* NGSPICE file created from nmos_10x10_flat.ext - technology: sky130A

.subckt nmos_10x10_flat
X0 S.t188 G D.t88 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1 D.t87 G S.t187 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 S.t186 G D.t50 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D.t131 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 S.t184 G D.t49 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 D.t78 G S.t183 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 S.t182 G D.t77 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 D.t58 G S.t181 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 S.t180 G D.t57 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 D.t90 G S.t179 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 S.t178 G D.t89 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 D.t130 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 D.t134 G S.t176 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D.t133 G S.t175 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 S.t174 G D.t60 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D.t59 G S.t173 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 S.t0 G D.t129 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 D.t62 G S.t171 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 S.t0 G D.t128 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 D.t61 G S.t169 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 D.t64 G S.t168 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 D.t63 G S.t167 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 D.t136 G S.t166 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 S.t165 G D.t135 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 S.t164 G D.t163 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 D.t162 G S.t163 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D.t142 G S.t162 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 S.t161 G D.t141 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D.t173 G S.t160 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 S.t159 G D.t172 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 S.t158 G D.t138 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 D.t137 G S.t157 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 S.t156 G D.t165 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 D.t164 G S.t155 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 S.t154 G D.t144 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 S.t153 G D.t143 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 D.t175 G S.t152 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 D.t174 G S.t151 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 D.t177 G S.t150 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 S.t149 G D.t176 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D.t179 G S.t148 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 S.t0 G D.t127 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 D.t178 G S.t146 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 S.t145 G D.t148 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 D.t147 G S.t144 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 S.t143 G D.t32 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 D.t31 G S.t142 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 D.t20 G S.t141 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 D.t19 G S.t140 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 S.t139 G D.t24 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 S.t138 G D.t23 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D.t85 G S.t137 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 S.t136 G D.t84 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 S.t135 G D.t154 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 D.t153 G S.t134 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 S.t133 G D.t152 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 D.t151 G S.t132 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 D.t126 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 S.t130 G D.t101 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D.t100 G S.t129 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 S.t128 G D.t103 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 S.t127 G D.t102 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 D.t105 G S.t126 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 D.t125 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 S.t124 G D.t104 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 D.t22 G S.t123 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 D.t21 G S.t122 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 S.t121 G D.t26 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 D.t25 G S.t120 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 D.t28 G S.t119 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 S.t118 G D.t27 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D.t92 G S.t117 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 D.t91 G S.t116 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 S.t115 G D.t66 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 D.t65 G S.t114 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 S.t113 G D.t80 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 S.t0 G D.t124 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 D.t79 G S.t111 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 S.t110 G D.t46 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 D.t123 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 S.t108 G D.t45 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 D.t94 G S.t107 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 S.t106 G D.t93 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 D.t12 G S.t105 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 S.t104 G D.t11 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 D.t8 G S.t103 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 S.t102 G D.t7 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 D.t52 G S.t101 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 D.t51 G S.t100 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 D.t54 G S.t99 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 S.t98 G D.t53 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 S.t97 G D.t70 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 S.t0 G D.t122 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 S.t95 G D.t69 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 S.t0 G D.t121 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 D.t96 G S.t93 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 S.t92 G D.t95 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 D.t98 G S.t91 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 S.t90 G D.t97 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 S.t89 G D.t82 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 D.t81 G S.t88 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 S.t87 G D.t48 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 D.t47 G S.t86 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 S.t85 G D.t56 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 D.t120 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 S.t83 G D.t55 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 D.t72 G S.t82 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 S.t81 G D.t71 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 D.t74 G S.t80 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 S.t79 G D.t73 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D.t30 G S.t78 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 S.t77 G D.t29 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t76 G D.t107 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 S.t75 G D.t106 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 D.t109 G S.t74 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 D.t108 G S.t73 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 S.t72 G D.t150 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 D.t119 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 S.t70 G D.t149 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 S.t0 G D.t118 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 D.t40 G S.t68 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 S.t67 G D.t39 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 D.t42 G S.t66 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 S.t65 G D.t41 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 S.t64 G D.t159 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 D.t158 G S.t63 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 S.t62 G D.t157 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 D.t156 G S.t61 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 S.t60 G D.t161 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 S.t0 G D.t117 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 S.t58 G D.t160 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 S.t57 G D.t169 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 D.t168 G S.t56 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t55 G D.t167 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 D.t166 G S.t54 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t53 G D.t171 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 D.t170 G S.t52 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 S.t51 G D.t146 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 S.t0 G D.t116 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 S.t49 G D.t145 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 S.t48 G D.t140 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 D.t139 G S.t47 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 D.t34 G S.t46 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 D.t33 G S.t45 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 S.t44 G D.t36 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 D.t35 G S.t43 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 D.t38 G S.t42 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 S.t41 G D.t37 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 D.t44 G S.t40 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 S.t39 G D.t43 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 D.t68 G S.t38 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 D.t67 G S.t37 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 S.t36 G D.t16 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 S.t35 G D.t15 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 D.t18 G S.t34 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 S.t33 G D.t17 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 S.t32 G D.t111 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 D.t110 G S.t31 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 D.t115 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 S.t29 G D.t14 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 D.t13 G S.t28 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 S.t27 G D.t1 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 D.t0 G S.t26 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 S.t24 G D.t112 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 D.t4 G S.t22 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 S.t20 G D.t2 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 D.t3 G S.t18 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 D.t10 G S.t16 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 D.t9 G S.t15 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 S.t14 G D.t132 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 D.t76 G S.t12 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 S.t0 G D.t114 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 D.t113 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 S.t8 G D.t83 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 S.t7 G D.t6 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 D.t99 G S.t6 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 S.t5 G D.t155 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 D.t5 G S.t4 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 D.t86 G S.t2 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 S.t1 G D.t75 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 D.n273 D.n272 41.943
R1 D.n272 D.n271 8.553
R2 D.n17 D.t140 4.386
R3 D.n21 D.t91 4.386
R4 D.n20 D.t84 4.386
R5 D.n3 D.t35 4.386
R6 D.n22 D.t51 4.386
R7 D.n23 D.t172 4.386
R8 D.n16 D.t122 4.386
R9 D.n15 D.t41 4.386
R10 D.n24 D.t162 4.386
R11 D.n25 D.t132 4.386
R12 D.n27 D.t85 4.386
R13 D.n26 D.t2 4.386
R14 D.n29 D.t31 4.386
R15 D.n28 D.t112 4.386
R16 D.n31 D.t147 4.386
R17 D.n30 D.t1 4.386
R18 D.n33 D.t179 4.386
R19 D.n32 D.t111 4.386
R20 D.n35 D.t120 4.386
R21 D.n34 D.t127 4.386
R22 D.n14 D.t146 4.386
R23 D.n36 D.t20 4.386
R24 D.n37 D.t107 4.386
R25 D.n38 D.t76 4.386
R26 D.n39 D.t71 4.386
R27 D.n40 D.t3 4.386
R28 D.n41 D.t56 4.386
R29 D.n42 D.t126 4.386
R30 D.n43 D.t114 4.386
R31 D.n45 D.t64 4.386
R32 D.n44 D.t23 4.386
R33 D.n47 D.t74 4.386
R34 D.n46 D.t32 4.386
R35 D.n49 D.t72 4.386
R36 D.n48 D.t148 4.386
R37 D.n51 D.t47 4.386
R38 D.n50 D.t176 4.386
R39 D.n53 D.t81 4.386
R40 D.n52 D.t143 4.386
R41 D.n55 D.t96 4.386
R42 D.n54 D.t165 4.386
R43 D.n57 D.t54 4.386
R44 D.n56 D.t138 4.386
R45 D.n58 D.t115 4.386
R46 D.n59 D.t121 4.386
R47 D.n61 D.t4 4.386
R48 D.n60 D.t48 4.386
R49 D.n63 D.t0 4.386
R50 D.n62 D.t82 4.386
R51 D.n13 D.t38 4.386
R52 D.n65 D.t44 4.386
R53 D.n64 D.t11 4.386
R54 D.n67 D.t67 4.386
R55 D.n66 D.t7 4.386
R56 D.n69 D.t110 4.386
R57 D.n68 D.t53 4.386
R58 D.n71 D.t13 4.386
R59 D.n70 D.t95 4.386
R60 D.n73 D.t177 4.386
R61 D.n72 D.t15 4.386
R62 D.n75 D.t175 4.386
R63 D.n74 D.t16 4.386
R64 D.n12 D.t142 4.386
R65 D.n77 D.t173 4.386
R66 D.n76 D.t36 4.386
R67 D.n79 D.t164 4.386
R68 D.n78 D.t43 4.386
R69 D.n2 D.t8 4.386
R70 D.n80 D.t52 4.386
R71 D.n81 D.t141 4.386
R72 D.n19 D.t118 4.386
R73 D.n18 D.t131 4.386
R74 D.n261 D.t17 4.327
R75 D.n260 D.t123 4.327
R76 D.n85 D.t116 4.327
R77 D.n232 D.t103 4.327
R78 D.n231 D.t108 4.327
R79 D.n88 D.t128 4.327
R80 D.n319 D.t160 4.327
R81 D.n318 D.t174 4.327
R82 D.n325 D.t60 4.327
R83 D.n324 D.t65 4.327
R84 D.n329 D.t89 4.327
R85 D.n328 D.t92 4.327
R86 D.n333 D.t57 4.327
R87 D.n332 D.t25 4.327
R88 D.n337 D.t49 4.327
R89 D.n336 D.t125 4.327
R90 D.n341 D.t88 4.327
R91 D.n340 D.t170 4.327
R92 D.n84 D.t124 4.327
R93 D.n286 D.t145 4.327
R94 D.n285 D.t28 4.327
R95 D.n291 D.t171 4.327
R96 D.n290 D.t59 4.327
R97 D.n295 D.t167 4.327
R98 D.n294 D.t130 4.327
R99 D.n299 D.t161 4.327
R100 D.n298 D.t79 4.327
R101 D.n86 D.t129 4.327
R102 D.n96 D.t97 4.327
R103 D.n95 D.t63 4.327
R104 D.n100 D.t66 4.327
R105 D.n99 D.t166 4.327
R106 D.n104 D.t27 4.327
R107 D.n103 D.t168 4.327
R108 D.n108 D.t26 4.327
R109 D.n107 D.t156 4.327
R110 D.n112 D.t104 4.327
R111 D.n111 D.t158 4.327
R112 D.n116 D.t102 4.327
R113 D.n115 D.t40 4.327
R114 D.n120 D.t101 4.327
R115 D.n119 D.t119 4.327
R116 D.n128 D.t152 4.327
R117 D.n127 D.t134 4.327
R118 D.n11 D.t133 4.327
R119 D.n163 D.t169 4.327
R120 D.n162 D.t90 4.327
R121 D.n167 D.t157 4.327
R122 D.n166 D.t58 4.327
R123 D.n191 D.t106 4.327
R124 D.n190 D.t99 4.327
R125 D.n185 D.t149 4.327
R126 D.n184 D.t86 4.327
R127 D.n179 D.t39 4.327
R128 D.n178 D.t87 4.327
R129 D.n173 D.t159 4.327
R130 D.n172 D.t78 4.327
R131 D.n10 D.t21 4.327
R132 D.n204 D.t77 4.327
R133 D.n203 D.t22 4.327
R134 D.n208 D.t50 4.327
R135 D.n207 D.t105 4.327
R136 D.n220 D.t155 4.327
R137 D.n219 D.t151 4.327
R138 D.n214 D.t75 4.327
R139 D.n213 D.t100 4.327
R140 D.n235 D.t154 4.327
R141 D.n234 D.t109 4.327
R142 D.n9 D.t42 4.327
R143 D.n8 D.t5 4.327
R144 D.n273 D.t80 4.327
R145 D.n274 D.t61 4.327
R146 D.n7 D.t37 4.091
R147 D.n89 D.t18 4.091
R148 D.n6 D.t45 4.091
R149 D.n87 D.t163 4.091
R150 D.n11 D.t9 4.091
R151 D.n10 D.t178 4.091
R152 D.n9 D.t144 4.091
R153 D.n8 D.t93 4.091
R154 D.n90 D.t117 4.084
R155 D.n17 D.t46 4.083
R156 D.n3 D.t29 4.083
R157 D.n16 D.t150 4.083
R158 D.n15 D.t6 4.083
R159 D.n14 D.t135 4.083
R160 D.n93 D.t139 4.083
R161 D.n13 D.t73 4.083
R162 D.n12 D.t83 4.083
R163 D.n2 D.t24 4.083
R164 D.n93 D.t70 4.06
R165 D.n90 D.t136 4.06
R166 D.n275 D.t137 4.057
R167 D.n253 D.t69 4.057
R168 D.n344 D.t34 4.057
R169 D.n308 D.t12 4.057
R170 D.n160 D.t55 4.057
R171 D.n201 D.t14 4.057
R172 D.n229 D.t98 4.057
R173 D.n243 D.t68 4.057
R174 D.n267 D.t94 4.031
R175 D.n241 D.t10 4.031
R176 D.n254 D.t33 4.031
R177 D.n321 D.t62 4.031
R178 D.n281 D.t153 4.031
R179 D.n152 D.t113 4.031
R180 D.n198 D.t19 4.031
R181 D.n228 D.t30 4.031
R182 D.n239 D.n237 0.345
R183 D.n255 D.n16 0.24
R184 D.n227 D.n226 0.225
R185 D.n159 D.n158 0.225
R186 D.n200 D.n199 0.225
R187 D.n239 D.n238 0.225
R188 D.n233 D.n9 0.203
R189 D.n251 D.n250 0.184
R190 D.n131 D.n129 0.174
R191 D.n131 D.n130 0.156
R192 D.n5 D.n89 0.152
R193 D.n91 D.n304 0.156
R194 D.n89 D.n248 0.143
R195 D.n6 D.n312 0.143
R196 D.n87 D.n309 0.143
R197 D.n87 D.n277 0.143
R198 D.n7 D.n257 0.143
R199 D.n59 D.n132 0.143
R200 D.n244 D.n3 0.143
R201 D.n252 D.n249 0.133
R202 D.n157 D.n156 0.125
R203 D.n25 D.n15 0.123
R204 D.n310 D.n87 0.122
R205 D.n21 D.n17 0.122
R206 D.n45 D.n93 0.122
R207 D.n244 D.n2 0.114
R208 D.n307 D.n301 0.113
R209 D.n245 D.n12 0.111
R210 D.n246 D.n13 0.111
R211 D.n4 D.n0 0.216
R212 D.n5 D.n1 0.216
R213 D.n0 D.n6 0.1
R214 D.n1 D.n7 0.1
R215 D.n157 D.n155 0.092
R216 D.n142 D.n141 0.092
R217 D.n90 D.n149 0.091
R218 D.n247 D.n150 0.085
R219 D.n266 D.n265 0.083
R220 D.n3 D.n8 0.079
R221 D.n61 D.n11 0.078
R222 D.n73 D.n10 0.078
R223 D.n138 D.n137 0.075
R224 D.n92 D.n123 0.075
R225 D.n317 D.n316 0.075
R226 D.n288 D.n284 0.075
R227 D.n148 D.n83 0.072
R228 D.n292 D.n288 0.072
R229 D.n296 D.n292 0.072
R230 D.n300 D.n296 0.072
R231 D.n237 D.n233 0.072
R232 D.n155 D.n154 0.064
R233 D.n142 D.n138 0.064
R234 D.n150 D.n90 0.061
R235 D.n90 D.n144 0.06
R236 D.n347 D.n346 0.058
R237 D.n16 D.n254 0.055
R238 D.n144 D.n142 0.055
R239 D.n155 D.n153 0.055
R240 D.n82 D.n221 0.055
R241 D.n252 D.n251 0.053
R242 D.n270 D.n269 0.053
R243 D.n82 D.n222 0.053
R244 D.n35 D.n33 0.053
R245 D.n19 D.n21 0.053
R246 D.n122 D.n121 0.053
R247 D.n343 D.n342 0.053
R248 D.n301 D.n300 0.053
R249 D.n280 D.n278 0.052
R250 D.n146 D.n145 0.052
R251 D.n21 D.n260 0.052
R252 D.n21 D.n261 0.052
R253 D.n23 D.n231 0.052
R254 D.n23 D.n232 0.052
R255 D.n25 D.n319 0.052
R256 D.n25 D.n318 0.052
R257 D.n27 D.n324 0.052
R258 D.n27 D.n325 0.052
R259 D.n29 D.n328 0.052
R260 D.n29 D.n329 0.052
R261 D.n31 D.n332 0.052
R262 D.n31 D.n333 0.052
R263 D.n33 D.n336 0.052
R264 D.n33 D.n337 0.052
R265 D.n35 D.n340 0.052
R266 D.n35 D.n341 0.052
R267 D.n37 D.n286 0.052
R268 D.n37 D.n285 0.052
R269 D.n39 D.n290 0.052
R270 D.n39 D.n291 0.052
R271 D.n41 D.n294 0.052
R272 D.n41 D.n295 0.052
R273 D.n43 D.n298 0.052
R274 D.n43 D.n299 0.052
R275 D.n45 D.n95 0.052
R276 D.n45 D.n96 0.052
R277 D.n47 D.n99 0.052
R278 D.n47 D.n100 0.052
R279 D.n49 D.n103 0.052
R280 D.n49 D.n104 0.052
R281 D.n51 D.n107 0.052
R282 D.n51 D.n108 0.052
R283 D.n53 D.n111 0.052
R284 D.n53 D.n112 0.052
R285 D.n55 D.n115 0.052
R286 D.n55 D.n116 0.052
R287 D.n57 D.n119 0.052
R288 D.n57 D.n120 0.052
R289 D.n59 D.n128 0.052
R290 D.n59 D.n127 0.052
R291 D.n61 D.n162 0.052
R292 D.n61 D.n163 0.052
R293 D.n63 D.n166 0.052
R294 D.n63 D.n167 0.052
R295 D.n65 D.n190 0.052
R296 D.n65 D.n191 0.052
R297 D.n67 D.n184 0.052
R298 D.n67 D.n185 0.052
R299 D.n69 D.n178 0.052
R300 D.n69 D.n179 0.052
R301 D.n71 D.n172 0.052
R302 D.n71 D.n173 0.052
R303 D.n73 D.n203 0.052
R304 D.n73 D.n204 0.052
R305 D.n75 D.n207 0.052
R306 D.n75 D.n208 0.052
R307 D.n77 D.n219 0.052
R308 D.n77 D.n220 0.052
R309 D.n79 D.n213 0.052
R310 D.n79 D.n214 0.052
R311 D.n81 D.n235 0.052
R312 D.n81 D.n234 0.052
R313 D.n19 D.n273 0.052
R314 D.n19 D.n274 0.052
R315 D.n17 D.n267 0.051
R316 D.n3 D.n241 0.051
R317 D.n15 D.n321 0.051
R318 D.n14 D.n281 0.051
R319 D.n13 D.n152 0.051
R320 D.n12 D.n198 0.051
R321 D.n2 D.n228 0.051
R322 D.n140 D.n139 0.051
R323 D.n141 D.n140 0.051
R324 D.n158 D.n157 0.051
R325 D.n144 D.n143 0.049
R326 D.n27 D.n25 0.049
R327 D.n33 D.n31 0.049
R328 D.n31 D.n29 0.049
R329 D.n29 D.n27 0.049
R330 D.n59 D.n57 0.049
R331 D.n57 D.n55 0.049
R332 D.n55 D.n53 0.049
R333 D.n53 D.n51 0.049
R334 D.n51 D.n49 0.049
R335 D.n49 D.n47 0.049
R336 D.n47 D.n45 0.049
R337 D.n65 D.n67 0.049
R338 D.n67 D.n69 0.049
R339 D.n69 D.n71 0.049
R340 D.n71 D.n63 0.049
R341 D.n63 D.n61 0.049
R342 D.n77 D.n79 0.049
R343 D.n79 D.n75 0.049
R344 D.n75 D.n73 0.049
R345 D.n13 D.n65 0.046
R346 D.n12 D.n77 0.046
R347 D.n6 D.n35 0.046
R348 D.n90 D.n59 0.045
R349 D.n303 D.n302 0.045
R350 D.n7 D.n19 0.045
R351 D D.n247 0.044
R352 D.n63 D.n170 0.042
R353 D.n71 D.n176 0.042
R354 D.n69 D.n182 0.042
R355 D.n67 D.n188 0.042
R356 D.n65 D.n194 0.042
R357 D.n75 D.n211 0.042
R358 D.n79 D.n217 0.042
R359 D.n77 D.n225 0.042
R360 D.n306 D.n305 0.039
R361 D.n59 D.n131 0.039
R362 D.n59 D.n125 0.039
R363 D.n6 D.n345 0.035
R364 D.n7 D.n276 0.035
R365 D.n89 D.n255 0.035
R366 D.n7 D.n275 0.034
R367 D.n89 D.n253 0.034
R368 D.n6 D.n344 0.034
R369 D.n87 D.n308 0.034
R370 D.n136 D.n135 0.034
R371 D D.n347 0.032
R372 D.n245 D.n244 0.031
R373 D.n246 D.n245 0.031
R374 D.n247 D.n246 0.031
R375 D.n4 D.n310 0.029
R376 D.n265 D.n264 0.029
R377 D.n316 D.n315 0.029
R378 D.n284 D.n283 0.029
R379 D.n316 D.n313 0.028
R380 D.n265 D.n263 0.028
R381 D.n89 D.n252 0.027
R382 D.n87 D.n307 0.027
R383 D.n59 D.n126 0.027
R384 D.n138 D.n133 0.026
R385 D.n315 D.n314 0.025
R386 D.n283 D.n282 0.025
R387 D.n263 D.n262 0.025
R388 D.n149 D.n148 0.024
R389 D.n305 D.n91 0.024
R390 D.n125 D.n92 0.023
R391 D.n91 D.n303 0.023
R392 D.n13 D.n196 0.023
R393 D.n63 D.n169 0.023
R394 D.n71 D.n175 0.023
R395 D.n69 D.n181 0.023
R396 D.n67 D.n187 0.023
R397 D.n65 D.n193 0.023
R398 D.n75 D.n210 0.023
R399 D.n79 D.n216 0.023
R400 D.n77 D.n224 0.023
R401 D.n284 D.n280 0.02
R402 D.n13 D.n151 0.019
R403 D.n3 D.n242 0.016
R404 D.n81 D.n236 0.016
R405 D.n65 D.n189 0.016
R406 D.n67 D.n183 0.016
R407 D.n69 D.n177 0.016
R408 D.n71 D.n171 0.016
R409 D.n77 D.n218 0.016
R410 D.n79 D.n212 0.016
R411 D.n12 D.n200 0.016
R412 D.n2 D.n239 0.016
R413 D.n92 D.n124 0.041
R414 D.n279 D.n14 0.04
R415 D.n11 D.n160 0.038
R416 D.n10 D.n201 0.038
R417 D.n9 D.n229 0.038
R418 D.n8 D.n243 0.038
R419 D.n310 D.n5 0.034
R420 D.n347 D.n4 0.033
R421 D.n77 D.n82 0.028
R422 D.n2 D.n227 0.021
R423 D.n3 D.n240 0.02
R424 D.n13 D.n159 0.02
R425 D.n1 D.n256 0.019
R426 D.n0 D.n311 0.019
R427 D.n83 D.n146 0.016
R428 D.n12 D.n197 0.015
R429 D.n169 D.n168 0.013
R430 D.n175 D.n174 0.013
R431 D.n181 D.n180 0.013
R432 D.n187 D.n186 0.013
R433 D.n193 D.n192 0.013
R434 D.n196 D.n195 0.013
R435 D.n210 D.n209 0.013
R436 D.n216 D.n215 0.013
R437 D.n224 D.n223 0.013
R438 D.n307 D.n306 0.012
R439 D.n45 D.n97 0.011
R440 D.n21 D.n266 0.011
R441 D.n27 D.n326 0.011
R442 D.n29 D.n330 0.011
R443 D.n31 D.n334 0.011
R444 D.n33 D.n338 0.011
R445 D.n35 D.n343 0.011
R446 D.n292 D.n39 0.011
R447 D.n296 D.n41 0.011
R448 D.n300 D.n43 0.011
R449 D.n47 D.n101 0.011
R450 D.n49 D.n105 0.011
R451 D.n51 D.n109 0.011
R452 D.n53 D.n113 0.011
R453 D.n55 D.n117 0.011
R454 D.n57 D.n122 0.011
R455 D.n233 D.n23 0.011
R456 D.n137 D.n136 0.01
R457 D.n237 D.n81 0.01
R458 D.n19 D.n270 0.01
R459 D.n135 D.n134 0.01
R460 D.n61 D.n164 0.01
R461 D.n73 D.n205 0.01
R462 D.n25 D.n320 0.009
R463 D.n37 D.n287 0.009
R464 D.n280 D.n279 0.008
R465 D.n25 D.n317 0.008
R466 D.n288 D.n37 0.008
R467 D.n45 D.n94 0.006
R468 D.n21 D.n259 0.006
R469 D.n83 D.n147 0.015
R470 D.n17 D.n268 0.015
R471 D.n15 D.n322 0.015
R472 D.n7 D.n85 0.01
R473 D.n6 D.n84 0.01
R474 D.n79 D.n78 0.009
R475 D.n77 D.n76 0.009
R476 D.n75 D.n74 0.009
R477 D.n73 D.n72 0.009
R478 D.n71 D.n70 0.009
R479 D.n69 D.n68 0.009
R480 D.n67 D.n66 0.009
R481 D.n65 D.n64 0.009
R482 D.n63 D.n62 0.009
R483 D.n61 D.n60 0.009
R484 D.n59 D.n58 0.009
R485 D.n57 D.n56 0.009
R486 D.n55 D.n54 0.009
R487 D.n53 D.n52 0.009
R488 D.n51 D.n50 0.009
R489 D.n49 D.n48 0.009
R490 D.n47 D.n46 0.009
R491 D.n45 D.n44 0.009
R492 D.n33 D.n32 0.009
R493 D.n31 D.n30 0.009
R494 D.n29 D.n28 0.009
R495 D.n27 D.n26 0.009
R496 D.n25 D.n24 0.009
R497 D.n21 D.n20 0.009
R498 D.n35 D.n34 0.008
R499 D.n19 D.n18 0.008
R500 D.n81 D.n80 0.007
R501 D.n43 D.n42 0.007
R502 D.n41 D.n40 0.007
R503 D.n39 D.n38 0.007
R504 D.n37 D.n36 0.007
R505 D.n23 D.n22 0.007
R506 D.n61 D.n161 0.006
R507 D.n73 D.n202 0.006
R508 D.n89 D.n88 0.006
R509 D.n87 D.n86 0.006
R510 D.n23 D.n230 0.006
R511 D.n35 D.n339 0.006
R512 D.n33 D.n335 0.006
R513 D.n31 D.n331 0.006
R514 D.n29 D.n327 0.006
R515 D.n27 D.n323 0.006
R516 D.n43 D.n297 0.006
R517 D.n41 D.n293 0.006
R518 D.n39 D.n289 0.006
R519 D.n57 D.n118 0.006
R520 D.n55 D.n114 0.006
R521 D.n53 D.n110 0.006
R522 D.n51 D.n106 0.006
R523 D.n49 D.n102 0.006
R524 D.n47 D.n98 0.006
R525 D.n63 D.n165 0.006
R526 D.n75 D.n206 0.006
R527 D.n19 D.n258 0.006
R528 S.n533 S.n532 91.519
R529 S.n754 S.n753 91.519
R530 S.n159 S.n158 91.519
R531 S.n358 S.n357 91.519
R532 S.n659 S.n658 91.519
R533 S.n264 S.n263 91.519
R534 S.n450 S.n449 91.519
R535 S.n557 S.n556 87.091
R536 S.n31 S.n30 87.091
R537 S.n61 S.n60 87.091
R538 S.n42 S.n41 87.091
R539 S.n52 S.n51 87.091
R540 S.n549 S.n548 87.091
R541 S.n553 S.n552 87.091
R542 S.n544 S.n543 87.091
R543 S.n470 S.t99 3.773
R544 S.n470 S.n469 3.773
R545 S.n472 S.n471 3.773
R546 S.n472 S.t32 3.773
R547 S.n541 S.t34 3.773
R548 S.n540 S.t45 3.773
R549 S.n533 S.t116 3.773
R550 S.n461 S.t72 3.773
R551 S.n512 S.t107 3.773
R552 S.n557 S.t111 3.773
R553 S.n554 S.t41 3.773
R554 S.n555 S.t105 3.773
R555 S.n480 S.n479 3.773
R556 S.n480 S.t136 3.773
R557 S.n491 S.t18 3.773
R558 S.n491 S.n490 3.773
R559 S.n488 S.t173 3.773
R560 S.n488 S.n487 3.773
R561 S.n483 S.n482 3.773
R562 S.n483 S.t113 3.773
R563 S.n685 S.n684 3.773
R564 S.n685 S.t48 3.773
R565 S.n703 S.t12 3.773
R566 S.n703 S.n702 3.773
R567 S.n700 S.t119 3.773
R568 S.n700 S.n699 3.773
R569 S.n688 S.n687 3.773
R570 S.n688 S.t33 3.773
R571 S.n754 S.t141 3.773
R572 S.n756 S.t134 3.773
R573 S.n758 S.t110 3.773
R574 S.n159 S.t161 3.773
R575 S.n160 S.t16 3.773
R576 S.n152 S.t139 3.773
R577 S.n243 S.n242 3.773
R578 S.n243 S.t159 3.773
R579 S.n258 S.t43 3.773
R580 S.n258 S.n257 3.773
R581 S.n261 S.t4 3.773
R582 S.n261 S.n260 3.773
R583 S.n246 S.n245 3.773
R584 S.n246 S.t135 3.773
R585 S.n31 S.t128 3.773
R586 S.n28 S.t154 3.773
R587 S.n29 S.t38 3.773
R588 S.n61 S.t90 3.773
R589 S.n57 S.t97 3.773
R590 S.n58 S.t15 3.773
R591 S.n141 S.n140 3.773
R592 S.n141 S.t138 3.773
R593 S.n231 S.t22 3.773
R594 S.n231 S.n230 3.773
R595 S.n228 S.t175 3.773
R596 S.n228 S.n227 3.773
R597 S.n144 S.n143 3.773
R598 S.n144 S.t115 3.773
R599 S.n309 S.n308 3.773
R600 S.n309 S.t145 3.773
R601 S.n326 S.t28 3.773
R602 S.n326 S.n325 3.773
R603 S.n323 S.t181 3.773
R604 S.n323 S.n322 3.773
R605 S.n306 S.n305 3.773
R606 S.n306 S.t121 3.773
R607 S.n499 S.n498 3.773
R608 S.n499 S.t158 3.773
R609 S.n507 S.t42 3.773
R610 S.n507 S.n506 3.773
R611 S.n510 S.t6 3.773
R612 S.n510 S.n509 3.773
R613 S.n496 S.n495 3.773
R614 S.n496 S.t133 3.773
R615 S.n668 S.n667 3.773
R616 S.n668 S.t156 3.773
R617 S.n679 S.t40 3.773
R618 S.n679 S.n678 3.773
R619 S.n676 S.t2 3.773
R620 S.n676 S.n675 3.773
R621 S.n665 S.n664 3.773
R622 S.n665 S.t130 3.773
R623 S.n577 S.n576 3.773
R624 S.n577 S.t153 3.773
R625 S.n594 S.t37 3.773
R626 S.n594 S.n593 3.773
R627 S.n591 S.t187 3.773
R628 S.n591 S.n590 3.773
R629 S.n574 S.n573 3.773
R630 S.n574 S.t127 3.773
R631 S.n386 S.n385 3.773
R632 S.n386 S.t149 3.773
R633 S.n395 S.t31 3.773
R634 S.n395 S.n394 3.773
R635 S.n392 S.t183 3.773
R636 S.n392 S.n391 3.773
R637 S.n383 S.n382 3.773
R638 S.n383 S.t124 3.773
R639 S.n150 S.n149 3.773
R640 S.n150 S.t143 3.773
R641 S.n215 S.t26 3.773
R642 S.n215 S.n214 3.773
R643 S.n218 S.t179 3.773
R644 S.n218 S.n217 3.773
R645 S.n221 S.n220 3.773
R646 S.n221 S.t118 3.773
R647 S.n42 S.t182 3.773
R648 S.n39 S.t29 3.773
R649 S.n40 S.t91 3.773
R650 S.n86 S.n85 3.773
R651 S.n86 S.t35 3.773
R652 S.n103 S.t100 3.773
R653 S.n103 S.n102 3.773
R654 S.n100 S.t66 3.773
R655 S.n100 S.n99 3.773
R656 S.n89 S.n88 3.773
R657 S.n89 S.t186 3.773
R658 S.n165 S.n164 3.773
R659 S.n165 S.t36 3.773
R660 S.n178 S.t101 3.773
R661 S.n178 S.n177 3.773
R662 S.n175 S.t73 3.773
R663 S.n175 S.n174 3.773
R664 S.n168 S.n167 3.773
R665 S.n168 S.t1 3.773
R666 S.n334 S.n333 3.773
R667 S.n334 S.t39 3.773
R668 S.n343 S.t103 3.773
R669 S.n343 S.n342 3.773
R670 S.n346 S.t74 3.773
R671 S.n346 S.n345 3.773
R672 S.n337 S.n336 3.773
R673 S.n337 S.t5 3.773
R674 S.n358 S.t44 3.773
R675 S.n359 S.t78 3.773
R676 S.n352 S.t8 3.773
R677 S.n187 S.n186 3.773
R678 S.n187 S.t89 3.773
R679 S.n195 S.t152 3.773
R680 S.n195 S.n194 3.773
R681 S.n192 S.t123 3.773
R682 S.n192 S.n191 3.773
R683 S.n184 S.n183 3.773
R684 S.n184 S.t64 3.773
R685 S.n289 S.n288 3.773
R686 S.n289 S.t92 3.773
R687 S.n301 S.t155 3.773
R688 S.n301 S.n300 3.773
R689 S.n298 S.t126 3.773
R690 S.n298 S.n297 3.773
R691 S.n292 S.n291 3.773
R692 S.n292 S.t67 3.773
R693 S.n365 S.n364 3.773
R694 S.n365 S.t98 3.773
R695 S.n378 S.t160 3.773
R696 S.n378 S.n377 3.773
R697 S.n375 S.t129 3.773
R698 S.n375 S.n374 3.773
R699 S.n368 S.n367 3.773
R700 S.n368 S.t70 3.773
R701 S.n607 S.n606 3.773
R702 S.n607 S.t102 3.773
R703 S.n616 S.t162 3.773
R704 S.n616 S.n615 3.773
R705 S.n619 S.t132 3.773
R706 S.n619 S.n618 3.773
R707 S.n610 S.n609 3.773
R708 S.n610 S.t75 3.773
R709 S.n659 S.t104 3.773
R710 S.n660 S.t140 3.773
R711 S.n650 S.t79 3.773
R712 S.n52 S.t57 3.773
R713 S.n47 S.t83 3.773
R714 S.n48 S.t146 3.773
R715 S.n113 S.n112 3.773
R716 S.n113 S.t87 3.773
R717 S.n131 S.t150 3.773
R718 S.n131 S.n130 3.773
R719 S.n128 S.t122 3.773
R720 S.n128 S.n127 3.773
R721 S.n116 S.n115 3.773
R722 S.n116 S.t62 3.773
R723 S.n16 S.t106 3.773
R724 S.n0 S.t77 3.773
R725 S.n264 S.t168 3.773
R726 S.n266 S.t47 3.773
R727 S.n268 S.t7 3.773
R728 S.n200 S.n199 3.773
R729 S.n200 S.t65 3.773
R730 S.n209 S.t80 3.773
R731 S.n209 S.n208 3.773
R732 S.n212 S.t167 3.773
R733 S.n212 S.n211 3.773
R734 S.n203 S.n202 3.773
R735 S.n203 S.t58 3.773
R736 S.n435 S.n434 3.773
R737 S.n435 S.t14 3.773
R738 S.n444 S.t82 3.773
R739 S.n444 S.n443 3.773
R740 S.n447 S.t54 3.773
R741 S.n447 S.n446 3.773
R742 S.n438 S.n437 3.773
R743 S.n438 S.t174 3.773
R744 S.n350 S.n349 3.773
R745 S.n350 S.t20 3.773
R746 S.n421 S.t86 3.773
R747 S.n421 S.n420 3.773
R748 S.n424 S.t56 3.773
R749 S.n424 S.n423 3.773
R750 S.n427 S.n426 3.773
R751 S.n427 S.t178 3.773
R752 S.n624 S.n623 3.773
R753 S.n624 S.t24 3.773
R754 S.n636 S.t88 3.773
R755 S.n636 S.n635 3.773
R756 S.n639 S.t61 3.773
R757 S.n639 S.n638 3.773
R758 S.n627 S.n626 3.773
R759 S.n627 S.t180 3.773
R760 S.n707 S.n706 3.773
R761 S.n707 S.t27 3.773
R762 S.n717 S.t93 3.773
R763 S.n717 S.n716 3.773
R764 S.n720 S.t63 3.773
R765 S.n720 S.n719 3.773
R766 S.n710 S.n709 3.773
R767 S.n710 S.t184 3.773
R768 S.n549 S.t176 3.773
R769 S.n546 S.t108 3.773
R770 S.n547 S.t166 3.773
R771 S.n450 S.t163 3.773
R772 S.n452 S.t171 3.773
R773 S.n454 S.t165 3.773
R774 S.n398 S.n397 3.773
R775 S.n398 S.t51 3.773
R776 S.n415 S.t137 3.773
R777 S.n415 S.n414 3.773
R778 S.n418 S.t151 3.773
R779 S.n418 S.n417 3.773
R780 S.n401 S.n400 3.773
R781 S.n401 S.t49 3.773
R782 S.n739 S.n738 3.773
R783 S.n739 S.t76 3.773
R784 S.n748 S.t142 3.773
R785 S.n748 S.n747 3.773
R786 S.n751 S.t114 3.773
R787 S.n751 S.n750 3.773
R788 S.n742 S.n741 3.773
R789 S.n742 S.t53 3.773
R790 S.n553 S.t52 3.773
R791 S.n550 S.t164 3.773
R792 S.n551 S.t46 3.773
R793 S.n519 S.n518 3.773
R794 S.n519 S.t85 3.773
R795 S.n527 S.t148 3.773
R796 S.n527 S.n526 3.773
R797 S.n530 S.t120 3.773
R798 S.n530 S.n529 3.773
R799 S.n522 S.n521 3.773
R800 S.n522 S.t60 3.773
R801 S.n648 S.n647 3.773
R802 S.n648 S.t81 3.773
R803 S.n723 S.t144 3.773
R804 S.n723 S.n722 3.773
R805 S.n726 S.t117 3.773
R806 S.n726 S.n725 3.773
R807 S.n729 S.n728 3.773
R808 S.n729 S.t55 3.773
R809 S.n544 S.t169 3.773
R810 S.n545 S.t95 3.773
R811 S.n542 S.t157 3.773
R812 S.n463 S.t68 3.773
R813 S.n463 S.n462 3.773
R814 S.n535 S.n534 3.773
R815 S.n535 S.t188 3.773
R816 S.n272 S.n271 0.172
R817 S.n5 S.n2 0.164
R818 S.n560 S.n559 0.143
R819 S.n340 S.n339 0.133
R820 S.n613 S.n612 0.133
R821 S.n295 S.n294 0.133
R822 S.n441 S.n440 0.133
R823 S.n66 S.n62 0.123
R824 S.n777 S.n460 0.114
R825 S.n778 S.n277 0.111
R826 S.n776 S.n775 0.11
R827 S.n560 S.n539 0.11
R828 S.n696 S.n691 0.106
R829 S.n768 S.n767 0.095
R830 S.n653 S.n652 0.093
R831 S.n694 S.n693 0.07
R832 S.n55 S.n53 0.067
R833 S.n55 S.n54 0.067
R834 S.n36 S.n34 0.067
R835 S.n45 S.n43 0.067
R836 S.n45 S.n44 0.067
R837 S.n36 S.n35 0.067
R838 S.n25 S.n24 0.067
R839 S.n25 S.n23 0.067
R840 S.n274 S.n273 0.067
R841 S.n274 S.n270 0.067
R842 S.n12 S.n11 0.067
R843 S.n98 S.n97 0.066
R844 S.n276 S.n275 0.065
R845 S.n225 S.n224 0.064
R846 S.n458 S.n457 0.063
R847 S.n321 S.n320 0.063
R848 S.n589 S.n588 0.063
R849 S.n674 S.n673 0.063
R850 S.n226 S.n134 0.063
R851 S.n296 S.n283 0.063
R852 S.n126 S.n107 0.063
R853 S.n256 S.n255 0.063
R854 S.n56 S.n55 0.062
R855 S.n46 S.n45 0.062
R856 S.n37 S.n36 0.061
R857 S.n597 S.n596 0.059
R858 S.n412 S.n411 0.059
R859 S.n26 S.n25 0.059
R860 S.n276 S.n274 0.058
R861 S S.n778 0.056
R862 S.n15 S.n0 0.055
R863 S.n536 S.n461 0.054
R864 S.n157 S.n152 0.054
R865 S.n356 S.n352 0.054
R866 S.n657 S.n650 0.054
R867 S.n757 S.n756 0.054
R868 S.n267 S.n266 0.054
R869 S.n453 S.n452 0.054
R870 S.n489 S.n488 0.053
R871 S.n701 S.n700 0.053
R872 S.n262 S.n261 0.053
R873 S.n229 S.n228 0.053
R874 S.n324 S.n323 0.053
R875 S.n511 S.n510 0.053
R876 S.n677 S.n676 0.053
R877 S.n592 S.n591 0.053
R878 S.n393 S.n392 0.053
R879 S.n219 S.n218 0.053
R880 S.n101 S.n100 0.053
R881 S.n176 S.n175 0.053
R882 S.n347 S.n346 0.053
R883 S.n193 S.n192 0.053
R884 S.n299 S.n298 0.053
R885 S.n376 S.n375 0.053
R886 S.n620 S.n619 0.053
R887 S.n129 S.n128 0.053
R888 S.n213 S.n212 0.053
R889 S.n448 S.n447 0.053
R890 S.n425 S.n424 0.053
R891 S.n640 S.n639 0.053
R892 S.n721 S.n720 0.053
R893 S.n419 S.n418 0.053
R894 S.n752 S.n751 0.053
R895 S.n531 S.n530 0.053
R896 S.n727 S.n726 0.053
R897 S.n281 S.n280 0.052
R898 S.n773 S.n772 0.052
R899 S.n693 S.n692 0.052
R900 S.n558 S.n540 0.052
R901 S.t17 S.n535 0.051
R902 S.t17 S.n463 0.051
R903 S.n235 S.n234 0.051
R904 S S.n66 0.051
R905 S.n614 S.n600 0.05
R906 S.n256 S.n237 0.05
R907 S.n137 S.n136 0.05
R908 S.n486 S.n484 0.047
R909 S.n698 S.n689 0.047
R910 S.n775 S.n759 0.047
R911 S.n256 S.n247 0.047
R912 S.n226 S.n145 0.047
R913 S.n321 S.n307 0.047
R914 S.n505 S.n497 0.047
R915 S.n674 S.n666 0.047
R916 S.n589 S.n575 0.047
R917 S.n390 S.n384 0.047
R918 S.n223 S.n222 0.047
R919 S.n98 S.n90 0.047
R920 S.n173 S.n169 0.047
R921 S.n341 S.n338 0.047
R922 S.n190 S.n185 0.047
R923 S.n296 S.n293 0.047
R924 S.n373 S.n369 0.047
R925 S.n614 S.n611 0.047
R926 S.n126 S.n117 0.047
R927 S.n277 S.n269 0.047
R928 S.n207 S.n204 0.047
R929 S.n442 S.n439 0.047
R930 S.n432 S.n428 0.047
R931 S.n634 S.n628 0.047
R932 S.n715 S.n711 0.047
R933 S.n459 S.n455 0.047
R934 S.n413 S.n402 0.047
R935 S.n746 S.n743 0.047
R936 S.n525 S.n523 0.047
R937 S.n732 S.n730 0.047
R938 S.n33 S.n32 0.046
R939 S.t3 S.n27 0.046
R940 S.n442 S.n432 0.046
R941 S.n19 S.n17 0.045
R942 S.n745 S.n744 0.045
R943 S.n82 S.n81 0.045
R944 S.n746 S.n732 0.045
R945 S.n634 S.n621 0.044
R946 S.n600 S.n599 0.043
R947 S.n94 S.n93 0.043
R948 S.n585 S.n580 0.042
R949 S.n317 S.n312 0.042
R950 S.n285 S.n284 0.042
R951 S.n110 S.n109 0.041
R952 S.n70 S.n69 0.041
R953 S.n13 S.n5 0.04
R954 S.n4 S.n3 0.039
R955 S.n764 S.n763 0.039
R956 S.n653 S.n651 0.038
R957 S.n571 S.n570 0.038
R958 S.n250 S.n249 0.038
R959 S.n331 S.n329 0.037
R960 S.n764 S.n761 0.037
R961 S.n763 S.n762 0.037
R962 S.n516 S.n515 0.037
R963 S.n736 S.n735 0.037
R964 S.n277 S.n70 0.036
R965 S.n362 S.n361 0.036
R966 S.n477 S.n476 0.035
R967 S.n765 S.n764 0.035
R968 S.n571 S.n566 0.035
R969 S.n513 S.n512 0.034
R970 S.n161 S.n160 0.034
R971 S.n360 S.n359 0.034
R972 S.n661 S.n660 0.034
R973 S.n26 S.n22 0.034
R974 S.t17 S.n465 0.034
R975 S.n715 S.n712 0.034
R976 S.n634 S.n630 0.034
R977 S.n432 S.n429 0.034
R978 S.n459 S.n278 0.034
R979 S.n775 S.n774 0.034
R980 S.n155 S.n154 0.034
R981 S.t0 S.n555 0.034
R982 S.t0 S.n554 0.034
R983 S.t3 S.n29 0.034
R984 S.t3 S.n28 0.034
R985 S.t3 S.n58 0.034
R986 S.t3 S.n57 0.034
R987 S.t3 S.n40 0.034
R988 S.t3 S.n39 0.034
R989 S.t3 S.n48 0.034
R990 S.t3 S.n47 0.034
R991 S.t0 S.n547 0.034
R992 S.t0 S.n546 0.034
R993 S.t0 S.n551 0.034
R994 S.t0 S.n550 0.034
R995 S.t0 S.n542 0.034
R996 S.t0 S.n545 0.034
R997 S.n13 S.n12 0.033
R998 S.n654 S.n653 0.032
R999 S.t17 S.n513 0.031
R1000 S.t25 S.n161 0.031
R1001 S.t19 S.n360 0.031
R1002 S.t11 S.n661 0.031
R1003 S.n566 S.n565 0.031
R1004 S.n64 S.n63 0.031
R1005 S.n65 S.n64 0.031
R1006 S.n66 S.n65 0.031
R1007 S.n778 S.n777 0.031
R1008 S.n777 S.n776 0.031
R1009 S.n776 S.n560 0.031
R1010 S.n68 S.n67 0.031
R1011 S.n467 S.n466 0.031
R1012 S.n632 S.n631 0.031
R1013 S.n75 S.n74 0.03
R1014 S.n239 S.n238 0.03
R1015 S.n317 S.n316 0.029
R1016 S.n585 S.n584 0.029
R1017 S.n74 S.n73 0.029
R1018 S.n566 S.n563 0.028
R1019 S.n503 S.n502 0.028
R1020 S.n516 S.n514 0.027
R1021 S.n736 S.n734 0.027
R1022 S.n119 S.n118 0.027
R1023 S.n98 S.n95 0.027
R1024 S.n630 S.n629 0.027
R1025 S.n321 S.n318 0.026
R1026 S.n390 S.n389 0.026
R1027 S.n589 S.n586 0.026
R1028 S.n674 S.n671 0.026
R1029 S.n505 S.n504 0.026
R1030 S.n223 S.n148 0.026
R1031 S.n372 S.n371 0.026
R1032 S.n296 S.n286 0.026
R1033 S.n614 S.n604 0.026
R1034 S.n126 S.n111 0.026
R1035 S.n256 S.n251 0.026
R1036 S.n256 S.n240 0.026
R1037 S.n698 S.n682 0.026
R1038 S.n691 S.n690 0.023
R1039 S.n773 S.n760 0.023
R1040 S.n251 S.n248 0.023
R1041 S.n171 S.n170 0.023
R1042 S.n120 S.n119 0.023
R1043 S.n95 S.n91 0.023
R1044 S.n281 S.n279 0.023
R1045 S.n76 S.n72 0.022
R1046 S.n599 S.n598 0.022
R1047 S.n235 S.n233 0.022
R1048 S.n603 S.n602 0.022
R1049 S.n316 S.n315 0.021
R1050 S.n312 S.n311 0.021
R1051 S.n584 S.n583 0.021
R1052 S.n580 S.n579 0.021
R1053 S.n502 S.n501 0.021
R1054 S.n136 S.n135 0.021
R1055 S.n565 S.n564 0.021
R1056 S.n134 S.n133 0.021
R1057 S.n331 S.n330 0.021
R1058 S.n237 S.n235 0.021
R1059 S.n93 S.n92 0.021
R1060 S.n109 S.n108 0.02
R1061 S.n254 S.n253 0.02
R1062 S.n476 S.n475 0.02
R1063 S.n600 S.n597 0.02
R1064 S.n237 S.n236 0.02
R1065 S.n125 S.n124 0.02
R1066 S.n83 S.n82 0.019
R1067 S.t3 S.n19 0.019
R1068 S.n645 S.n644 0.019
R1069 S.n19 S.n18 0.018
R1070 S.n409 S.n408 0.018
R1071 S.n407 S.n406 0.017
R1072 S.n413 S.n410 0.017
R1073 S.n770 S.n769 0.017
R1074 S.n769 S.n768 0.017
R1075 S.n734 S.n733 0.015
R1076 S.n77 S.n76 0.015
R1077 S.n76 S.n75 0.015
R1078 S.n602 S.n601 0.015
R1079 S.n123 S.n122 0.015
R1080 S.n643 S.n642 0.015
R1081 S.n642 S.n641 0.015
R1082 S.n568 S.n567 0.015
R1083 S.n80 S.n79 0.014
R1084 S.n459 S.n458 0.014
R1085 S.n525 S.n516 0.014
R1086 S.n746 S.n736 0.014
R1087 S.n697 S.n696 0.014
R1088 S.n572 S.n571 0.013
R1089 S.n329 S.n328 0.013
R1090 S.n696 S.n695 0.013
R1091 S.n766 S.n765 0.012
R1092 S.n569 S.n568 0.012
R1093 S.n226 S.n138 0.012
R1094 S.n695 S.n694 0.012
R1095 S.n413 S.n407 0.01
R1096 S.n173 S.n171 0.01
R1097 S.n373 S.n370 0.01
R1098 S.n190 S.n182 0.01
R1099 S.n126 S.n125 0.01
R1100 S.n207 S.n205 0.01
R1101 S.n459 S.n281 0.01
R1102 S.n775 S.n773 0.01
R1103 S.n98 S.n80 0.01
R1104 S.n768 S.n766 0.01
R1105 S.n539 S.n537 0.009
R1106 S.n771 S.n770 0.009
R1107 S.n341 S.n331 0.009
R1108 S.n775 S.n561 0.009
R1109 S.n570 S.n569 0.008
R1110 S.n320 S.n319 0.008
R1111 S.n582 S.n581 0.008
R1112 S.n588 S.n587 0.008
R1113 S.n673 S.n672 0.008
R1114 S.n314 S.n313 0.008
R1115 S.n173 S.n172 0.008
R1116 S.n373 S.n372 0.008
R1117 S.n190 S.n181 0.008
R1118 S.n283 S.n282 0.008
R1119 S.n107 S.n106 0.008
R1120 S.n122 S.n120 0.008
R1121 S.n122 S.n121 0.008
R1122 S.n255 S.n252 0.008
R1123 S.n207 S.n206 0.008
R1124 S.n277 S.n68 0.008
R1125 S.n413 S.n412 0.008
R1126 S.n474 S.n473 0.008
R1127 S.n97 S.n96 0.008
R1128 S.t3 S.n26 0.007
R1129 S.n79 S.n78 0.007
R1130 S.n406 S.n405 0.007
R1131 S.n315 S.n314 0.006
R1132 S.n583 S.n582 0.006
R1133 S.n255 S.n254 0.006
R1134 S.n475 S.n474 0.006
R1135 S.t3 S.n20 0.005
R1136 S.t3 S.n37 0.005
R1137 S.n484 S.n483 0.004
R1138 S.n689 S.n688 0.004
R1139 S.n759 S.n758 0.004
R1140 S.n247 S.n246 0.004
R1141 S.n145 S.n144 0.004
R1142 S.n307 S.n306 0.004
R1143 S.n497 S.n496 0.004
R1144 S.n666 S.n665 0.004
R1145 S.n575 S.n574 0.004
R1146 S.n384 S.n383 0.004
R1147 S.n222 S.n221 0.004
R1148 S.n90 S.n89 0.004
R1149 S.n169 S.n168 0.004
R1150 S.n338 S.n337 0.004
R1151 S.n185 S.n184 0.004
R1152 S.n293 S.n292 0.004
R1153 S.n369 S.n368 0.004
R1154 S.n611 S.n610 0.004
R1155 S.n117 S.n116 0.004
R1156 S.n269 S.n268 0.004
R1157 S.n204 S.n203 0.004
R1158 S.n439 S.n438 0.004
R1159 S.n428 S.n427 0.004
R1160 S.n628 S.n627 0.004
R1161 S.n711 S.n710 0.004
R1162 S.n455 S.n454 0.004
R1163 S.n402 S.n401 0.004
R1164 S.n743 S.n742 0.004
R1165 S.n523 S.n522 0.004
R1166 S.n730 S.n729 0.004
R1167 S.n226 S.n225 0.004
R1168 S.t3 S.n46 0.004
R1169 S.n156 S.n153 0.004
R1170 S.n72 S.n71 0.004
R1171 S.n190 S.n189 0.004
R1172 S.n373 S.n362 0.004
R1173 S.n656 S.n654 0.004
R1174 S.n156 S.n155 0.004
R1175 S.n645 S.n643 0.004
R1176 S.t0 S.n557 0.004
R1177 S.t25 S.n159 0.004
R1178 S.t3 S.n31 0.004
R1179 S.t3 S.n61 0.004
R1180 S.t3 S.n42 0.004
R1181 S.t19 S.n358 0.004
R1182 S.t11 S.n659 0.004
R1183 S.t3 S.n52 0.004
R1184 S.t3 S.n16 0.004
R1185 S.t0 S.n549 0.004
R1186 S.t0 S.n553 0.004
R1187 S.t0 S.n544 0.004
R1188 S.t3 S.n59 0.004
R1189 S.t17 S.n533 0.004
R1190 S.t3 S.n56 0.004
R1191 S.n355 S.n354 0.004
R1192 S.n656 S.n655 0.004
R1193 S.n492 S.n491 0.003
R1194 S.n704 S.n703 0.003
R1195 S.n755 S.n754 0.003
R1196 S.n259 S.n258 0.003
R1197 S.n232 S.n231 0.003
R1198 S.n327 S.n326 0.003
R1199 S.n508 S.n507 0.003
R1200 S.n680 S.n679 0.003
R1201 S.n595 S.n594 0.003
R1202 S.n396 S.n395 0.003
R1203 S.n216 S.n215 0.003
R1204 S.n104 S.n103 0.003
R1205 S.n179 S.n178 0.003
R1206 S.n344 S.n343 0.003
R1207 S.n196 S.n195 0.003
R1208 S.n302 S.n301 0.003
R1209 S.n379 S.n378 0.003
R1210 S.n617 S.n616 0.003
R1211 S.n132 S.n131 0.003
R1212 S.n265 S.n264 0.003
R1213 S.n210 S.n209 0.003
R1214 S.n445 S.n444 0.003
R1215 S.n422 S.n421 0.003
R1216 S.n637 S.n636 0.003
R1217 S.n718 S.n717 0.003
R1218 S.n451 S.n450 0.003
R1219 S.n416 S.n415 0.003
R1220 S.n749 S.n748 0.003
R1221 S.n528 S.n527 0.003
R1222 S.n724 S.n723 0.003
R1223 S.n486 S.n481 0.003
R1224 S.n698 S.n686 0.003
R1225 S.n256 S.n244 0.003
R1226 S.n226 S.n142 0.003
R1227 S.n321 S.n310 0.003
R1228 S.n505 S.n500 0.003
R1229 S.n674 S.n669 0.003
R1230 S.n589 S.n578 0.003
R1231 S.n390 S.n387 0.003
R1232 S.n223 S.n151 0.003
R1233 S.n98 S.n87 0.003
R1234 S.n173 S.n166 0.003
R1235 S.n341 S.n335 0.003
R1236 S.n190 S.n188 0.003
R1237 S.n296 S.n290 0.003
R1238 S.n373 S.n366 0.003
R1239 S.n614 S.n608 0.003
R1240 S.n126 S.n114 0.003
R1241 S.n207 S.n201 0.003
R1242 S.n442 S.n436 0.003
R1243 S.n432 S.n351 0.003
R1244 S.n634 S.n625 0.003
R1245 S.n715 S.n708 0.003
R1246 S.n413 S.n399 0.003
R1247 S.n746 S.n740 0.003
R1248 S.n525 S.n520 0.003
R1249 S.n732 S.n649 0.003
R1250 S.n277 S.n276 0.003
R1251 S.n355 S.n353 0.003
R1252 S.n251 S.n250 0.003
R1253 S.n732 S.n645 0.003
R1254 S.n539 S.n538 0.003
R1255 S.t17 S.n472 0.003
R1256 S.t17 S.n470 0.003
R1257 S.t0 S.n541 0.003
R1258 S.n604 S.n603 0.003
R1259 S.n486 S.n477 0.003
R1260 S.n138 S.n137 0.003
R1261 S.n78 S.n77 0.003
R1262 S.n405 S.n404 0.003
R1263 S.n98 S.n84 0.002
R1264 S.n173 S.n163 0.002
R1265 S.n373 S.n363 0.002
R1266 S.n296 S.n287 0.002
R1267 S.n190 S.n180 0.002
R1268 S.n126 S.n105 0.002
R1269 S.n442 S.n433 0.002
R1270 S.n432 S.n348 0.002
R1271 S.n634 S.n622 0.002
R1272 S.n715 S.n705 0.002
R1273 S.t17 S.n464 0.002
R1274 S.n732 S.n646 0.002
R1275 S.n525 S.n517 0.002
R1276 S.n413 S.n403 0.002
R1277 S.n746 S.n737 0.002
R1278 S.n698 S.n683 0.002
R1279 S.n486 S.n478 0.002
R1280 S.n341 S.n332 0.002
R1281 S.n614 S.n605 0.002
R1282 S.t3 S.n33 0.002
R1283 S.t3 S.n50 0.002
R1284 S.n442 S.n441 0.002
R1285 S.n240 S.n239 0.002
R1286 S.n504 S.n503 0.002
R1287 S.n321 S.n304 0.002
R1288 S.n732 S.n731 0.002
R1289 S.n525 S.n524 0.002
R1290 S.n698 S.n697 0.002
R1291 S.n486 S.n485 0.002
R1292 S.n10 S.n9 0.002
R1293 S.n674 S.n663 0.002
R1294 S.n589 S.n572 0.002
R1295 S.n390 S.n381 0.002
R1296 S.n224 S.n223 0.002
R1297 S.n746 S.n745 0.002
R1298 S.n98 S.n83 0.002
R1299 S.n126 S.n123 0.002
R1300 S.n413 S.n409 0.002
R1301 S.n505 S.n494 0.002
R1302 S.n14 S.n13 0.002
R1303 S.n341 S.n340 0.002
R1304 S.n614 S.n613 0.002
R1305 S.n296 S.n295 0.002
R1306 S.n173 S.n162 0.002
R1307 S.n207 S.n197 0.002
R1308 S.n256 S.n241 0.002
R1309 S.n505 S.n493 0.002
R1310 S.n674 S.n662 0.002
R1311 S.n589 S.n562 0.002
R1312 S.n390 S.n380 0.002
R1313 S.n321 S.n303 0.002
R1314 S.n223 S.n146 0.002
R1315 S.n226 S.n139 0.002
R1316 S.n559 S.n558 0.002
R1317 S.n111 S.n110 0.002
R1318 S.n15 S.n14 0.001
R1319 S.t3 S.n15 0.001
R1320 S.n286 S.n285 0.001
R1321 S.n558 S.t0 0.001
R1322 S.t3 S.n21 0.001
R1323 S.t3 S.n38 0.001
R1324 S.n772 S.n771 0.001
R1325 S.n318 S.n317 0.001
R1326 S.n389 S.n388 0.001
R1327 S.n586 S.n585 0.001
R1328 S.n671 S.n670 0.001
R1329 S.n148 S.n147 0.001
R1330 S.n207 S.n198 0.001
R1331 S.n62 S.t3 0.001
R1332 S.t3 S.n49 0.001
R1333 S.n356 S.n355 0.001
R1334 S.n657 S.n656 0.001
R1335 S.n157 S.n156 0.001
R1336 S.n539 S.n536 0.001
R1337 S.n10 S.n8 0.001
R1338 S.t17 S.n468 0.001
R1339 S.n715 S.n714 0.001
R1340 S.n634 S.n633 0.001
R1341 S.n432 S.n431 0.001
R1342 S.n536 S.t17 0.001
R1343 S.t25 S.n157 0.001
R1344 S.t19 S.n356 0.001
R1345 S.t11 S.n657 0.001
R1346 S.n460 S.n459 0.001
R1347 S.n682 S.n681 0.001
R1348 S.n11 S.n10 0.001
R1349 S.n95 S.n94 0.001
R1350 S.n10 S.n6 0.001
R1351 S.n481 S.n480 0.001
R1352 S.n686 S.n685 0.001
R1353 S.n244 S.n243 0.001
R1354 S.n142 S.n141 0.001
R1355 S.n310 S.n309 0.001
R1356 S.n500 S.n499 0.001
R1357 S.n669 S.n668 0.001
R1358 S.n578 S.n577 0.001
R1359 S.n387 S.n386 0.001
R1360 S.n151 S.n150 0.001
R1361 S.n87 S.n86 0.001
R1362 S.n166 S.n165 0.001
R1363 S.n335 S.n334 0.001
R1364 S.n188 S.n187 0.001
R1365 S.n290 S.n289 0.001
R1366 S.n366 S.n365 0.001
R1367 S.n608 S.n607 0.001
R1368 S.n114 S.n113 0.001
R1369 S.n201 S.n200 0.001
R1370 S.n436 S.n435 0.001
R1371 S.n351 S.n350 0.001
R1372 S.n625 S.n624 0.001
R1373 S.n708 S.n707 0.001
R1374 S.n399 S.n398 0.001
R1375 S.n740 S.n739 0.001
R1376 S.n520 S.n519 0.001
R1377 S.n649 S.n648 0.001
R1378 S.n10 S.n7 0.001
R1379 S.t17 S.n492 0.001
R1380 S.t17 S.n489 0.001
R1381 S.n489 S.n486 0.001
R1382 S.t11 S.n704 0.001
R1383 S.t11 S.n701 0.001
R1384 S.n701 S.n698 0.001
R1385 S.n755 S.t23 0.001
R1386 S.n775 S.n757 0.001
R1387 S.t21 S.n259 0.001
R1388 S.t21 S.n262 0.001
R1389 S.t21 S.n232 0.001
R1390 S.t21 S.n229 0.001
R1391 S.n229 S.n226 0.001
R1392 S.t13 S.n327 0.001
R1393 S.t13 S.n324 0.001
R1394 S.n324 S.n321 0.001
R1395 S.t17 S.n508 0.001
R1396 S.t17 S.n511 0.001
R1397 S.t11 S.n680 0.001
R1398 S.t11 S.n677 0.001
R1399 S.n677 S.n674 0.001
R1400 S.t23 S.n595 0.001
R1401 S.t23 S.n592 0.001
R1402 S.n592 S.n589 0.001
R1403 S.t19 S.n396 0.001
R1404 S.t19 S.n393 0.001
R1405 S.n393 S.n390 0.001
R1406 S.n216 S.t25 0.001
R1407 S.n223 S.n219 0.001
R1408 S.t21 S.n104 0.001
R1409 S.t21 S.n101 0.001
R1410 S.n101 S.n98 0.001
R1411 S.t25 S.n179 0.001
R1412 S.t25 S.n176 0.001
R1413 S.n176 S.n173 0.001
R1414 S.t13 S.n344 0.001
R1415 S.t13 S.n347 0.001
R1416 S.t25 S.n196 0.001
R1417 S.t25 S.n193 0.001
R1418 S.n193 S.n190 0.001
R1419 S.t13 S.n302 0.001
R1420 S.t13 S.n299 0.001
R1421 S.n299 S.n296 0.001
R1422 S.t19 S.n379 0.001
R1423 S.t19 S.n376 0.001
R1424 S.n376 S.n373 0.001
R1425 S.t23 S.n617 0.001
R1426 S.t23 S.n620 0.001
R1427 S.t21 S.n132 0.001
R1428 S.t21 S.n129 0.001
R1429 S.n129 S.n126 0.001
R1430 S.n265 S.t21 0.001
R1431 S.n277 S.n267 0.001
R1432 S.t25 S.n210 0.001
R1433 S.t25 S.n213 0.001
R1434 S.t13 S.n445 0.001
R1435 S.t13 S.n448 0.001
R1436 S.n422 S.t19 0.001
R1437 S.n432 S.n425 0.001
R1438 S.t23 S.n637 0.001
R1439 S.t23 S.n640 0.001
R1440 S.t11 S.n718 0.001
R1441 S.t11 S.n721 0.001
R1442 S.n468 S.n467 0.001
R1443 S.n714 S.n713 0.001
R1444 S.n633 S.n632 0.001
R1445 S.n431 S.n430 0.001
R1446 S.n451 S.t13 0.001
R1447 S.n459 S.n453 0.001
R1448 S.t19 S.n416 0.001
R1449 S.t19 S.n419 0.001
R1450 S.t23 S.n749 0.001
R1451 S.t23 S.n752 0.001
R1452 S.t17 S.n528 0.001
R1453 S.t17 S.n531 0.001
R1454 S.n724 S.t11 0.001
R1455 S.n732 S.n727 0.001
R1456 S.n2 S.n1 0.001
R1457 S.n5 S.n4 0.001
R1458 S.n274 S.n272 0.001
R1459 S.n457 S.n456 0.001
R1460 S.n775 S.n755 0.001
R1461 S.n223 S.n216 0.001
R1462 S.n508 S.n505 0.001
R1463 S.n617 S.n614 0.001
R1464 S.n344 S.n341 0.001
R1465 S.n259 S.n256 0.001
R1466 S.n277 S.n265 0.001
R1467 S.n718 S.n715 0.001
R1468 S.n637 S.n634 0.001
R1469 S.n432 S.n422 0.001
R1470 S.n445 S.n442 0.001
R1471 S.n210 S.n207 0.001
R1472 S.n459 S.n451 0.001
R1473 S.n528 S.n525 0.001
R1474 S.n732 S.n724 0.001
R1475 S.n749 S.n746 0.001
R1476 S.n416 S.n413 0.001
C0 D DNW 165.20fF
C1 G S 291.31fF
C2 D S 442.22fF
C3 G D 190.00fF
C4 DNW S 749.93fF
C5 G DNW 2.66fF
C6 D VSUBS -10.06fF $ **FLOATING
C7 G VSUBS -18.93fF
C8 S VSUBS 49.04fF $ **FLOATING
C9 DNW VSUBS 3204.16fF $ **FLOATING
C10 S.t77 VSUBS 0.02fF
C11 S.n0 VSUBS 1.24fF $ **FLOATING
C12 S.n1 VSUBS 20.83fF $ **FLOATING
C13 S.n2 VSUBS 2.11fF $ **FLOATING
C14 S.n3 VSUBS 0.59fF $ **FLOATING
C15 S.n4 VSUBS 0.50fF $ **FLOATING
C16 S.n5 VSUBS 3.49fF $ **FLOATING
C17 S.n6 VSUBS 4.04fF $ **FLOATING
C18 S.n7 VSUBS 4.08fF $ **FLOATING
C19 S.n8 VSUBS 4.06fF $ **FLOATING
C20 S.n9 VSUBS 4.46fF $ **FLOATING
C21 S.n10 VSUBS 32.46fF $ **FLOATING
C22 S.n11 VSUBS 2.09fF $ **FLOATING
C23 S.n12 VSUBS 12.26fF $ **FLOATING
C24 S.n13 VSUBS 1.79fF $ **FLOATING
C25 S.n14 VSUBS 8.93fF $ **FLOATING
C26 S.n15 VSUBS 0.24fF $ **FLOATING
C27 S.t106 VSUBS 0.02fF
C28 S.n16 VSUBS 0.42fF $ **FLOATING
C29 S.n17 VSUBS 1.00fF $ **FLOATING
C30 S.n18 VSUBS 0.99fF $ **FLOATING
C31 S.n19 VSUBS 0.40fF $ **FLOATING
C32 S.n20 VSUBS 0.26fF $ **FLOATING
C33 S.n21 VSUBS 3.22fF $ **FLOATING
C34 S.n22 VSUBS 0.29fF $ **FLOATING
C35 S.n23 VSUBS 12.93fF $ **FLOATING
C36 S.n24 VSUBS 12.93fF $ **FLOATING
C37 S.n25 VSUBS 4.96fF $ **FLOATING
C38 S.n26 VSUBS 0.95fF $ **FLOATING
C39 S.n27 VSUBS 0.34fF $ **FLOATING
C40 S.t154 VSUBS 0.02fF
C41 S.n28 VSUBS 0.84fF $ **FLOATING
C42 S.t38 VSUBS 0.02fF
C43 S.n29 VSUBS 0.84fF $ **FLOATING
C44 S.n30 VSUBS 0.02fF $ **FLOATING
C45 S.t128 VSUBS 0.02fF
C46 S.n31 VSUBS 0.35fF $ **FLOATING
C47 S.n32 VSUBS 0.76fF $ **FLOATING
C48 S.n33 VSUBS 1.76fF $ **FLOATING
C49 S.n34 VSUBS 8.52fF $ **FLOATING
C50 S.n35 VSUBS 8.52fF $ **FLOATING
C51 S.n36 VSUBS 5.42fF $ **FLOATING
C52 S.n37 VSUBS 1.69fF $ **FLOATING
C53 S.n38 VSUBS 2.51fF $ **FLOATING
C54 S.t29 VSUBS 0.02fF
C55 S.n39 VSUBS 0.84fF $ **FLOATING
C56 S.t91 VSUBS 0.02fF
C57 S.n40 VSUBS 0.84fF $ **FLOATING
C58 S.n41 VSUBS 0.02fF $ **FLOATING
C59 S.t182 VSUBS 0.02fF
C60 S.n42 VSUBS 0.35fF $ **FLOATING
C61 S.n43 VSUBS 8.52fF $ **FLOATING
C62 S.n44 VSUBS 8.52fF $ **FLOATING
C63 S.n45 VSUBS 5.27fF $ **FLOATING
C64 S.n46 VSUBS 1.53fF $ **FLOATING
C65 S.t83 VSUBS 0.02fF
C66 S.n47 VSUBS 0.84fF $ **FLOATING
C67 S.t146 VSUBS 0.02fF
C68 S.n48 VSUBS 0.84fF $ **FLOATING
C69 S.n49 VSUBS 2.51fF $ **FLOATING
C70 S.n50 VSUBS 1.44fF $ **FLOATING
C71 S.n51 VSUBS 0.02fF $ **FLOATING
C72 S.t57 VSUBS 0.02fF
C73 S.n52 VSUBS 0.35fF $ **FLOATING
C74 S.n53 VSUBS 19.76fF $ **FLOATING
C75 S.n54 VSUBS 19.76fF $ **FLOATING
C76 S.n55 VSUBS 5.50fF $ **FLOATING
C77 S.n56 VSUBS 1.86fF $ **FLOATING
C78 S.t97 VSUBS 0.02fF
C79 S.n57 VSUBS 0.84fF $ **FLOATING
C80 S.t15 VSUBS 0.02fF
C81 S.n58 VSUBS 0.84fF $ **FLOATING
C82 S.n59 VSUBS 1.54fF $ **FLOATING
C83 S.n60 VSUBS 0.02fF $ **FLOATING
C84 S.t90 VSUBS 0.02fF
C85 S.n61 VSUBS 0.35fF $ **FLOATING
C86 S.t3 VSUBS 46.64fF
C87 S.n62 VSUBS 3.12fF $ **FLOATING
C88 S.n63 VSUBS 15.59fF $ **FLOATING
C89 S.n64 VSUBS 8.90fF $ **FLOATING
C90 S.n65 VSUBS 8.96fF $ **FLOATING
C91 S.n66 VSUBS 11.51fF $ **FLOATING
C92 S.n67 VSUBS 1.11fF $ **FLOATING
C93 S.n68 VSUBS 0.36fF $ **FLOATING
C94 S.n69 VSUBS 1.15fF $ **FLOATING
C95 S.n70 VSUBS 0.35fF $ **FLOATING
C96 S.n71 VSUBS 0.03fF $ **FLOATING
C97 S.n72 VSUBS 0.03fF $ **FLOATING
C98 S.n73 VSUBS 0.10fF $ **FLOATING
C99 S.n74 VSUBS 0.34fF $ **FLOATING
C100 S.n75 VSUBS 0.36fF $ **FLOATING
C101 S.n76 VSUBS 0.10fF $ **FLOATING
C102 S.n77 VSUBS 0.11fF $ **FLOATING
C103 S.n78 VSUBS 0.03fF $ **FLOATING
C104 S.n79 VSUBS 0.07fF $ **FLOATING
C105 S.n80 VSUBS 1.33fF $ **FLOATING
C106 S.n81 VSUBS 0.04fF $ **FLOATING
C107 S.n82 VSUBS 0.46fF $ **FLOATING
C108 S.n83 VSUBS 0.36fF $ **FLOATING
C109 S.n84 VSUBS 1.54fF $ **FLOATING
C110 S.n85 VSUBS 0.11fF $ **FLOATING
C111 S.t35 VSUBS 0.02fF
C112 S.n86 VSUBS 0.13fF $ **FLOATING
C113 S.t186 VSUBS 0.02fF
C114 S.n88 VSUBS 0.23fF $ **FLOATING
C115 S.n89 VSUBS 0.34fF $ **FLOATING
C116 S.n90 VSUBS 0.58fF $ **FLOATING
C117 S.n91 VSUBS 0.60fF $ **FLOATING
C118 S.n92 VSUBS 0.40fF $ **FLOATING
C119 S.n93 VSUBS 0.19fF $ **FLOATING
C120 S.n94 VSUBS 0.29fF $ **FLOATING
C121 S.n95 VSUBS 0.25fF $ **FLOATING
C122 S.n96 VSUBS 0.24fF $ **FLOATING
C123 S.n97 VSUBS 0.08fF $ **FLOATING
C124 S.n98 VSUBS 1.86fF $ **FLOATING
C125 S.t66 VSUBS 0.02fF
C126 S.n99 VSUBS 0.23fF $ **FLOATING
C127 S.n100 VSUBS 0.87fF $ **FLOATING
C128 S.n101 VSUBS 0.05fF $ **FLOATING
C129 S.t100 VSUBS 0.02fF
C130 S.n102 VSUBS 0.11fF $ **FLOATING
C131 S.n103 VSUBS 0.13fF $ **FLOATING
C132 S.n105 VSUBS 1.43fF $ **FLOATING
C133 S.n106 VSUBS 0.24fF $ **FLOATING
C134 S.n107 VSUBS 0.08fF $ **FLOATING
C135 S.n108 VSUBS 0.74fF $ **FLOATING
C136 S.n109 VSUBS 0.20fF $ **FLOATING
C137 S.n110 VSUBS 1.65fF $ **FLOATING
C138 S.n111 VSUBS 0.42fF $ **FLOATING
C139 S.n112 VSUBS 0.11fF $ **FLOATING
C140 S.t87 VSUBS 0.02fF
C141 S.n113 VSUBS 0.13fF $ **FLOATING
C142 S.t62 VSUBS 0.02fF
C143 S.n115 VSUBS 0.23fF $ **FLOATING
C144 S.n116 VSUBS 0.34fF $ **FLOATING
C145 S.n117 VSUBS 0.58fF $ **FLOATING
C146 S.n118 VSUBS 0.35fF $ **FLOATING
C147 S.n119 VSUBS 0.24fF $ **FLOATING
C148 S.n120 VSUBS 0.60fF $ **FLOATING
C149 S.n121 VSUBS 0.21fF $ **FLOATING
C150 S.n122 VSUBS 0.57fF $ **FLOATING
C151 S.n123 VSUBS 0.26fF $ **FLOATING
C152 S.n124 VSUBS 0.13fF $ **FLOATING
C153 S.n125 VSUBS 1.65fF $ **FLOATING
C154 S.n126 VSUBS 1.84fF $ **FLOATING
C155 S.t122 VSUBS 0.02fF
C156 S.n127 VSUBS 0.23fF $ **FLOATING
C157 S.n128 VSUBS 0.87fF $ **FLOATING
C158 S.n129 VSUBS 0.05fF $ **FLOATING
C159 S.t150 VSUBS 0.02fF
C160 S.n130 VSUBS 0.11fF $ **FLOATING
C161 S.n131 VSUBS 0.13fF $ **FLOATING
C162 S.n133 VSUBS 0.18fF $ **FLOATING
C163 S.n134 VSUBS 0.09fF $ **FLOATING
C164 S.n135 VSUBS 0.65fF $ **FLOATING
C165 S.n136 VSUBS 0.26fF $ **FLOATING
C166 S.n137 VSUBS 1.65fF $ **FLOATING
C167 S.n138 VSUBS 0.20fF $ **FLOATING
C168 S.n139 VSUBS 1.75fF $ **FLOATING
C169 S.n140 VSUBS 0.11fF $ **FLOATING
C170 S.t138 VSUBS 0.02fF
C171 S.n141 VSUBS 0.13fF $ **FLOATING
C172 S.t115 VSUBS 0.02fF
C173 S.n143 VSUBS 0.23fF $ **FLOATING
C174 S.n144 VSUBS 0.34fF $ **FLOATING
C175 S.n145 VSUBS 0.58fF $ **FLOATING
C176 S.n146 VSUBS 1.79fF $ **FLOATING
C177 S.n147 VSUBS 1.10fF $ **FLOATING
C178 S.n148 VSUBS 0.21fF $ **FLOATING
C179 S.n149 VSUBS 0.11fF $ **FLOATING
C180 S.t143 VSUBS 0.02fF
C181 S.n150 VSUBS 0.13fF $ **FLOATING
C182 S.t139 VSUBS 0.02fF
C183 S.n152 VSUBS 1.16fF $ **FLOATING
C184 S.n153 VSUBS 2.18fF $ **FLOATING
C185 S.n154 VSUBS 0.58fF $ **FLOATING
C186 S.n155 VSUBS 2.33fF $ **FLOATING
C187 S.n156 VSUBS 3.74fF $ **FLOATING
C188 S.n157 VSUBS 0.24fF $ **FLOATING
C189 S.n158 VSUBS 0.01fF $ **FLOATING
C190 S.t161 VSUBS 0.02fF
C191 S.n159 VSUBS 0.24fF $ **FLOATING
C192 S.t16 VSUBS 0.02fF
C193 S.n160 VSUBS 0.90fF $ **FLOATING
C194 S.n161 VSUBS 0.67fF $ **FLOATING
C195 S.n162 VSUBS 1.37fF $ **FLOATING
C196 S.n163 VSUBS 1.78fF $ **FLOATING
C197 S.n164 VSUBS 0.11fF $ **FLOATING
C198 S.t36 VSUBS 0.02fF
C199 S.n165 VSUBS 0.13fF $ **FLOATING
C200 S.t1 VSUBS 0.02fF
C201 S.n167 VSUBS 0.23fF $ **FLOATING
C202 S.n168 VSUBS 0.34fF $ **FLOATING
C203 S.n169 VSUBS 0.58fF $ **FLOATING
C204 S.n170 VSUBS 0.86fF $ **FLOATING
C205 S.n171 VSUBS 1.57fF $ **FLOATING
C206 S.n172 VSUBS 0.33fF $ **FLOATING
C207 S.n173 VSUBS 2.05fF $ **FLOATING
C208 S.t73 VSUBS 0.02fF
C209 S.n174 VSUBS 0.23fF $ **FLOATING
C210 S.n175 VSUBS 0.87fF $ **FLOATING
C211 S.n176 VSUBS 0.05fF $ **FLOATING
C212 S.t101 VSUBS 0.02fF
C213 S.n177 VSUBS 0.11fF $ **FLOATING
C214 S.n178 VSUBS 0.13fF $ **FLOATING
C215 S.n180 VSUBS 1.78fF $ **FLOATING
C216 S.n181 VSUBS 0.33fF $ **FLOATING
C217 S.n182 VSUBS 1.18fF $ **FLOATING
C218 S.t64 VSUBS 0.02fF
C219 S.n183 VSUBS 0.23fF $ **FLOATING
C220 S.n184 VSUBS 0.34fF $ **FLOATING
C221 S.n185 VSUBS 0.58fF $ **FLOATING
C222 S.n186 VSUBS 0.11fF $ **FLOATING
C223 S.t89 VSUBS 0.02fF
C224 S.n187 VSUBS 0.13fF $ **FLOATING
C225 S.n189 VSUBS 2.18fF $ **FLOATING
C226 S.n190 VSUBS 1.92fF $ **FLOATING
C227 S.t123 VSUBS 0.02fF
C228 S.n191 VSUBS 0.23fF $ **FLOATING
C229 S.n192 VSUBS 0.87fF $ **FLOATING
C230 S.n193 VSUBS 0.05fF $ **FLOATING
C231 S.t152 VSUBS 0.02fF
C232 S.n194 VSUBS 0.11fF $ **FLOATING
C233 S.n195 VSUBS 0.13fF $ **FLOATING
C234 S.n197 VSUBS 2.60fF $ **FLOATING
C235 S.n198 VSUBS 1.84fF $ **FLOATING
C236 S.n199 VSUBS 0.11fF $ **FLOATING
C237 S.t65 VSUBS 0.02fF
C238 S.n200 VSUBS 0.13fF $ **FLOATING
C239 S.t58 VSUBS 0.02fF
C240 S.n202 VSUBS 0.23fF $ **FLOATING
C241 S.n203 VSUBS 0.34fF $ **FLOATING
C242 S.n204 VSUBS 0.58fF $ **FLOATING
C243 S.n205 VSUBS 1.48fF $ **FLOATING
C244 S.n206 VSUBS 0.27fF $ **FLOATING
C245 S.n207 VSUBS 2.00fF $ **FLOATING
C246 S.t80 VSUBS 0.02fF
C247 S.n208 VSUBS 0.11fF $ **FLOATING
C248 S.n209 VSUBS 0.13fF $ **FLOATING
C249 S.t167 VSUBS 0.02fF
C250 S.n211 VSUBS 0.23fF $ **FLOATING
C251 S.n212 VSUBS 0.87fF $ **FLOATING
C252 S.n213 VSUBS 0.05fF $ **FLOATING
C253 S.t25 VSUBS 13.78fF
C254 S.t26 VSUBS 0.02fF
C255 S.n214 VSUBS 0.11fF $ **FLOATING
C256 S.n215 VSUBS 0.13fF $ **FLOATING
C257 S.t179 VSUBS 0.02fF
C258 S.n217 VSUBS 0.23fF $ **FLOATING
C259 S.n218 VSUBS 0.87fF $ **FLOATING
C260 S.n219 VSUBS 0.05fF $ **FLOATING
C261 S.t118 VSUBS 0.02fF
C262 S.n220 VSUBS 0.23fF $ **FLOATING
C263 S.n221 VSUBS 0.34fF $ **FLOATING
C264 S.n222 VSUBS 0.58fF $ **FLOATING
C265 S.n223 VSUBS 1.78fF $ **FLOATING
C266 S.n224 VSUBS 2.60fF $ **FLOATING
C267 S.n225 VSUBS 2.37fF $ **FLOATING
C268 S.n226 VSUBS 1.76fF $ **FLOATING
C269 S.t175 VSUBS 0.02fF
C270 S.n227 VSUBS 0.23fF $ **FLOATING
C271 S.n228 VSUBS 0.87fF $ **FLOATING
C272 S.n229 VSUBS 0.05fF $ **FLOATING
C273 S.t22 VSUBS 0.02fF
C274 S.n230 VSUBS 0.11fF $ **FLOATING
C275 S.n231 VSUBS 0.13fF $ **FLOATING
C276 S.n233 VSUBS 0.06fF $ **FLOATING
C277 S.n234 VSUBS 0.19fF $ **FLOATING
C278 S.n235 VSUBS 0.09fF $ **FLOATING
C279 S.n236 VSUBS 0.20fF $ **FLOATING
C280 S.n237 VSUBS 0.09fF $ **FLOATING
C281 S.n238 VSUBS 0.29fF $ **FLOATING
C282 S.n239 VSUBS 0.71fF $ **FLOATING
C283 S.n240 VSUBS 0.43fF $ **FLOATING
C284 S.n241 VSUBS 1.61fF $ **FLOATING
C285 S.n242 VSUBS 0.11fF $ **FLOATING
C286 S.t159 VSUBS 0.02fF
C287 S.n243 VSUBS 0.13fF $ **FLOATING
C288 S.t135 VSUBS 0.02fF
C289 S.n245 VSUBS 0.23fF $ **FLOATING
C290 S.n246 VSUBS 0.34fF $ **FLOATING
C291 S.n247 VSUBS 0.58fF $ **FLOATING
C292 S.n248 VSUBS 0.38fF $ **FLOATING
C293 S.n249 VSUBS 0.64fF $ **FLOATING
C294 S.n250 VSUBS 0.37fF $ **FLOATING
C295 S.n251 VSUBS 0.42fF $ **FLOATING
C296 S.n252 VSUBS 0.24fF $ **FLOATING
C297 S.n253 VSUBS 0.75fF $ **FLOATING
C298 S.n254 VSUBS 0.18fF $ **FLOATING
C299 S.n255 VSUBS 0.08fF $ **FLOATING
C300 S.n256 VSUBS 1.62fF $ **FLOATING
C301 S.t43 VSUBS 0.02fF
C302 S.n257 VSUBS 0.11fF $ **FLOATING
C303 S.n258 VSUBS 0.13fF $ **FLOATING
C304 S.t4 VSUBS 0.02fF
C305 S.n260 VSUBS 0.23fF $ **FLOATING
C306 S.n261 VSUBS 0.87fF $ **FLOATING
C307 S.n262 VSUBS 0.05fF $ **FLOATING
C308 S.t21 VSUBS 13.41fF
C309 S.t168 VSUBS 0.02fF
C310 S.n263 VSUBS 0.01fF $ **FLOATING
C311 S.n264 VSUBS 0.24fF $ **FLOATING
C312 S.t47 VSUBS 0.02fF
C313 S.n266 VSUBS 1.14fF $ **FLOATING
C314 S.n267 VSUBS 0.05fF $ **FLOATING
C315 S.t7 VSUBS 0.02fF
C316 S.n268 VSUBS 0.61fF $ **FLOATING
C317 S.n269 VSUBS 0.58fF $ **FLOATING
C318 S.n270 VSUBS 19.35fF $ **FLOATING
C319 S.n271 VSUBS 0.20fF $ **FLOATING
C320 S.n272 VSUBS 1.35fF $ **FLOATING
C321 S.n273 VSUBS 19.35fF $ **FLOATING
C322 S.n274 VSUBS 4.03fF $ **FLOATING
C323 S.n275 VSUBS 1.08fF $ **FLOATING
C324 S.n276 VSUBS 1.71fF $ **FLOATING
C325 S.n277 VSUBS 4.03fF $ **FLOATING
C326 S.n278 VSUBS 0.23fF $ **FLOATING
C327 S.n279 VSUBS 1.42fF $ **FLOATING
C328 S.n280 VSUBS 1.19fF $ **FLOATING
C329 S.n281 VSUBS 0.26fF $ **FLOATING
C330 S.n282 VSUBS 0.24fF $ **FLOATING
C331 S.n283 VSUBS 0.08fF $ **FLOATING
C332 S.n284 VSUBS 0.20fF $ **FLOATING
C333 S.n285 VSUBS 1.22fF $ **FLOATING
C334 S.n286 VSUBS 0.50fF $ **FLOATING
C335 S.n287 VSUBS 1.78fF $ **FLOATING
C336 S.n288 VSUBS 0.11fF $ **FLOATING
C337 S.t92 VSUBS 0.02fF
C338 S.n289 VSUBS 0.13fF $ **FLOATING
C339 S.t67 VSUBS 0.02fF
C340 S.n291 VSUBS 0.23fF $ **FLOATING
C341 S.n292 VSUBS 0.34fF $ **FLOATING
C342 S.n293 VSUBS 0.58fF $ **FLOATING
C343 S.n294 VSUBS 0.68fF $ **FLOATING
C344 S.n295 VSUBS 1.50fF $ **FLOATING
C345 S.n296 VSUBS 2.32fF $ **FLOATING
C346 S.t126 VSUBS 0.02fF
C347 S.n297 VSUBS 0.23fF $ **FLOATING
C348 S.n298 VSUBS 0.87fF $ **FLOATING
C349 S.n299 VSUBS 0.05fF $ **FLOATING
C350 S.t155 VSUBS 0.02fF
C351 S.n300 VSUBS 0.11fF $ **FLOATING
C352 S.n301 VSUBS 0.13fF $ **FLOATING
C353 S.n303 VSUBS 1.79fF $ **FLOATING
C354 S.n304 VSUBS 2.54fF $ **FLOATING
C355 S.t121 VSUBS 0.02fF
C356 S.n305 VSUBS 0.23fF $ **FLOATING
C357 S.n306 VSUBS 0.34fF $ **FLOATING
C358 S.n307 VSUBS 0.58fF $ **FLOATING
C359 S.n308 VSUBS 0.11fF $ **FLOATING
C360 S.t145 VSUBS 0.02fF
C361 S.n309 VSUBS 0.13fF $ **FLOATING
C362 S.n311 VSUBS 0.66fF $ **FLOATING
C363 S.n312 VSUBS 0.21fF $ **FLOATING
C364 S.n313 VSUBS 0.24fF $ **FLOATING
C365 S.n314 VSUBS 0.08fF $ **FLOATING
C366 S.n315 VSUBS 0.21fF $ **FLOATING
C367 S.n316 VSUBS 0.66fF $ **FLOATING
C368 S.n317 VSUBS 1.10fF $ **FLOATING
C369 S.n318 VSUBS 0.21fF $ **FLOATING
C370 S.n319 VSUBS 0.24fF $ **FLOATING
C371 S.n320 VSUBS 0.08fF $ **FLOATING
C372 S.n321 VSUBS 1.79fF $ **FLOATING
C373 S.t181 VSUBS 0.02fF
C374 S.n322 VSUBS 0.23fF $ **FLOATING
C375 S.n323 VSUBS 0.87fF $ **FLOATING
C376 S.n324 VSUBS 0.05fF $ **FLOATING
C377 S.t28 VSUBS 0.02fF
C378 S.n325 VSUBS 0.11fF $ **FLOATING
C379 S.n326 VSUBS 0.13fF $ **FLOATING
C380 S.n328 VSUBS 0.18fF $ **FLOATING
C381 S.n329 VSUBS 1.50fF $ **FLOATING
C382 S.n330 VSUBS 2.10fF $ **FLOATING
C383 S.n331 VSUBS 0.31fF $ **FLOATING
C384 S.n332 VSUBS 2.27fF $ **FLOATING
C385 S.n333 VSUBS 0.11fF $ **FLOATING
C386 S.t39 VSUBS 0.02fF
C387 S.n334 VSUBS 0.13fF $ **FLOATING
C388 S.t5 VSUBS 0.02fF
C389 S.n336 VSUBS 0.23fF $ **FLOATING
C390 S.n337 VSUBS 0.34fF $ **FLOATING
C391 S.n338 VSUBS 0.58fF $ **FLOATING
C392 S.n339 VSUBS 0.68fF $ **FLOATING
C393 S.n340 VSUBS 1.64fF $ **FLOATING
C394 S.n341 VSUBS 2.29fF $ **FLOATING
C395 S.t103 VSUBS 0.02fF
C396 S.n342 VSUBS 0.11fF $ **FLOATING
C397 S.n343 VSUBS 0.13fF $ **FLOATING
C398 S.t74 VSUBS 0.02fF
C399 S.n345 VSUBS 0.23fF $ **FLOATING
C400 S.n346 VSUBS 0.87fF $ **FLOATING
C401 S.n347 VSUBS 0.05fF $ **FLOATING
C402 S.n348 VSUBS 1.78fF $ **FLOATING
C403 S.n349 VSUBS 0.11fF $ **FLOATING
C404 S.t20 VSUBS 0.02fF
C405 S.n350 VSUBS 0.13fF $ **FLOATING
C406 S.t8 VSUBS 0.02fF
C407 S.n352 VSUBS 1.16fF $ **FLOATING
C408 S.n353 VSUBS 1.90fF $ **FLOATING
C409 S.n354 VSUBS 2.35fF $ **FLOATING
C410 S.n355 VSUBS 4.15fF $ **FLOATING
C411 S.n356 VSUBS 0.24fF $ **FLOATING
C412 S.n357 VSUBS 0.01fF $ **FLOATING
C413 S.t44 VSUBS 0.02fF
C414 S.n358 VSUBS 0.24fF $ **FLOATING
C415 S.t78 VSUBS 0.02fF
C416 S.n359 VSUBS 0.90fF $ **FLOATING
C417 S.n360 VSUBS 0.67fF $ **FLOATING
C418 S.n361 VSUBS 0.74fF $ **FLOATING
C419 S.n362 VSUBS 2.15fF $ **FLOATING
C420 S.n363 VSUBS 1.78fF $ **FLOATING
C421 S.n364 VSUBS 0.11fF $ **FLOATING
C422 S.t98 VSUBS 0.02fF
C423 S.n365 VSUBS 0.13fF $ **FLOATING
C424 S.t70 VSUBS 0.02fF
C425 S.n367 VSUBS 0.23fF $ **FLOATING
C426 S.n368 VSUBS 0.34fF $ **FLOATING
C427 S.n369 VSUBS 0.58fF $ **FLOATING
C428 S.n370 VSUBS 1.32fF $ **FLOATING
C429 S.n371 VSUBS 1.08fF $ **FLOATING
C430 S.n372 VSUBS 0.33fF $ **FLOATING
C431 S.n373 VSUBS 1.92fF $ **FLOATING
C432 S.t129 VSUBS 0.02fF
C433 S.n374 VSUBS 0.23fF $ **FLOATING
C434 S.n375 VSUBS 0.87fF $ **FLOATING
C435 S.n376 VSUBS 0.05fF $ **FLOATING
C436 S.t160 VSUBS 0.02fF
C437 S.n377 VSUBS 0.11fF $ **FLOATING
C438 S.n378 VSUBS 0.13fF $ **FLOATING
C439 S.n380 VSUBS 1.79fF $ **FLOATING
C440 S.n381 VSUBS 2.55fF $ **FLOATING
C441 S.t124 VSUBS 0.02fF
C442 S.n382 VSUBS 0.23fF $ **FLOATING
C443 S.n383 VSUBS 0.34fF $ **FLOATING
C444 S.n384 VSUBS 0.58fF $ **FLOATING
C445 S.n385 VSUBS 0.11fF $ **FLOATING
C446 S.t149 VSUBS 0.02fF
C447 S.n386 VSUBS 0.13fF $ **FLOATING
C448 S.n388 VSUBS 1.10fF $ **FLOATING
C449 S.n389 VSUBS 0.21fF $ **FLOATING
C450 S.n390 VSUBS 1.79fF $ **FLOATING
C451 S.t183 VSUBS 0.02fF
C452 S.n391 VSUBS 0.23fF $ **FLOATING
C453 S.n392 VSUBS 0.87fF $ **FLOATING
C454 S.n393 VSUBS 0.05fF $ **FLOATING
C455 S.t31 VSUBS 0.02fF
C456 S.n394 VSUBS 0.11fF $ **FLOATING
C457 S.n395 VSUBS 0.13fF $ **FLOATING
C458 S.n397 VSUBS 0.11fF $ **FLOATING
C459 S.t51 VSUBS 0.02fF
C460 S.n398 VSUBS 0.13fF $ **FLOATING
C461 S.t49 VSUBS 0.02fF
C462 S.n400 VSUBS 0.23fF $ **FLOATING
C463 S.n401 VSUBS 0.34fF $ **FLOATING
C464 S.n402 VSUBS 0.58fF $ **FLOATING
C465 S.n403 VSUBS 1.51fF $ **FLOATING
C466 S.n404 VSUBS 0.11fF $ **FLOATING
C467 S.n405 VSUBS 0.03fF $ **FLOATING
C468 S.n406 VSUBS 0.13fF $ **FLOATING
C469 S.n407 VSUBS 0.55fF $ **FLOATING
C470 S.n408 VSUBS 0.51fF $ **FLOATING
C471 S.n409 VSUBS 0.39fF $ **FLOATING
C472 S.n410 VSUBS 0.24fF $ **FLOATING
C473 S.n411 VSUBS 0.49fF $ **FLOATING
C474 S.n412 VSUBS 0.66fF $ **FLOATING
C475 S.n413 VSUBS 1.87fF $ **FLOATING
C476 S.t137 VSUBS 0.02fF
C477 S.n414 VSUBS 0.11fF $ **FLOATING
C478 S.n415 VSUBS 0.13fF $ **FLOATING
C479 S.t151 VSUBS 0.02fF
C480 S.n417 VSUBS 0.23fF $ **FLOATING
C481 S.n418 VSUBS 0.87fF $ **FLOATING
C482 S.n419 VSUBS 0.05fF $ **FLOATING
C483 S.t19 VSUBS 13.78fF
C484 S.t86 VSUBS 0.02fF
C485 S.n420 VSUBS 0.11fF $ **FLOATING
C486 S.n421 VSUBS 0.13fF $ **FLOATING
C487 S.t56 VSUBS 0.02fF
C488 S.n423 VSUBS 0.23fF $ **FLOATING
C489 S.n424 VSUBS 0.87fF $ **FLOATING
C490 S.n425 VSUBS 0.05fF $ **FLOATING
C491 S.t178 VSUBS 0.02fF
C492 S.n426 VSUBS 0.23fF $ **FLOATING
C493 S.n427 VSUBS 0.34fF $ **FLOATING
C494 S.n428 VSUBS 0.58fF $ **FLOATING
C495 S.n429 VSUBS 0.30fF $ **FLOATING
C496 S.n430 VSUBS 1.47fF $ **FLOATING
C497 S.n431 VSUBS 0.15fF $ **FLOATING
C498 S.n432 VSUBS 4.72fF $ **FLOATING
C499 S.n433 VSUBS 1.78fF $ **FLOATING
C500 S.n434 VSUBS 0.11fF $ **FLOATING
C501 S.t14 VSUBS 0.02fF
C502 S.n435 VSUBS 0.13fF $ **FLOATING
C503 S.t174 VSUBS 0.02fF
C504 S.n437 VSUBS 0.23fF $ **FLOATING
C505 S.n438 VSUBS 0.34fF $ **FLOATING
C506 S.n439 VSUBS 0.58fF $ **FLOATING
C507 S.n440 VSUBS 0.67fF $ **FLOATING
C508 S.n441 VSUBS 1.21fF $ **FLOATING
C509 S.n442 VSUBS 5.67fF $ **FLOATING
C510 S.t82 VSUBS 0.02fF
C511 S.n443 VSUBS 0.11fF $ **FLOATING
C512 S.n444 VSUBS 0.13fF $ **FLOATING
C513 S.t54 VSUBS 0.02fF
C514 S.n446 VSUBS 0.23fF $ **FLOATING
C515 S.n447 VSUBS 0.87fF $ **FLOATING
C516 S.n448 VSUBS 0.05fF $ **FLOATING
C517 S.t13 VSUBS 13.41fF
C518 S.t163 VSUBS 0.02fF
C519 S.n449 VSUBS 0.01fF $ **FLOATING
C520 S.n450 VSUBS 0.24fF $ **FLOATING
C521 S.t171 VSUBS 0.02fF
C522 S.n452 VSUBS 1.14fF $ **FLOATING
C523 S.n453 VSUBS 0.05fF $ **FLOATING
C524 S.t165 VSUBS 0.02fF
C525 S.n454 VSUBS 0.61fF $ **FLOATING
C526 S.n455 VSUBS 0.58fF $ **FLOATING
C527 S.n456 VSUBS 0.26fF $ **FLOATING
C528 S.n457 VSUBS 4.05fF $ **FLOATING
C529 S.n458 VSUBS 2.84fF $ **FLOATING
C530 S.n459 VSUBS 1.72fF $ **FLOATING
C531 S.n460 VSUBS 2.51fF $ **FLOATING
C532 S.t72 VSUBS 0.02fF
C533 S.n461 VSUBS 1.16fF $ **FLOATING
C534 S.t68 VSUBS 0.02fF
C535 S.n462 VSUBS 0.23fF $ **FLOATING
C536 S.n463 VSUBS 0.88fF $ **FLOATING
C537 S.n464 VSUBS 1.79fF $ **FLOATING
C538 S.n465 VSUBS 0.30fF $ **FLOATING
C539 S.n466 VSUBS 0.88fF $ **FLOATING
C540 S.n467 VSUBS 1.03fF $ **FLOATING
C541 S.n468 VSUBS 0.15fF $ **FLOATING
C542 S.t99 VSUBS 0.02fF
C543 S.n469 VSUBS 0.11fF $ **FLOATING
C544 S.n470 VSUBS 0.13fF $ **FLOATING
C545 S.n471 VSUBS 0.11fF $ **FLOATING
C546 S.t32 VSUBS 0.02fF
C547 S.n472 VSUBS 0.13fF $ **FLOATING
C548 S.n473 VSUBS 0.24fF $ **FLOATING
C549 S.n474 VSUBS 0.08fF $ **FLOATING
C550 S.n475 VSUBS 0.19fF $ **FLOATING
C551 S.n476 VSUBS 0.74fF $ **FLOATING
C552 S.n477 VSUBS 1.84fF $ **FLOATING
C553 S.n478 VSUBS 1.78fF $ **FLOATING
C554 S.n479 VSUBS 0.11fF $ **FLOATING
C555 S.t136 VSUBS 0.02fF
C556 S.n480 VSUBS 0.13fF $ **FLOATING
C557 S.t113 VSUBS 0.02fF
C558 S.n482 VSUBS 0.23fF $ **FLOATING
C559 S.n483 VSUBS 0.34fF $ **FLOATING
C560 S.n484 VSUBS 0.58fF $ **FLOATING
C561 S.n485 VSUBS 2.53fF $ **FLOATING
C562 S.n486 VSUBS 2.84fF $ **FLOATING
C563 S.t173 VSUBS 0.02fF
C564 S.n487 VSUBS 0.23fF $ **FLOATING
C565 S.n488 VSUBS 0.87fF $ **FLOATING
C566 S.n489 VSUBS 0.05fF $ **FLOATING
C567 S.t18 VSUBS 0.02fF
C568 S.n490 VSUBS 0.11fF $ **FLOATING
C569 S.n491 VSUBS 0.13fF $ **FLOATING
C570 S.n493 VSUBS 1.69fF $ **FLOATING
C571 S.n494 VSUBS 2.89fF $ **FLOATING
C572 S.t133 VSUBS 0.02fF
C573 S.n495 VSUBS 0.23fF $ **FLOATING
C574 S.n496 VSUBS 0.34fF $ **FLOATING
C575 S.n497 VSUBS 0.58fF $ **FLOATING
C576 S.n498 VSUBS 0.11fF $ **FLOATING
C577 S.t158 VSUBS 0.02fF
C578 S.n499 VSUBS 0.13fF $ **FLOATING
C579 S.n501 VSUBS 0.21fF $ **FLOATING
C580 S.n502 VSUBS 0.63fF $ **FLOATING
C581 S.n503 VSUBS 0.86fF $ **FLOATING
C582 S.n504 VSUBS 0.21fF $ **FLOATING
C583 S.n505 VSUBS 1.89fF $ **FLOATING
C584 S.t42 VSUBS 0.02fF
C585 S.n506 VSUBS 0.11fF $ **FLOATING
C586 S.n507 VSUBS 0.13fF $ **FLOATING
C587 S.t6 VSUBS 0.02fF
C588 S.n509 VSUBS 0.23fF $ **FLOATING
C589 S.n510 VSUBS 0.87fF $ **FLOATING
C590 S.n511 VSUBS 0.05fF $ **FLOATING
C591 S.t107 VSUBS 0.02fF
C592 S.n512 VSUBS 0.90fF $ **FLOATING
C593 S.n513 VSUBS 0.67fF $ **FLOATING
C594 S.n514 VSUBS 0.34fF $ **FLOATING
C595 S.n515 VSUBS 0.44fF $ **FLOATING
C596 S.n516 VSUBS 1.08fF $ **FLOATING
C597 S.n517 VSUBS 1.78fF $ **FLOATING
C598 S.n518 VSUBS 0.11fF $ **FLOATING
C599 S.t85 VSUBS 0.02fF
C600 S.n519 VSUBS 0.13fF $ **FLOATING
C601 S.t60 VSUBS 0.02fF
C602 S.n521 VSUBS 0.23fF $ **FLOATING
C603 S.n522 VSUBS 0.34fF $ **FLOATING
C604 S.n523 VSUBS 0.58fF $ **FLOATING
C605 S.n524 VSUBS 2.53fF $ **FLOATING
C606 S.n525 VSUBS 3.71fF $ **FLOATING
C607 S.t148 VSUBS 0.02fF
C608 S.n526 VSUBS 0.11fF $ **FLOATING
C609 S.n527 VSUBS 0.13fF $ **FLOATING
C610 S.t120 VSUBS 0.02fF
C611 S.n529 VSUBS 0.23fF $ **FLOATING
C612 S.n530 VSUBS 0.87fF $ **FLOATING
C613 S.n531 VSUBS 0.05fF $ **FLOATING
C614 S.t116 VSUBS 0.02fF
C615 S.n532 VSUBS 0.01fF $ **FLOATING
C616 S.n533 VSUBS 0.24fF $ **FLOATING
C617 S.n534 VSUBS 0.23fF $ **FLOATING
C618 S.t188 VSUBS 0.02fF
C619 S.n535 VSUBS 0.87fF $ **FLOATING
C620 S.t17 VSUBS 18.57fF
C621 S.n536 VSUBS 0.24fF $ **FLOATING
C622 S.n537 VSUBS 2.77fF $ **FLOATING
C623 S.n538 VSUBS 2.21fF $ **FLOATING
C624 S.n539 VSUBS 4.34fF $ **FLOATING
C625 S.t45 VSUBS 0.02fF
C626 S.n540 VSUBS 1.21fF $ **FLOATING
C627 S.t34 VSUBS 0.02fF
C628 S.n541 VSUBS 0.42fF $ **FLOATING
C629 S.t157 VSUBS 0.02fF
C630 S.n542 VSUBS 0.84fF $ **FLOATING
C631 S.t169 VSUBS 0.02fF
C632 S.n543 VSUBS 0.02fF $ **FLOATING
C633 S.n544 VSUBS 0.35fF $ **FLOATING
C634 S.t95 VSUBS 0.02fF
C635 S.n545 VSUBS 0.84fF $ **FLOATING
C636 S.t108 VSUBS 0.02fF
C637 S.n546 VSUBS 0.84fF $ **FLOATING
C638 S.t166 VSUBS 0.02fF
C639 S.n547 VSUBS 0.84fF $ **FLOATING
C640 S.t176 VSUBS 0.02fF
C641 S.n548 VSUBS 0.02fF $ **FLOATING
C642 S.n549 VSUBS 0.35fF $ **FLOATING
C643 S.t164 VSUBS 0.02fF
C644 S.n550 VSUBS 0.84fF $ **FLOATING
C645 S.t46 VSUBS 0.02fF
C646 S.n551 VSUBS 0.84fF $ **FLOATING
C647 S.t52 VSUBS 0.02fF
C648 S.n552 VSUBS 0.02fF $ **FLOATING
C649 S.n553 VSUBS 0.35fF $ **FLOATING
C650 S.t41 VSUBS 0.02fF
C651 S.n554 VSUBS 0.84fF $ **FLOATING
C652 S.t105 VSUBS 0.02fF
C653 S.n555 VSUBS 0.84fF $ **FLOATING
C654 S.t111 VSUBS 0.02fF
C655 S.n556 VSUBS 0.02fF $ **FLOATING
C656 S.n557 VSUBS 0.35fF $ **FLOATING
C657 S.t0 VSUBS 530.76fF
C658 S.n558 VSUBS 0.44fF $ **FLOATING
C659 S.n559 VSUBS 6.58fF $ **FLOATING
C660 S.n560 VSUBS 15.33fF $ **FLOATING
C661 S.n561 VSUBS 2.67fF $ **FLOATING
C662 S.n562 VSUBS 1.79fF $ **FLOATING
C663 S.n563 VSUBS 0.06fF $ **FLOATING
C664 S.n564 VSUBS 0.03fF $ **FLOATING
C665 S.n565 VSUBS 0.03fF $ **FLOATING
C666 S.n566 VSUBS 0.94fF $ **FLOATING
C667 S.n567 VSUBS 0.02fF $ **FLOATING
C668 S.n568 VSUBS 0.01fF $ **FLOATING
C669 S.n569 VSUBS 0.01fF $ **FLOATING
C670 S.n570 VSUBS 0.08fF $ **FLOATING
C671 S.n571 VSUBS 0.34fF $ **FLOATING
C672 S.n572 VSUBS 1.76fF $ **FLOATING
C673 S.t127 VSUBS 0.02fF
C674 S.n573 VSUBS 0.23fF $ **FLOATING
C675 S.n574 VSUBS 0.34fF $ **FLOATING
C676 S.n575 VSUBS 0.58fF $ **FLOATING
C677 S.n576 VSUBS 0.11fF $ **FLOATING
C678 S.t153 VSUBS 0.02fF
C679 S.n577 VSUBS 0.13fF $ **FLOATING
C680 S.n579 VSUBS 0.66fF $ **FLOATING
C681 S.n580 VSUBS 0.21fF $ **FLOATING
C682 S.n581 VSUBS 0.24fF $ **FLOATING
C683 S.n582 VSUBS 0.08fF $ **FLOATING
C684 S.n583 VSUBS 0.21fF $ **FLOATING
C685 S.n584 VSUBS 0.66fF $ **FLOATING
C686 S.n585 VSUBS 1.10fF $ **FLOATING
C687 S.n586 VSUBS 0.21fF $ **FLOATING
C688 S.n587 VSUBS 0.24fF $ **FLOATING
C689 S.n588 VSUBS 0.08fF $ **FLOATING
C690 S.n589 VSUBS 1.79fF $ **FLOATING
C691 S.t187 VSUBS 0.02fF
C692 S.n590 VSUBS 0.23fF $ **FLOATING
C693 S.n591 VSUBS 0.87fF $ **FLOATING
C694 S.n592 VSUBS 0.05fF $ **FLOATING
C695 S.t37 VSUBS 0.02fF
C696 S.n593 VSUBS 0.11fF $ **FLOATING
C697 S.n594 VSUBS 0.13fF $ **FLOATING
C698 S.n596 VSUBS 0.09fF $ **FLOATING
C699 S.n597 VSUBS 0.20fF $ **FLOATING
C700 S.n598 VSUBS 0.06fF $ **FLOATING
C701 S.n599 VSUBS 0.06fF $ **FLOATING
C702 S.n600 VSUBS 0.06fF $ **FLOATING
C703 S.n601 VSUBS 0.17fF $ **FLOATING
C704 S.n602 VSUBS 0.19fF $ **FLOATING
C705 S.n603 VSUBS 0.98fF $ **FLOATING
C706 S.n604 VSUBS 0.51fF $ **FLOATING
C707 S.n605 VSUBS 2.22fF $ **FLOATING
C708 S.n606 VSUBS 0.11fF $ **FLOATING
C709 S.t102 VSUBS 0.02fF
C710 S.n607 VSUBS 0.13fF $ **FLOATING
C711 S.t75 VSUBS 0.02fF
C712 S.n609 VSUBS 0.23fF $ **FLOATING
C713 S.n610 VSUBS 0.34fF $ **FLOATING
C714 S.n611 VSUBS 0.58fF $ **FLOATING
C715 S.n612 VSUBS 0.68fF $ **FLOATING
C716 S.n613 VSUBS 1.64fF $ **FLOATING
C717 S.n614 VSUBS 2.32fF $ **FLOATING
C718 S.t162 VSUBS 0.02fF
C719 S.n615 VSUBS 0.11fF $ **FLOATING
C720 S.n616 VSUBS 0.13fF $ **FLOATING
C721 S.t132 VSUBS 0.02fF
C722 S.n618 VSUBS 0.23fF $ **FLOATING
C723 S.n619 VSUBS 0.87fF $ **FLOATING
C724 S.n620 VSUBS 0.05fF $ **FLOATING
C725 S.n621 VSUBS 2.79fF $ **FLOATING
C726 S.n622 VSUBS 1.78fF $ **FLOATING
C727 S.n623 VSUBS 0.11fF $ **FLOATING
C728 S.t24 VSUBS 0.02fF
C729 S.n624 VSUBS 0.13fF $ **FLOATING
C730 S.t180 VSUBS 0.02fF
C731 S.n626 VSUBS 0.23fF $ **FLOATING
C732 S.n627 VSUBS 0.34fF $ **FLOATING
C733 S.n628 VSUBS 0.58fF $ **FLOATING
C734 S.n629 VSUBS 0.88fF $ **FLOATING
C735 S.n630 VSUBS 0.30fF $ **FLOATING
C736 S.n631 VSUBS 0.88fF $ **FLOATING
C737 S.n632 VSUBS 1.03fF $ **FLOATING
C738 S.n633 VSUBS 0.15fF $ **FLOATING
C739 S.n634 VSUBS 4.45fF $ **FLOATING
C740 S.t88 VSUBS 0.02fF
C741 S.n635 VSUBS 0.11fF $ **FLOATING
C742 S.n636 VSUBS 0.13fF $ **FLOATING
C743 S.t61 VSUBS 0.02fF
C744 S.n638 VSUBS 0.23fF $ **FLOATING
C745 S.n639 VSUBS 0.87fF $ **FLOATING
C746 S.n640 VSUBS 0.05fF $ **FLOATING
C747 S.n641 VSUBS 0.10fF $ **FLOATING
C748 S.n642 VSUBS 0.11fF $ **FLOATING
C749 S.n643 VSUBS 0.09fF $ **FLOATING
C750 S.n644 VSUBS 0.11fF $ **FLOATING
C751 S.n645 VSUBS 0.17fF $ **FLOATING
C752 S.n646 VSUBS 1.78fF $ **FLOATING
C753 S.n647 VSUBS 0.11fF $ **FLOATING
C754 S.t81 VSUBS 0.02fF
C755 S.n648 VSUBS 0.13fF $ **FLOATING
C756 S.t79 VSUBS 0.02fF
C757 S.n650 VSUBS 1.16fF $ **FLOATING
C758 S.n651 VSUBS 0.06fF $ **FLOATING
C759 S.n652 VSUBS 0.09fF $ **FLOATING
C760 S.n653 VSUBS 0.57fF $ **FLOATING
C761 S.n654 VSUBS 2.30fF $ **FLOATING
C762 S.n655 VSUBS 2.35fF $ **FLOATING
C763 S.n656 VSUBS 4.07fF $ **FLOATING
C764 S.n657 VSUBS 0.24fF $ **FLOATING
C765 S.n658 VSUBS 0.01fF $ **FLOATING
C766 S.t104 VSUBS 0.02fF
C767 S.n659 VSUBS 0.24fF $ **FLOATING
C768 S.t140 VSUBS 0.02fF
C769 S.n660 VSUBS 0.90fF $ **FLOATING
C770 S.n661 VSUBS 0.67fF $ **FLOATING
C771 S.n662 VSUBS 1.79fF $ **FLOATING
C772 S.n663 VSUBS 1.78fF $ **FLOATING
C773 S.t130 VSUBS 0.02fF
C774 S.n664 VSUBS 0.23fF $ **FLOATING
C775 S.n665 VSUBS 0.34fF $ **FLOATING
C776 S.n666 VSUBS 0.58fF $ **FLOATING
C777 S.n667 VSUBS 0.11fF $ **FLOATING
C778 S.t156 VSUBS 0.02fF
C779 S.n668 VSUBS 0.13fF $ **FLOATING
C780 S.n670 VSUBS 1.10fF $ **FLOATING
C781 S.n671 VSUBS 0.21fF $ **FLOATING
C782 S.n672 VSUBS 0.24fF $ **FLOATING
C783 S.n673 VSUBS 0.08fF $ **FLOATING
C784 S.n674 VSUBS 1.79fF $ **FLOATING
C785 S.t2 VSUBS 0.02fF
C786 S.n675 VSUBS 0.23fF $ **FLOATING
C787 S.n676 VSUBS 0.87fF $ **FLOATING
C788 S.n677 VSUBS 0.05fF $ **FLOATING
C789 S.t40 VSUBS 0.02fF
C790 S.n678 VSUBS 0.11fF $ **FLOATING
C791 S.n679 VSUBS 0.13fF $ **FLOATING
C792 S.n681 VSUBS 0.73fF $ **FLOATING
C793 S.n682 VSUBS 0.42fF $ **FLOATING
C794 S.n683 VSUBS 1.50fF $ **FLOATING
C795 S.n684 VSUBS 0.11fF $ **FLOATING
C796 S.t48 VSUBS 0.02fF
C797 S.n685 VSUBS 0.13fF $ **FLOATING
C798 S.t33 VSUBS 0.02fF
C799 S.n687 VSUBS 0.23fF $ **FLOATING
C800 S.n688 VSUBS 0.34fF $ **FLOATING
C801 S.n689 VSUBS 0.58fF $ **FLOATING
C802 S.n690 VSUBS 0.01fF $ **FLOATING
C803 S.n691 VSUBS 0.06fF $ **FLOATING
C804 S.n692 VSUBS 0.01fF $ **FLOATING
C805 S.n693 VSUBS 0.01fF $ **FLOATING
C806 S.n694 VSUBS 0.01fF $ **FLOATING
C807 S.n695 VSUBS 0.23fF $ **FLOATING
C808 S.n696 VSUBS 1.10fF $ **FLOATING
C809 S.n697 VSUBS 1.27fF $ **FLOATING
C810 S.n698 VSUBS 1.89fF $ **FLOATING
C811 S.t119 VSUBS 0.02fF
C812 S.n699 VSUBS 0.23fF $ **FLOATING
C813 S.n700 VSUBS 0.87fF $ **FLOATING
C814 S.n701 VSUBS 0.05fF $ **FLOATING
C815 S.t12 VSUBS 0.02fF
C816 S.n702 VSUBS 0.11fF $ **FLOATING
C817 S.n703 VSUBS 0.13fF $ **FLOATING
C818 S.n705 VSUBS 1.78fF $ **FLOATING
C819 S.n706 VSUBS 0.11fF $ **FLOATING
C820 S.t27 VSUBS 0.02fF
C821 S.n707 VSUBS 0.13fF $ **FLOATING
C822 S.t184 VSUBS 0.02fF
C823 S.n709 VSUBS 0.23fF $ **FLOATING
C824 S.n710 VSUBS 0.34fF $ **FLOATING
C825 S.n711 VSUBS 0.58fF $ **FLOATING
C826 S.n712 VSUBS 0.30fF $ **FLOATING
C827 S.n713 VSUBS 1.03fF $ **FLOATING
C828 S.n714 VSUBS 0.15fF $ **FLOATING
C829 S.n715 VSUBS 1.99fF $ **FLOATING
C830 S.t93 VSUBS 0.02fF
C831 S.n716 VSUBS 0.11fF $ **FLOATING
C832 S.n717 VSUBS 0.13fF $ **FLOATING
C833 S.t63 VSUBS 0.02fF
C834 S.n719 VSUBS 0.23fF $ **FLOATING
C835 S.n720 VSUBS 0.87fF $ **FLOATING
C836 S.n721 VSUBS 0.05fF $ **FLOATING
C837 S.t11 VSUBS 13.78fF
C838 S.t144 VSUBS 0.02fF
C839 S.n722 VSUBS 0.11fF $ **FLOATING
C840 S.n723 VSUBS 0.13fF $ **FLOATING
C841 S.t117 VSUBS 0.02fF
C842 S.n725 VSUBS 0.23fF $ **FLOATING
C843 S.n726 VSUBS 0.87fF $ **FLOATING
C844 S.n727 VSUBS 0.05fF $ **FLOATING
C845 S.t55 VSUBS 0.02fF
C846 S.n728 VSUBS 0.23fF $ **FLOATING
C847 S.n729 VSUBS 0.34fF $ **FLOATING
C848 S.n730 VSUBS 0.58fF $ **FLOATING
C849 S.n731 VSUBS 2.52fF $ **FLOATING
C850 S.n732 VSUBS 3.12fF $ **FLOATING
C851 S.n733 VSUBS 0.10fF $ **FLOATING
C852 S.n734 VSUBS 0.34fF $ **FLOATING
C853 S.n735 VSUBS 0.44fF $ **FLOATING
C854 S.n736 VSUBS 1.08fF $ **FLOATING
C855 S.n737 VSUBS 1.78fF $ **FLOATING
C856 S.n738 VSUBS 0.11fF $ **FLOATING
C857 S.t76 VSUBS 0.02fF
C858 S.n739 VSUBS 0.13fF $ **FLOATING
C859 S.t53 VSUBS 0.02fF
C860 S.n741 VSUBS 0.23fF $ **FLOATING
C861 S.n742 VSUBS 0.34fF $ **FLOATING
C862 S.n743 VSUBS 0.58fF $ **FLOATING
C863 S.n744 VSUBS 1.21fF $ **FLOATING
C864 S.n745 VSUBS 2.26fF $ **FLOATING
C865 S.n746 VSUBS 3.99fF $ **FLOATING
C866 S.t142 VSUBS 0.02fF
C867 S.n747 VSUBS 0.11fF $ **FLOATING
C868 S.n748 VSUBS 0.13fF $ **FLOATING
C869 S.t114 VSUBS 0.02fF
C870 S.n750 VSUBS 0.23fF $ **FLOATING
C871 S.n751 VSUBS 0.87fF $ **FLOATING
C872 S.n752 VSUBS 0.05fF $ **FLOATING
C873 S.t23 VSUBS 13.41fF
C874 S.t141 VSUBS 0.02fF
C875 S.n753 VSUBS 0.01fF $ **FLOATING
C876 S.n754 VSUBS 0.24fF $ **FLOATING
C877 S.t134 VSUBS 0.02fF
C878 S.n756 VSUBS 1.14fF $ **FLOATING
C879 S.n757 VSUBS 0.05fF $ **FLOATING
C880 S.t110 VSUBS 0.02fF
C881 S.n758 VSUBS 0.61fF $ **FLOATING
C882 S.n759 VSUBS 0.58fF $ **FLOATING
C883 S.n760 VSUBS 1.42fF $ **FLOATING
C884 S.n761 VSUBS 0.02fF $ **FLOATING
C885 S.n762 VSUBS 0.01fF $ **FLOATING
C886 S.n763 VSUBS 0.01fF $ **FLOATING
C887 S.n764 VSUBS 0.01fF $ **FLOATING
C888 S.n765 VSUBS 0.01fF $ **FLOATING
C889 S.n766 VSUBS 0.02fF $ **FLOATING
C890 S.n767 VSUBS 0.02fF $ **FLOATING
C891 S.n768 VSUBS 0.03fF $ **FLOATING
C892 S.n769 VSUBS 0.15fF $ **FLOATING
C893 S.n770 VSUBS 0.10fF $ **FLOATING
C894 S.n771 VSUBS 0.16fF $ **FLOATING
C895 S.n772 VSUBS 0.14fF $ **FLOATING
C896 S.n773 VSUBS 0.26fF $ **FLOATING
C897 S.n774 VSUBS 0.23fF $ **FLOATING
C898 S.n775 VSUBS 4.45fF $ **FLOATING
C899 S.n776 VSUBS 8.82fF $ **FLOATING
C900 S.n777 VSUBS 8.88fF $ **FLOATING
C901 S.n778 VSUBS 11.78fF $ **FLOATING
C902 D.n0 VSUBS 1.26fF $ **FLOATING
C903 D.n1 VSUBS 1.26fF $ **FLOATING
C904 D.n2 VSUBS 3.86fF $ **FLOATING
C905 D.n3 VSUBS 7.00fF $ **FLOATING
C906 D.n4 VSUBS 8.26fF $ **FLOATING
C907 D.n5 VSUBS 16.73fF $ **FLOATING
C908 D.n6 VSUBS 6.03fF $ **FLOATING
C909 D.n7 VSUBS 4.47fF $ **FLOATING
C910 D.n8 VSUBS 10.52fF $ **FLOATING
C911 D.n9 VSUBS 11.39fF $ **FLOATING
C912 D.n10 VSUBS 10.37fF $ **FLOATING
C913 D.n11 VSUBS 10.37fF $ **FLOATING
C914 D.n12 VSUBS 5.27fF $ **FLOATING
C915 D.n13 VSUBS 5.11fF $ **FLOATING
C916 D.n14 VSUBS 8.38fF $ **FLOATING
C917 D.n15 VSUBS 7.56fF $ **FLOATING
C918 D.n16 VSUBS 12.28fF $ **FLOATING
C919 D.n17 VSUBS 7.64fF $ **FLOATING
C920 D.n18 VSUBS 0.19fF $ **FLOATING
C921 D.n19 VSUBS 3.91fF $ **FLOATING
C922 D.n20 VSUBS 0.20fF $ **FLOATING
C923 D.n21 VSUBS 4.36fF $ **FLOATING
C924 D.n22 VSUBS 0.20fF $ **FLOATING
C925 D.n23 VSUBS 4.11fF $ **FLOATING
C926 D.n24 VSUBS 0.20fF $ **FLOATING
C927 D.n25 VSUBS 4.42fF $ **FLOATING
C928 D.n26 VSUBS 0.20fF $ **FLOATING
C929 D.n27 VSUBS 4.00fF $ **FLOATING
C930 D.n28 VSUBS 0.20fF $ **FLOATING
C931 D.n29 VSUBS 4.00fF $ **FLOATING
C932 D.n30 VSUBS 0.20fF $ **FLOATING
C933 D.n31 VSUBS 4.00fF $ **FLOATING
C934 D.n32 VSUBS 0.20fF $ **FLOATING
C935 D.n33 VSUBS 4.01fF $ **FLOATING
C936 D.n34 VSUBS 0.20fF $ **FLOATING
C937 D.n35 VSUBS 3.92fF $ **FLOATING
C938 D.n36 VSUBS 0.20fF $ **FLOATING
C939 D.n37 VSUBS 4.22fF $ **FLOATING
C940 D.n38 VSUBS 0.20fF $ **FLOATING
C941 D.n39 VSUBS 4.02fF $ **FLOATING
C942 D.n40 VSUBS 0.20fF $ **FLOATING
C943 D.n41 VSUBS 4.02fF $ **FLOATING
C944 D.n42 VSUBS 0.20fF $ **FLOATING
C945 D.n43 VSUBS 4.02fF $ **FLOATING
C946 D.n44 VSUBS 0.20fF $ **FLOATING
C947 D.n45 VSUBS 4.22fF $ **FLOATING
C948 D.n46 VSUBS 0.20fF $ **FLOATING
C949 D.n47 VSUBS 4.00fF $ **FLOATING
C950 D.n48 VSUBS 0.20fF $ **FLOATING
C951 D.n49 VSUBS 4.00fF $ **FLOATING
C952 D.n50 VSUBS 0.20fF $ **FLOATING
C953 D.n51 VSUBS 4.00fF $ **FLOATING
C954 D.n52 VSUBS 0.20fF $ **FLOATING
C955 D.n53 VSUBS 4.00fF $ **FLOATING
C956 D.n54 VSUBS 0.20fF $ **FLOATING
C957 D.n55 VSUBS 4.00fF $ **FLOATING
C958 D.n56 VSUBS 0.20fF $ **FLOATING
C959 D.n57 VSUBS 4.00fF $ **FLOATING
C960 D.n58 VSUBS 0.20fF $ **FLOATING
C961 D.n59 VSUBS 3.22fF $ **FLOATING
C962 D.n60 VSUBS 0.20fF $ **FLOATING
C963 D.n61 VSUBS 5.48fF $ **FLOATING
C964 D.n62 VSUBS 0.20fF $ **FLOATING
C965 D.n63 VSUBS 4.97fF $ **FLOATING
C966 D.n64 VSUBS 0.20fF $ **FLOATING
C967 D.n65 VSUBS 4.41fF $ **FLOATING
C968 D.n66 VSUBS 0.20fF $ **FLOATING
C969 D.n67 VSUBS 4.48fF $ **FLOATING
C970 D.n68 VSUBS 0.20fF $ **FLOATING
C971 D.n69 VSUBS 4.48fF $ **FLOATING
C972 D.n70 VSUBS 0.20fF $ **FLOATING
C973 D.n71 VSUBS 4.48fF $ **FLOATING
C974 D.n72 VSUBS 0.20fF $ **FLOATING
C975 D.n73 VSUBS 5.48fF $ **FLOATING
C976 D.n74 VSUBS 0.20fF $ **FLOATING
C977 D.n75 VSUBS 4.97fF $ **FLOATING
C978 D.n76 VSUBS 0.20fF $ **FLOATING
C979 D.n77 VSUBS 3.85fF $ **FLOATING
C980 D.n78 VSUBS 0.20fF $ **FLOATING
C981 D.n79 VSUBS 4.48fF $ **FLOATING
C982 D.n80 VSUBS 0.20fF $ **FLOATING
C983 D.n81 VSUBS 3.53fF $ **FLOATING
C984 D.n82 VSUBS 0.59fF $ **FLOATING
C985 D.n83 VSUBS 0.75fF $ **FLOATING
C986 D.n84 VSUBS 0.25fF $ **FLOATING
C987 D.n85 VSUBS 0.25fF $ **FLOATING
C988 D.n86 VSUBS 0.25fF $ **FLOATING
C989 D.n87 VSUBS 26.03fF $ **FLOATING
C990 D.n88 VSUBS 0.25fF $ **FLOATING
C991 D.n89 VSUBS 6.06fF $ **FLOATING
C992 D.n90 VSUBS 4.31fF $ **FLOATING
C993 D.n91 VSUBS 3.16fF $ **FLOATING
C994 D.n92 VSUBS 1.34fF $ **FLOATING
C995 D.n93 VSUBS 8.80fF $ **FLOATING
C996 D.t139 VSUBS -0.01fF
C997 D.t70 VSUBS 0.00fF
C998 D.n94 VSUBS 1.69fF $ **FLOATING
C999 D.t63 VSUBS -0.06fF
C1000 D.n95 VSUBS 0.59fF $ **FLOATING
C1001 D.t23 VSUBS -0.02fF
C1002 D.t64 VSUBS -0.02fF
C1003 D.t97 VSUBS -0.06fF
C1004 D.n96 VSUBS 0.59fF $ **FLOATING
C1005 D.n97 VSUBS 2.09fF $ **FLOATING
C1006 D.n98 VSUBS 1.80fF $ **FLOATING
C1007 D.t166 VSUBS -0.06fF
C1008 D.n99 VSUBS 0.59fF $ **FLOATING
C1009 D.t32 VSUBS -0.02fF
C1010 D.t74 VSUBS -0.02fF
C1011 D.t66 VSUBS -0.06fF
C1012 D.n100 VSUBS 0.59fF $ **FLOATING
C1013 D.n101 VSUBS 2.20fF $ **FLOATING
C1014 D.n102 VSUBS 1.80fF $ **FLOATING
C1015 D.t168 VSUBS -0.06fF
C1016 D.n103 VSUBS 0.59fF $ **FLOATING
C1017 D.t148 VSUBS -0.02fF
C1018 D.t72 VSUBS -0.02fF
C1019 D.t27 VSUBS -0.06fF
C1020 D.n104 VSUBS 0.59fF $ **FLOATING
C1021 D.n105 VSUBS 2.20fF $ **FLOATING
C1022 D.n106 VSUBS 1.80fF $ **FLOATING
C1023 D.t156 VSUBS -0.06fF
C1024 D.n107 VSUBS 0.59fF $ **FLOATING
C1025 D.t176 VSUBS -0.02fF
C1026 D.t47 VSUBS -0.02fF
C1027 D.t26 VSUBS -0.06fF
C1028 D.n108 VSUBS 0.59fF $ **FLOATING
C1029 D.n109 VSUBS 2.20fF $ **FLOATING
C1030 D.n110 VSUBS 1.80fF $ **FLOATING
C1031 D.t158 VSUBS -0.06fF
C1032 D.n111 VSUBS 0.59fF $ **FLOATING
C1033 D.t143 VSUBS -0.02fF
C1034 D.t81 VSUBS -0.02fF
C1035 D.t104 VSUBS -0.06fF
C1036 D.n112 VSUBS 0.59fF $ **FLOATING
C1037 D.n113 VSUBS 2.20fF $ **FLOATING
C1038 D.n114 VSUBS 1.80fF $ **FLOATING
C1039 D.t40 VSUBS -0.06fF
C1040 D.n115 VSUBS 0.59fF $ **FLOATING
C1041 D.t165 VSUBS -0.02fF
C1042 D.t96 VSUBS -0.02fF
C1043 D.t102 VSUBS -0.06fF
C1044 D.n116 VSUBS 0.59fF $ **FLOATING
C1045 D.n117 VSUBS 2.20fF $ **FLOATING
C1046 D.n118 VSUBS 2.27fF $ **FLOATING
C1047 D.t119 VSUBS -0.06fF
C1048 D.n119 VSUBS 0.59fF $ **FLOATING
C1049 D.t138 VSUBS -0.02fF
C1050 D.t54 VSUBS -0.02fF
C1051 D.t101 VSUBS -0.06fF
C1052 D.n120 VSUBS 0.59fF $ **FLOATING
C1053 D.n121 VSUBS 1.19fF $ **FLOATING
C1054 D.n122 VSUBS 1.88fF $ **FLOATING
C1055 D.n123 VSUBS 0.07fF $ **FLOATING
C1056 D.n124 VSUBS 0.43fF $ **FLOATING
C1057 D.n125 VSUBS 0.18fF $ **FLOATING
C1058 D.n126 VSUBS 0.13fF $ **FLOATING
C1059 D.t121 VSUBS -0.02fF
C1060 D.t134 VSUBS -0.06fF
C1061 D.n127 VSUBS 0.59fF $ **FLOATING
C1062 D.t115 VSUBS -0.02fF
C1063 D.t152 VSUBS -0.06fF
C1064 D.n128 VSUBS 0.59fF $ **FLOATING
C1065 D.n129 VSUBS 0.11fF $ **FLOATING
C1066 D.n130 VSUBS 0.09fF $ **FLOATING
C1067 D.n131 VSUBS 0.10fF $ **FLOATING
C1068 D.n132 VSUBS 0.61fF $ **FLOATING
C1069 D.n133 VSUBS 0.32fF $ **FLOATING
C1070 D.n134 VSUBS 4.03fF $ **FLOATING
C1071 D.n135 VSUBS 2.89fF $ **FLOATING
C1072 D.n136 VSUBS 3.16fF $ **FLOATING
C1073 D.n137 VSUBS 11.17fF $ **FLOATING
C1074 D.n138 VSUBS 1.28fF $ **FLOATING
C1075 D.n139 VSUBS 9.41fF $ **FLOATING
C1076 D.n140 VSUBS 9.33fF $ **FLOATING
C1077 D.n141 VSUBS 13.94fF $ **FLOATING
C1078 D.n142 VSUBS 1.96fF $ **FLOATING
C1079 D.n143 VSUBS 0.07fF $ **FLOATING
C1080 D.n144 VSUBS 0.23fF $ **FLOATING
C1081 D.t136 VSUBS 0.00fF
C1082 D.t117 VSUBS -0.01fF
C1083 D.n145 VSUBS 0.07fF $ **FLOATING
C1084 D.n146 VSUBS 0.10fF $ **FLOATING
C1085 D.n147 VSUBS 0.75fF $ **FLOATING
C1086 D.n148 VSUBS 0.05fF $ **FLOATING
C1087 D.n149 VSUBS 0.05fF $ **FLOATING
C1088 D.n150 VSUBS 1.59fF $ **FLOATING
C1089 D.n151 VSUBS 0.77fF $ **FLOATING
C1090 D.t38 VSUBS -0.02fF
C1091 D.t73 VSUBS -0.01fF
C1092 D.t113 VSUBS -0.02fF
C1093 D.n152 VSUBS 0.54fF $ **FLOATING
C1094 D.n153 VSUBS 0.19fF $ **FLOATING
C1095 D.n154 VSUBS 1.09fF $ **FLOATING
C1096 D.n155 VSUBS 1.96fF $ **FLOATING
C1097 D.n156 VSUBS 11.05fF $ **FLOATING
C1098 D.n157 VSUBS 13.78fF $ **FLOATING
C1099 D.n158 VSUBS 9.02fF $ **FLOATING
C1100 D.n159 VSUBS 2.09fF $ **FLOATING
C1101 D.t9 VSUBS 0.00fF
C1102 D.t133 VSUBS -0.06fF
C1103 D.t55 VSUBS 0.00fF
C1104 D.n160 VSUBS 0.32fF $ **FLOATING
C1105 D.n161 VSUBS 2.13fF $ **FLOATING
C1106 D.t90 VSUBS -0.06fF
C1107 D.n162 VSUBS 0.59fF $ **FLOATING
C1108 D.t48 VSUBS -0.02fF
C1109 D.t4 VSUBS -0.02fF
C1110 D.t169 VSUBS -0.06fF
C1111 D.n163 VSUBS 0.59fF $ **FLOATING
C1112 D.n164 VSUBS 1.29fF $ **FLOATING
C1113 D.n165 VSUBS 2.23fF $ **FLOATING
C1114 D.t58 VSUBS -0.06fF
C1115 D.n166 VSUBS 0.59fF $ **FLOATING
C1116 D.t82 VSUBS -0.02fF
C1117 D.t0 VSUBS -0.02fF
C1118 D.t157 VSUBS -0.06fF
C1119 D.n167 VSUBS 0.59fF $ **FLOATING
C1120 D.n168 VSUBS 0.73fF $ **FLOATING
C1121 D.n169 VSUBS 0.43fF $ **FLOATING
C1122 D.n170 VSUBS 0.24fF $ **FLOATING
C1123 D.n171 VSUBS 2.02fF $ **FLOATING
C1124 D.t78 VSUBS -0.06fF
C1125 D.n172 VSUBS 0.59fF $ **FLOATING
C1126 D.t95 VSUBS -0.02fF
C1127 D.t13 VSUBS -0.02fF
C1128 D.t159 VSUBS -0.06fF
C1129 D.n173 VSUBS 0.59fF $ **FLOATING
C1130 D.n174 VSUBS 0.73fF $ **FLOATING
C1131 D.n175 VSUBS 0.43fF $ **FLOATING
C1132 D.n176 VSUBS 0.24fF $ **FLOATING
C1133 D.n177 VSUBS 2.28fF $ **FLOATING
C1134 D.t87 VSUBS -0.06fF
C1135 D.n178 VSUBS 0.59fF $ **FLOATING
C1136 D.t53 VSUBS -0.02fF
C1137 D.t110 VSUBS -0.02fF
C1138 D.t39 VSUBS -0.06fF
C1139 D.n179 VSUBS 0.59fF $ **FLOATING
C1140 D.n180 VSUBS 0.73fF $ **FLOATING
C1141 D.n181 VSUBS 0.43fF $ **FLOATING
C1142 D.n182 VSUBS 0.24fF $ **FLOATING
C1143 D.n183 VSUBS 2.28fF $ **FLOATING
C1144 D.t86 VSUBS -0.06fF
C1145 D.n184 VSUBS 0.59fF $ **FLOATING
C1146 D.t7 VSUBS -0.02fF
C1147 D.t67 VSUBS -0.02fF
C1148 D.t149 VSUBS -0.06fF
C1149 D.n185 VSUBS 0.59fF $ **FLOATING
C1150 D.n186 VSUBS 0.73fF $ **FLOATING
C1151 D.n187 VSUBS 0.43fF $ **FLOATING
C1152 D.n188 VSUBS 0.24fF $ **FLOATING
C1153 D.n189 VSUBS 2.28fF $ **FLOATING
C1154 D.t99 VSUBS -0.06fF
C1155 D.n190 VSUBS 0.59fF $ **FLOATING
C1156 D.t11 VSUBS -0.02fF
C1157 D.t44 VSUBS -0.02fF
C1158 D.t106 VSUBS -0.06fF
C1159 D.n191 VSUBS 0.59fF $ **FLOATING
C1160 D.n192 VSUBS 0.73fF $ **FLOATING
C1161 D.n193 VSUBS 0.43fF $ **FLOATING
C1162 D.n194 VSUBS 0.24fF $ **FLOATING
C1163 D.n195 VSUBS 0.80fF $ **FLOATING
C1164 D.n196 VSUBS 0.43fF $ **FLOATING
C1165 D.n197 VSUBS 0.65fF $ **FLOATING
C1166 D.t142 VSUBS -0.02fF
C1167 D.t83 VSUBS -0.01fF
C1168 D.t19 VSUBS -0.02fF
C1169 D.n198 VSUBS 0.54fF $ **FLOATING
C1170 D.n199 VSUBS 9.02fF $ **FLOATING
C1171 D.n200 VSUBS 2.09fF $ **FLOATING
C1172 D.t178 VSUBS 0.00fF
C1173 D.t21 VSUBS -0.06fF
C1174 D.t14 VSUBS 0.00fF
C1175 D.n201 VSUBS 0.32fF $ **FLOATING
C1176 D.n202 VSUBS 2.13fF $ **FLOATING
C1177 D.t22 VSUBS -0.06fF
C1178 D.n203 VSUBS 0.59fF $ **FLOATING
C1179 D.t15 VSUBS -0.02fF
C1180 D.t177 VSUBS -0.02fF
C1181 D.t77 VSUBS -0.06fF
C1182 D.n204 VSUBS 0.59fF $ **FLOATING
C1183 D.n205 VSUBS 1.29fF $ **FLOATING
C1184 D.n206 VSUBS 2.23fF $ **FLOATING
C1185 D.t105 VSUBS -0.06fF
C1186 D.n207 VSUBS 0.59fF $ **FLOATING
C1187 D.t16 VSUBS -0.02fF
C1188 D.t175 VSUBS -0.02fF
C1189 D.t50 VSUBS -0.06fF
C1190 D.n208 VSUBS 0.59fF $ **FLOATING
C1191 D.n209 VSUBS 0.73fF $ **FLOATING
C1192 D.n210 VSUBS 0.43fF $ **FLOATING
C1193 D.n211 VSUBS 0.24fF $ **FLOATING
C1194 D.n212 VSUBS 2.02fF $ **FLOATING
C1195 D.t100 VSUBS -0.06fF
C1196 D.n213 VSUBS 0.59fF $ **FLOATING
C1197 D.t43 VSUBS -0.02fF
C1198 D.t164 VSUBS -0.02fF
C1199 D.t75 VSUBS -0.06fF
C1200 D.n214 VSUBS 0.59fF $ **FLOATING
C1201 D.n215 VSUBS 0.73fF $ **FLOATING
C1202 D.n216 VSUBS 0.43fF $ **FLOATING
C1203 D.n217 VSUBS 0.24fF $ **FLOATING
C1204 D.n218 VSUBS 2.28fF $ **FLOATING
C1205 D.t151 VSUBS -0.06fF
C1206 D.n219 VSUBS 0.59fF $ **FLOATING
C1207 D.t36 VSUBS -0.02fF
C1208 D.t173 VSUBS -0.02fF
C1209 D.t155 VSUBS -0.06fF
C1210 D.n220 VSUBS 0.59fF $ **FLOATING
C1211 D.n221 VSUBS 0.94fF $ **FLOATING
C1212 D.n222 VSUBS 0.13fF $ **FLOATING
C1213 D.n223 VSUBS 0.73fF $ **FLOATING
C1214 D.n224 VSUBS 0.43fF $ **FLOATING
C1215 D.n225 VSUBS 0.24fF $ **FLOATING
C1216 D.n226 VSUBS 18.51fF $ **FLOATING
C1217 D.n227 VSUBS 2.10fF $ **FLOATING
C1218 D.t30 VSUBS -0.02fF
C1219 D.n228 VSUBS 0.54fF $ **FLOATING
C1220 D.t8 VSUBS -0.02fF
C1221 D.t24 VSUBS -0.01fF
C1222 D.t42 VSUBS -0.06fF
C1223 D.t144 VSUBS 0.00fF
C1224 D.t98 VSUBS 0.00fF
C1225 D.n229 VSUBS 0.32fF $ **FLOATING
C1226 D.n230 VSUBS 2.59fF $ **FLOATING
C1227 D.t108 VSUBS -0.06fF
C1228 D.n231 VSUBS 0.59fF $ **FLOATING
C1229 D.t172 VSUBS -0.02fF
C1230 D.t51 VSUBS -0.02fF
C1231 D.t103 VSUBS -0.06fF
C1232 D.n232 VSUBS 0.59fF $ **FLOATING
C1233 D.n233 VSUBS 2.66fF $ **FLOATING
C1234 D.t141 VSUBS -0.02fF
C1235 D.t109 VSUBS -0.06fF
C1236 D.n234 VSUBS 0.59fF $ **FLOATING
C1237 D.t52 VSUBS -0.02fF
C1238 D.t154 VSUBS -0.06fF
C1239 D.n235 VSUBS 0.59fF $ **FLOATING
C1240 D.n236 VSUBS 2.01fF $ **FLOATING
C1241 D.n237 VSUBS 2.58fF $ **FLOATING
C1242 D.n238 VSUBS 18.52fF $ **FLOATING
C1243 D.n239 VSUBS 1.81fF $ **FLOATING
C1244 D.n240 VSUBS 4.83fF $ **FLOATING
C1245 D.t35 VSUBS -0.02fF
C1246 D.t29 VSUBS -0.01fF
C1247 D.t10 VSUBS -0.02fF
C1248 D.n241 VSUBS 0.54fF $ **FLOATING
C1249 D.n242 VSUBS 4.80fF $ **FLOATING
C1250 D.t5 VSUBS -0.06fF
C1251 D.t93 VSUBS 0.00fF
C1252 D.t68 VSUBS 0.00fF
C1253 D.n243 VSUBS 0.32fF $ **FLOATING
C1254 D.n244 VSUBS 16.11fF $ **FLOATING
C1255 D.n245 VSUBS 7.77fF $ **FLOATING
C1256 D.n246 VSUBS 7.77fF $ **FLOATING
C1257 D.n247 VSUBS 8.80fF $ **FLOATING
C1258 D.n248 VSUBS 0.12fF $ **FLOATING
C1259 D.n249 VSUBS 0.67fF $ **FLOATING
C1260 D.n250 VSUBS 16.34fF $ **FLOATING
C1261 D.n251 VSUBS 4.69fF $ **FLOATING
C1262 D.n252 VSUBS 0.23fF $ **FLOATING
C1263 D.t18 VSUBS 0.00fF
C1264 D.t128 VSUBS -0.06fF
C1265 D.t69 VSUBS 0.00fF
C1266 D.n253 VSUBS 0.32fF $ **FLOATING
C1267 D.t122 VSUBS -0.02fF
C1268 D.t150 VSUBS -0.01fF
C1269 D.t33 VSUBS -0.02fF
C1270 D.n254 VSUBS 0.54fF $ **FLOATING
C1271 D.n255 VSUBS 4.62fF $ **FLOATING
C1272 D.n256 VSUBS 0.04fF $ **FLOATING
C1273 D.n257 VSUBS 0.09fF $ **FLOATING
C1274 D.n258 VSUBS 2.43fF $ **FLOATING
C1275 D.n259 VSUBS 1.83fF $ **FLOATING
C1276 D.t123 VSUBS -0.06fF
C1277 D.n260 VSUBS 0.59fF $ **FLOATING
C1278 D.t84 VSUBS -0.02fF
C1279 D.t91 VSUBS -0.02fF
C1280 D.t17 VSUBS -0.06fF
C1281 D.n261 VSUBS 0.59fF $ **FLOATING
C1282 D.n262 VSUBS 0.26fF $ **FLOATING
C1283 D.n263 VSUBS 0.13fF $ **FLOATING
C1284 D.n264 VSUBS 0.71fF $ **FLOATING
C1285 D.n265 VSUBS 1.10fF $ **FLOATING
C1286 D.n266 VSUBS 1.73fF $ **FLOATING
C1287 D.t94 VSUBS -0.02fF
C1288 D.n267 VSUBS 0.54fF $ **FLOATING
C1289 D.t140 VSUBS -0.02fF
C1290 D.t46 VSUBS -0.01fF
C1291 D.n268 VSUBS 1.71fF $ **FLOATING
C1292 D.n269 VSUBS 1.16fF $ **FLOATING
C1293 D.n270 VSUBS 1.87fF $ **FLOATING
C1294 D.t118 VSUBS -0.02fF
C1295 D.n271 VSUBS 0.01fF $ **FLOATING
C1296 D.t80 VSUBS -0.06fF
C1297 D.n273 VSUBS 0.58fF $ **FLOATING
C1298 D.t61 VSUBS -0.06fF
C1299 D.n274 VSUBS 0.59fF $ **FLOATING
C1300 D.t131 VSUBS -0.02fF
C1301 D.t116 VSUBS -0.06fF
C1302 D.t37 VSUBS 0.00fF
C1303 D.t137 VSUBS 0.00fF
C1304 D.n275 VSUBS 0.32fF $ **FLOATING
C1305 D.n276 VSUBS 1.85fF $ **FLOATING
C1306 D.n277 VSUBS 0.09fF $ **FLOATING
C1307 D.n278 VSUBS 1.71fF $ **FLOATING
C1308 D.n279 VSUBS 0.09fF $ **FLOATING
C1309 D.n280 VSUBS 0.81fF $ **FLOATING
C1310 D.t153 VSUBS -0.02fF
C1311 D.n281 VSUBS 0.54fF $ **FLOATING
C1312 D.t146 VSUBS -0.02fF
C1313 D.t135 VSUBS -0.01fF
C1314 D.n282 VSUBS 0.26fF $ **FLOATING
C1315 D.n283 VSUBS 0.13fF $ **FLOATING
C1316 D.n284 VSUBS 0.88fF $ **FLOATING
C1317 D.t107 VSUBS -0.02fF
C1318 D.t28 VSUBS -0.06fF
C1319 D.n285 VSUBS 0.59fF $ **FLOATING
C1320 D.t20 VSUBS -0.02fF
C1321 D.t145 VSUBS -0.06fF
C1322 D.n286 VSUBS 0.59fF $ **FLOATING
C1323 D.n287 VSUBS 2.06fF $ **FLOATING
C1324 D.n288 VSUBS 1.70fF $ **FLOATING
C1325 D.n289 VSUBS 1.67fF $ **FLOATING
C1326 D.t59 VSUBS -0.06fF
C1327 D.n290 VSUBS 0.59fF $ **FLOATING
C1328 D.t71 VSUBS -0.02fF
C1329 D.t76 VSUBS -0.02fF
C1330 D.t171 VSUBS -0.06fF
C1331 D.n291 VSUBS 0.59fF $ **FLOATING
C1332 D.n292 VSUBS 2.20fF $ **FLOATING
C1333 D.n293 VSUBS 1.80fF $ **FLOATING
C1334 D.t130 VSUBS -0.06fF
C1335 D.n294 VSUBS 0.59fF $ **FLOATING
C1336 D.t56 VSUBS -0.02fF
C1337 D.t3 VSUBS -0.02fF
C1338 D.t167 VSUBS -0.06fF
C1339 D.n295 VSUBS 0.59fF $ **FLOATING
C1340 D.n296 VSUBS 2.20fF $ **FLOATING
C1341 D.n297 VSUBS 2.32fF $ **FLOATING
C1342 D.t79 VSUBS -0.06fF
C1343 D.n298 VSUBS 0.59fF $ **FLOATING
C1344 D.t114 VSUBS -0.02fF
C1345 D.t126 VSUBS -0.02fF
C1346 D.t161 VSUBS -0.06fF
C1347 D.n299 VSUBS 0.59fF $ **FLOATING
C1348 D.n300 VSUBS 1.88fF $ **FLOATING
C1349 D.n301 VSUBS 1.15fF $ **FLOATING
C1350 D.n302 VSUBS 0.03fF $ **FLOATING
C1351 D.n303 VSUBS 0.04fF $ **FLOATING
C1352 D.n304 VSUBS 24.73fF $ **FLOATING
C1353 D.n305 VSUBS 0.07fF $ **FLOATING
C1354 D.n306 VSUBS 0.10fF $ **FLOATING
C1355 D.n307 VSUBS 0.11fF $ **FLOATING
C1356 D.t129 VSUBS -0.06fF
C1357 D.t163 VSUBS 0.00fF
C1358 D.t12 VSUBS 0.00fF
C1359 D.n308 VSUBS 0.32fF $ **FLOATING
C1360 D.n309 VSUBS 0.55fF $ **FLOATING
C1361 D.n310 VSUBS 7.24fF $ **FLOATING
C1362 D.n311 VSUBS 0.04fF $ **FLOATING
C1363 D.n312 VSUBS 0.09fF $ **FLOATING
C1364 D.n313 VSUBS 0.67fF $ **FLOATING
C1365 D.n314 VSUBS 0.26fF $ **FLOATING
C1366 D.n315 VSUBS 0.13fF $ **FLOATING
C1367 D.n316 VSUBS 1.11fF $ **FLOATING
C1368 D.n317 VSUBS 1.70fF $ **FLOATING
C1369 D.t132 VSUBS -0.02fF
C1370 D.t174 VSUBS -0.06fF
C1371 D.n318 VSUBS 0.59fF $ **FLOATING
C1372 D.t162 VSUBS -0.02fF
C1373 D.t160 VSUBS -0.06fF
C1374 D.n319 VSUBS 0.59fF $ **FLOATING
C1375 D.n320 VSUBS 2.06fF $ **FLOATING
C1376 D.t62 VSUBS -0.02fF
C1377 D.n321 VSUBS 0.54fF $ **FLOATING
C1378 D.t41 VSUBS -0.02fF
C1379 D.t6 VSUBS -0.01fF
C1380 D.n322 VSUBS 1.71fF $ **FLOATING
C1381 D.n323 VSUBS 1.67fF $ **FLOATING
C1382 D.t65 VSUBS -0.06fF
C1383 D.n324 VSUBS 0.59fF $ **FLOATING
C1384 D.t2 VSUBS -0.02fF
C1385 D.t85 VSUBS -0.02fF
C1386 D.t60 VSUBS -0.06fF
C1387 D.n325 VSUBS 0.59fF $ **FLOATING
C1388 D.n326 VSUBS 2.20fF $ **FLOATING
C1389 D.n327 VSUBS 1.80fF $ **FLOATING
C1390 D.t92 VSUBS -0.06fF
C1391 D.n328 VSUBS 0.59fF $ **FLOATING
C1392 D.t112 VSUBS -0.02fF
C1393 D.t31 VSUBS -0.02fF
C1394 D.t89 VSUBS -0.06fF
C1395 D.n329 VSUBS 0.59fF $ **FLOATING
C1396 D.n330 VSUBS 2.20fF $ **FLOATING
C1397 D.n331 VSUBS 1.80fF $ **FLOATING
C1398 D.t25 VSUBS -0.06fF
C1399 D.n332 VSUBS 0.59fF $ **FLOATING
C1400 D.t1 VSUBS -0.02fF
C1401 D.t147 VSUBS -0.02fF
C1402 D.t57 VSUBS -0.06fF
C1403 D.n333 VSUBS 0.59fF $ **FLOATING
C1404 D.n334 VSUBS 2.20fF $ **FLOATING
C1405 D.n335 VSUBS 1.80fF $ **FLOATING
C1406 D.t125 VSUBS -0.06fF
C1407 D.n336 VSUBS 0.59fF $ **FLOATING
C1408 D.t111 VSUBS -0.02fF
C1409 D.t179 VSUBS -0.02fF
C1410 D.t49 VSUBS -0.06fF
C1411 D.n337 VSUBS 0.59fF $ **FLOATING
C1412 D.n338 VSUBS 2.20fF $ **FLOATING
C1413 D.n339 VSUBS 2.44fF $ **FLOATING
C1414 D.t170 VSUBS -0.06fF
C1415 D.n340 VSUBS 0.59fF $ **FLOATING
C1416 D.t127 VSUBS -0.02fF
C1417 D.t120 VSUBS -0.02fF
C1418 D.t88 VSUBS -0.06fF
C1419 D.n341 VSUBS 0.59fF $ **FLOATING
C1420 D.n342 VSUBS 1.15fF $ **FLOATING
C1421 D.n343 VSUBS 1.88fF $ **FLOATING
C1422 D.t124 VSUBS -0.06fF
C1423 D.t45 VSUBS 0.00fF
C1424 D.t34 VSUBS 0.00fF
C1425 D.n344 VSUBS 0.32fF $ **FLOATING
C1426 D.n345 VSUBS 1.85fF $ **FLOATING
C1427 D.n346 VSUBS 1.02fF $ **FLOATING
C1428 D.n347 VSUBS 7.05fF $ **FLOATING
.ends

