* NGSPICE file created from mag_files/POSTLAYOUT/nmos_flat_4x4.ext - technology: sky130A

.subckt nmos_flat_4x4 G S D DNW VSUBS
X0 S.t30 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1 S.t29 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2 S.t28 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3 D G S.t27 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X4 S.t26 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5 D G S.t25 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6 D G S.t24 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7 D G S.t23 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X8 D G S.t21 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9 S.t20 G D S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10 S.t19 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X11 D G S.t18 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12 D G S.t17 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X13 S.t16 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X14 S.t14 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X15 S.t13 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X16 D G S.t12 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X17 D G S.t10 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X18 S.t8 G D S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X19 D G S.t7 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X20 S.t6 G D S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X21 D G S.t4 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X22 S.t2 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X23 D G S.t1 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
R0 S.t15 S.t0 355.882
R1 S.n2 S.t3 310.588
R2 S.n1 S.t9 310.588
R3 S.t5 S.n111 300.235
R4 S.t11 S.n73 300.235
R5 S.t22 S.n30 300.235
R6 S.n52 S.n51 169.353
R7 S.n54 S.n53 137.98
R8 S.n70 S.n69 135.611
R9 S.n50 S.n49 129.387
R10 S.n64 S.n63 91.65
R11 S.n113 S.n112 91.389
R12 S.n19 S.n18 87.222
R13 S.n32 S.n31 86.961
R14 S.n43 S.t23 3.904
R15 S.n29 S.t17 3.904
R16 S.n86 S.n85 3.904
R17 S.n108 S.t21 3.904
R18 S.n105 S.n104 3.904
R19 S.n88 S.t1 3.904
R20 S.n21 S.t25 3.904
R21 S.n113 S.t24 3.904
R22 S.n109 S.t7 3.904
R23 S.n62 S.n61 3.904
R24 S.n80 S.t12 3.904
R25 S.n82 S.n81 3.904
R26 S.n76 S.t18 3.904
R27 S.n33 S.t27 3.904
R28 S.n32 S.t10 3.904
R29 S.n65 S.t4 3.904
R30 S.n74 S.t14 3.643
R31 S.n17 S.t16 3.643
R32 S.n16 S.t2 3.643
R33 S.n86 S.t6 3.643
R34 S.n108 S.n107 3.643
R35 S.n105 S.t20 3.643
R36 S.n88 S.n87 3.643
R37 S.n19 S.t29 3.643
R38 S.n20 S.t19 3.643
R39 S.n84 S.t8 3.643
R40 S.n62 S.t26 3.643
R41 S.n80 S.n79 3.643
R42 S.n82 S.t13 3.643
R43 S.n76 S.n75 3.643
R44 S.n42 S.t28 3.643
R45 S.n64 S.t30 3.643
R46 S.n1 S.n70 2.799
R47 S.n52 S.n50 2.511
R48 S.n7 S.n44 0.218
R49 S.n6 S.n55 0.172
R50 S.n118 S.n47 0.141
R51 S.n26 S.t15 0.123
R52 S.n118 S.n4 0.11
R53 S S.n118 0.09
R54 S.n3 S.n8 0.129
R55 S.n6 S.n2 0.083
R56 S.n28 S.n27 0.079
R57 S.n25 S.n23 0.076
R58 S.n71 S.n1 0.126
R59 S.n39 S.n38 0.071
R60 S.n4 S.n0 0.071
R61 S.t22 S.n34 0.068
R62 S.n6 S.n48 0.067
R63 S.n11 S.n10 0.067
R64 S.n6 S.n56 0.067
R65 S.n11 S.n9 0.067
R66 S.n98 S.n97 0.066
R67 S.n5 S.n92 0.063
R68 S.n99 S.n98 0.059
R69 S.n3 S.n16 0.055
R70 S.n4 S.n84 0.054
R71 S.n46 S.n7 0.054
R72 S.t22 S.n29 0.053
R73 S.t11 S.n65 0.052
R74 S.t11 S.n74 0.051
R75 S.n5 S.n103 0.05
R76 S.n5 S.n106 0.05
R77 S.n0 S.n83 0.05
R78 S.n58 S.n6 0.049
R79 S.n12 S.n11 0.048
R80 S.n14 S.n12 0.044
R81 S.n103 S.n102 0.043
R82 S.n1 S.n68 0.039
R83 S.n41 S.n39 0.039
R84 S.n2 S.n52 0.039
R85 S.t22 S.n33 0.036
R86 S.n110 S.n109 0.035
R87 S.t15 S.n21 0.035
R88 S.n37 S.n36 0.035
R89 S.t15 S.n20 0.034
R90 S.t22 S.n42 0.034
R91 S.n71 S.n66 0.032
R92 S.t5 S.n110 0.031
R93 S.n5 S.n90 0.031
R94 S.n0 S.n78 0.031
R95 S.n90 S.n89 0.031
R96 S.n78 S.n77 0.031
R97 S.n25 S.n24 0.029
R98 S.n4 S.n117 0.027
R99 S.n60 S.n59 0.026
R100 S.n58 S.n57 0.026
R101 S.n5 S.n96 0.026
R102 S.n7 S.n45 0.025
R103 S.n117 S.n116 0.024
R104 S.n60 S.n58 0.023
R105 S.n37 S.n35 0.023
R106 S.n115 S.n114 0.023
R107 S.n14 S.n13 0.022
R108 S.n102 S.n101 0.022
R109 S.n95 S.n94 0.021
R110 S.n103 S.n99 0.02
R111 S.t15 S.n14 0.019
R112 S S.n26 0.018
R113 S.n101 S.n100 0.018
R114 S.t15 S.n22 0.016
R115 S.n94 S.n93 0.015
R116 S.t22 S.n37 0.015
R117 S.n4 S.n60 0.01
R118 S.n4 S.n115 0.01
R119 S.n92 S.n91 0.008
R120 S.t15 S.n25 0.008
R121 S.t15 S.n15 0.005
R122 S.n106 S.n105 0.004
R123 S.n83 S.n82 0.004
R124 S.n89 S.n88 0.004
R125 S.n77 S.n76 0.004
R126 S.t11 S.n72 0.004
R127 S.t11 S.n71 0.004
R128 S.t5 S.n86 0.004
R129 S.t11 S.n62 0.004
R130 S.t22 S.n41 0.167
R131 S.n1 S.n67 0.041
R132 S.n2 S.n54 0.03
R133 S.n0 S.t11 0.005
R134 S.t11 S.n64 0.004
R135 S.t15 S.n19 0.004
R136 S.t5 S.n113 0.004
R137 S.n41 S.n40 0.003
R138 S.t5 S.n108 0.003
R139 S.n0 S.n80 0.003
R140 S.n47 S.n46 0.003
R141 S.n47 S.n28 0.003
R142 S.t5 S.n5 0.003
R143 S.t15 S.n17 0.003
R144 S.t22 S.n43 0.003
R145 S.t22 S.n32 0.003
R146 S.n47 S.t22 0.003
R147 S.t15 S.n3 0.003
R148 S.n4 S.t5 0.002
R149 S.n96 S.n95 0.002
C0 G S 225.81fF
C1 G DNW 1.44fF
C2 D S 55.77fF
C3 D DNW 82.22fF
C4 G D 56.67fF
C5 S DNW 240.69fF
C6 D SUB 1.96fF
C7 G SUB -26.44fF
C8 S SUB -68.86fF
C9 DNW SUB 1993.74fF $ **FLOATING
C10 S.n0 SUB 8.60fF
C11 S.n1 SUB 10.35fF
C12 S.n2 SUB 7.03fF
C13 S.t22 SUB 22.18fF
C14 S.n3 SUB 61.92fF
C15 S.t15 SUB 17.65fF
C16 S.t5 SUB 7.38fF
C17 S.n4 SUB 3.49fF
C18 S.t11 SUB 12.46fF
C19 S.n5 SUB 5.90fF
C20 S.n6 SUB 5.97fF
C21 S.n7 SUB 15.91fF
C22 S.n8 SUB 17.57fF
C23 S.n9 SUB 27.97fF
C24 S.n10 SUB 27.97fF
C25 S.n11 SUB 5.83fF
C26 S.n12 SUB 1.16fF
C27 S.n13 SUB 0.77fF
C28 S.n14 SUB 0.50fF
C29 S.n15 SUB 0.33fF
C30 S.t2 SUB 0.02fF
C31 S.n16 SUB 1.44fF
C32 S.t16 SUB 0.02fF
C33 S.n17 SUB 0.48fF
C34 S.n18 SUB 0.02fF
C35 S.t29 SUB 0.02fF
C36 S.n19 SUB 0.40fF
C37 S.t0 SUB 4.28fF
C38 S.t19 SUB 0.02fF
C39 S.n20 SUB 0.98fF
C40 S.t25 SUB 0.03fF
C41 S.n21 SUB 0.98fF
C42 S.n22 SUB 0.29fF
C43 S.n23 SUB 0.97fF
C44 S.n24 SUB 1.23fF
C45 S.n25 SUB 0.68fF
C46 S.n26 SUB 16.25fF
C47 S.n27 SUB 4.87fF
C48 S.n28 SUB 2.77fF
C49 S.t17 SUB 0.03fF
C50 S.n29 SUB 1.40fF
C51 S.n30 SUB 3.70fF
C52 S.t10 SUB 0.03fF
C53 S.n31 SUB 0.02fF
C54 S.n32 SUB 0.41fF
C55 S.t27 SUB 0.03fF
C56 S.n33 SUB 0.98fF
C57 S.n34 SUB 0.34fF
C58 S.n35 SUB 2.33fF
C59 S.n36 SUB 1.31fF
C60 S.n37 SUB 0.36fF
C61 S.n38 SUB 0.62fF
C62 S.n39 SUB 0.97fF
C63 S.n40 SUB 8.65fF
C64 S.n41 SUB 20.67fF
C65 S.t28 SUB 0.02fF
C66 S.n42 SUB 0.98fF
C67 S.t23 SUB 0.03fF
C68 S.n43 SUB 0.48fF
C69 S.n44 SUB 16.21fF
C70 S.n45 SUB 0.84fF
C71 S.n46 SUB 2.76fF
C72 S.n47 SUB 7.67fF
C73 S.n48 SUB 27.49fF
C74 S.t3 SUB 3.81fF
C75 S.n49 SUB 0.97fF
C76 S.n50 SUB 0.09fF
C77 S.n51 SUB 0.97fF
C78 S.n52 SUB 1.66fF
C79 S.n53 SUB 0.66fF
C80 S.n54 SUB 0.24fF
C81 S.n55 SUB 0.23fF
C82 S.n56 SUB 27.49fF
C83 S.n57 SUB 0.15fF
C84 S.n58 SUB 1.63fF
C85 S.n59 SUB 1.51fF
C86 S.n60 SUB 0.29fF
C87 S.n61 SUB 0.13fF
C88 S.t26 SUB 0.02fF
C89 S.n62 SUB 0.15fF
C90 S.n63 SUB 0.01fF
C91 S.t30 SUB 0.02fF
C92 S.n64 SUB 0.28fF
C93 S.t4 SUB 0.03fF
C94 S.n65 SUB 1.33fF
C95 S.n66 SUB 0.67fF
C96 S.n67 SUB 1.27fF
C97 S.n68 SUB 0.90fF
C98 S.n69 SUB 0.93fF
C99 S.n70 SUB 0.02fF
C100 S.t9 SUB 3.81fF
C101 S.n71 SUB 4.64fF
C102 S.n72 SUB 2.52fF
C103 S.n73 SUB 3.70fF
C104 S.t14 SUB 0.02fF
C105 S.n74 SUB 1.31fF
C106 S.n75 SUB 0.26fF
C107 S.t18 SUB 0.03fF
C108 S.n76 SUB 0.39fF
C109 S.n77 SUB 0.40fF
C110 S.n78 SUB 0.74fF
C111 S.t12 SUB 0.03fF
C112 S.n79 SUB 0.13fF
C113 S.n80 SUB 0.16fF
C114 S.n81 SUB 0.26fF
C115 S.t13 SUB 0.02fF
C116 S.n82 SUB 0.39fF
C117 S.n83 SUB 0.69fF
C118 S.t8 SUB 0.02fF
C119 S.n84 SUB 1.34fF
C120 S.n85 SUB 0.13fF
C121 S.t6 SUB 0.02fF
C122 S.n86 SUB 0.15fF
C123 S.n87 SUB 0.26fF
C124 S.t1 SUB 0.03fF
C125 S.n88 SUB 0.39fF
C126 S.n89 SUB 0.40fF
C127 S.n90 SUB 0.74fF
C128 S.n91 SUB 0.27fF
C129 S.n92 SUB 0.10fF
C130 S.n93 SUB 0.20fF
C131 S.n94 SUB 0.22fF
C132 S.n95 SUB 1.33fF
C133 S.n96 SUB 0.25fF
C134 S.n97 SUB 0.11fF
C135 S.n98 SUB 0.10fF
C136 S.n99 SUB 0.23fF
C137 S.n100 SUB 0.07fF
C138 S.n101 SUB 0.07fF
C139 S.n102 SUB 0.06fF
C140 S.n103 SUB 0.08fF
C141 S.n104 SUB 0.26fF
C142 S.t20 SUB 0.02fF
C143 S.n105 SUB 0.39fF
C144 S.n106 SUB 0.69fF
C145 S.t21 SUB 0.03fF
C146 S.n107 SUB 0.13fF
C147 S.n108 SUB 0.16fF
C148 S.t7 SUB 0.03fF
C149 S.n109 SUB 1.05fF
C150 S.n110 SUB 0.77fF
C151 S.n111 SUB 3.70fF
C152 S.t24 SUB 0.03fF
C153 S.n112 SUB 0.01fF
C154 S.n113 SUB 0.28fF
C155 S.n114 SUB 1.65fF
C156 S.n115 SUB 0.39fF
C157 S.n116 SUB 1.44fF
C158 S.n117 SUB 0.17fF
C159 S.n118 SUB 27.02fF
.ends

