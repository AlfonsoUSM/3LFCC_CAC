magic
tech sky130A
timestamp 1675431308
<< error_p >>
rect 507 575 610 663
rect 81 560 610 575
rect 81 553 519 560
rect 345 550 385 553
rect -463 547 -187 550
rect 610 507 663 560
rect 550 345 571 433
rect -975 53 156 160
rect 396 156 550 160
rect 103 0 156 53
rect 117 -21 205 0
rect -10 -113 43 -60
<< pwell >>
rect -575 0 550 550
<< mvnmos >>
rect 81 500 519 550
<< mvndiff >>
rect 81 550 519 553
rect 81 494 519 500
rect 81 477 87 494
rect 513 477 519 494
rect 81 471 519 477
rect 79 469 521 471
rect 79 463 550 469
rect 79 415 527 463
rect 79 85 135 415
rect 465 85 527 415
rect 79 37 527 85
rect 544 37 550 463
rect 79 31 550 37
rect 79 29 521 31
rect 81 23 519 29
rect 81 6 87 23
rect 513 6 519 23
rect 81 0 519 6
<< mvndiffc >>
rect 87 477 513 494
rect 527 37 544 463
rect 87 6 513 23
<< mvpsubdiff >>
rect -475 17 -463 550
rect -187 17 -175 550
rect -475 0 -175 17
rect 135 403 465 415
rect 135 97 147 403
rect 453 97 465 403
rect 135 85 465 97
<< mvpsubdiffcont >>
rect -463 17 -187 550
rect 147 97 453 403
<< poly >>
rect 0 542 81 550
rect 0 508 8 542
rect 42 508 81 542
rect 0 500 81 508
rect 519 500 550 550
rect 0 0 50 500
<< polycont >>
rect 8 508 42 542
<< locali >>
rect -475 17 -463 550
rect -187 17 -175 550
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 79 477 87 494
rect 513 477 521 494
rect 73 471 527 477
rect 73 463 544 471
rect 73 415 527 463
rect 73 85 135 415
rect 465 85 527 415
rect 73 37 527 85
rect 73 29 544 37
rect 73 23 527 29
rect -475 0 -175 17
rect 79 6 87 23
rect 513 6 521 23
<< viali >>
rect -463 19 -187 550
rect 8 508 42 542
rect 87 477 513 494
rect 135 403 465 415
rect 135 97 147 403
rect 147 97 453 403
rect 453 97 465 403
rect 135 85 465 97
rect 527 37 544 463
rect 87 6 513 23
<< metal1 >>
rect -475 19 -463 550
rect -187 19 -175 550
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 81 494 519 497
rect 81 477 87 494
rect 513 477 519 494
rect 81 474 519 477
rect 76 469 524 474
rect 76 463 547 469
rect 76 415 527 463
rect 76 85 135 415
rect 465 85 527 415
rect 76 37 527 85
rect 544 37 547 463
rect 76 31 547 37
rect 76 26 524 31
rect -475 0 -175 19
rect 81 23 519 26
rect 81 6 87 23
rect 513 6 519 23
rect 81 3 519 6
<< via1 >>
rect -375 362 -275 462
rect 8 508 42 542
rect 135 85 465 415
<< metal2 >>
rect -175 542 550 550
rect -175 508 8 542
rect 42 508 550 542
rect -175 500 550 508
rect -385 462 -265 472
rect -385 362 -375 462
rect -275 362 -265 462
rect -385 352 -265 362
rect -175 0 50 500
rect 125 415 475 425
rect 125 85 135 415
rect 465 85 475 415
rect 125 75 475 85
<< via2 >>
rect -375 362 -275 462
rect 240 190 360 310
<< metal3 >>
rect -475 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 550 550
rect -475 462 266 510
rect -475 362 -375 462
rect -275 412 266 462
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 550 510
rect -275 362 364 412
rect -475 314 364 362
tri 364 314 462 412 sw
tri 462 324 550 412 ne
rect -475 310 462 314
rect -475 190 240 310
rect 360 226 462 310
tri 462 226 550 314 sw
rect 360 190 550 226
rect -475 186 550 190
tri 138 88 236 186 ne
rect 236 88 550 186
rect -975 0 138 88
tri 138 0 226 88 sw
tri 236 0 324 88 ne
rect 324 0 550 88
<< via3 >>
rect -375 362 -275 462
rect 240 190 360 310
<< metal4 >>
rect -475 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 550 550
rect -475 462 266 510
rect -475 362 -375 462
rect -275 412 266 462
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 550 510
rect -275 362 364 412
rect -475 314 364 362
tri 364 314 462 412 sw
tri 462 324 550 412 ne
rect -475 310 462 314
rect -475 190 240 310
rect 360 226 462 310
tri 462 226 550 314 sw
rect 360 190 550 226
rect -475 186 550 190
tri 138 88 236 186 ne
rect 236 88 550 186
rect -975 0 138 88
tri 138 0 226 88 sw
tri 236 0 324 88 ne
rect 324 0 550 88
<< via4 >>
rect 240 190 360 310
<< metal5 >>
rect -475 447 156 550
tri 156 447 259 550 sw
tri 394 447 497 550 ne
rect 497 447 550 550
rect -475 310 259 447
tri 259 310 396 447 sw
tri 497 394 550 447 ne
rect -475 292 240 310
tri 102 190 204 292 ne
rect 204 190 240 292
rect 360 190 396 310
rect -975 0 103 53
tri 103 0 156 53 sw
tri 204 0 394 190 ne
rect 394 156 396 190
tri 396 156 550 310 sw
rect 394 0 550 156
<< properties >>
string MASKHINTS_HVI 880 0 1100 220 960 960 1100 1100
string MASKHINTS_HVNTM 93 21 121 979
<< end >>
