**.subckt PMOS_RONcalc
VGS G VDD {VGS}
VDS D VDD -5
XM1 D G VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='mul' m='mul'
VDD VDD GND 5
**** begin user architecture code


.param VGS = -5
.param mul = 264
.option temp=70
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.control
compose voltage values -5 (-2.5)
foreach volt $&voltage
alterparam VGS=$volt
reset
save i(VDS)
dc VDS -3 0 0.0001
wrdata SPICE_files/PMOS/PRELAYOUT/PMOS_R_on_calc_PRELAYOUT.txt i(VDS)
set appendwrite
end

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
.control
quit
.endc