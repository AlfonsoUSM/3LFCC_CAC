* NGSPICE file created from nmos_6x6_flat.ext - technology: sky130A

.subckt nmos_6x6_flat
X0 S.t69 G D.t37 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1 D.t36 G S S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.31847e+14p ps=5.9064e+08u w=4.38e+06u l=500000u
X2 S.t66 G D.t20 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D.t35 G S S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 S.t64 G D.t22 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 D.t6 G S.t63 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 S G D.t34 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 D.t1 G S.t61 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 S G D.t33 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 D.t0 G S.t59 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 D.t3 G S.t58 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 S.t57 G D.t43 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 D.t54 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D.t16 G S.t55 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 S.t54 G D.t15 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D.t57 G S.t53 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 D.t55 G S.t52 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 D.t32 G S S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 D.t44 G S.t49 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 D.t31 G S S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 S.t47 G D.t5 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 D.t58 G S.t46 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 D.t53 G S.t0 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D.t52 G S.t0 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 S.t43 G D.t8 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 D.t9 G S.t42 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D.t13 G S.t41 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 D.t7 G S.t40 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 S.t39 G D.t17 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 D.t30 G S S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 D.t23 G S.t37 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 D.t41 G S.t36 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 S.t35 G D.t4 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 S G D.t29 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 D.t38 G S.t32 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 S.t31 G D.t12 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 D.t42 G S.t30 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t0 G D.t51 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 S.t28 G D.t18 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 S G D.t28 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 S.t25 G D.t59 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 D.t50 G S.t0 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 S.t23 G D.t24 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 D.t10 G S.t21 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 S.t0 G D.t49 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 S.t19 G D.t19 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 S G D.t27 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 S.t17 G D.t14 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 S.t16 G D.t56 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 S.t0 G D.t48 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 S.t14 G D.t39 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D.t11 G S.t13 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 S.t0 G D.t47 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 D.t25 G S.t10 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 S.t0 G D.t46 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 S.t8 G D.t40 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 D.t21 G S.t6 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 S.t4 G D.t2 S.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 S G D.t26 S sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D.t45 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 D.n39 D.n38 41.943
R1 D.n38 D.n37 8.553
R2 D.n15 D.t48 4.386
R3 D.n11 D.t38 4.386
R4 D.n14 D.t29 4.386
R5 D.n10 D.t45 4.386
R6 D.n10 D.t51 4.386
R7 D.n3 D.t32 4.386
R8 D.n3 D.t26 4.386
R9 D.n2 D.t21 4.386
R10 D.n2 D.t12 4.386
R11 D.n1 D.t55 4.386
R12 D.n1 D.t18 4.386
R13 D.n6 D.t3 4.386
R14 D.n17 D.t54 4.386
R15 D.n16 D.t46 4.386
R16 D.n5 D.t16 4.386
R17 D.n5 D.t40 4.386
R18 D.n0 D.t13 4.386
R19 D.n0 D.t15 4.386
R20 D.n4 D.t28 4.386
R21 D.n4 D.t36 4.386
R22 D.n7 D.t27 4.327
R23 D.n8 D.t33 4.327
R24 D.n60 D.t19 4.327
R25 D.n59 D.t6 4.327
R26 D.n72 D.t24 4.327
R27 D.n71 D.t7 4.327
R28 D.n65 D.t49 4.327
R29 D.n64 D.t35 4.327
R30 D.n57 D.t56 4.327
R31 D.n56 D.t53 4.327
R32 D.n13 D.t9 4.327
R33 D.n101 D.t20 4.327
R34 D.n100 D.t58 4.327
R35 D.n96 D.t22 4.327
R36 D.n95 D.t52 4.327
R37 D.n12 D.t10 4.327
R38 D.n33 D.t47 4.327
R39 D.n32 D.t30 4.327
R40 D.n39 D.t8 4.327
R41 D.n40 D.t1 4.327
R42 D.n7 D.t39 4.091
R43 D.n8 D.t25 4.091
R44 D.n13 D.t57 4.091
R45 D.n12 D.t43 4.091
R46 D.n18 D.t34 4.084
R47 D.n15 D.t17 4.083
R48 D.n11 D.t5 4.083
R49 D.n14 D.t59 4.083
R50 D.n21 D.t44 4.083
R51 D.n6 D.t37 4.083
R52 D.n21 D.t14 4.06
R53 D.n18 D.t23 4.06
R54 D.n49 D.t0 4.057
R55 D.n26 D.t4 4.057
R56 D.n94 D.t2 4.057
R57 D.n106 D.t42 4.057
R58 D.n35 D.t41 4.031
R59 D.n104 D.t50 4.031
R60 D.n27 D.t11 4.031
R61 D.n88 D.t31 4.031
R62 D.n28 D.n14 0.24
R63 D.n87 D.n86 0.225
R64 D.n93 D.n92 0.225
R65 D.n75 D.n73 0.174
R66 D.n98 D.n13 0.166
R67 D.n52 D.n8 0.16
R68 D.n75 D.n74 0.156
R69 D.n19 D.n45 0.298
R70 D.n8 D.n22 0.143
R71 D.n7 D.n29 0.143
R72 D.n3 D.n76 0.143
R73 D.n107 D.n11 0.143
R74 D.n25 D.n23 0.133
R75 D.n52 D.n7 0.127
R76 D.n107 D.n6 0.118
R77 D.n48 D.n42 0.113
R78 D.n51 D.n50 0.096
R79 D.n85 D.n84 0.092
R80 D.n91 D.n90 0.092
R81 D.n18 D.n78 0.091
R82 D.n108 D.n82 0.085
R83 D.n31 D.n30 0.083
R84 D.n11 D.n12 0.079
R85 D.n20 D.n67 0.075
R86 D.n99 D.n98 0.072
R87 D.n41 D.n31 0.072
R88 D.n1 D.n21 0.066
R89 D.n82 D.n18 0.061
R90 D.n54 D.n53 0.058
R91 D.n6 D.n17 0.057
R92 D.n90 D.n89 0.055
R93 D.n84 D.n83 0.055
R94 D.n68 D.n109 0.055
R95 D.n25 D.n24 0.053
R96 D.n42 D.n41 0.053
R97 D.n4 D.n0 0.053
R98 D.n63 D.n62 0.053
R99 D.n10 D.n59 0.052
R100 D.n10 D.n60 0.052
R101 D.n3 D.n72 0.052
R102 D.n3 D.n71 0.052
R103 D.n2 D.n65 0.052
R104 D.n2 D.n64 0.052
R105 D.n1 D.n57 0.052
R106 D.n1 D.n56 0.052
R107 D.n17 D.n101 0.052
R108 D.n17 D.n100 0.052
R109 D.n5 D.n96 0.052
R110 D.n5 D.n95 0.052
R111 D.n0 D.n33 0.052
R112 D.n0 D.n32 0.052
R113 D.n4 D.n39 0.052
R114 D.n4 D.n40 0.052
R115 D.n15 D.n35 0.051
R116 D.n11 D.n104 0.051
R117 D.n6 D.n88 0.051
R118 D.n68 D.n110 0.051
R119 D.n92 D.n91 0.051
R120 D.n86 D.n85 0.051
R121 D.n10 D.n1 0.049
R122 D.n3 D.n2 0.049
R123 D.n2 D.n10 0.049
R124 D.n44 D.n43 0.045
R125 D D.n108 0.045
R126 D.n18 D.n81 0.192
R127 D.n0 D.n15 0.04
R128 D.n47 D.n46 0.039
R129 D.n3 D.n75 0.039
R130 D.n3 D.n69 0.039
R131 D.n7 D.n51 0.245
R132 D.n8 D.n28 0.035
R133 D.n7 D.n49 0.034
R134 D.n8 D.n26 0.034
R135 D.n54 D.n52 0.032
R136 D.n108 D.n107 0.031
R137 D D.n54 0.031
R138 D.n78 D.n77 0.024
R139 D.n19 D.n44 0.023
R140 D.n69 D.n20 0.023
R141 D.n81 D.n80 0.019
R142 D.n6 D.n93 0.016
R143 D.n11 D.n105 0.016
R144 D.n17 D.n102 0.016
R145 D.n5 D.n97 0.016
R146 D.n2 D.n66 0.016
R147 D.n1 D.n58 0.015
R148 D.n20 D.n68 0.014
R149 D.n48 D.n47 0.012
R150 D.n17 D.n99 0.011
R151 D.n10 D.n61 0.011
R152 D.n81 D.n79 0.057
R153 D.n14 D.n27 0.055
R154 D.n18 D.n3 0.045
R155 D.n13 D.n94 0.038
R156 D.n12 D.n106 0.038
R157 D.n3 D.n70 0.036
R158 D.n8 D.n25 0.033
R159 D.n7 D.n48 0.033
R160 D.n46 D.n19 0.024
R161 D.n0 D.n34 0.024
R162 D.n6 D.n87 0.023
R163 D.n11 D.n103 0.02
R164 D.n1 D.n55 0.02
R165 D.n2 D.n63 0.02
R166 D.n41 D.n4 0.018
R167 D.n98 D.n5 0.018
R168 D.n15 D.n36 0.015
R169 D.n10 D.n9 0.013
R170 D.n17 D.n16 0.01
R171 S.n65 S.n64 91.519
R172 S.n124 S.n123 91.519
R173 S S.n78 87.091
R174 S S.n77 87.091
R175 S.n30 S.n29 87.091
R176 S.n21 S.n20 87.091
R177 S S.t59 3.773
R178 S S.t61 3.773
R179 S S.t35 3.773
R180 S.n65 S.t41 3.773
R181 S.n35 S.t25 3.773
R182 S.n62 S.t36 3.773
R183 S S.t10 3.773
R184 S S.t13 3.773
R185 S.n124 S.t52 3.773
R186 S.n1 S.n37 3.773
R187 S.n1 S.t54 3.773
R188 S.n46 S.t6 3.773
R189 S.n46 S.n45 3.773
R190 S.n44 S.t63 3.773
R191 S.n44 S.n43 3.773
R192 S.n39 S.n38 3.773
R193 S.n39 S.t43 3.773
R194 S S.t40 3.773
R195 S S.t14 3.773
R196 S S.t37 3.773
R197 S.n28 S.t57 3.773
R198 S.n23 S.t47 3.773
R199 S.n30 S.t64 3.773
R200 S.n32 S.t4 3.773
R201 S.n31 S.t30 3.773
R202 S.n2 S.n114 3.773
R203 S.n2 S.t8 3.773
R204 S.n120 S.t32 3.773
R205 S.n120 S.n119 3.773
R206 S.n122 S.t21 3.773
R207 S.n122 S.n121 3.773
R208 S.n116 S.n115 3.773
R209 S.n116 S.t66 3.773
R210 S.n3 S.n92 3.773
R211 S.n3 S.t28 3.773
R212 S.n107 S.t55 3.773
R213 S.n107 S.n106 3.773
R214 S.n105 S.t42 3.773
R215 S.n105 S.n104 3.773
R216 S.n94 S.n93 3.773
R217 S.n94 S.t19 3.773
R218 S.n21 S.t16 3.773
R219 S.n22 S.t17 3.773
R220 S.n19 S.t53 3.773
R221 S.n4 S.n55 3.773
R222 S.n4 S.t31 3.773
R223 S.n59 S.t58 3.773
R224 S.n59 S.n58 3.773
R225 S.n61 S.t46 3.773
R226 S.n61 S.n60 3.773
R227 S.n53 S.n52 3.773
R228 S.n53 S.t23 3.773
R229 S.n125 S.t39 3.773
R230 S.n127 S.t49 3.773
R231 S.n72 S.t69 3.773
R232 S S.t12 0.178
R233 S S.n34 0.12
R234 S.t22 S.n75 0.118
R235 S.t12 S.n76 0.118
R236 S S.n71 0.112
R237 S S.n9 0.11
R238 S.n76 S.t22 0.068
R239 S.n6 S.n87 0.063
R240 S.n27 S.n23 0.055
R241 S.n66 S.n35 0.054
R242 S.n9 S.n127 0.054
R243 S.n5 S.n44 0.053
R244 S.t7 S.n122 0.053
R245 S.n6 S.n105 0.053
R246 S.t5 S.n61 0.053
R247 S.n85 S.n84 0.052
R248 S.t0 S.n72 0.051
R249 S.n0 S.n108 0.05
R250 S.n89 S.n88 0.05
R251 S.n5 S.n40 0.047
R252 S.n0 S.n117 0.047
R253 S.n6 S.n95 0.047
R254 S.n7 S.n54 0.047
R255 S.n9 S.n126 0.047
R256 S.n18 S.n17 0.038
R257 S.n101 S.n100 0.038
R258 S.n103 S.n96 0.036
R259 S.n63 S.n62 0.034
R260 S.n9 S.n86 0.034
R261 S.t3 S.n31 0.034
R262 S.t3 S.n32 0.034
R263 S.t3 S.n19 0.034
R264 S.t3 S.n22 0.034
R265 S.t5 S.n63 0.031
R266 S.n16 S.n15 0.029
R267 S.n101 S.n99 0.028
R268 S.n75 S.t11 0.028
R269 S.n0 S.n118 0.028
R270 S.n9 S.n80 0.027
R271 S.n7 S.n57 0.026
R272 S.n70 S.n67 0.026
R273 S.n0 S.n112 0.026
R274 S.n80 S.n79 0.024
R275 S.n85 S.n83 0.023
R276 S.n102 S.n97 0.023
R277 S.n82 S.n81 0.023
R278 S.n13 S.n12 0.022
R279 S.n111 S.n110 0.021
R280 S.t3 S.n13 0.019
R281 S.n7 S.n51 0.016
R282 S.t3 S.n16 0.016
R283 S.n110 S.n109 0.015
R284 S.n6 S.n90 0.012
R285 S.n103 S.n102 0.012
R286 S.n6 S.n103 0.011
R287 S.n70 S.n68 0.01
R288 S.n5 S.n41 0.01
R289 S.n9 S.n82 0.01
R290 S.n9 S.n85 0.01
R291 S.n70 S.n69 0.01
R292 S.n50 S.n48 0.008
R293 S.t3 S.n18 0.008
R294 S.n99 S.n98 0.008
R295 S.n5 S.n42 0.008
R296 S.t3 S.n14 0.005
R297 S.n26 S.n24 0.005
R298 S.t3 S.n33 0.005
R299 S.n40 S.n39 0.004
R300 S.n117 S.n116 0.004
R301 S.n95 S.n94 0.004
R302 S.n54 S.n53 0.004
R303 S.n126 S.n125 0.004
R304 S.n73 S.t0 0.131
R305 S.n7 S.n50 0.004
R306 S.n7 S.n4 0.004
R307 S.n6 S.n3 0.004
R308 S.n0 S.n2 0.004
R309 S.n5 S.n1 0.004
R310 S.t3 S.n28 0.004
R311 S.t3 S.n30 0.004
R312 S.t3 S.n21 0.004
R313 S.t5 S.n65 0.004
R314 S.n8 S.n124 0.003
R315 S.t5 S.n46 0.003
R316 S.n0 S.n120 0.003
R317 S.t7 S.n107 0.003
R318 S.n7 S.n59 0.003
R319 S.n112 S.n111 0.003
R320 S.n102 S.n101 0.003
R321 S.n26 S.n25 0.003
R322 S.n90 S.n89 0.003
R323 S.n5 S.n36 0.002
R324 S.n0 S.n113 0.002
R325 S.t3 S.n10 0.002
R326 S.n57 S.n56 0.002
R327 S.n71 S.n70 0.002
R328 S.t7 S.n0 0.002
R329 S.n6 S.n91 0.002
R330 S.n7 S.n47 0.002
R331 S.t7 S.n6 0.002
R332 S.t5 S.n5 0.002
R333 S.n66 S.t5 0.001
R334 S.n27 S.n26 0.001
R335 S.t3 S.n27 0.001
R336 S.n34 S.t3 0.001
R337 S.t3 S.n11 0.001
R338 S.n50 S.n49 0.001
R339 S.n74 S.n73 0.001
R340 S.n70 S.n66 0.001
R341 S.t5 S.n7 0.001
R342 S.n9 S.n8 0.001
R343 S.n8 S.t7 0.001
R344 S.t11 S.n74 0.001
C0 D S 180.22fF
C1 DNW S 386.59fF
C2 DNW D 110.79fF
C3 G S 125.11fF
C4 G D 73.67fF
C5 DNW G 1.64fF
C6 D VSUBS -2.71fF $ **FLOATING
C7 G VSUBS -5.46fF
C8 S VSUBS 239.92fF
C9 DNW VSUBS 2400.13fF $ **FLOATING
C10 S.n0 VSUBS 3.88fF $ **FLOATING
C11 S.n1 VSUBS 0.13fF $ **FLOATING
C12 S.n2 VSUBS 0.13fF $ **FLOATING
C13 S.n3 VSUBS 0.13fF $ **FLOATING
C14 S.n4 VSUBS 0.13fF $ **FLOATING
C15 S.t5 VSUBS 8.52fF
C16 S.n5 VSUBS 4.87fF $ **FLOATING
C17 S.t7 VSUBS 8.17fF
C18 S.n6 VSUBS 1.60fF $ **FLOATING
C19 S.n7 VSUBS 1.66fF $ **FLOATING
C20 S.n9 VSUBS 3.62fF $ **FLOATING
C21 S.t22 VSUBS 19.71fF
C22 S.n10 VSUBS 1.34fF $ **FLOATING
C23 S.n11 VSUBS 2.40fF $ **FLOATING
C24 S.n12 VSUBS 0.73fF $ **FLOATING
C25 S.n13 VSUBS 0.42fF $ **FLOATING
C26 S.n14 VSUBS 0.27fF $ **FLOATING
C27 S.n15 VSUBS 0.28fF $ **FLOATING
C28 S.n16 VSUBS 0.20fF $ **FLOATING
C29 S.n17 VSUBS 0.31fF $ **FLOATING
C30 S.n18 VSUBS 0.59fF $ **FLOATING
C31 S.t53 VSUBS 0.02fF
C32 S.n19 VSUBS 0.81fF $ **FLOATING
C33 S.n20 VSUBS 0.01fF $ **FLOATING
C34 S.t16 VSUBS 0.02fF
C35 S.n21 VSUBS 0.34fF $ **FLOATING
C36 S.t17 VSUBS 0.02fF
C37 S.n22 VSUBS 0.81fF $ **FLOATING
C38 S.t47 VSUBS 0.02fF
C39 S.n23 VSUBS 1.19fF $ **FLOATING
C40 S.n24 VSUBS 1.89fF $ **FLOATING
C41 S.n25 VSUBS 1.73fF $ **FLOATING
C42 S.n26 VSUBS 7.19fF $ **FLOATING
C43 S.n27 VSUBS 0.23fF $ **FLOATING
C44 S.t57 VSUBS 0.02fF
C45 S.n28 VSUBS 0.40fF $ **FLOATING
C46 S.n29 VSUBS 0.01fF $ **FLOATING
C47 S.t64 VSUBS 0.02fF
C48 S.n30 VSUBS 0.34fF $ **FLOATING
C49 S.t30 VSUBS 0.02fF
C50 S.n31 VSUBS 0.81fF $ **FLOATING
C51 S.t4 VSUBS 0.02fF
C52 S.n32 VSUBS 0.81fF $ **FLOATING
C53 S.n33 VSUBS 1.14fF $ **FLOATING
C54 S.t3 VSUBS 26.84fF
C55 S.n34 VSUBS 3.08fF $ **FLOATING
C56 S.t25 VSUBS 0.02fF
C57 S.n35 VSUBS 1.11fF $ **FLOATING
C58 S.n36 VSUBS 1.71fF $ **FLOATING
C59 S.n37 VSUBS 0.11fF $ **FLOATING
C60 S.t54 VSUBS 0.02fF
C61 S.t43 VSUBS 0.02fF
C62 S.n38 VSUBS 0.22fF $ **FLOATING
C63 S.n39 VSUBS 0.32fF $ **FLOATING
C64 S.n40 VSUBS 0.55fF $ **FLOATING
C65 S.n41 VSUBS 1.13fF $ **FLOATING
C66 S.n42 VSUBS 0.32fF $ **FLOATING
C67 S.t63 VSUBS 0.02fF
C68 S.n43 VSUBS 0.22fF $ **FLOATING
C69 S.n44 VSUBS 0.83fF $ **FLOATING
C70 S.t6 VSUBS 0.02fF
C71 S.n45 VSUBS 0.11fF $ **FLOATING
C72 S.n46 VSUBS 0.13fF $ **FLOATING
C73 S.n47 VSUBS 1.73fF $ **FLOATING
C74 S.n48 VSUBS 0.29fF $ **FLOATING
C75 S.n49 VSUBS 0.42fF $ **FLOATING
C76 S.n50 VSUBS 0.15fF $ **FLOATING
C77 S.n51 VSUBS 1.96fF $ **FLOATING
C78 S.t23 VSUBS 0.02fF
C79 S.n52 VSUBS 0.22fF $ **FLOATING
C80 S.n53 VSUBS 0.32fF $ **FLOATING
C81 S.n54 VSUBS 0.55fF $ **FLOATING
C82 S.n55 VSUBS 0.11fF $ **FLOATING
C83 S.t31 VSUBS 0.02fF
C84 S.n56 VSUBS 0.82fF $ **FLOATING
C85 S.n57 VSUBS 0.21fF $ **FLOATING
C86 S.t58 VSUBS 0.02fF
C87 S.n58 VSUBS 0.11fF $ **FLOATING
C88 S.n59 VSUBS 0.13fF $ **FLOATING
C89 S.t46 VSUBS 0.02fF
C90 S.n60 VSUBS 0.22fF $ **FLOATING
C91 S.n61 VSUBS 0.83fF $ **FLOATING
C92 S.t36 VSUBS 0.02fF
C93 S.n62 VSUBS 0.86fF $ **FLOATING
C94 S.n63 VSUBS 0.64fF $ **FLOATING
C95 S.t41 VSUBS 0.02fF
C96 S.n64 VSUBS 0.01fF $ **FLOATING
C97 S.n65 VSUBS 0.23fF $ **FLOATING
C98 S.n66 VSUBS 0.23fF $ **FLOATING
C99 S.n67 VSUBS 0.17fF $ **FLOATING
C100 S.n68 VSUBS 0.31fF $ **FLOATING
C101 S.n69 VSUBS 2.06fF $ **FLOATING
C102 S.n70 VSUBS 1.05fF $ **FLOATING
C103 S.n71 VSUBS 1.87fF $ **FLOATING
C104 S.t13 VSUBS 0.02fF
C105 S.t69 VSUBS 0.02fF
C106 S.n72 VSUBS 1.09fF $ **FLOATING
C107 S.t0 VSUBS 47.18fF
C108 S.n73 VSUBS 2.94fF $ **FLOATING
C109 S.n74 VSUBS 1.41fF $ **FLOATING
C110 S.t11 VSUBS 14.54fF
C111 S.n75 VSUBS 0.70fF $ **FLOATING
C112 S.n76 VSUBS 74.05fF $ **FLOATING
C113 S.t12 VSUBS 183.29fF
C114 S.t37 VSUBS 0.02fF
C115 S.t40 VSUBS 0.02fF
C116 S.n77 VSUBS 0.01fF $ **FLOATING
C117 S.t14 VSUBS 0.02fF
C118 S.t10 VSUBS 0.02fF
C119 S.t61 VSUBS 0.02fF
C120 S.n78 VSUBS 0.01fF $ **FLOATING
C121 S.t35 VSUBS 0.02fF
C122 S.t59 VSUBS 0.02fF
C123 S.n79 VSUBS 1.19fF $ **FLOATING
C124 S.n80 VSUBS 0.14fF $ **FLOATING
C125 S.n81 VSUBS 1.37fF $ **FLOATING
C126 S.n82 VSUBS 0.32fF $ **FLOATING
C127 S.n83 VSUBS 1.36fF $ **FLOATING
C128 S.n84 VSUBS 1.19fF $ **FLOATING
C129 S.n85 VSUBS 0.25fF $ **FLOATING
C130 S.n86 VSUBS 0.22fF $ **FLOATING
C131 S.n87 VSUBS 0.09fF $ **FLOATING
C132 S.n88 VSUBS 0.25fF $ **FLOATING
C133 S.n89 VSUBS 1.35fF $ **FLOATING
C134 S.n90 VSUBS 0.19fF $ **FLOATING
C135 S.n91 VSUBS 1.70fF $ **FLOATING
C136 S.n92 VSUBS 0.11fF $ **FLOATING
C137 S.t28 VSUBS 0.02fF
C138 S.t19 VSUBS 0.02fF
C139 S.n93 VSUBS 0.22fF $ **FLOATING
C140 S.n94 VSUBS 0.32fF $ **FLOATING
C141 S.n95 VSUBS 0.55fF $ **FLOATING
C142 S.n96 VSUBS 0.33fF $ **FLOATING
C143 S.n97 VSUBS 0.37fF $ **FLOATING
C144 S.n98 VSUBS 0.53fF $ **FLOATING
C145 S.n99 VSUBS 0.20fF $ **FLOATING
C146 S.n100 VSUBS 0.62fF $ **FLOATING
C147 S.n101 VSUBS 0.33fF $ **FLOATING
C148 S.n102 VSUBS 0.42fF $ **FLOATING
C149 S.n103 VSUBS 0.07fF $ **FLOATING
C150 S.t42 VSUBS 0.02fF
C151 S.n104 VSUBS 0.22fF $ **FLOATING
C152 S.n105 VSUBS 0.83fF $ **FLOATING
C153 S.t55 VSUBS 0.02fF
C154 S.n106 VSUBS 0.11fF $ **FLOATING
C155 S.n107 VSUBS 0.13fF $ **FLOATING
C156 S.n108 VSUBS 0.06fF $ **FLOATING
C157 S.n109 VSUBS 0.16fF $ **FLOATING
C158 S.n110 VSUBS 0.20fF $ **FLOATING
C159 S.n111 VSUBS 1.33fF $ **FLOATING
C160 S.n112 VSUBS 0.41fF $ **FLOATING
C161 S.n113 VSUBS 2.29fF $ **FLOATING
C162 S.n114 VSUBS 0.11fF $ **FLOATING
C163 S.t8 VSUBS 0.02fF
C164 S.t66 VSUBS 0.02fF
C165 S.n115 VSUBS 0.22fF $ **FLOATING
C166 S.n116 VSUBS 0.32fF $ **FLOATING
C167 S.n117 VSUBS 0.55fF $ **FLOATING
C168 S.n118 VSUBS 1.71fF $ **FLOATING
C169 S.t32 VSUBS 0.02fF
C170 S.n119 VSUBS 0.11fF $ **FLOATING
C171 S.n120 VSUBS 0.13fF $ **FLOATING
C172 S.t21 VSUBS 0.02fF
C173 S.n121 VSUBS 0.22fF $ **FLOATING
C174 S.n122 VSUBS 0.83fF $ **FLOATING
C175 S.t52 VSUBS 0.02fF
C176 S.n123 VSUBS 0.01fF $ **FLOATING
C177 S.n124 VSUBS 0.23fF $ **FLOATING
C178 S.t39 VSUBS 0.02fF
C179 S.n125 VSUBS 0.58fF $ **FLOATING
C180 S.n126 VSUBS 0.55fF $ **FLOATING
C181 S.t49 VSUBS 0.02fF
C182 S.n127 VSUBS 1.09fF $ **FLOATING
C183 D.n0 VSUBS 3.57fF $ **FLOATING
C184 D.n1 VSUBS 3.95fF $ **FLOATING
C185 D.n2 VSUBS 3.50fF $ **FLOATING
C186 D.n3 VSUBS 3.23fF $ **FLOATING
C187 D.n4 VSUBS 7.27fF $ **FLOATING
C188 D.n5 VSUBS 3.62fF $ **FLOATING
C189 D.n6 VSUBS 4.14fF $ **FLOATING
C190 D.n7 VSUBS 8.66fF $ **FLOATING
C191 D.n8 VSUBS 6.05fF $ **FLOATING
C192 D.n9 VSUBS 2.70fF $ **FLOATING
C193 D.n10 VSUBS 3.86fF $ **FLOATING
C194 D.n11 VSUBS 6.79fF $ **FLOATING
C195 D.n12 VSUBS 10.45fF $ **FLOATING
C196 D.n13 VSUBS 10.99fF $ **FLOATING
C197 D.n14 VSUBS 11.60fF $ **FLOATING
C198 D.n15 VSUBS 9.23fF $ **FLOATING
C199 D.n16 VSUBS 0.19fF $ **FLOATING
C200 D.n17 VSUBS 2.98fF $ **FLOATING
C201 D.n18 VSUBS 4.67fF $ **FLOATING
C202 D.n19 VSUBS 14.09fF $ **FLOATING
C203 D.n20 VSUBS 0.67fF $ **FLOATING
C204 D.n21 VSUBS 8.45fF $ **FLOATING
C205 D.n22 VSUBS 0.11fF $ **FLOATING
C206 D.n23 VSUBS 0.64fF $ **FLOATING
C207 D.n24 VSUBS 4.43fF $ **FLOATING
C208 D.n25 VSUBS 0.22fF $ **FLOATING
C209 D.t25 VSUBS 0.00fF
C210 D.t33 VSUBS -0.05fF
C211 D.t4 VSUBS 0.00fF
C212 D.n26 VSUBS 0.31fF $ **FLOATING
C213 D.t29 VSUBS -0.02fF
C214 D.t59 VSUBS -0.01fF
C215 D.t11 VSUBS -0.02fF
C216 D.n27 VSUBS 0.51fF $ **FLOATING
C217 D.n28 VSUBS 4.36fF $ **FLOATING
C218 D.n29 VSUBS 0.09fF $ **FLOATING
C219 D.n30 VSUBS 0.82fF $ **FLOATING
C220 D.n31 VSUBS 1.63fF $ **FLOATING
C221 D.t15 VSUBS -0.02fF
C222 D.t30 VSUBS -0.05fF
C223 D.n32 VSUBS 0.56fF $ **FLOATING
C224 D.t13 VSUBS -0.02fF
C225 D.t47 VSUBS -0.05fF
C226 D.n33 VSUBS 0.56fF $ **FLOATING
C227 D.n34 VSUBS 1.30fF $ **FLOATING
C228 D.t41 VSUBS -0.02fF
C229 D.n35 VSUBS 0.51fF $ **FLOATING
C230 D.t48 VSUBS -0.02fF
C231 D.t17 VSUBS -0.01fF
C232 D.n36 VSUBS 1.61fF $ **FLOATING
C233 D.t28 VSUBS -0.02fF
C234 D.n37 VSUBS 0.01fF $ **FLOATING
C235 D.t8 VSUBS -0.05fF
C236 D.n39 VSUBS 0.55fF $ **FLOATING
C237 D.t1 VSUBS -0.05fF
C238 D.n40 VSUBS 0.56fF $ **FLOATING
C239 D.t36 VSUBS -0.02fF
C240 D.n41 VSUBS 1.77fF $ **FLOATING
C241 D.n42 VSUBS 1.10fF $ **FLOATING
C242 D.n43 VSUBS 0.03fF $ **FLOATING
C243 D.n44 VSUBS 0.04fF $ **FLOATING
C244 D.n45 VSUBS 18.02fF $ **FLOATING
C245 D.n46 VSUBS 0.07fF $ **FLOATING
C246 D.n47 VSUBS 0.09fF $ **FLOATING
C247 D.n48 VSUBS 0.10fF $ **FLOATING
C248 D.t27 VSUBS -0.05fF
C249 D.t39 VSUBS 0.00fF
C250 D.t0 VSUBS 0.00fF
C251 D.n49 VSUBS 0.31fF $ **FLOATING
C252 D.n50 VSUBS 1.03fF $ **FLOATING
C253 D.n51 VSUBS 26.07fF $ **FLOATING
C254 D.n52 VSUBS 15.54fF $ **FLOATING
C255 D.n53 VSUBS 0.96fF $ **FLOATING
C256 D.n54 VSUBS 6.74fF $ **FLOATING
C257 D.n55 VSUBS 1.98fF $ **FLOATING
C258 D.t18 VSUBS -0.02fF
C259 D.t53 VSUBS -0.05fF
C260 D.n56 VSUBS 0.56fF $ **FLOATING
C261 D.t55 VSUBS -0.02fF
C262 D.t56 VSUBS -0.05fF
C263 D.n57 VSUBS 0.56fF $ **FLOATING
C264 D.n58 VSUBS 1.26fF $ **FLOATING
C265 D.t44 VSUBS -0.01fF
C266 D.t14 VSUBS 0.00fF
C267 D.t6 VSUBS -0.05fF
C268 D.n59 VSUBS 0.56fF $ **FLOATING
C269 D.t51 VSUBS -0.02fF
C270 D.t45 VSUBS -0.02fF
C271 D.t19 VSUBS -0.05fF
C272 D.n60 VSUBS 0.56fF $ **FLOATING
C273 D.n61 VSUBS 2.08fF $ **FLOATING
C274 D.n62 VSUBS 1.12fF $ **FLOATING
C275 D.n63 VSUBS 1.78fF $ **FLOATING
C276 D.t12 VSUBS -0.02fF
C277 D.t35 VSUBS -0.05fF
C278 D.n64 VSUBS 0.56fF $ **FLOATING
C279 D.t21 VSUBS -0.02fF
C280 D.t49 VSUBS -0.05fF
C281 D.n65 VSUBS 0.56fF $ **FLOATING
C282 D.n66 VSUBS 1.71fF $ **FLOATING
C283 D.n67 VSUBS 0.07fF $ **FLOATING
C284 D.n68 VSUBS 0.39fF $ **FLOATING
C285 D.n69 VSUBS 0.17fF $ **FLOATING
C286 D.n70 VSUBS 0.12fF $ **FLOATING
C287 D.t26 VSUBS -0.02fF
C288 D.t7 VSUBS -0.05fF
C289 D.n71 VSUBS 0.56fF $ **FLOATING
C290 D.t32 VSUBS -0.02fF
C291 D.t24 VSUBS -0.05fF
C292 D.n72 VSUBS 0.56fF $ **FLOATING
C293 D.n73 VSUBS 0.10fF $ **FLOATING
C294 D.n74 VSUBS 0.09fF $ **FLOATING
C295 D.n75 VSUBS 0.10fF $ **FLOATING
C296 D.n76 VSUBS 1.06fF $ **FLOATING
C297 D.n77 VSUBS 0.06fF $ **FLOATING
C298 D.n78 VSUBS 0.05fF $ **FLOATING
C299 D.t23 VSUBS 0.00fF
C300 D.t34 VSUBS -0.01fF
C301 D.n79 VSUBS 0.17fF $ **FLOATING
C302 D.n80 VSUBS 0.37fF $ **FLOATING
C303 D.n81 VSUBS 0.99fF $ **FLOATING
C304 D.n82 VSUBS 1.50fF $ **FLOATING
C305 D.n83 VSUBS 0.18fF $ **FLOATING
C306 D.n84 VSUBS 1.85fF $ **FLOATING
C307 D.n85 VSUBS 13.00fF $ **FLOATING
C308 D.n86 VSUBS 17.47fF $ **FLOATING
C309 D.n87 VSUBS 1.98fF $ **FLOATING
C310 D.t31 VSUBS -0.02fF
C311 D.n88 VSUBS 0.51fF $ **FLOATING
C312 D.t3 VSUBS -0.02fF
C313 D.t37 VSUBS -0.01fF
C314 D.n89 VSUBS 0.18fF $ **FLOATING
C315 D.n90 VSUBS 1.85fF $ **FLOATING
C316 D.n91 VSUBS 13.00fF $ **FLOATING
C317 D.n92 VSUBS 17.47fF $ **FLOATING
C318 D.n93 VSUBS 1.71fF $ **FLOATING
C319 D.t57 VSUBS 0.00fF
C320 D.t9 VSUBS -0.05fF
C321 D.t2 VSUBS 0.00fF
C322 D.n94 VSUBS 0.31fF $ **FLOATING
C323 D.t40 VSUBS -0.02fF
C324 D.t52 VSUBS -0.05fF
C325 D.n95 VSUBS 0.56fF $ **FLOATING
C326 D.t16 VSUBS -0.02fF
C327 D.t22 VSUBS -0.05fF
C328 D.n96 VSUBS 0.56fF $ **FLOATING
C329 D.n97 VSUBS 2.30fF $ **FLOATING
C330 D.n98 VSUBS 2.59fF $ **FLOATING
C331 D.n99 VSUBS 2.44fF $ **FLOATING
C332 D.t46 VSUBS -0.02fF
C333 D.t58 VSUBS -0.05fF
C334 D.n100 VSUBS 0.56fF $ **FLOATING
C335 D.t54 VSUBS -0.02fF
C336 D.t20 VSUBS -0.05fF
C337 D.n101 VSUBS 0.56fF $ **FLOATING
C338 D.n102 VSUBS 2.15fF $ **FLOATING
C339 D.n103 VSUBS 4.03fF $ **FLOATING
C340 D.t38 VSUBS -0.02fF
C341 D.t5 VSUBS -0.01fF
C342 D.t50 VSUBS -0.02fF
C343 D.n104 VSUBS 0.51fF $ **FLOATING
C344 D.n105 VSUBS 4.53fF $ **FLOATING
C345 D.t10 VSUBS -0.05fF
C346 D.t43 VSUBS 0.00fF
C347 D.t42 VSUBS 0.00fF
C348 D.n106 VSUBS 0.31fF $ **FLOATING
C349 D.n107 VSUBS 15.29fF $ **FLOATING
C350 D.n108 VSUBS 8.35fF $ **FLOATING
C351 D.n109 VSUBS 0.46fF $ **FLOATING
C352 D.n110 VSUBS 0.13fF $ **FLOATING
.ends

