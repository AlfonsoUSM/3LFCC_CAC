* NGSPICE file created from mag_files/POSTLAYOUT/nmos_flat_24x24.ext - technology: sky130A

.subckt mag_files/POSTLAYOUT/nmos_flat_24x24
X0 D G S.t1150 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=1.53148e+15p pd=1.0396e+10u as=0p ps=0u w=4.38e+06u l=500000u
X1 D G S.t1149 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 S.t1148 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D G S.t1147 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 D G S.t1146 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 D G S.t1145 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 D G S.t1144 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 S.t1143 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 S.t1142 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 D G S.t1141 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 S.t1140 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 S.t1139 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 S.t1138 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D G S.t1137 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 D G S.t1136 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D G S.t1135 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 D G S.t1134 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 D G S.t1133 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 D G S.t1132 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 D G S.t1131 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 D G S.t1130 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 D G S.t1129 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 D G S.t1128 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D G S.t1127 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 D G S.t1126 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 D G S.t1125 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D G S.t1124 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 D G S.t1123 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D G S.t1122 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 D G S.t1121 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 D G S.t1120 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 S.t1119 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 D G S.t1118 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 D G S.t1117 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 D G S.t1116 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 D G S.t1115 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 D G S.t1114 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t1113 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 S.t1112 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 D G S.t1111 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D G S.t1110 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 D G S.t1109 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 D G S.t1108 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 D G S.t1107 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 D G S.t1106 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 S.t1105 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 D G S.t1104 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 S.t1103 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 D G S.t1102 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 D G S.t1101 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 S.t1100 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D G S.t1099 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 D G S.t1098 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 D G S.t1097 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 S.t1096 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 D G S.t1095 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 D G S.t1094 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 S.t1093 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 S.t1092 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D G S.t1091 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 S.t1090 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 S.t1089 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 S.t1088 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 S.t1087 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 D G S.t1086 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 S.t1085 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 S.t1084 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 D G S.t1083 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 D G S.t1082 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 D G S.t1081 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 S.t1080 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D G S.t1079 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 S.t1078 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 D G S.t1077 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 D G S.t1076 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 S.t1075 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 S.t1074 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 S.t1073 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 D G S.t1072 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 S.t1071 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 S.t1070 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 S.t1069 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 S.t1068 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 D G S.t1067 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 S.t1066 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 S.t1065 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 S.t1064 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 S.t1063 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 S.t1062 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 S.t1061 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D G S.t1060 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 S.t1059 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 D G S.t1058 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 S.t1057 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 S.t1056 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 S.t1055 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D G S.t1054 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 S.t1053 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 S.t1052 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 D G S.t1051 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 S.t1050 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 D G S.t1049 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 S.t1048 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 S.t1047 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 S.t1046 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 D G S.t1045 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 S.t1044 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 D G S.t1043 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 D G S.t1042 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 S.t1041 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D G S.t1040 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 S.t1039 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t1038 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 S.t1037 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 S.t1036 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 D G S.t1035 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 S.t1034 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 S.t1033 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 S.t1032 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 S.t1031 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 S.t1030 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 D G S.t1029 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 D G S.t1028 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 S.t1027 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 S.t1026 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 D G S.t1025 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 S.t1024 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 D G S.t1023 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 D G S.t1022 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 S.t1021 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 S.t1020 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 D G S.t1019 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 D G S.t1018 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 D G S.t1017 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 D G S.t1016 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t1015 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 S.t1014 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 D G S.t1013 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 S.t1012 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 D G S.t1011 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 S.t1010 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 D G S.t1009 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 S.t1008 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 S.t1007 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 D G S.t1006 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 S.t1005 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 S.t1004 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 D G S.t1003 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 S.t1002 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 S.t1001 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 D G S.t1000 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 S.t999 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 S.t998 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 D G S.t997 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 D G S.t996 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 D G S.t995 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 S.t994 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 S.t993 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 S.t992 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 S.t991 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 S.t990 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 S.t989 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 S.t988 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 S.t987 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 S.t986 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 D G S.t985 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 S.t984 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 D G S.t983 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 S.t982 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 D G S.t981 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 S.t980 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 D G S.t979 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 D G S.t978 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 S.t977 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 S.t976 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 S.t975 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 S.t974 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 S.t973 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 D G S.t972 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 S.t971 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 S.t970 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 S.t969 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 D G S.t968 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 S.t967 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 S.t966 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 S.t965 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 D G S.t964 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 S.t963 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 D G S.t962 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 D G S.t961 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 D G S.t960 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 D G S.t959 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 D G S.t958 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 S.t957 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 S.t956 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 D G S.t955 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 D G S.t954 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 D G S.t953 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 S.t952 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 S.t951 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 D G S.t950 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 D G S.t949 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 D G S.t948 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 S.t947 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 D G S.t946 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 D G S.t945 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 D G S.t944 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 D G S.t943 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 D G S.t942 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 D G S.t941 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 S.t940 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 D G S.t939 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 D G S.t938 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 D G S.t937 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 S.t936 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 D G S.t935 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 D G S.t934 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 D G S.t933 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 D G S.t932 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 D G S.t931 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 D G S.t930 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 S.t929 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 D G S.t928 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 S.t927 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 D G S.t926 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 S.t925 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 S.t924 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 D G S.t923 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 S.t922 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 S.t921 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 D G S.t920 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 S.t919 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 D G S.t918 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 S.t917 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 D G S.t916 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 D G S.t915 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 D G S.t914 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 D G S.t913 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 D G S.t912 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 S.t911 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 S.t910 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 D G S.t909 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 D G S.t908 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 D G S.t907 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 S.t906 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 D G S.t905 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 D G S.t904 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 S.t903 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 D G S.t902 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 D G S.t901 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 D G S.t900 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 D G S.t899 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 D G S.t898 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 D G S.t897 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 S.t896 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 S.t895 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 D G S.t894 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 S.t893 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 D G S.t892 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 S.t891 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 S.t890 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 D G S.t889 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 D G S.t888 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 D G S.t887 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 S.t886 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 S.t885 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 D G S.t884 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 S.t883 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 D G S.t882 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 S.t881 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 S.t880 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 D G S.t879 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 S.t878 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 S.t877 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 S.t876 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 S.t875 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 S.t874 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 D G S.t873 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 S.t872 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 D G S.t871 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 D G S.t870 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 D G S.t869 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 S.t868 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D G S.t867 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 D G S.t866 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 D G S.t865 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 D G S.t864 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 S.t863 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 S.t862 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 S.t861 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 S.t860 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 S.t859 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 S.t858 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 D G S.t857 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 D G S.t856 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 S.t855 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 S.t854 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 D G S.t853 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 S.t852 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 D G S.t851 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 S.t850 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 S.t849 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 S.t848 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 S.t847 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 S.t846 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 S.t845 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 S.t844 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 S.t843 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 S.t842 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 S.t841 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 S.t840 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 D G S.t839 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 S.t838 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 S.t837 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 S.t836 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 D G S.t835 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 D G S.t834 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 S.t833 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 S.t832 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 S.t831 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 D G S.t830 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 S.t829 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 D G S.t828 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 S.t827 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 S.t826 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 S.t825 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 S.t824 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 S.t823 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 S.t822 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 S.t821 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 D G S.t820 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 D G S.t819 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 S.t818 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 D G S.t817 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 S.t816 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 S.t815 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 S.t814 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 S.t813 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 D G S.t812 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 S.t811 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 D G S.t810 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 S.t809 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 S.t808 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 D G S.t807 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 S.t806 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 S.t805 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 S.t804 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 D G S.t803 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 S.t802 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t801 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 D G S.t800 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 D G S.t799 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 D G S.t798 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 D G S.t797 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 D G S.t796 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 D G S.t795 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 D G S.t794 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 S.t793 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 D G S.t792 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 D G S.t791 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 D G S.t790 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 S.t789 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 D G S.t788 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 D G S.t787 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 S.t786 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 D G S.t785 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 S.t784 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 D G S.t783 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 S.t782 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 S.t781 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 D G S.t780 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 S.t779 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 D G S.t778 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 D G S.t777 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 D G S.t776 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 D G S.t775 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 D G S.t774 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 S.t773 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 S.t772 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 D G S.t771 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 D G S.t770 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 S.t769 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 D G S.t768 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 S.t767 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 D G S.t766 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 D G S.t765 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 D G S.t764 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 D G S.t763 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 S.t762 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 S.t761 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 D G S.t760 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 D G S.t759 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 D G S.t758 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 D G S.t757 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 D G S.t756 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 D G S.t755 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 S.t754 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 D G S.t753 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 D G S.t752 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 S.t751 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 S.t750 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 D G S.t749 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 D G S.t748 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 D G S.t747 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 D G S.t746 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 D G S.t745 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 D G S.t744 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 D G S.t743 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 S.t742 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 D G S.t741 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 D G S.t740 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 D G S.t739 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 D G S.t738 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 S.t737 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 D G S.t736 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 D G S.t735 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 S.t734 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 D G S.t733 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 D G S.t732 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 D G S.t731 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 S.t730 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 S.t729 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 S.t728 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 D G S.t727 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 S.t726 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 D G S.t725 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 S.t724 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 D G S.t723 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 S.t722 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 D G S.t721 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 D G S.t720 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 S.t719 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 S.t718 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 D G S.t717 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 S.t716 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 S.t715 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 D G S.t714 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 D G S.t713 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 S.t712 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 D G S.t711 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 D G S.t710 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 D G S.t709 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 S.t708 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 S.t707 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 D G S.t706 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 D G S.t705 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 S.t704 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 S.t703 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 D G S.t702 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 S.t701 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 S.t700 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 S.t699 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 D G S.t698 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 S.t697 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 S.t696 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 D G S.t695 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 S.t694 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 S.t693 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 S.t692 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 S.t691 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 D G S.t690 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 S.t689 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 D G S.t688 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t687 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 S.t686 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 S.t685 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 D G S.t684 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 S.t683 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 S.t682 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 S.t681 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 S.t680 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 S.t679 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 D G S.t678 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 D G S.t677 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 S.t676 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 S.t675 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 S.t674 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 S.t673 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 D G S.t672 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 S.t671 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 S.t670 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 S.t669 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 D G S.t668 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 S.t667 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 D G S.t666 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 D G S.t665 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 D G S.t664 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 S.t663 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 S.t662 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 D G S.t661 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 S.t660 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 D G S.t659 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 D G S.t658 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 S.t657 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t656 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 S.t655 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 D G S.t654 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 S.t653 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 D G S.t652 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 D G S.t651 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 D G S.t650 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 D G S.t649 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 S.t648 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 S.t647 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 S.t646 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 D G S.t645 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 D G S.t644 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 D G S.t643 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 S.t642 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 S.t641 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t640 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 S.t639 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 D G S.t638 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 S.t637 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 D G S.t636 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 S.t635 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 S.t634 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 S.t633 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 S.t632 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 S.t631 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 S.t630 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 D G S.t629 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 D G S.t628 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 S.t627 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 D G S.t626 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 S.t625 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 S.t624 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 D G S.t623 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 D G S.t622 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 S.t621 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 D G S.t620 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D G S.t619 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 D G S.t618 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 S.t617 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 S.t616 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 D G S.t615 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 S.t614 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 S.t613 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 D G S.t612 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 S.t611 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 D G S.t610 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 S.t609 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 S.t608 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 S.t607 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 D G S.t606 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t605 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 D G S.t604 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 S.t603 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 D G S.t602 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 S.t601 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 S.t600 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 D G S.t599 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 D G S.t598 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 S.t597 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 D G S.t596 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 S.t595 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 D G S.t594 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 D G S.t593 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 D G S.t592 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 D G S.t591 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 D G S.t590 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 S.t589 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 D G S.t588 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 S.t587 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 D G S.t586 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 D G S.t585 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 D G S.t584 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 D G S.t583 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 D G S.t582 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 D G S.t581 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 D G S.t580 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 S.t579 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 D G S.t578 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 D G S.t577 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 D G S.t576 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 S.t575 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 D G S.t574 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 D G S.t573 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 S.t572 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 D G S.t571 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 D G S.t570 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 S.t569 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 S.t568 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 D G S.t567 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 S.t566 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 D G S.t565 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 D G S.t564 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 D G S.t563 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 S.t562 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 D G S.t561 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 S.t560 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 S.t559 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 D G S.t558 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 D G S.t557 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 D G S.t556 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 D G S.t555 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 D G S.t554 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 D G S.t553 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 D G S.t552 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 D G S.t551 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 S.t550 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D G S.t549 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 D G S.t548 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 S.t547 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 S.t546 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 D G S.t545 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 S.t544 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 D G S.t543 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 D G S.t542 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 S.t541 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 S.t540 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 D G S.t539 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 D G S.t538 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 D G S.t537 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 D G S.t536 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 D G S.t535 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 D G S.t534 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 D G S.t533 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 S.t532 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 D G S.t531 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 S.t530 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 D G S.t529 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 S.t528 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 D G S.t527 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 S.t526 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 D G S.t525 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 D G S.t524 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 S.t523 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 S.t522 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 S.t521 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 D G S.t520 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 S.t519 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 D G S.t518 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 D G S.t517 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 D G S.t516 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 S.t515 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 D G S.t514 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 S.t513 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 S.t512 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 S.t511 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 S.t510 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 S.t509 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 S.t508 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 D G S.t507 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 D G S.t506 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 S.t505 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 S.t504 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 D G S.t503 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 D G S.t502 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 S.t501 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 D G S.t500 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 S.t499 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 S.t498 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 S.t497 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 S.t496 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 S.t495 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 S.t494 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 D G S.t493 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 D G S.t492 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 S.t491 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 D G S.t490 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 D G S.t489 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 S.t488 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 D G S.t487 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 S.t486 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 S.t485 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 S.t484 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 S.t483 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 S.t482 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 D G S.t481 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 D G S.t480 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 S.t479 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 S.t478 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 D G S.t477 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 S.t476 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 S.t475 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 S.t474 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 S.t473 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 D G S.t472 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 S.t471 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 S.t470 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 S.t469 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 S.t468 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 D G S.t467 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 S.t466 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 S.t465 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 S.t464 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 S.t463 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 S.t462 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 S.t461 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 D G S.t460 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 S.t459 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 S.t458 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 S.t457 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 D G S.t456 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 S.t455 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 D G S.t454 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 D G S.t453 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 S.t452 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 S.t451 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 S.t450 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 D G S.t449 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 S.t448 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 D G S.t447 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 D G S.t446 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 D G S.t445 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 S.t444 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 S.t443 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 S.t442 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 D G S.t441 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 S.t440 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 D G S.t439 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 S.t438 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 S.t437 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 S.t436 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 D G S.t435 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 D G S.t434 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 S.t433 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 D G S.t432 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 D G S.t431 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 D G S.t430 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 S.t429 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 S.t428 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 D G S.t427 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 D G S.t426 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 S.t425 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 D G S.t424 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 S.t423 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 S.t422 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 S.t421 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 D G S.t420 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 D G S.t419 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 D G S.t418 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 D G S.t417 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 D G S.t416 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 D G S.t415 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 S.t414 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 D G S.t413 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 D G S.t412 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 D G S.t411 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 D G S.t410 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 D G S.t409 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 S.t408 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 S.t407 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 D G S.t406 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 D G S.t405 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 S.t404 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 D G S.t403 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 D G S.t402 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 S.t401 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 D G S.t400 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 D G S.t399 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 D G S.t398 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 D G S.t397 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 D G S.t396 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 D G S.t395 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 D G S.t394 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 D G S.t393 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 S.t392 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 S.t391 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 D G S.t390 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 D G S.t389 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 D G S.t388 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 D G S.t387 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 D G S.t386 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 D G S.t385 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 S.t384 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 D G S.t383 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 D G S.t382 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 D G S.t381 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 D G S.t380 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 D G S.t379 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 D G S.t378 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 S.t377 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 D G S.t376 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 D G S.t375 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 D G S.t374 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 D G S.t373 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 D G S.t372 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 D G S.t371 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 D G S.t370 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 S.t369 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 S.t368 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 D G S.t367 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 D G S.t366 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 S.t365 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 S.t364 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 D G S.t363 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 S.t362 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 S.t361 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 D G S.t360 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 S.t359 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 D G S.t358 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 S.t357 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 D G S.t356 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 D G S.t355 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 S.t354 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 S.t353 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 D G S.t352 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 D G S.t351 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 D G S.t350 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 S.t349 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 S.t348 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 S.t347 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 D G S.t346 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 S.t345 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 S.t344 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 S.t343 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 D G S.t342 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 D G S.t341 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 D G S.t340 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 D G S.t339 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 S.t338 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 D G S.t337 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 S.t336 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 S.t335 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 S.t334 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 S.t333 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 D G S.t332 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 S.t331 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 S.t330 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 S.t329 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 D G S.t328 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 D G S.t327 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 S.t326 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 S.t325 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 S.t324 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 S.t323 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 S.t322 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 D G S.t321 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 S.t320 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 S.t319 G D S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 S.t318 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 S.t317 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 S.t316 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 D G S.t315 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 S.t314 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 D G S.t313 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 S.t312 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 S.t311 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 D G S.t310 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 S.t309 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 S.t308 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 D G S.t307 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 S.t306 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 S.t305 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 S.t304 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 S.t303 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 S.t302 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 S.t301 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 S.t300 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 S.t299 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 D G S.t298 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 D G S.t297 S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 S.t296 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 S.t295 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 D G S.t294 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 S.t293 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 S.t292 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 D G S.t291 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 D G S.t290 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 S.t289 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 D G S.t288 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 S.t287 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 S.t286 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 S.t285 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 S.t284 G D S.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 D G S.t282 S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 D G S.t281 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 D G S.t280 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 D G S.t279 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 D G S.t278 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 D G S.t277 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 S.t276 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 S.t275 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 D G S.t274 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 S.t273 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 S.t272 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 S.t271 G D S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 D G S.t270 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 S.t269 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 S.t268 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 S.t267 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 S.t266 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 D G S.t265 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 S.t264 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 D G S.t263 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 S.t262 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 S.t261 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 D G S.t260 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 S.t258 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 S.t257 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 D G S.t256 S.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 S.t254 G D S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 S.t253 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 D G S.t252 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 S.t251 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 D G S.t250 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 S.t249 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 D G S.t248 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 S.t247 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 D G S.t246 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 S.t245 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 D G S.t244 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 D G S.t243 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 D G S.t242 S.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 S.t240 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 S.t239 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 S.t238 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 S.t237 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 S.t236 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 D G S.t235 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 S.t234 G D S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 S.t233 G D S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 D G S.t232 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 D G S.t231 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 S.t230 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 D G S.t229 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 S.t228 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 D G S.t227 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 S.t226 G D S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 S.t225 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 D G S.t224 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 S.t223 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 S.t222 G D S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 D G S.t221 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 S.t220 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 D G S.t219 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 S.t218 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 S.t217 G D S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 D G S.t216 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 D G S.t215 S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 S.t214 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 D G S.t213 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 D G S.t212 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 S.t211 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 D G S.t210 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 D G S.t209 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 D G S.t208 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 D G S.t207 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 D G S.t206 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 D G S.t205 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 S.t204 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 D G S.t203 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 D G S.t202 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 D G S.t201 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 D G S.t200 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 S.t199 G D S.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 D G S.t197 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 D G S.t196 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 D G S.t195 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 D G S.t194 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 D G S.t193 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 S.t192 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 S.t191 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 D G S.t190 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 D G S.t189 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 S.t188 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 S.t187 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 D G S.t186 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 D G S.t185 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 S.t184 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 D G S.t183 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 D G S.t182 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 S.t181 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 S.t180 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 D G S.t179 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 S.t178 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 D G S.t177 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 D G S.t176 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 D G S.t175 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 D G S.t174 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 S.t173 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 D G S.t172 S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 D G S.t171 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 S.t170 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 D G S.t169 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 S.t168 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 D G S.t167 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 D G S.t166 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 S.t165 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 D G S.t164 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 D G S.t163 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 D G S.t162 S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 D G S.t161 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 D G S.t160 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 D G S.t159 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 S.t158 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 D G S.t157 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 D G S.t155 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 S.t154 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 S.t153 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 D G S.t152 S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 S.t151 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 D G S.t150 S.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 D G S.t148 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 S.t147 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 S.t146 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 S.t145 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 D G S.t144 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 S.t143 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 D G S.t142 S.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 D G S.t140 S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 D G S.t139 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 S.t138 G D S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 D G S.t137 S.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 S.t135 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 D G S.t134 S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 S.t133 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 S.t132 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 S.t131 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 S.t130 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 S.t129 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 S.t128 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 D G S.t127 S.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 D G S.t125 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 D G S.t124 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 S.t123 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 D G S.t122 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 S.t121 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 D G S.t120 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 S.t119 G D S.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 S.t117 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 S.t116 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 S.t115 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 S.t114 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 S.t113 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 S.t112 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 S.t110 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 S.t109 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 S.t108 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 S.t107 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 S.t105 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 S.t104 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 D G S.t102 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 S.t101 G D S.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 D G S.t99 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 S.t98 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 S.t97 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 D G S.t96 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 S.t95 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 S.t94 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 S.t93 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 S.t92 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 S.t90 G D S.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 D G S.t88 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 S.t86 G D S.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 D G S.t84 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 S.t83 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 D G S.t82 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 D G S.t81 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 S.t80 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 D G S.t79 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 S.t78 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 S.t77 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 S.t76 G D S.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 D G S.t74 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 S.t73 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 D G S.t72 S.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 S.t70 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 S.t69 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 S.t68 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 D G S.t67 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 S.t65 G D S.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 S.t63 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 S.t61 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 S.t60 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 S.t58 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 D G S.t56 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 D G S.t55 S.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 D G S.t53 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 D G S.t51 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 S.t50 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 D G S.t49 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 D G S.t48 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 S.t46 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 D G S.t45 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 D G S.t43 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 S.t41 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 D G S.t40 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 D G S.t39 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 S.t38 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 S.t37 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 S.t36 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 S.t34 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 D G S.t32 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 S.t31 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 S.t30 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 D G S.t28 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 D G S.t27 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 D G S.t26 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 D G S.t24 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 S.t22 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 S.t20 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 S.t18 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 D G S.t17 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 D G S.t15 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 S.t13 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 D G S.t11 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 S.t9 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 D G S.t7 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 D G S.t5 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 S.t3 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 D G S.t1 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 S.n365 S.n363 169.353
R1 S.n1212 S.n1211 169.353
R2 S.n1248 S.n1247 169.353
R3 S.n1834 S.n1833 169.353
R4 S.n2875 S.n2874 169.353
R5 S.n2925 S.n2924 169.353
R6 S.n3440 S.n3439 169.353
R7 S.n3946 S.n3945 169.353
R8 S.n4417 S.n4416 169.353
R9 S.n5452 S.n5451 169.353
R10 S.n5272 S.n5271 169.353
R11 S.n365 S.n364 169.353
R12 S.n5270 S.n5269 137.98
R13 S.n5450 S.n5449 137.98
R14 S.n4415 S.n4414 137.98
R15 S.n3944 S.n3943 137.98
R16 S.n3438 S.n3437 137.98
R17 S.n2923 S.n2922 137.98
R18 S.n2873 S.n2872 137.98
R19 S.n1832 S.n1831 137.98
R20 S.n1246 S.n1245 137.98
R21 S.n1210 S.n1209 137.98
R22 S.n362 S.n361 137.98
R23 S.n89 S.n88 135.611
R24 S.n977 S.n976 135.611
R25 S.n1551 S.n1550 135.611
R26 S.n2165 S.n2164 135.611
R27 S.n2679 S.n2678 135.611
R28 S.n3216 S.n3215 135.611
R29 S.n3611 S.n3610 135.611
R30 S.n4218 S.n4217 135.611
R31 S.n4673 S.n4672 135.611
R32 S.n5660 S.n5659 135.611
R33 S.n5037 S.n5036 135.611
R34 S.n100 S.n99 91.65
R35 S.n5028 S.n5027 91.65
R36 S.n3228 S.n3227 91.65
R37 S.n3622 S.n3621 91.65
R38 S.n4230 S.n4229 91.65
R39 S.n4684 S.n4683 91.65
R40 S.n5672 S.n5671 91.65
R41 S.n2177 S.n2176 91.65
R42 S.n2690 S.n2689 91.65
R43 S.n989 S.n988 91.65
R44 S.n1562 S.n1561 91.65
R45 S.n5265 S.n5264 91.389
R46 S.n5879 S.n5878 91.389
R47 S.n380 S.n379 91.389
R48 S.n1203 S.n1202 91.389
R49 S.n1803 S.n1802 91.389
R50 S.n2353 S.n2352 91.389
R51 S.n2863 S.n2862 91.389
R52 S.n3409 S.n3408 91.389
R53 S.n3915 S.n3914 91.389
R54 S.n4396 S.n4395 91.389
R55 S.n4850 S.n4849 91.389
R56 S.n650 S.n649 87.222
R57 S.n647 S.n646 87.222
R58 S.n559 S.n558 87.222
R59 S.n662 S.n661 87.222
R60 S.n574 S.n573 87.222
R61 S.n621 S.n620 87.222
R62 S.n638 S.n637 87.222
R63 S.n547 S.n546 87.222
R64 S.n658 S.n657 87.222
R65 S.n535 S.n534 87.222
R66 S.n654 S.n653 87.222
R67 S.n5441 S.n5440 86.961
R68 S.n5359 S.n5358 86.961
R69 S.n5369 S.n5368 86.961
R70 S.n5377 S.n5376 86.961
R71 S.n5385 S.n5384 86.961
R72 S.n5393 S.n5392 86.961
R73 S.n5401 S.n5400 86.961
R74 S.n5409 S.n5408 86.961
R75 S.n5417 S.n5416 86.961
R76 S.n5425 S.n5424 86.961
R77 S.n5347 S.n5346 86.961
R78 S.t241 S.t111 84.027
R79 S.n367 S.t2 73.333
R80 S.n91 S.t259 73.333
R81 S.n1214 S.t33 73.333
R82 S.n979 S.t91 73.333
R83 S.n1250 S.t141 73.333
R84 S.n1553 S.t106 73.333
R85 S.n1836 S.t149 73.333
R86 S.n2167 S.t75 73.333
R87 S.n2877 S.t44 73.333
R88 S.n2681 S.t89 73.333
R89 S.n2927 S.t136 73.333
R90 S.n3218 S.t103 73.333
R91 S.n3442 S.t52 73.333
R92 S.n3613 S.t19 73.333
R93 S.n3948 S.t156 73.333
R94 S.n4220 S.t85 73.333
R95 S.n4419 S.t126 73.333
R96 S.n4675 S.t100 73.333
R97 S.n5454 S.t118 73.333
R98 S.n5662 S.t29 73.333
R99 S.n5274 S.t87 73.333
R100 S.n5039 S.t62 73.333
R101 S.t198 S.n355 70.888
R102 S.t255 S.n261 70.888
R103 S.t59 S.n942 70.888
R104 S.t6 S.n1157 70.888
R105 S.t23 S.n1507 70.888
R106 S.t21 S.n1716 70.888
R107 S.t47 S.n2051 70.888
R108 S.t16 S.n2312 70.888
R109 S.t66 S.n2543 70.888
R110 S.t0 S.n2808 70.888
R111 S.t14 S.n3081 70.888
R112 S.t12 S.n3327 70.888
R113 S.t42 S.n3567 70.888
R114 S.t10 S.n3704 70.888
R115 S.t54 S.n4041 70.888
R116 S.t57 S.n4293 70.888
R117 S.t71 S.n4478 70.888
R118 S.t8 S.n4726 70.888
R119 S.t25 S.n5491 70.888
R120 S.t4 S.n5718 70.888
R121 S.t35 S.n5243 70.888
R122 S.t64 S.n5001 70.888
R123 S.t283 S.n5292 70.888
R124 S.n5291 S.t725 3.904
R125 S.n5290 S.t503 3.904
R126 S.n5265 S.t913 3.904
R127 S.n5215 S.t200 3.904
R128 S.n5441 S.t477 3.904
R129 S.n5439 S.t297 3.904
R130 S.n5012 S.n5011 3.904
R131 S.n5020 S.t332 3.904
R132 S.n5023 S.t88 3.904
R133 S.n5015 S.n5014 3.904
R134 S.n5251 S.n5250 3.904
R135 S.n5259 S.t678 3.904
R136 S.n5262 S.t39 3.904
R137 S.n5254 S.n5253 3.904
R138 S.n5698 S.n5697 3.904
R139 S.n5716 S.t894 3.904
R140 S.n5713 S.t402 3.904
R141 S.n5701 S.n5700 3.904
R142 S.n5879 S.t1130 3.904
R143 S.n5881 S.t580 3.904
R144 S.n101 S.t705 3.904
R145 S.n477 S.n476 3.904
R146 S.n480 S.t252 3.904
R147 S.n483 S.t931 3.904
R148 S.n486 S.n485 3.904
R149 S.n648 S.t1049 3.904
R150 S.n644 S.t581 3.904
R151 S.n342 S.n341 3.904
R152 S.n353 S.t215 3.904
R153 S.n350 S.t839 3.904
R154 S.n345 S.n344 3.904
R155 S.n926 S.n925 3.904
R156 S.n940 S.t232 3.904
R157 S.n937 S.t1094 3.904
R158 S.n923 S.n922 3.904
R159 S.n5025 S.t612 3.904
R160 S.n5223 S.n5222 3.904
R161 S.n5241 S.t82 3.904
R162 S.n5238 S.t870 3.904
R163 S.n5220 S.n5219 3.904
R164 S.n5681 S.n5680 3.904
R165 S.n5692 S.t1023 3.904
R166 S.n5689 S.t420 3.904
R167 S.n5678 S.n5677 3.904
R168 S.n5474 S.n5473 3.904
R169 S.n5489 S.t1060 3.904
R170 S.n5486 S.t636 3.904
R171 S.n5471 S.n5470 3.904
R172 S.n4713 S.n4712 3.904
R173 S.n4724 S.t743 3.904
R174 S.n4721 S.t981 3.904
R175 S.n4710 S.n4709 3.904
R176 S.n4461 S.n4460 3.904
R177 S.n4476 S.t472 3.904
R178 S.n4473 S.t205 3.904
R179 S.n4458 S.n4457 3.904
R180 S.n4280 S.n4279 3.904
R181 S.n4291 S.t785 3.904
R182 S.n4288 S.t972 3.904
R183 S.n4277 S.n4276 3.904
R184 S.n4024 S.n4023 3.904
R185 S.n4039 S.t460 3.904
R186 S.n4036 S.t190 3.904
R187 S.n4021 S.n4020 3.904
R188 S.n3691 S.n3690 3.904
R189 S.n3702 S.t768 3.904
R190 S.n3699 S.t959 3.904
R191 S.n3688 S.n3687 3.904
R192 S.n3550 S.n3549 3.904
R193 S.n3565 S.t43 3.904
R194 S.n3562 S.t175 3.904
R195 S.n3547 S.n3546 3.904
R196 S.n3317 S.n3316 3.904
R197 S.n3325 S.t753 3.904
R198 S.n3309 S.t570 3.904
R199 S.n3314 S.n3313 3.904
R200 S.n3064 S.n3063 3.904
R201 S.n3079 S.t15 3.904
R202 S.n3076 S.t162 3.904
R203 S.n3061 S.n3060 3.904
R204 S.n2795 S.n2794 3.904
R205 S.n2806 S.t735 3.904
R206 S.n2803 S.t551 3.904
R207 S.n2792 S.n2791 3.904
R208 S.n2526 S.n2525 3.904
R209 S.n2541 S.t1145 3.904
R210 S.n2538 S.t221 3.904
R211 S.n2523 S.n2522 3.904
R212 S.n2299 S.n2298 3.904
R213 S.n2310 S.t798 3.904
R214 S.n2307 S.t538 3.904
R215 S.n2296 S.n2295 3.904
R216 S.n2034 S.n2033 3.904
R217 S.n2049 S.t1124 3.904
R218 S.n2046 S.t202 3.904
R219 S.n2031 S.n2030 3.904
R220 S.n1703 S.n1702 3.904
R221 S.n1714 S.t783 3.904
R222 S.n1711 S.t527 3.904
R223 S.n1700 S.n1699 3.904
R224 S.n1488 S.n1487 3.904
R225 S.n1505 S.t1110 3.904
R226 S.n1502 S.t189 3.904
R227 S.n1485 S.n1484 3.904
R228 S.n1146 S.n1145 3.904
R229 S.n1155 S.t764 3.904
R230 S.n1152 S.t698 3.904
R231 S.n1143 S.n1142 3.904
R232 S.n248 S.n247 3.904
R233 S.n259 S.t622 3.904
R234 S.n256 S.t684 3.904
R235 S.n251 S.n250 3.904
R236 S.n553 S.t242 3.904
R237 S.n64 S.n63 3.904
R238 S.n75 S.t1017 3.904
R239 S.n72 S.t713 3.904
R240 S.n67 S.n66 3.904
R241 S.n781 S.n780 3.904
R242 S.n794 S.t1025 3.904
R243 S.n791 S.t727 3.904
R244 S.n778 S.n777 3.904
R245 S.n3229 S.t310 3.904
R246 S.n3088 S.n3087 3.904
R247 S.n3102 S.t937 3.904
R248 S.n3105 S.t378 3.904
R249 S.n3085 S.n3084 3.904
R250 S.n2699 S.n2698 3.904
R251 S.n2710 S.t537 3.904
R252 S.n2707 S.t45 3.904
R253 S.n2696 S.n2695 3.904
R254 S.n2379 S.n2378 3.904
R255 S.n2394 S.t702 3.904
R256 S.n2391 S.t134 3.904
R257 S.n2376 S.n2375 3.904
R258 S.n2203 S.n2202 3.904
R259 S.n2214 S.t288 3.904
R260 S.n2211 S.t243 3.904
R261 S.n2200 S.n2199 3.904
R262 S.n1887 S.n1886 3.904
R263 S.n1902 S.t830 3.904
R264 S.n1899 S.t950 3.904
R265 S.n1884 S.n1883 3.904
R266 S.n1607 S.n1606 3.904
R267 S.n1618 S.t427 3.904
R268 S.n1615 S.t229 3.904
R269 S.n1604 S.n1603 3.904
R270 S.n1335 S.n1334 3.904
R271 S.n1352 S.t819 3.904
R272 S.n1349 S.t934 3.904
R273 S.n1332 S.n1331 3.904
R274 S.n1049 S.n1048 3.904
R275 S.n1058 S.t412 3.904
R276 S.n1055 S.t411 3.904
R277 S.n1046 S.n1045 3.904
R278 S.n660 S.t1018 3.904
R279 S.n12 S.n11 3.904
R280 S.n385 S.t643 3.904
R281 S.n388 S.t409 3.904
R282 S.n391 S.n390 3.904
R283 S.n3623 S.t53 3.904
R284 S.n3578 S.n3577 3.904
R285 S.n3593 S.t803 3.904
R286 S.n3596 S.t281 3.904
R287 S.n3581 S.n3580 3.904
R288 S.n3235 S.n3234 3.904
R289 S.n3246 S.t400 3.904
R290 S.n3243 S.t1040 3.904
R291 S.n3238 S.n3237 3.904
R292 S.n2941 S.n2940 3.904
R293 S.n2961 S.t626 3.904
R294 S.n2958 S.t1099 3.904
R295 S.n2944 S.n2943 3.904
R296 S.n2716 S.n2715 3.904
R297 S.n2727 S.t148 3.904
R298 S.n2724 S.t979 3.904
R299 S.n2719 S.n2718 3.904
R300 S.n2403 S.n2402 3.904
R301 S.n2423 S.t467 3.904
R302 S.n2420 S.t590 3.904
R303 S.n2406 S.n2405 3.904
R304 S.n2220 S.n2219 3.904
R305 S.n2231 S.t17 3.904
R306 S.n2228 S.t968 3.904
R307 S.n2223 S.n2222 3.904
R308 S.n1911 S.n1910 3.904
R309 S.n1931 S.t456 3.904
R310 S.n1928 S.t571 3.904
R311 S.n1914 S.n1913 3.904
R312 S.n1624 S.n1623 3.904
R313 S.n1635 S.t1146 3.904
R314 S.n1632 S.t953 3.904
R315 S.n1627 S.n1626 3.904
R316 S.n1361 S.n1360 3.904
R317 S.n1381 S.t446 3.904
R318 S.n1378 S.t555 3.904
R319 S.n1364 S.n1363 3.904
R320 S.n1064 S.n1063 3.904
R321 S.n1077 S.t1131 3.904
R322 S.n1074 S.t1125 3.904
R323 S.n1067 S.n1066 3.904
R324 S.n1083 S.n1082 3.904
R325 S.n1097 S.t741 3.904
R326 S.n1094 S.t740 3.904
R327 S.n1086 S.n1085 3.904
R328 S.n832 S.n831 3.904
R329 S.n856 S.t277 3.904
R330 S.n853 S.t1144 3.904
R331 S.n835 S.n834 3.904
R332 S.n79 S.n78 3.904
R333 S.n281 S.t652 3.904
R334 S.n284 S.t721 3.904
R335 S.n287 S.n286 3.904
R336 S.n295 S.n294 3.904
R337 S.n310 S.t263 3.904
R338 S.n307 S.t1128 3.904
R339 S.n298 S.n297 3.904
R340 S.n567 S.t644 3.904
R341 S.n1399 S.n1398 3.904
R342 S.n1416 S.t24 3.904
R343 S.n1413 S.t163 3.904
R344 S.n1396 S.n1395 3.904
R345 S.n1948 S.n1947 3.904
R346 S.n1963 S.t48 3.904
R347 S.n1960 S.t177 3.904
R348 S.n1945 S.n1944 3.904
R349 S.n2440 S.n2439 3.904
R350 S.n2455 S.t67 3.904
R351 S.n2452 S.t193 3.904
R352 S.n2437 S.n2436 3.904
R353 S.n2978 S.n2977 3.904
R354 S.n2993 S.t79 3.904
R355 S.n2990 S.t208 3.904
R356 S.n2975 S.n2974 3.904
R357 S.n3464 S.n3463 3.904
R358 S.n3479 S.t481 3.904
R359 S.n3476 S.t1009 3.904
R360 S.n3461 S.n3460 3.904
R361 S.n4051 S.n4050 3.904
R362 S.n4065 S.t563 3.904
R363 S.n4068 S.t139 3.904
R364 S.n4048 S.n4047 3.904
R365 S.n4231 S.t1042 3.904
R366 S.n3631 S.n3630 3.904
R367 S.n3642 S.t291 3.904
R368 S.n3639 S.t796 3.904
R369 S.n3628 S.n3627 3.904
R370 S.n3254 S.n3253 3.904
R371 S.n3265 S.t1121 3.904
R372 S.n3262 S.t615 3.904
R373 S.n3251 S.n3250 3.904
R374 S.n2735 S.n2734 3.904
R375 S.n2746 S.t788 3.904
R376 S.n2743 S.t602 3.904
R377 S.n2732 S.n2731 3.904
R378 S.n2239 S.n2238 3.904
R379 S.n2250 S.t771 3.904
R380 S.n2247 S.t591 3.904
R381 S.n2236 S.n2235 3.904
R382 S.n1643 S.n1642 3.904
R383 S.n1654 S.t757 3.904
R384 S.n1651 S.t573 3.904
R385 S.n1640 S.n1639 3.904
R386 S.n871 S.n870 3.904
R387 S.n890 S.t995 3.904
R388 S.n887 S.t756 3.904
R389 S.n874 S.n873 3.904
R390 S.n205 S.n204 3.904
R391 S.n220 S.t278 3.904
R392 S.n217 S.t339 3.904
R393 S.n208 S.n207 3.904
R394 S.n583 S.n582 3.904
R395 S.n586 S.t983 3.904
R396 S.n589 S.t744 3.904
R397 S.n592 S.n591 3.904
R398 S.n578 S.t265 3.904
R399 S.n4685 S.t932 3.904
R400 S.n4492 S.n4491 3.904
R401 S.n4500 S.t432 3.904
R402 S.n4503 S.t1107 3.904
R403 S.n4489 S.n4488 3.904
R404 S.n4244 S.n4243 3.904
R405 S.n4252 S.t155 3.904
R406 S.n4249 S.t666 3.904
R407 S.n4241 S.n4240 3.904
R408 S.n3969 S.n3968 3.904
R409 S.n3987 S.t246 3.904
R410 S.n3984 S.t864 3.904
R411 S.n3966 S.n3965 3.904
R412 S.n3655 S.n3654 3.904
R413 S.n3663 S.t1019 3.904
R414 S.n3660 S.t623 3.904
R415 S.n3652 S.n3651 3.904
R416 S.n3495 S.n3494 3.904
R417 S.n3513 S.t828 3.904
R418 S.n3510 S.t945 3.904
R419 S.n3492 S.n3491 3.904
R420 S.n3278 S.n3277 3.904
R421 S.n3286 S.t424 3.904
R422 S.n3283 S.t227 3.904
R423 S.n3275 S.n3274 3.904
R424 S.n3009 S.n3008 3.904
R425 S.n3027 S.t817 3.904
R426 S.n3024 S.t930 3.904
R427 S.n3006 S.n3005 3.904
R428 S.n2759 S.n2758 3.904
R429 S.n2767 S.t406 3.904
R430 S.n2764 S.t209 3.904
R431 S.n2756 S.n2755 3.904
R432 S.n2471 S.n2470 3.904
R433 S.n2489 S.t807 3.904
R434 S.n2486 S.t916 3.904
R435 S.n2468 S.n2467 3.904
R436 S.n2263 S.n2262 3.904
R437 S.n2271 S.t390 3.904
R438 S.n2268 S.t194 3.904
R439 S.n2260 S.n2259 3.904
R440 S.n1979 S.n1978 3.904
R441 S.n1997 S.t790 3.904
R442 S.n1994 S.t901 3.904
R443 S.n1976 S.n1975 3.904
R444 S.n1667 S.n1666 3.904
R445 S.n1675 S.t370 3.904
R446 S.n1672 S.t176 3.904
R447 S.n1664 S.n1663 3.904
R448 S.n1432 S.n1431 3.904
R449 S.n1450 S.t774 3.904
R450 S.n1447 S.t964 3.904
R451 S.n1429 S.n1428 3.904
R452 S.n1110 S.n1109 3.904
R453 S.n1118 S.t439 3.904
R454 S.n1115 S.t356 3.904
R455 S.n1107 S.n1106 3.904
R456 S.n899 S.n898 3.904
R457 S.n918 S.t620 3.904
R458 S.n915 S.t372 3.904
R459 S.n902 S.n901 3.904
R460 S.n225 S.n224 3.904
R461 S.n239 S.t997 3.904
R462 S.n236 S.t1067 3.904
R463 S.n228 S.n227 3.904
R464 S.n1129 S.n1128 3.904
R465 S.n1138 S.t7 3.904
R466 S.n1135 S.t1081 3.904
R467 S.n1126 S.n1125 3.904
R468 S.n1459 S.n1458 3.904
R469 S.n1471 S.t388 3.904
R470 S.n1468 S.t583 3.904
R471 S.n1462 S.n1461 3.904
R472 S.n1681 S.n1680 3.904
R473 S.n1695 S.t40 3.904
R474 S.n1692 S.t900 3.904
R475 S.n1684 S.n1683 3.904
R476 S.n2006 S.n2005 3.904
R477 S.n2017 S.t410 3.904
R478 S.n2014 S.t599 3.904
R479 S.n2009 S.n2008 3.904
R480 S.n2277 S.n2276 3.904
R481 S.n2291 S.t1109 3.904
R482 S.n2288 S.t915 3.904
R483 S.n2280 S.n2279 3.904
R484 S.n2498 S.n2497 3.904
R485 S.n2509 S.t426 3.904
R486 S.n2506 S.t539 3.904
R487 S.n2501 S.n2500 3.904
R488 S.n2773 S.n2772 3.904
R489 S.n2787 S.t1126 3.904
R490 S.n2784 S.t933 3.904
R491 S.n2776 S.n2775 3.904
R492 S.n3036 S.n3035 3.904
R493 S.n3047 S.t441 3.904
R494 S.n3044 S.t552 3.904
R495 S.n3039 S.n3038 3.904
R496 S.n3292 S.n3291 3.904
R497 S.n3306 S.t1141 3.904
R498 S.n3303 S.t949 3.904
R499 S.n3295 S.n3294 3.904
R500 S.n3522 S.n3521 3.904
R501 S.n3533 S.t453 3.904
R502 S.n3530 S.t567 3.904
R503 S.n3525 S.n3524 3.904
R504 S.n3669 S.n3668 3.904
R505 S.n3683 S.t11 3.904
R506 S.n3680 S.t235 3.904
R507 S.n3672 S.n3671 3.904
R508 S.n3996 S.n3995 3.904
R509 S.n4007 S.t835 3.904
R510 S.n4004 S.t585 3.904
R511 S.n3999 S.n3998 3.904
R512 S.n4258 S.n4257 3.904
R513 S.n4272 S.t884 3.904
R514 S.n4269 S.t248 3.904
R515 S.n4261 S.n4260 3.904
R516 S.n4433 S.n4432 3.904
R517 S.n4444 S.t96 3.904
R518 S.n4441 S.t714 3.904
R519 S.n4436 S.n4435 3.904
R520 S.n4691 S.n4690 3.904
R521 S.n4705 S.t1127 3.904
R522 S.n4702 S.t554 3.904
R523 S.n4694 S.n4693 3.904
R524 S.n5503 S.n5502 3.904
R525 S.n5511 S.t298 3.904
R526 S.n5514 S.t1013 3.904
R527 S.n5506 S.n5505 3.904
R528 S.n5673 S.t800 3.904
R529 S.n626 S.t985 3.904
R530 S.n315 S.n314 3.904
R531 S.n332 S.t606 3.904
R532 S.n329 S.t358 3.904
R533 S.n318 S.n317 3.904
R534 S.n803 S.n802 3.904
R535 S.n822 S.t651 3.904
R536 S.n819 S.t346 3.904
R537 S.n806 S.n805 3.904
R538 S.n189 S.n188 3.904
R539 S.n200 S.t978 3.904
R540 S.n197 S.t1111 3.904
R541 S.n192 S.n191 3.904
R542 S.n172 S.n171 3.904
R543 S.n183 S.t256 3.904
R544 S.n180 S.t389 3.904
R545 S.n175 S.n174 3.904
R546 S.n541 S.t1003 3.904
R547 S.n43 S.n42 3.904
R548 S.n54 S.t659 3.904
R549 S.n51 S.t381 3.904
R550 S.n46 S.n45 3.904
R551 S.n722 S.n721 3.904
R552 S.n735 S.t665 3.904
R553 S.n732 S.t399 3.904
R554 S.n719 S.n718 3.904
R555 S.n2178 S.t592 3.904
R556 S.n2058 S.n2057 3.904
R557 S.n2072 S.t56 3.904
R558 S.n2075 S.t654 3.904
R559 S.n2055 S.n2054 3.904
R560 S.n1571 S.n1570 3.904
R561 S.n1582 S.t777 3.904
R562 S.n1579 S.t307 3.904
R563 S.n1568 S.n1567 3.904
R564 S.n1272 S.n1271 3.904
R565 S.n1289 S.t996 3.904
R566 S.n1286 S.t371 3.904
R567 S.n1269 S.n1268 3.904
R568 S.n1015 S.n1014 3.904
R569 S.n1024 S.t533 3.904
R570 S.n1021 S.t49 3.904
R571 S.n1012 S.n1011 3.904
R572 S.n656 S.t628 3.904
R573 S.n413 S.n412 3.904
R574 S.n416 S.t290 3.904
R575 S.n419 S.t1102 3.904
R576 S.n422 S.n421 3.904
R577 S.n2691 S.t454 3.904
R578 S.n2554 S.n2553 3.904
R579 S.n2569 S.t1043 3.904
R580 S.n2572 S.t524 3.904
R581 S.n2557 S.n2556 3.904
R582 S.n2184 S.n2183 3.904
R583 S.n2195 S.t658 3.904
R584 S.n2192 S.t195 3.904
R585 S.n2187 S.n2186 3.904
R586 S.n1850 S.n1849 3.904
R587 S.n1870 S.t856 3.904
R588 S.n1867 S.t280 3.904
R589 S.n1853 S.n1852 3.904
R590 S.n1588 S.n1587 3.904
R591 S.n1599 S.t395 3.904
R592 S.n1596 S.t618 3.904
R593 S.n1591 S.n1590 3.904
R594 S.n1298 S.n1297 3.904
R595 S.n1318 S.t81 3.904
R596 S.n1315 S.t210 3.904
R597 S.n1301 S.n1300 3.904
R598 S.n1030 S.n1029 3.904
R599 S.n1041 S.t792 3.904
R600 S.n1038 S.t791 3.904
R601 S.n1033 S.n1032 3.904
R602 S.n744 S.n743 3.904
R603 S.n764 S.t294 3.904
R604 S.n761 S.t1118 3.904
R605 S.n747 S.n746 3.904
R606 S.n156 S.n155 3.904
R607 S.n167 S.t638 3.904
R608 S.n164 S.t776 3.904
R609 S.n159 S.n158 3.904
R610 S.n139 S.n138 3.904
R611 S.n150 S.t1011 3.904
R612 S.n147 S.t27 3.904
R613 S.n142 S.n141 3.904
R614 S.n528 S.t672 3.904
R615 S.n22 S.n21 3.904
R616 S.n33 S.t1022 3.904
R617 S.n30 S.t553 3.904
R618 S.n25 S.n24 3.904
R619 S.n949 S.n948 3.904
R620 S.n961 S.t99 3.904
R621 S.n964 S.t799 3.904
R622 S.n946 S.n945 3.904
R623 S.n990 S.t629 3.904
R624 S.n652 S.t279 3.904
R625 S.n444 S.n443 3.904
R626 S.n447 S.t1035 3.904
R627 S.n450 S.t766 3.904
R628 S.n453 S.n452 3.904
R629 S.n1563 S.t677 3.904
R630 S.n1518 S.n1517 3.904
R631 S.n1533 S.t206 3.904
R632 S.n1536 S.t755 3.904
R633 S.n1521 S.n1520 3.904
R634 S.n996 S.n995 3.904
R635 S.n1007 S.t907 3.904
R636 S.n1004 S.t244 3.904
R637 S.n999 S.n998 3.904
R638 S.n685 S.n684 3.904
R639 S.n705 S.t887 3.904
R640 S.n702 S.t419 3.904
R641 S.n688 S.n687 3.904
R642 S.n123 S.n122 3.904
R643 S.n134 S.t578 3.904
R644 S.n131 S.t447 3.904
R645 S.n126 S.n125 3.904
R646 S.n106 S.n105 3.904
R647 S.n117 S.t961 3.904
R648 S.n114 S.t327 3.904
R649 S.n109 S.n108 3.904
R650 S.n380 S.t219 3.904
R651 S.n382 S.t397 3.904
R652 S.n265 S.n264 3.904
R653 S.n275 S.t1051 3.904
R654 S.n278 S.t1117 3.904
R655 S.n268 S.n267 3.904
R656 S.n1189 S.n1188 3.904
R657 S.n1197 S.t954 3.904
R658 S.n1200 S.t260 3.904
R659 S.n1192 S.n1191 3.904
R660 S.n968 S.n967 3.904
R661 S.n1175 S.t382 3.904
R662 S.n1178 S.t315 3.904
R663 S.n1181 S.n1180 3.904
R664 S.n1753 S.n1752 3.904
R665 S.n1765 S.t720 3.904
R666 S.n1768 S.t912 3.904
R667 S.n1756 S.n1755 3.904
R668 S.n1540 S.n1539 3.904
R669 S.n1738 S.t398 3.904
R670 S.n1741 S.t142 3.904
R671 S.n1744 S.n1743 3.904
R672 S.n2097 S.n2096 3.904
R673 S.n2109 S.t738 3.904
R674 S.n2112 S.t926 3.904
R675 S.n2100 S.n2099 3.904
R676 S.n2079 S.n2078 3.904
R677 S.n2082 S.t417 3.904
R678 S.n2085 S.t150 3.904
R679 S.n2088 S.n2087 3.904
R680 S.n2594 S.n2593 3.904
R681 S.n2606 S.t752 3.904
R682 S.n2609 S.t943 3.904
R683 S.n2597 S.n2596 3.904
R684 S.n2576 S.n2575 3.904
R685 S.n2579 S.t435 3.904
R686 S.n2582 S.t161 3.904
R687 S.n2585 S.n2584 3.904
R688 S.n3127 S.n3126 3.904
R689 S.n3139 S.t770 3.904
R690 S.n3142 S.t962 3.904
R691 S.n3130 S.n3129 3.904
R692 S.n3109 S.n3108 3.904
R693 S.n3112 S.t366 3.904
R694 S.n3115 S.t174 3.904
R695 S.n3118 S.n3117 3.904
R696 S.n3804 S.n3803 3.904
R697 S.n3816 S.t787 3.904
R698 S.n3819 S.t899 3.904
R699 S.n3807 S.n3806 3.904
R700 S.n3600 S.n3599 3.904
R701 S.n3789 S.t387 3.904
R702 S.n3792 S.t577 3.904
R703 S.n3795 S.n3794 3.904
R704 S.n4090 S.n4089 3.904
R705 S.n4102 S.t55 3.904
R706 S.n4105 S.t914 3.904
R707 S.n4093 S.n4092 3.904
R708 S.n4072 S.n4071 3.904
R709 S.n4075 S.t403 3.904
R710 S.n4078 S.t594 3.904
R711 S.n4081 S.n4080 3.904
R712 S.n4525 S.n4524 3.904
R713 S.n4537 S.t72 3.904
R714 S.n4540 S.t928 3.904
R715 S.n4528 S.n4527 3.904
R716 S.n4507 S.n4506 3.904
R717 S.n4510 S.t418 3.904
R718 S.n4513 S.t604 3.904
R719 S.n4516 S.n4515 3.904
R720 S.n5519 S.n5518 3.904
R721 S.n5531 S.t84 3.904
R722 S.n5534 S.t946 3.904
R723 S.n5522 S.n5521 3.904
R724 S.n5721 S.n5720 3.904
R725 S.n5731 S.t649 3.904
R726 S.n5734 S.t619 3.904
R727 S.n5724 S.n5723 3.904
R728 S.n5198 S.n5197 3.904
R729 S.n5213 S.t873 3.904
R730 S.n5210 S.t493 3.904
R731 S.n5201 S.n5200 3.904
R732 S.n4999 S.n4998 3.904
R733 S.n5183 S.t385 3.904
R734 S.n5186 S.t224 3.904
R735 S.n5189 S.n5188 3.904
R736 S.n5359 S.t645 3.904
R737 S.n5353 S.t812 3.904
R738 S.n1203 S.t688 3.904
R739 S.n1205 S.t1133 3.904
R740 S.n1161 S.n1160 3.904
R741 S.n1169 S.t160 3.904
R742 S.n1172 S.t520 3.904
R743 S.n1164 S.n1163 3.904
R744 S.n1776 S.n1775 3.904
R745 S.n1795 S.t341 3.904
R746 S.n1798 S.t445 3.904
R747 S.n1773 S.n1772 3.904
R748 S.n5369 S.t270 3.904
R749 S.n5364 S.t489 3.904
R750 S.n4986 S.n4985 3.904
R751 S.n4983 S.t1106 3.904
R752 S.n4980 S.t935 3.904
R753 S.n4977 S.n4976 3.904
R754 S.n4972 S.n4971 3.904
R755 S.n4995 S.t431 3.904
R756 S.n4992 S.t586 3.904
R757 S.n4969 S.n4968 3.904
R758 S.n5742 S.n5741 3.904
R759 S.n5746 S.t5 3.904
R760 S.n5749 S.t231 3.904
R761 S.n5739 S.n5738 3.904
R762 S.n5542 S.n5541 3.904
R763 S.n5547 S.t820 3.904
R764 S.n5550 S.t565 3.904
R765 S.n5539 S.n5538 3.904
R766 S.n4562 S.n4561 3.904
R767 S.n4559 S.t1137 3.904
R768 S.n4556 S.t213 3.904
R769 S.n4553 S.n4552 3.904
R770 S.n4548 S.n4547 3.904
R771 S.n4568 S.t810 3.904
R772 S.n4571 S.t549 3.904
R773 S.n4545 S.n4544 3.904
R774 S.n4127 S.n4126 3.904
R775 S.n4124 S.t1123 3.904
R776 S.n4121 S.t197 3.904
R777 S.n4118 S.n4117 3.904
R778 S.n4113 S.n4112 3.904
R779 S.n4133 S.t795 3.904
R780 S.n4136 S.t536 3.904
R781 S.n4110 S.n4109 3.904
R782 S.n3841 S.n3840 3.904
R783 S.n3838 S.t1104 3.904
R784 S.n3835 S.t183 3.904
R785 S.n3832 S.n3831 3.904
R786 S.n3827 S.n3826 3.904
R787 S.n3847 S.t405 3.904
R788 S.n3850 S.t596 3.904
R789 S.n3824 S.n3823 3.904
R790 S.n3164 S.n3163 3.904
R791 S.n3161 S.t32 3.904
R792 S.n3158 S.t898 3.904
R793 S.n3155 S.n3154 3.904
R794 S.n3150 S.n3149 3.904
R795 S.n3170 S.t386 3.904
R796 S.n3173 S.t582 3.904
R797 S.n3147 S.n3146 3.904
R798 S.n2631 S.n2630 3.904
R799 S.n2628 S.t1 3.904
R800 S.n2625 S.t888 3.904
R801 S.n2622 S.n2621 3.904
R802 S.n2617 S.n2616 3.904
R803 S.n2637 S.t367 3.904
R804 S.n2640 S.t564 3.904
R805 S.n2614 S.n2613 3.904
R806 S.n2137 S.n2136 3.904
R807 S.n2134 S.t1135 3.904
R808 S.n2131 S.t879 3.904
R809 S.n2128 S.n2127 3.904
R810 S.n2123 S.n2122 3.904
R811 S.n2120 S.t355 3.904
R812 S.n2143 S.t548 3.904
R813 S.n2117 S.n2116 3.904
R814 S.n1790 S.n1789 3.904
R815 S.n1787 S.t1120 3.904
R816 S.n1784 S.t867 3.904
R817 S.n1781 S.n1780 3.904
R818 S.n1803 S.t74 3.904
R819 S.n1800 S.t948 3.904
R820 S.n1720 S.n1719 3.904
R821 S.n1732 S.t664 3.904
R822 S.n1735 S.t1083 3.904
R823 S.n1723 S.n1722 3.904
R824 S.n2151 S.n2150 3.904
R825 S.n2345 S.t1082 3.904
R826 S.n2348 S.t955 3.904
R827 S.n2148 S.n2147 3.904
R828 S.n5377 S.t869 3.904
R829 S.n5371 S.t732 3.904
R830 S.n5053 S.n5052 3.904
R831 S.n5058 S.t736 3.904
R832 S.n5061 S.t556 3.904
R833 S.n5050 S.n5049 3.904
R834 S.n4957 S.n4956 3.904
R835 S.n4964 S.t1147 3.904
R836 S.n4961 S.t186 3.904
R837 S.n4954 S.n4953 3.904
R838 S.n5757 S.n5756 3.904
R839 S.n5762 S.t765 3.904
R840 S.n5765 S.t960 3.904
R841 S.n5754 S.n5753 3.904
R842 S.n5558 S.n5557 3.904
R843 S.n5562 S.t449 3.904
R844 S.n5565 S.t172 3.904
R845 S.n5555 S.n5554 3.904
R846 S.n4733 S.n4732 3.904
R847 S.n4738 S.t749 3.904
R848 S.n4741 S.t939 3.904
R849 S.n4730 S.n4729 3.904
R850 S.n4579 S.n4578 3.904
R851 S.n4583 S.t430 3.904
R852 S.n4586 S.t159 3.904
R853 S.n4576 S.n4575 3.904
R854 S.n4300 S.n4299 3.904
R855 S.n4305 S.t731 3.904
R856 S.n4308 S.t920 3.904
R857 S.n4297 S.n4296 3.904
R858 S.n4144 S.n4143 3.904
R859 S.n4148 S.t415 3.904
R860 S.n4151 S.t216 3.904
R861 S.n4141 S.n4140 3.904
R862 S.n3711 S.n3710 3.904
R863 S.n3716 S.t797 3.904
R864 S.n3719 S.t905 3.904
R865 S.n3708 S.n3707 3.904
R866 S.n3858 S.n3857 3.904
R867 S.n3862 S.t1122 3.904
R868 S.n3865 S.t201 3.904
R869 S.n3855 S.n3854 3.904
R870 S.n3334 S.n3333 3.904
R871 S.n3339 S.t780 3.904
R872 S.n3342 S.t525 3.904
R873 S.n3331 S.n3330 3.904
R874 S.n3181 S.n3180 3.904
R875 S.n3185 S.t1108 3.904
R876 S.n3188 S.t185 3.904
R877 S.n3178 S.n3177 3.904
R878 S.n2815 S.n2814 3.904
R879 S.n2820 S.t763 3.904
R880 S.n2823 S.t516 3.904
R881 S.n2812 S.n2811 3.904
R882 S.n2648 S.n2647 3.904
R883 S.n2652 S.t1091 3.904
R884 S.n2655 S.t171 3.904
R885 S.n2645 S.n2644 3.904
R886 S.n2340 S.n2339 3.904
R887 S.n2337 S.t748 3.904
R888 S.n2334 S.t502 3.904
R889 S.n2156 S.n2155 3.904
R890 S.n2353 S.t610 3.904
R891 S.n2350 S.t588 3.904
R892 S.n2316 S.n2315 3.904
R893 S.n2328 S.t51 3.904
R894 S.n2331 S.t490 3.904
R895 S.n2319 S.n2318 3.904
R896 S.n2663 S.n2662 3.904
R897 S.n2857 S.t706 3.904
R898 S.n2860 S.t321 3.904
R899 S.n2660 S.n2659 3.904
R900 S.n5385 S.t492 3.904
R901 S.n5379 S.t350 3.904
R902 S.n5069 S.n5068 3.904
R903 S.n5074 S.t352 3.904
R904 S.n5077 S.t164 3.904
R905 S.n5066 S.n5065 3.904
R906 S.n4942 S.n4941 3.904
R907 S.n4949 S.t758 3.904
R908 S.n4946 S.t909 3.904
R909 S.n4939 S.n4938 3.904
R910 S.n5773 S.n5772 3.904
R911 S.n5778 S.t383 3.904
R912 S.n5781 S.t574 3.904
R913 S.n5770 S.n5769 3.904
R914 S.n5573 S.n5572 3.904
R915 S.n5577 S.t26 3.904
R916 S.n5580 S.t897 3.904
R917 S.n5570 S.n5569 3.904
R918 S.n4749 S.n4748 3.904
R919 S.n4754 S.t363 3.904
R920 S.n4757 S.t558 3.904
R921 S.n4746 S.n4745 3.904
R922 S.n4594 S.n4593 3.904
R923 S.n4598 S.t1149 3.904
R924 S.n4601 S.t958 3.904
R925 S.n4591 S.n4590 3.904
R926 S.n4316 S.n4315 3.904
R927 S.n4321 S.t434 3.904
R928 S.n4324 S.t543 3.904
R929 S.n4313 S.n4312 3.904
R930 S.n4159 S.n4158 3.904
R931 S.n4163 S.t1134 3.904
R932 S.n4166 S.t941 3.904
R933 S.n4156 S.n4155 3.904
R934 S.n3727 S.n3726 3.904
R935 S.n3732 S.t416 3.904
R936 S.n3735 S.t531 3.904
R937 S.n3724 S.n3723 3.904
R938 S.n3873 S.n3872 3.904
R939 S.n3877 S.t733 3.904
R940 S.n3880 S.t923 3.904
R941 S.n3870 S.n3869 3.904
R942 S.n3350 S.n3349 3.904
R943 S.n3355 S.t396 3.904
R944 S.n3358 S.t137 3.904
R945 S.n3347 S.n3346 3.904
R946 S.n3196 S.n3195 3.904
R947 S.n3200 S.t717 3.904
R948 S.n3203 S.t908 3.904
R949 S.n3193 S.n3192 3.904
R950 S.n2852 S.n2851 3.904
R951 S.n2849 S.t379 3.904
R952 S.n2846 S.t124 3.904
R953 S.n2668 S.n2667 3.904
R954 S.n4609 S.n4608 3.904
R955 S.n4613 S.t760 3.904
R956 S.n4616 S.t576 3.904
R957 S.n4606 S.n4605 3.904
R958 S.n5393 S.t102 3.904
R959 S.n5387 S.t1077 3.904
R960 S.n5085 S.n5084 3.904
R961 S.n5090 S.t1076 3.904
R962 S.n5093 S.t889 3.904
R963 S.n5082 S.n5081 3.904
R964 S.n4927 S.n4926 3.904
R965 S.n4934 S.t374 3.904
R966 S.n4931 S.t534 3.904
R967 S.n4924 S.n4923 3.904
R968 S.n5789 S.n5788 3.904
R969 S.n5794 S.t1101 3.904
R970 S.n5797 S.t179 3.904
R971 S.n5786 S.n5785 3.904
R972 S.n5588 S.n5587 3.904
R973 S.n5592 S.t775 3.904
R974 S.n5595 S.t593 3.904
R975 S.n5585 S.n5584 3.904
R976 S.n4765 S.n4764 3.904
R977 S.n4770 S.t28 3.904
R978 S.n4773 S.t167 3.904
R979 S.n4762 S.n4761 3.904
R980 S.n4170 S.n4169 3.904
R981 S.n4178 S.t746 3.904
R982 S.n4181 S.t561 3.904
R983 S.n4173 S.n4172 3.904
R984 S.n3740 S.n3739 3.904
R985 S.n3748 S.t1132 3.904
R986 S.n3751 S.t144 3.904
R987 S.n3743 S.n3742 3.904
R988 S.n3884 S.n3883 3.904
R989 S.n3892 S.t351 3.904
R990 S.n3895 S.t545 3.904
R991 S.n3887 S.n3886 3.904
R992 S.n3207 S.n3206 3.904
R993 S.n3381 S.t1116 3.904
R994 S.n3384 S.t865 3.904
R995 S.n3387 S.n3386 3.904
R996 S.n3393 S.n3392 3.904
R997 S.n3401 S.t337 3.904
R998 S.n3404 S.t851 3.904
R999 S.n3396 S.n3395 3.904
R1000 S.n2828 S.n2827 3.904
R1001 S.n2840 S.t598 3.904
R1002 S.n2843 S.t1000 3.904
R1003 S.n2831 S.n2830 3.904
R1004 S.n2863 S.t1072 3.904
R1005 S.n2865 S.t207 3.904
R1006 S.n3409 S.t500 3.904
R1007 S.n3406 S.t944 3.904
R1008 S.n3363 S.n3362 3.904
R1009 S.n3375 S.t1058 3.904
R1010 S.n3378 S.t342 3.904
R1011 S.n3366 S.n3365 3.904
R1012 S.n3903 S.n3902 3.904
R1013 S.n3907 S.t1079 3.904
R1014 S.n3910 S.t274 3.904
R1015 S.n3900 S.n3899 3.904
R1016 S.n5401 S.t834 3.904
R1017 S.n5395 S.t690 3.904
R1018 S.n5101 S.n5100 3.904
R1019 S.n5106 S.t695 3.904
R1020 S.n5109 S.t518 3.904
R1021 S.n5098 S.n5097 3.904
R1022 S.n4912 S.n4911 3.904
R1023 S.n4919 S.t1095 3.904
R1024 S.n4916 S.t212 3.904
R1025 S.n4909 S.n4908 3.904
R1026 S.n5805 S.n5804 3.904
R1027 S.n5810 S.t794 3.904
R1028 S.n5813 S.t902 3.904
R1029 S.n5802 S.n5801 3.904
R1030 S.n5603 S.n5602 3.904
R1031 S.n5607 S.t394 3.904
R1032 S.n5610 S.t196 3.904
R1033 S.n5600 S.n5599 3.904
R1034 S.n4781 S.n4780 3.904
R1035 S.n4786 S.t778 3.904
R1036 S.n4789 S.t892 3.904
R1037 S.n4778 S.n4777 3.904
R1038 S.n4624 S.n4623 3.904
R1039 S.n4628 S.t375 3.904
R1040 S.n4631 S.t182 3.904
R1041 S.n4621 S.n4620 3.904
R1042 S.n4332 S.n4331 3.904
R1043 S.n4337 S.t759 3.904
R1044 S.n4340 S.t882 3.904
R1045 S.n4329 S.n4328 3.904
R1046 S.n4189 S.n4188 3.904
R1047 S.n4193 S.t360 3.904
R1048 S.n4196 S.t169 3.904
R1049 S.n4186 S.n4185 3.904
R1050 S.n3759 S.n3758 3.904
R1051 S.n3763 S.t747 3.904
R1052 S.n3766 S.t871 3.904
R1053 S.n3756 S.n3755 3.904
R1054 S.n3915 S.t1016 3.904
R1055 S.n3912 S.t584 3.904
R1056 S.n3771 S.n3770 3.904
R1057 S.n3783 S.t487 3.904
R1058 S.n3786 S.t1136 3.904
R1059 S.n3774 S.n3773 3.904
R1060 S.n4204 S.n4203 3.904
R1061 S.n4388 S.t1086 3.904
R1062 S.n4391 S.t739 3.904
R1063 S.n4201 S.n4200 3.904
R1064 S.n5409 S.t514 3.904
R1065 S.n5403 S.t313 3.904
R1066 S.n5117 S.n5116 3.904
R1067 S.n5122 S.t380 3.904
R1068 S.n5125 S.t125 3.904
R1069 S.n5114 S.n5113 3.904
R1070 S.n4897 S.n4896 3.904
R1071 S.n4904 S.t710 3.904
R1072 S.n4901 S.t938 3.904
R1073 S.n4894 S.n4893 3.904
R1074 S.n5821 S.n5820 3.904
R1075 S.n5826 S.t413 3.904
R1076 S.n5829 S.t529 3.904
R1077 S.n5818 S.n5817 3.904
R1078 S.n5618 S.n5617 3.904
R1079 S.n5622 S.t1114 3.904
R1080 S.n5625 S.t918 3.904
R1081 S.n5615 S.n5614 3.904
R1082 S.n4797 S.n4796 3.904
R1083 S.n4802 S.t393 3.904
R1084 S.n4805 S.t517 3.904
R1085 S.n4794 S.n4793 3.904
R1086 S.n4639 S.n4638 3.904
R1087 S.n4643 S.t1098 3.904
R1088 S.n4646 S.t904 3.904
R1089 S.n4636 S.n4635 3.904
R1090 S.n4383 S.n4382 3.904
R1091 S.n4380 S.t376 3.904
R1092 S.n4377 S.t506 3.904
R1093 S.n4209 S.n4208 3.904
R1094 S.n4396 S.t120 3.904
R1095 S.n4393 S.t203 3.904
R1096 S.n4345 S.n4344 3.904
R1097 S.n4357 S.t1006 3.904
R1098 S.n4360 S.t535 3.904
R1099 S.n4348 S.n4347 3.904
R1100 S.n4654 S.n4653 3.904
R1101 S.n4842 S.t709 3.904
R1102 S.n4845 S.t152 3.904
R1103 S.n4651 S.n4650 3.904
R1104 S.n5417 S.t122 3.904
R1105 S.n5411 S.t1045 3.904
R1106 S.n5133 S.n5132 3.904
R1107 S.n5138 S.t1097 3.904
R1108 S.n5141 S.t857 3.904
R1109 S.n5130 S.n5129 3.904
R1110 S.n4882 S.n4881 3.904
R1111 S.n4889 S.t328 3.904
R1112 S.n4886 S.t557 3.904
R1113 S.n4879 S.n4878 3.904
R1114 S.n5837 S.n5836 3.904
R1115 S.n5842 S.t1129 3.904
R1116 S.n5845 S.t140 3.904
R1117 S.n5834 S.n5833 3.904
R1118 S.n5633 S.n5632 3.904
R1119 S.n5637 S.t723 3.904
R1120 S.n5640 S.t542 3.904
R1121 S.n5630 S.n5629 3.904
R1122 S.n4837 S.n4836 3.904
R1123 S.n4834 S.t1115 3.904
R1124 S.n4831 S.t127 3.904
R1125 S.n4659 S.n4658 3.904
R1126 S.n4850 S.t650 3.904
R1127 S.n4847 S.t942 3.904
R1128 S.n4808 S.n4807 3.904
R1129 S.n4825 S.t373 3.904
R1130 S.n4828 S.t1029 3.904
R1131 S.n4811 S.n4810 3.904
R1132 S.n5864 S.n5863 3.904
R1133 S.n5873 S.t340 3.904
R1134 S.n5876 S.t661 3.904
R1135 S.n5867 S.n5866 3.904
R1136 S.n5425 S.t853 3.904
R1137 S.n5422 S.t668 3.904
R1138 S.n5146 S.n5145 3.904
R1139 S.n5154 S.t711 3.904
R1140 S.n5157 S.t480 3.904
R1141 S.n5149 S.n5148 3.904
R1142 S.n4863 S.n4862 3.904
R1143 S.n4874 S.t1054 3.904
R1144 S.n4871 S.t166 3.904
R1145 S.n4866 S.n4865 3.904
R1146 S.n5649 S.n5648 3.904
R1147 S.n5848 S.t745 3.904
R1148 S.n5851 S.t866 3.904
R1149 S.n5854 S.n5853 3.904
R1150 S.n5347 S.t250 3.904
R1151 S.n5345 S.t1028 3.904
R1152 S.n5169 S.n5168 3.904
R1153 S.n5177 S.t282 3.904
R1154 S.n5180 S.t507 3.904
R1155 S.n5172 S.n5171 3.904
R1156 S.n4370 S.n4369 3.904
R1157 S.n4374 S.t157 3.904
R1158 S.n4363 S.n4362 3.904
R1159 S.n4365 S.t1150 3.904
R1160 S.n4857 S.t218 3.643
R1161 S.n5438 S.t284 3.643
R1162 S.n5012 S.t1092 3.643
R1163 S.n5020 S.n5019 3.643
R1164 S.n5023 S.n5022 3.643
R1165 S.n5015 S.t369 3.643
R1166 S.n5251 S.t129 3.643
R1167 S.n5259 S.n5258 3.643
R1168 S.n5262 S.n5261 3.643
R1169 S.n5254 S.t676 3.643
R1170 S.n5698 S.t589 3.643
R1171 S.n5716 S.n5715 3.643
R1172 S.n5713 S.n5712 3.643
R1173 S.n5701 S.t1063 3.643
R1174 S.n5883 S.t999 3.643
R1175 S.n100 S.t991 3.643
R1176 S.n81 S.t1074 3.643
R1177 S.n477 S.t211 3.643
R1178 S.n480 S.n479 3.643
R1179 S.n483 S.n482 3.643
R1180 S.n486 S.t442 3.643
R1181 S.n650 S.t845 3.643
R1182 S.n651 S.t761 3.643
R1183 S.n647 S.t220 3.643
R1184 S.n643 S.t254 3.643
R1185 S.n342 S.t540 3.643
R1186 S.n353 S.n352 3.643
R1187 S.n350 S.n349 3.643
R1188 S.n345 S.t1073 3.643
R1189 S.n926 S.t192 3.643
R1190 S.n940 S.n939 3.643
R1191 S.n937 S.n936 3.643
R1192 S.n923 S.t429 3.643
R1193 S.n5028 S.t433 3.643
R1194 S.n5029 S.t929 3.643
R1195 S.n5223 S.t36 3.643
R1196 S.n5241 S.n5240 3.643
R1197 S.n5238 S.n5237 3.643
R1198 S.n5220 S.t296 3.643
R1199 S.n5681 S.t691 3.643
R1200 S.n5692 S.n5691 3.643
R1201 S.n5689 S.n5688 3.643
R1202 S.n5678 S.t779 3.643
R1203 S.n5474 S.t1012 3.643
R1204 S.n5489 S.n5488 3.643
R1205 S.n5486 S.n5485 3.643
R1206 S.n5471 S.t119 3.643
R1207 S.n4713 S.t510 3.643
R1208 S.n4724 S.n4723 3.643
R1209 S.n4721 S.n4720 3.643
R1210 S.n4710 S.t180 3.643
R1211 S.n4461 S.t359 3.643
R1212 S.n4476 S.n4475 3.643
R1213 S.n4473 S.n4472 3.643
R1214 S.n4458 S.t639 3.643
R1215 S.n4280 S.t497 3.643
R1216 S.n4291 S.n4290 3.643
R1217 S.n4288 S.n4287 3.643
R1218 S.n4277 S.t168 3.643
R1219 S.n4024 S.t344 3.643
R1220 S.n4039 S.n4038 3.643
R1221 S.n4036 S.n4035 3.643
R1222 S.n4021 S.t625 3.643
R1223 S.n3691 S.t486 3.643
R1224 S.n3702 S.n3701 3.643
R1225 S.n3699 S.n3698 3.643
R1226 S.n3688 S.t154 3.643
R1227 S.n3550 S.t1064 3.643
R1228 S.n3565 S.n3564 3.643
R1229 S.n3562 S.n3561 3.643
R1230 S.n3547 S.t614 3.643
R1231 S.n3317 S.t478 3.643
R1232 S.n3325 S.n3324 3.643
R1233 S.n3309 S.n3308 3.643
R1234 S.n3314 S.t145 3.643
R1235 S.n3064 S.t1052 3.643
R1236 S.n3079 S.n3078 3.643
R1237 S.n3076 S.n3075 3.643
R1238 S.n3061 S.t217 3.643
R1239 S.n2795 S.t469 3.643
R1240 S.n2806 S.n2805 3.643
R1241 S.n2803 S.n2802 3.643
R1242 S.n2792 S.t130 3.643
R1243 S.n2526 S.t1100 3.643
R1244 S.n2541 S.n2540 3.643
R1245 S.n2538 S.n2537 3.643
R1246 S.n2523 S.t275 3.643
R1247 S.n2299 S.t455 3.643
R1248 S.n2310 S.n2309 3.643
R1249 S.n2307 S.n2306 3.643
R1250 S.n2296 S.t116 3.643
R1251 S.n2034 S.t1088 3.643
R1252 S.n2049 S.n2048 3.643
R1253 S.n2046 S.n2045 3.643
R1254 S.n2031 S.t258 3.643
R1255 S.n1703 S.t444 3.643
R1256 S.n1714 S.n1713 3.643
R1257 S.n1711 S.n1710 3.643
R1258 S.n1700 S.t107 3.643
R1259 S.n1488 S.t1071 3.643
R1260 S.n1505 S.n1504 3.643
R1261 S.n1502 S.n1501 3.643
R1262 S.n1485 S.t245 3.643
R1263 S.n1146 S.t428 3.643
R1264 S.n1155 S.n1154 3.643
R1265 S.n1152 S.n1151 3.643
R1266 S.n1143 S.t92 3.643
R1267 S.n248 S.t271 3.643
R1268 S.n259 S.n258 3.643
R1269 S.n256 S.n255 3.643
R1270 S.n251 S.t1030 3.643
R1271 S.n559 S.t685 3.643
R1272 S.n552 S.t1032 3.643
R1273 S.n64 S.t921 3.643
R1274 S.n75 S.n74 3.643
R1275 S.n72 S.n71 3.643
R1276 S.n67 S.t3 3.643
R1277 S.n781 S.t940 3.643
R1278 S.n794 S.n793 3.643
R1279 S.n791 S.n790 3.643
R1280 S.n778 S.t34 3.643
R1281 S.n3228 S.t448 3.643
R1282 S.n3209 S.t575 3.643
R1283 S.n3088 S.t896 3.643
R1284 S.n3102 S.n3101 3.643
R1285 S.n3105 S.n3104 3.643
R1286 S.n3085 S.t1119 3.643
R1287 S.n2699 S.t257 3.643
R1288 S.n2710 S.n2709 3.643
R1289 S.n2707 S.n2706 3.643
R1290 S.n2696 S.t302 3.643
R1291 S.n2379 S.t653 3.643
R1292 S.n2394 S.n2393 3.643
R1293 S.n2391 S.n2390 3.643
R1294 S.n2376 S.t877 3.643
R1295 S.n2203 S.t135 3.643
R1296 S.n2214 S.n2213 3.643
R1297 S.n2211 S.n2210 3.643
R1298 S.n2200 S.t925 3.643
R1299 S.n1887 S.t719 3.643
R1300 S.n1902 S.n1901 3.643
R1301 S.n1899 S.n1898 3.643
R1302 S.n1884 S.t1001 3.643
R1303 S.n1607 S.t123 3.643
R1304 S.n1618 S.n1617 3.643
R1305 S.n1615 S.n1614 3.643
R1306 S.n1604 S.t910 3.643
R1307 S.n1335 S.t707 3.643
R1308 S.n1352 S.n1351 3.643
R1309 S.n1349 S.n1348 3.643
R1310 S.n1332 S.t987 3.643
R1311 S.n1049 S.t113 3.643
R1312 S.n1058 S.n1057 3.643
R1313 S.n1055 S.n1054 3.643
R1314 S.n1046 S.t895 3.643
R1315 S.n662 S.t312 3.643
R1316 S.n663 S.t657 3.643
R1317 S.n12 S.t613 3.643
R1318 S.n385 S.n384 3.643
R1319 S.n388 S.n387 3.643
R1320 S.n391 S.t831 3.643
R1321 S.n3622 S.t306 3.643
R1322 S.n3602 S.t443 3.643
R1323 S.n3578 S.t762 3.643
R1324 S.n3593 S.n3592 3.643
R1325 S.n3596 S.n3595 3.643
R1326 S.n3581 S.t885 3.643
R1327 S.n3235 S.t105 3.643
R1328 S.n3246 S.n3245 3.643
R1329 S.n3243 S.n3242 3.643
R1330 S.n3238 S.t181 3.643
R1331 S.n2941 S.t523 3.643
R1332 S.n2961 S.n2960 3.643
R1333 S.n2958 S.n2957 3.643
R1334 S.n2944 S.t728 3.643
R1335 S.n2716 S.t876 3.643
R1336 S.n2727 S.n2726 3.643
R1337 S.n2724 S.n2723 3.643
R1338 S.n2719 S.t562 3.643
R1339 S.n2403 S.t353 3.643
R1340 S.n2423 S.n2422 3.643
R1341 S.n2420 S.n2419 3.643
R1342 S.n2406 S.t634 3.643
R1343 S.n2220 S.t863 3.643
R1344 S.n2231 S.n2230 3.643
R1345 S.n2228 S.n2227 3.643
R1346 S.n2223 S.t547 3.643
R1347 S.n1911 S.t338 3.643
R1348 S.n1931 S.n1930 3.643
R1349 S.n1928 S.n1927 3.643
R1350 S.n1914 S.t624 3.643
R1351 S.n1624 S.t855 3.643
R1352 S.n1635 S.n1634 3.643
R1353 S.n1632 S.n1631 3.643
R1354 S.n1627 S.t532 3.643
R1355 S.n1361 S.t329 3.643
R1356 S.n1381 S.n1380 3.643
R1357 S.n1378 S.n1377 3.643
R1358 S.n1364 S.t608 3.643
R1359 S.n1064 S.t846 3.643
R1360 S.n1077 S.n1076 3.643
R1361 S.n1074 S.n1073 3.643
R1362 S.n1067 S.t522 3.643
R1363 S.n1083 S.t471 3.643
R1364 S.n1097 S.n1096 3.643
R1365 S.n1094 S.n1093 3.643
R1366 S.n1086 S.t132 3.643
R1367 S.n832 S.t236 3.643
R1368 S.n856 S.n855 3.643
R1369 S.n853 S.n852 3.643
R1370 S.n835 S.t468 3.643
R1371 S.n79 S.t292 3.643
R1372 S.n281 S.n280 3.643
R1373 S.n284 S.n283 3.643
R1374 S.n287 S.t1047 3.643
R1375 S.n295 S.t225 3.643
R1376 S.n310 S.n309 3.643
R1377 S.n307 S.n306 3.643
R1378 S.n298 S.t457 3.643
R1379 S.n574 S.t1044 3.643
R1380 S.n566 S.t286 3.643
R1381 S.n1399 S.t1053 3.643
R1382 S.n1416 S.n1415 3.643
R1383 S.n1413 S.n1412 3.643
R1384 S.n1396 S.t222 3.643
R1385 S.n1948 S.t1066 3.643
R1386 S.n1963 S.n1962 3.643
R1387 S.n1960 S.n1959 3.643
R1388 S.n1945 S.t234 3.643
R1389 S.n2440 S.t1080 3.643
R1390 S.n2455 S.n2454 3.643
R1391 S.n2452 S.n2451 3.643
R1392 S.n2437 S.t251 3.643
R1393 S.n2978 S.t1090 3.643
R1394 S.n2993 S.n2992 3.643
R1395 S.n2990 S.n2989 3.643
R1396 S.n2975 S.t264 3.643
R1397 S.n3464 S.t377 3.643
R1398 S.n3479 S.n3478 3.643
R1399 S.n3476 S.n3475 3.643
R1400 S.n3461 S.t505 3.643
R1401 S.n4051 S.t526 3.643
R1402 S.n4065 S.n4064 3.643
R1403 S.n4068 S.n4067 3.643
R1404 S.n4048 S.t737 3.643
R1405 S.n4230 S.t191 3.643
R1406 S.n4211 S.t305 3.643
R1407 S.n3631 S.t1069 3.643
R1408 S.n3642 S.n3641 3.643
R1409 S.n3639 S.n3638 3.643
R1410 S.n3628 S.t20 3.643
R1411 S.n3254 S.t512 3.643
R1412 S.n3265 S.n3264 3.643
R1413 S.n3262 S.n3261 3.643
R1414 S.n3251 S.t184 3.643
R1415 S.n2735 S.t499 3.643
R1416 S.n2746 S.n2745 3.643
R1417 S.n2743 S.n2742 3.643
R1418 S.n2732 S.t170 3.643
R1419 S.n2239 S.t488 3.643
R1420 S.n2250 S.n2249 3.643
R1421 S.n2247 S.n2246 3.643
R1422 S.n2236 S.t158 3.643
R1423 S.n1643 S.t479 3.643
R1424 S.n1654 S.n1653 3.643
R1425 S.n1651 S.n1650 3.643
R1426 S.n1640 S.t146 3.643
R1427 S.n871 S.t965 3.643
R1428 S.n890 S.n889 3.643
R1429 S.n887 S.n886 3.643
R1430 S.n874 S.t68 3.643
R1431 S.n205 S.t1020 3.643
R1432 S.n220 S.n219 3.643
R1433 S.n217 S.n216 3.643
R1434 S.n208 S.t670 3.643
R1435 S.n583 S.t947 3.643
R1436 S.n586 S.n585 3.643
R1437 S.n589 S.n588 3.643
R1438 S.n592 S.t50 3.643
R1439 S.n621 S.t667 3.643
R1440 S.n577 S.t1014 3.643
R1441 S.n4684 S.t37 3.643
R1442 S.n4661 S.t188 3.643
R1443 S.n4492 S.t384 3.643
R1444 S.n4500 S.n4499 3.643
R1445 S.n4503 S.n4502 3.643
R1446 S.n4489 S.t647 3.643
R1447 S.n4244 S.t982 3.643
R1448 S.n4252 S.n4251 3.643
R1449 S.n4249 S.n4248 3.643
R1450 S.n4241 S.t1034 3.643
R1451 S.n3969 S.t138 3.643
R1452 S.n3987 S.n3986 3.643
R1453 S.n3984 S.n3983 3.643
R1454 S.n3966 S.t354 3.643
R1455 S.n3655 S.t133 3.643
R1456 S.n3663 S.n3662 3.643
R1457 S.n3660 S.n3659 3.643
R1458 S.n3652 S.t922 3.643
R1459 S.n3495 S.t716 3.643
R1460 S.n3513 S.n3512 3.643
R1461 S.n3510 S.n3509 3.643
R1462 S.n3492 S.t268 3.643
R1463 S.n3278 S.t121 3.643
R1464 S.n3286 S.n3285 3.643
R1465 S.n3283 S.n3282 3.643
R1466 S.n3275 S.t906 3.643
R1467 S.n3009 S.t704 3.643
R1468 S.n3027 S.n3026 3.643
R1469 S.n3024 S.n3023 3.643
R1470 S.n3006 S.t986 3.643
R1471 S.n2759 S.t110 3.643
R1472 S.n2767 S.n2766 3.643
R1473 S.n2764 S.n2763 3.643
R1474 S.n2756 S.t893 3.643
R1475 S.n2471 S.t697 3.643
R1476 S.n2489 S.n2488 3.643
R1477 S.n2486 S.n2485 3.643
R1478 S.n2468 S.t971 3.643
R1479 S.n2263 S.t98 3.643
R1480 S.n2271 S.n2270 3.643
R1481 S.n2268 S.n2267 3.643
R1482 S.n2260 S.t886 3.643
R1483 S.n1979 S.t683 3.643
R1484 S.n1997 S.n1996 3.643
R1485 S.n1994 S.n1993 3.643
R1486 S.n1976 S.t963 3.643
R1487 S.n1667 S.t83 3.643
R1488 S.n1675 S.n1674 3.643
R1489 S.n1672 S.n1671 3.643
R1490 S.n1664 S.t874 3.643
R1491 S.n1432 S.t729 3.643
R1492 S.n1450 S.n1449 3.643
R1493 S.n1447 S.n1446 3.643
R1494 S.n1429 S.t1007 3.643
R1495 S.n1110 S.t69 3.643
R1496 S.n1118 S.n1117 3.643
R1497 S.n1115 S.n1114 3.643
R1498 S.n1107 S.t861 3.643
R1499 S.n899 S.t587 3.643
R1500 S.n918 S.n917 3.643
R1501 S.n915 S.n914 3.643
R1502 S.n902 S.t809 3.643
R1503 S.n225 S.t646 3.643
R1504 S.n239 S.n238 3.643
R1505 S.n236 S.n235 3.643
R1506 S.n228 S.t299 3.643
R1507 S.n1129 S.t808 3.643
R1508 S.n1138 S.n1137 3.643
R1509 S.n1135 S.n1134 3.643
R1510 S.n1126 S.t485 3.643
R1511 S.n1459 S.t348 3.643
R1512 S.n1471 S.n1470 3.643
R1513 S.n1468 S.n1467 3.643
R1514 S.n1462 S.t630 3.643
R1515 S.n1681 S.t818 3.643
R1516 S.n1695 S.n1694 3.643
R1517 S.n1692 S.n1691 3.643
R1518 S.n1684 S.t496 3.643
R1519 S.n2006 S.t362 3.643
R1520 S.n2017 S.n2016 3.643
R1521 S.n2014 S.n2013 3.643
R1522 S.n2009 S.t641 3.643
R1523 S.n2277 S.t832 3.643
R1524 S.n2291 S.n2290 3.643
R1525 S.n2288 S.n2287 3.643
R1526 S.n2280 S.t509 3.643
R1527 S.n2498 S.t314 3.643
R1528 S.n2509 S.n2508 3.643
R1529 S.n2506 S.n2505 3.643
R1530 S.n2501 S.t597 3.643
R1531 S.n2773 S.t843 3.643
R1532 S.n2787 S.n2786 3.643
R1533 S.n2784 S.n2783 3.643
R1534 S.n2776 S.t521 3.643
R1535 S.n3036 S.t326 3.643
R1536 S.n3047 S.n3046 3.643
R1537 S.n3044 S.n3043 3.643
R1538 S.n3039 S.t609 3.643
R1539 S.n3292 S.t854 3.643
R1540 S.n3306 S.n3305 3.643
R1541 S.n3303 S.n3302 3.643
R1542 S.n3295 S.t530 3.643
R1543 S.n3522 S.t335 3.643
R1544 S.n3533 S.n3532 3.643
R1545 S.n3530 S.n3529 3.643
R1546 S.n3525 S.t990 3.643
R1547 S.n3669 S.t862 3.643
R1548 S.n3683 S.n3682 3.643
R1549 S.n3680 S.n3679 3.643
R1550 S.n3672 S.t544 3.643
R1551 S.n3996 S.t724 3.643
R1552 S.n4007 S.n4006 3.643
R1553 S.n4004 S.n4003 3.643
R1554 S.n3999 S.t1004 3.643
R1555 S.n4258 S.t875 3.643
R1556 S.n4272 S.n4271 3.643
R1557 S.n4269 S.n4268 3.643
R1558 S.n4261 S.t560 3.643
R1559 S.n4433 S.t1105 3.643
R1560 S.n4444 S.n4443 3.643
R1561 S.n4441 S.n4440 3.643
R1562 S.n4436 S.t273 3.643
R1563 S.n4691 S.t844 3.643
R1564 S.n4705 S.n4704 3.643
R1565 S.n4702 S.n4701 3.643
R1566 S.n4694 S.t911 3.643
R1567 S.n5503 S.t285 3.643
R1568 S.n5511 S.n5510 3.643
R1569 S.n5514 S.n5513 3.643
R1570 S.n5506 S.t511 3.643
R1571 S.n5672 S.t1037 3.643
R1572 S.n5651 S.t30 3.643
R1573 S.n638 S.t295 3.643
R1574 S.n625 S.t640 3.643
R1575 S.n315 S.t569 3.643
R1576 S.n332 S.n331 3.643
R1577 S.n329 S.n328 3.643
R1578 S.n318 S.t793 3.643
R1579 S.n803 S.t559 3.643
R1580 S.n822 S.n821 3.643
R1581 S.n819 S.n818 3.643
R1582 S.n806 S.t781 3.643
R1583 S.n189 S.t662 3.643
R1584 S.n200 S.n199 3.643
R1585 S.n197 S.n196 3.643
R1586 S.n192 S.t316 3.643
R1587 S.n172 S.t1039 3.643
R1588 S.n183 S.n182 3.643
R1589 S.n180 S.n179 3.643
R1590 S.n175 S.t696 3.643
R1591 S.n547 S.t343 3.643
R1592 S.n540 S.t675 3.643
R1593 S.n43 S.t595 3.643
R1594 S.n54 S.n53 3.643
R1595 S.n51 S.n50 3.643
R1596 S.n46 S.t811 3.643
R1597 S.n722 S.t605 3.643
R1598 S.n735 S.n734 3.643
R1599 S.n732 S.n731 3.643
R1600 S.n719 S.t824 3.643
R1601 S.n2177 S.t673 3.643
R1602 S.n2158 S.t815 3.643
R1603 S.n2058 S.t1142 3.643
R1604 S.n2072 S.n2071 3.643
R1605 S.n2075 S.n2074 3.643
R1606 S.n2055 S.t287 3.643
R1607 S.n1571 S.t494 3.643
R1608 S.n1582 S.n1581 3.643
R1609 S.n1579 S.n1578 3.643
R1610 S.n1568 S.t568 3.643
R1611 S.n1272 S.t891 3.643
R1612 S.n1289 S.n1288 3.643
R1613 S.n1286 S.n1285 3.643
R1614 S.n1269 S.t1113 3.643
R1615 S.n1015 S.t878 3.643
R1616 S.n1024 S.n1023 3.643
R1617 S.n1021 S.n1020 3.643
R1618 S.n1012 S.t566 3.643
R1619 S.n658 S.t1065 3.643
R1620 S.n659 S.t303 3.643
R1621 S.n413 S.t199 3.643
R1622 S.n416 S.n415 3.643
R1623 S.n419 S.n418 3.643
R1624 S.n422 S.t436 3.643
R1625 S.n2690 S.t579 3.643
R1626 S.n2670 S.t674 3.643
R1627 S.n2554 S.t1027 3.643
R1628 S.n2569 S.n2568 3.643
R1629 S.n2572 S.n2571 3.643
R1630 S.n2557 S.t147 3.643
R1631 S.n2184 S.t336 3.643
R1632 S.n2195 S.n2194 3.643
R1633 S.n2192 S.n2191 3.643
R1634 S.n2187 S.t437 3.643
R1635 S.n1850 S.t754 3.643
R1636 S.n1870 S.n1869 3.643
R1637 S.n1867 S.n1866 3.643
R1638 S.n1853 S.t1015 3.643
R1639 S.n1588 S.t515 3.643
R1640 S.n1599 S.n1598 3.643
R1641 S.n1596 S.n1595 3.643
R1642 S.n1591 S.t187 3.643
R1643 S.n1298 S.t1093 3.643
R1644 S.n1318 S.n1317 3.643
R1645 S.n1315 S.n1314 3.643
R1646 S.n1301 S.t267 3.643
R1647 S.n1030 S.t501 3.643
R1648 S.n1041 S.n1040 3.643
R1649 S.n1038 S.n1037 3.643
R1650 S.n1033 S.t173 3.643
R1651 S.n744 S.t214 3.643
R1652 S.n764 S.n763 3.643
R1653 S.n761 S.n760 3.643
R1654 S.n747 S.t450 3.643
R1655 S.n156 S.t309 3.643
R1656 S.n167 S.n166 3.643
R1657 S.n164 S.n163 3.643
R1658 S.n159 S.t1084 3.643
R1659 S.n139 S.t680 3.643
R1660 S.n150 S.n149 3.643
R1661 S.n147 S.n146 3.643
R1662 S.n142 S.t357 3.643
R1663 S.n535 S.t1112 3.643
R1664 S.n527 S.t324 3.643
R1665 S.n22 S.t936 3.643
R1666 S.n33 S.n32 3.643
R1667 S.n30 S.n29 3.643
R1668 S.n25 S.t18 3.643
R1669 S.n949 S.t60 3.643
R1670 S.n961 S.n960 3.643
R1671 S.n964 S.n963 3.643
R1672 S.n946 S.t304 3.643
R1673 S.n989 S.t951 3.643
R1674 S.n970 S.t1046 3.643
R1675 S.n654 S.t722 3.643
R1676 S.n655 S.t1050 3.643
R1677 S.n444 S.t973 3.643
R1678 S.n447 S.n446 3.643
R1679 S.n450 S.n449 3.643
R1680 S.n453 S.t77 3.643
R1681 S.n1562 S.t814 3.643
R1682 S.n1542 S.t952 3.643
R1683 S.n1518 S.t165 3.643
R1684 S.n1533 S.n1532 3.643
R1685 S.n1536 S.n1535 3.643
R1686 S.n1521 S.t392 3.643
R1687 S.n996 S.t637 3.643
R1688 S.n1007 S.n1006 3.643
R1689 S.n1004 S.n1003 3.643
R1690 S.n999 S.t669 3.643
R1691 S.n685 S.t802 3.643
R1692 S.n705 S.n704 3.643
R1693 S.n702 S.n701 3.643
R1694 S.n688 S.t1033 3.643
R1695 S.n123 S.t1059 3.643
R1696 S.n134 S.n133 3.643
R1697 S.n131 S.n130 3.643
R1698 S.n126 S.t742 3.643
R1699 S.n106 S.t655 3.643
R1700 S.n117 S.n116 3.643
R1701 S.n114 S.n113 3.643
R1702 S.n109 S.t692 3.643
R1703 S.n522 S.t1078 3.643
R1704 S.n502 S.t112 3.643
R1705 S.n372 S.t822 3.643
R1706 S.n265 S.t718 3.643
R1707 S.n275 S.n274 3.643
R1708 S.n278 S.n277 3.643
R1709 S.n268 S.t679 3.643
R1710 S.n1189 S.t1036 3.643
R1711 S.n1197 S.n1196 3.643
R1712 S.n1200 S.n1199 3.643
R1713 S.n1192 S.t498 3.643
R1714 S.n968 S.t1148 3.643
R1715 S.n1175 S.n1174 3.643
R1716 S.n1178 S.n1177 3.643
R1717 S.n1181 S.t825 3.643
R1718 S.n1753 S.t689 3.643
R1719 S.n1765 S.n1764 3.643
R1720 S.n1768 S.n1767 3.643
R1721 S.n1756 S.t969 3.643
R1722 S.n1540 S.t22 3.643
R1723 S.n1738 S.n1737 3.643
R1724 S.n1741 S.n1740 3.643
R1725 S.n1744 S.t837 3.643
R1726 S.n2097 S.t701 3.643
R1727 S.n2109 S.n2108 3.643
R1728 S.n2112 S.n2111 3.643
R1729 S.n2100 S.t980 3.643
R1730 S.n2079 S.t46 3.643
R1731 S.n2082 S.n2081 3.643
R1732 S.n2085 S.n2084 3.643
R1733 S.n2088 S.t850 3.643
R1734 S.n2594 S.t712 3.643
R1735 S.n2606 S.n2605 3.643
R1736 S.n2609 S.n2608 3.643
R1737 S.n2597 S.t992 3.643
R1738 S.n2576 S.t61 3.643
R1739 S.n2579 S.n2578 3.643
R1740 S.n2582 S.n2581 3.643
R1741 S.n2585 S.t859 3.643
R1742 S.n3127 S.t726 3.643
R1743 S.n3139 S.n3138 3.643
R1744 S.n3142 S.n3141 3.643
R1745 S.n3130 S.t1005 3.643
R1746 S.n3109 S.t80 3.643
R1747 S.n3112 S.n3111 3.643
R1748 S.n3115 S.n3114 3.643
R1749 S.n3118 S.t872 3.643
R1750 S.n3804 S.t682 3.643
R1751 S.n3816 S.n3815 3.643
R1752 S.n3819 S.n3818 3.643
R1753 S.n3807 S.t226 3.643
R1754 S.n3600 S.t95 3.643
R1755 S.n3789 S.n3788 3.643
R1756 S.n3792 S.n3791 3.643
R1757 S.n3795 S.t883 3.643
R1758 S.n4090 S.t1068 3.643
R1759 S.n4102 S.n4101 3.643
R1760 S.n4105 S.n4104 3.643
R1761 S.n4093 S.t237 3.643
R1762 S.n4072 S.t108 3.643
R1763 S.n4075 S.n4074 3.643
R1764 S.n4078 S.n4077 3.643
R1765 S.n4081 S.t890 3.643
R1766 S.n4525 S.t1085 3.643
R1767 S.n4537 S.n4536 3.643
R1768 S.n4540 S.n4539 3.643
R1769 S.n4528 S.t253 3.643
R1770 S.n4507 S.t117 3.643
R1771 S.n4510 S.n4509 3.643
R1772 S.n4513 S.n4512 3.643
R1773 S.n4516 S.t903 3.643
R1774 S.n5519 S.t1096 3.643
R1775 S.n5531 S.n5530 3.643
R1776 S.n5534 S.n5533 3.643
R1777 S.n5522 S.t269 3.643
R1778 S.n5721 S.t131 3.643
R1779 S.n5731 S.n5730 3.643
R1780 S.n5734 S.n5733 3.643
R1781 S.n5724 S.t917 3.643
R1782 S.n5198 S.t782 3.643
R1783 S.n5213 S.n5212 3.643
R1784 S.n5210 S.n5209 3.643
R1785 S.n5201 S.t1026 3.643
R1786 S.n4999 S.t97 3.643
R1787 S.n5183 S.n5182 3.643
R1788 S.n5186 S.n5185 3.643
R1789 S.n5189 S.t550 3.643
R1790 S.n5352 S.t772 3.643
R1791 S.n1207 S.t459 3.643
R1792 S.n1161 S.t956 3.643
R1793 S.n1169 S.n1168 3.643
R1794 S.n1172 S.n1171 3.643
R1795 S.n1164 S.t475 3.643
R1796 S.n1776 S.t408 3.643
R1797 S.n1795 S.n1794 3.643
R1798 S.n1798 S.n1797 3.643
R1799 S.n1773 S.t989 3.643
R1800 S.n5365 S.t391 3.643
R1801 S.n4986 S.t842 3.643
R1802 S.n4983 S.n4982 3.643
R1803 S.n4980 S.n4979 3.643
R1804 S.n4977 S.t109 3.643
R1805 S.n4972 S.t317 3.643
R1806 S.n4995 S.n4994 3.643
R1807 S.n4992 S.n4991 3.643
R1808 S.n4969 S.t600 3.643
R1809 S.n5742 S.t860 3.643
R1810 S.n5746 S.n5745 3.643
R1811 S.n5749 S.n5748 3.643
R1812 S.n5739 S.t541 3.643
R1813 S.n5542 S.t708 3.643
R1814 S.n5547 S.n5546 3.643
R1815 S.n5550 S.n5549 3.643
R1816 S.n5539 S.t988 3.643
R1817 S.n4562 S.t852 3.643
R1818 S.n4559 S.n4558 3.643
R1819 S.n4556 S.n4555 3.643
R1820 S.n4553 S.t528 3.643
R1821 S.n4548 S.t699 3.643
R1822 S.n4568 S.n4567 3.643
R1823 S.n4571 S.n4570 3.643
R1824 S.n4545 S.t976 3.643
R1825 S.n4127 S.t840 3.643
R1826 S.n4124 S.n4123 3.643
R1827 S.n4121 S.n4120 3.643
R1828 S.n4118 S.t519 3.643
R1829 S.n4113 S.t686 3.643
R1830 S.n4133 S.n4132 3.643
R1831 S.n4136 S.n4135 3.643
R1832 S.n4110 S.t966 3.643
R1833 S.n3841 S.t829 3.643
R1834 S.n3838 S.n3837 3.643
R1835 S.n3835 S.n3834 3.643
R1836 S.n3832 S.t508 3.643
R1837 S.n3827 S.t361 3.643
R1838 S.n3847 S.n3846 3.643
R1839 S.n3850 S.n3849 3.643
R1840 S.n3824 S.t1010 3.643
R1841 S.n3164 S.t816 3.643
R1842 S.n3161 S.n3160 3.643
R1843 S.n3158 S.n3157 3.643
R1844 S.n3155 S.t495 3.643
R1845 S.n3150 S.t345 3.643
R1846 S.n3170 S.n3169 3.643
R1847 S.n3173 S.n3172 3.643
R1848 S.n3147 S.t627 3.643
R1849 S.n2631 S.t804 3.643
R1850 S.n2628 S.n2627 3.643
R1851 S.n2625 S.n2624 3.643
R1852 S.n2622 S.t483 3.643
R1853 S.n2617 S.t331 3.643
R1854 S.n2637 S.n2636 3.643
R1855 S.n2640 S.n2639 3.643
R1856 S.n2614 S.t616 3.643
R1857 S.n2137 S.t789 3.643
R1858 S.n2134 S.n2133 3.643
R1859 S.n2131 S.n2130 3.643
R1860 S.n2128 S.t474 3.643
R1861 S.n2123 S.t322 3.643
R1862 S.n2120 S.n2119 3.643
R1863 S.n2143 S.n2142 3.643
R1864 S.n2117 S.t603 3.643
R1865 S.n1790 S.t773 3.643
R1866 S.n1787 S.n1786 3.643
R1867 S.n1784 S.n1783 3.643
R1868 S.n1781 S.t463 3.643
R1869 S.n1255 S.t998 3.643
R1870 S.n1720 S.t318 3.643
R1871 S.n1732 S.n1731 3.643
R1872 S.n1735 S.n1734 3.643
R1873 S.n1723 S.t975 3.643
R1874 S.n2151 S.t919 3.643
R1875 S.n2345 S.n2344 3.643
R1876 S.n2348 S.n2347 3.643
R1877 S.n2148 S.t349 3.643
R1878 S.n5372 S.t663 3.643
R1879 S.n5053 S.t466 3.643
R1880 S.n5058 S.n5057 3.643
R1881 S.n5061 S.n5060 3.643
R1882 S.n5050 S.t841 3.643
R1883 S.n4957 S.t1048 3.643
R1884 S.n4964 S.n4963 3.643
R1885 S.n4961 S.n4960 3.643
R1886 S.n4954 S.t204 3.643
R1887 S.n5757 S.t484 3.643
R1888 S.n5762 S.n5761 3.643
R1889 S.n5765 S.n5764 3.643
R1890 S.n5754 S.t151 3.643
R1891 S.n5558 S.t330 3.643
R1892 S.n5562 S.n5561 3.643
R1893 S.n5565 S.n5564 3.643
R1894 S.n5555 S.t611 3.643
R1895 S.n4733 S.t476 3.643
R1896 S.n4738 S.n4737 3.643
R1897 S.n4741 S.n4740 3.643
R1898 S.n4730 S.t143 3.643
R1899 S.n4579 S.t319 3.643
R1900 S.n4583 S.n4582 3.643
R1901 S.n4586 S.n4585 3.643
R1902 S.n4576 S.t601 3.643
R1903 S.n4300 S.t464 3.643
R1904 S.n4305 S.n4304 3.643
R1905 S.n4308 S.n4307 3.643
R1906 S.n4297 S.t128 3.643
R1907 S.n4144 S.t365 3.643
R1908 S.n4148 S.n4147 3.643
R1909 S.n4151 S.n4150 3.643
R1910 S.n4141 S.t642 3.643
R1911 S.n3711 S.t452 3.643
R1912 S.n3716 S.n3715 3.643
R1913 S.n3719 S.n3718 3.643
R1914 S.n3708 S.t115 3.643
R1915 S.n3858 S.t1087 3.643
R1916 S.n3862 S.n3861 3.643
R1917 S.n3865 S.n3864 3.643
R1918 S.n3855 S.t633 3.643
R1919 S.n3334 S.t440 3.643
R1920 S.n3339 S.n3338 3.643
R1921 S.n3342 S.n3341 3.643
R1922 S.n3331 S.t104 3.643
R1923 S.n3181 S.t1070 3.643
R1924 S.n3185 S.n3184 3.643
R1925 S.n3188 S.n3187 3.643
R1926 S.n3178 S.t238 3.643
R1927 S.n2815 S.t425 3.643
R1928 S.n2820 S.n2819 3.643
R1929 S.n2823 S.n2822 3.643
R1930 S.n2812 S.t90 3.643
R1931 S.n2648 S.t1057 3.643
R1932 S.n2652 S.n2651 3.643
R1933 S.n2655 S.n2654 3.643
R1934 S.n2645 S.t228 3.643
R1935 S.n2340 S.t407 3.643
R1936 S.n2337 S.n2336 3.643
R1937 S.n2334 S.n2333 3.643
R1938 S.n2156 S.t76 3.643
R1939 S.n1841 S.t632 3.643
R1940 S.n2316 S.t849 3.643
R1941 S.n2328 S.n2327 3.643
R1942 S.n2331 S.n2330 3.643
R1943 S.n2319 S.t323 3.643
R1944 S.n2663 S.t308 3.643
R1945 S.n2857 S.n2856 3.643
R1946 S.n2860 S.n2859 3.643
R1947 S.n2660 S.t880 3.643
R1948 S.n5380 S.t293 3.643
R1949 S.n5069 S.t65 3.643
R1950 S.n5074 S.n5073 3.643
R1951 S.n5077 S.n5076 3.643
R1952 S.n5066 S.t465 3.643
R1953 S.n4942 S.t671 3.643
R1954 S.n4949 S.n4948 3.643
R1955 S.n4946 S.n4945 3.643
R1956 S.n4939 S.t927 3.643
R1957 S.n5773 S.t93 3.643
R1958 S.n5778 S.n5777 3.643
R1959 S.n5781 S.n5780 3.643
R1960 S.n5770 S.t881 3.643
R1961 S.n5573 S.t1056 3.643
R1962 S.n5577 S.n5576 3.643
R1963 S.n5580 S.n5579 3.643
R1964 S.n5570 S.t223 3.643
R1965 S.n4749 S.t78 3.643
R1966 S.n4754 S.n4753 3.643
R1967 S.n4757 S.n4756 3.643
R1968 S.n4746 S.t868 3.643
R1969 S.n4594 S.t1103 3.643
R1970 S.n4598 S.n4597 3.643
R1971 S.n4601 S.n4600 3.643
R1972 S.n4591 S.t276 3.643
R1973 S.n4316 S.t58 3.643
R1974 S.n4321 S.n4320 3.643
R1975 S.n4324 S.n4323 3.643
R1976 S.n4313 S.t858 3.643
R1977 S.n4159 S.t1089 3.643
R1978 S.n4163 S.n4162 3.643
R1979 S.n4166 S.n4165 3.643
R1980 S.n4156 S.t262 3.643
R1981 S.n3727 S.t41 3.643
R1982 S.n3732 S.n3731 3.643
R1983 S.n3735 S.n3734 3.643
R1984 S.n3724 S.t848 3.643
R1985 S.n3873 S.t700 3.643
R1986 S.n3877 S.n3876 3.643
R1987 S.n3880 S.n3879 3.643
R1988 S.n3870 S.t249 3.643
R1989 S.n3350 S.t13 3.643
R1990 S.n3355 S.n3354 3.643
R1991 S.n3358 S.n3357 3.643
R1992 S.n3347 S.t836 3.643
R1993 S.n3196 S.t687 3.643
R1994 S.n3200 S.n3199 3.643
R1995 S.n3203 S.n3202 3.643
R1996 S.n3193 S.t967 3.643
R1997 S.n2852 S.t1143 3.643
R1998 S.n2849 S.n2848 3.643
R1999 S.n2846 S.n2845 3.643
R2000 S.n2668 S.t823 3.643
R2001 S.n4609 S.t715 3.643
R2002 S.n4613 S.n4612 3.643
R2003 S.n4616 S.n4615 3.643
R2004 S.n4606 S.t994 3.643
R2005 S.n5388 S.t1021 3.643
R2006 S.n5085 S.t806 3.643
R2007 S.n5090 S.n5089 3.643
R2008 S.n5093 S.n5092 3.643
R2009 S.n5082 S.t63 3.643
R2010 S.n4927 S.t301 3.643
R2011 S.n4934 S.n4933 3.643
R2012 S.n4931 S.n4930 3.643
R2013 S.n4924 S.t546 3.643
R2014 S.n5789 S.t827 3.643
R2015 S.n5794 S.n5793 3.643
R2016 S.n5797 S.n5796 3.643
R2017 S.n5786 S.t504 3.643
R2018 S.n5588 S.t730 3.643
R2019 S.n5592 S.n5591 3.643
R2020 S.n5595 S.n5594 3.643
R2021 S.n5585 S.t1008 3.643
R2022 S.n4765 S.t813 3.643
R2023 S.n4770 S.n4769 3.643
R2024 S.n4773 S.n4772 3.643
R2025 S.n4762 S.t491 3.643
R2026 S.n4170 S.t703 3.643
R2027 S.n4178 S.n4177 3.643
R2028 S.n4181 S.n4180 3.643
R2029 S.n4173 S.t984 3.643
R2030 S.n3740 S.t786 3.643
R2031 S.n3748 S.n3747 3.643
R2032 S.n3751 S.n3750 3.643
R2033 S.n3743 S.t473 3.643
R2034 S.n3884 S.t320 3.643
R2035 S.n3892 S.n3891 3.643
R2036 S.n3895 S.n3894 3.643
R2037 S.n3887 S.t974 3.643
R2038 S.n3207 S.t769 3.643
R2039 S.n3381 S.n3380 3.643
R2040 S.n3384 S.n3383 3.643
R2041 S.n3387 S.t461 3.643
R2042 S.n3393 S.t826 3.643
R2043 S.n3401 S.n3400 3.643
R2044 S.n3404 S.n3403 3.643
R2045 S.n3396 S.t289 3.643
R2046 S.n2828 S.t272 3.643
R2047 S.n2840 S.n2839 3.643
R2048 S.n2843 S.n2842 3.643
R2049 S.n2831 S.t838 3.643
R2050 S.n2867 S.t261 3.643
R2051 S.n2932 S.t993 3.643
R2052 S.n3363 S.t734 3.643
R2053 S.n3375 S.n3374 3.643
R2054 S.n3378 S.n3377 3.643
R2055 S.n3366 S.t239 3.643
R2056 S.n3903 S.t240 3.643
R2057 S.n3907 S.n3906 3.643
R2058 S.n3910 S.n3909 3.643
R2059 S.n3900 S.t513 3.643
R2060 S.n5396 S.t648 3.643
R2061 S.n5101 S.t423 3.643
R2062 S.n5106 S.n5105 3.643
R2063 S.n5109 S.n5108 3.643
R2064 S.n5098 S.t805 3.643
R2065 S.n4912 S.t1061 3.643
R2066 S.n4919 S.n4918 3.643
R2067 S.n4916 S.n4915 3.643
R2068 S.n4909 S.t230 3.643
R2069 S.n5805 S.t451 3.643
R2070 S.n5810 S.n5809 3.643
R2071 S.n5813 S.n5812 3.643
R2072 S.n5802 S.t114 3.643
R2073 S.n5603 S.t347 3.643
R2074 S.n5607 S.n5606 3.643
R2075 S.n5610 S.n5609 3.643
R2076 S.n5600 S.t631 3.643
R2077 S.n4781 S.t438 3.643
R2078 S.n4786 S.n4785 3.643
R2079 S.n4789 S.n4788 3.643
R2080 S.n4778 S.t101 3.643
R2081 S.n4624 S.t333 3.643
R2082 S.n4628 S.n4627 3.643
R2083 S.n4631 S.n4630 3.643
R2084 S.n4621 S.t621 3.643
R2085 S.n4332 S.t421 3.643
R2086 S.n4337 S.n4336 3.643
R2087 S.n4340 S.n4339 3.643
R2088 S.n4329 S.t86 3.643
R2089 S.n4189 S.t325 3.643
R2090 S.n4193 S.n4192 3.643
R2091 S.n4196 S.n4195 3.643
R2092 S.n4186 S.t607 3.643
R2093 S.n3759 S.t404 3.643
R2094 S.n3763 S.n3762 3.643
R2095 S.n3766 S.n3765 3.643
R2096 S.n3756 S.t73 3.643
R2097 S.n3447 S.t1002 3.643
R2098 S.n3771 S.t153 3.643
R2099 S.n3783 S.n3782 3.643
R2100 S.n3786 S.n3785 3.643
R2101 S.n3774 S.t694 3.643
R2102 S.n4204 S.t462 3.643
R2103 S.n4388 S.n4387 3.643
R2104 S.n4391 S.n4390 3.643
R2105 S.n4201 S.t1024 3.643
R2106 S.n5404 S.t300 3.643
R2107 S.n5117 S.t1140 3.643
R2108 S.n5122 S.n5121 3.643
R2109 S.n5125 S.n5124 3.643
R2110 S.n5114 S.t422 3.643
R2111 S.n4897 S.t681 3.643
R2112 S.n4904 S.n4903 3.643
R2113 S.n4901 S.n4900 3.643
R2114 S.n4894 S.t957 3.643
R2115 S.n5821 S.t38 3.643
R2116 S.n5826 S.n5825 3.643
R2117 S.n5829 S.n5828 3.643
R2118 S.n5818 S.t847 3.643
R2119 S.n5618 S.t1075 3.643
R2120 S.n5622 S.n5621 3.643
R2121 S.n5625 S.n5624 3.643
R2122 S.n5615 S.t247 3.643
R2123 S.n4797 S.t9 3.643
R2124 S.n4802 S.n4801 3.643
R2125 S.n4805 S.n4804 3.643
R2126 S.n4794 S.t833 3.643
R2127 S.n4639 S.t1062 3.643
R2128 S.n4643 S.n4642 3.643
R2129 S.n4646 S.n4645 3.643
R2130 S.n4636 S.t233 3.643
R2131 S.n4383 S.t1139 3.643
R2132 S.n4380 S.n4379 3.643
R2133 S.n4377 S.n4376 3.643
R2134 S.n4209 S.t821 3.643
R2135 S.n3953 S.t635 3.643
R2136 S.n4345 S.t660 3.643
R2137 S.n4357 S.n4356 3.643
R2138 S.n4360 S.n4359 3.643
R2139 S.n4348 S.t94 3.643
R2140 S.n4654 S.t977 3.643
R2141 S.n4842 S.n4841 3.643
R2142 S.n4845 S.n4844 3.643
R2143 S.n4651 S.t414 3.643
R2144 S.n5412 S.t1031 3.643
R2145 S.n5133 S.t750 3.643
R2146 S.n5138 S.n5137 3.643
R2147 S.n5141 S.n5140 3.643
R2148 S.n5130 S.t1138 3.643
R2149 S.n4882 S.t311 3.643
R2150 S.n4889 S.n4888 3.643
R2151 S.n4886 S.n4885 3.643
R2152 S.n4879 S.t572 3.643
R2153 S.n5837 S.t784 3.643
R2154 S.n5842 S.n5841 3.643
R2155 S.n5845 S.n5844 3.643
R2156 S.n5834 S.t470 3.643
R2157 S.n5633 S.t693 3.643
R2158 S.n5637 S.n5636 3.643
R2159 S.n5640 S.n5639 3.643
R2160 S.n5630 S.t970 3.643
R2161 S.n4837 S.t767 3.643
R2162 S.n4834 S.n4833 3.643
R2163 S.n4831 S.n4830 3.643
R2164 S.n4659 S.t458 3.643
R2165 S.n4424 S.t266 3.643
R2166 S.n4808 S.t31 3.643
R2167 S.n4825 S.n4824 3.643
R2168 S.n4828 S.n4827 3.643
R2169 S.n4811 S.t617 3.643
R2170 S.n5864 S.t334 3.643
R2171 S.n5873 S.n5872 3.643
R2172 S.n5876 S.n5875 3.643
R2173 S.n5867 S.t924 3.643
R2174 S.n5421 S.t656 3.643
R2175 S.n5146 S.t368 3.643
R2176 S.n5154 S.n5153 3.643
R2177 S.n5157 S.n5156 3.643
R2178 S.n5149 S.t751 3.643
R2179 S.n4863 S.t1041 3.643
R2180 S.n4874 S.n4873 3.643
R2181 S.n4871 S.n4870 3.643
R2182 S.n4866 S.t178 3.643
R2183 S.n5649 S.t401 3.643
R2184 S.n5848 S.n5847 3.643
R2185 S.n5851 S.n5850 3.643
R2186 S.n5854 S.t70 3.643
R2187 S.n5348 S.t1055 3.643
R2188 S.n5169 S.t1038 3.643
R2189 S.n5177 S.n5176 3.643
R2190 S.n5180 S.n5179 3.643
R2191 S.n5172 S.t364 3.643
R2192 S.n4370 S.t482 3.643
R2193 S.n4374 S.n4373 3.643
R2194 S.n4363 S.t801 3.643
R2195 S.n4365 S.n4364 3.643
R2196 S.n91 S.n89 2.799
R2197 S.n979 S.n977 2.799
R2198 S.n1553 S.n1551 2.799
R2199 S.n2167 S.n2165 2.799
R2200 S.n2681 S.n2679 2.799
R2201 S.n3218 S.n3216 2.799
R2202 S.n3613 S.n3611 2.799
R2203 S.n4220 S.n4218 2.799
R2204 S.n4675 S.n4673 2.799
R2205 S.n5662 S.n5660 2.799
R2206 S.n5039 S.n5037 2.799
R2207 S.n506 S.n505 2.645
R2208 S.n85 S.n84 2.645
R2209 S.n973 S.n972 2.645
R2210 S.n1547 S.n1546 2.645
R2211 S.n2161 S.n2160 2.645
R2212 S.n2675 S.n2674 2.645
R2213 S.n3212 S.n3211 2.645
R2214 S.n3607 S.n3606 2.645
R2215 S.n4214 S.n4213 2.645
R2216 S.n4669 S.n4668 2.645
R2217 S.n5656 S.n5655 2.645
R2218 S.n4405 S.n4404 0.21
R2219 S.n5288 S.n5285 0.178
R2220 S.n369 S.n368 0.172
R2221 S.n508 S.n504 0.164
R2222 S.n5446 S.n5445 0.141
R2223 S.n1465 S.n1464 0.133
R2224 S.n496 S.n467 0.123
R2225 S.n673 S.n664 0.123
R2226 S.n530 S.n529 0.123
R2227 S.n5909 S.n1223 0.116
R2228 S.n5908 S.n1809 0.111
R2229 S.n5907 S.n2359 0.111
R2230 S.n5905 S.n3415 0.111
R2231 S.n5904 S.n3921 0.111
R2232 S.n5903 S.n4402 0.111
R2233 S.n5902 S.n4856 0.111
R2234 S.n5351 S.n5350 0.11
R2235 S.n5901 S.n5900 0.11
R2236 S.n5906 S.n2900 0.11
R2237 S.n5446 S.n5280 0.11
R2238 S.n4699 S.n4697 0.109
R2239 S.n4266 S.n4264 0.109
R2240 S.n3677 S.n3675 0.109
R2241 S.n3300 S.n3298 0.109
R2242 S.n2781 S.n2779 0.109
R2243 S.n2285 S.n2283 0.109
R2244 S.n1689 S.n1687 0.109
R2245 S.n272 S.n271 0.109
R2246 S.n1728 S.n1725 0.106
R2247 S.n2324 S.n2321 0.106
R2248 S.n2836 S.n2833 0.106
R2249 S.n3371 S.n3368 0.106
R2250 S.n3779 S.n3776 0.106
R2251 S.n4353 S.n4350 0.106
R2252 S.n5709 S.n5704 0.106
R2253 S.n1425 S.n1424 0.097
R2254 S.n1972 S.n1971 0.097
R2255 S.n2464 S.n2463 0.097
R2256 S.n3002 S.n3001 0.097
R2257 S.n3488 S.n3487 0.097
R2258 S.n3962 S.n3961 0.097
R2259 S.n4486 S.n4485 0.097
R2260 S.n881 S.n880 0.097
R2261 S.n909 S.n908 0.097
R2262 S.n5893 S.n5892 0.095
R2263 S.n5363 S.n5362 0.093
R2264 S.n5033 S.n5032 0.093
R2265 S.n5654 S.n5653 0.093
R2266 S.n5160 S.n5159 0.092
R2267 S.n5003 S.n5002 0.092
R2268 S S.n5910 0.09
R2269 S.n838 S.n837 0.087
R2270 S.n5344 S.n5343 0.087
R2271 S.n5361 S.n5360 0.085
R2272 S.n370 S.n367 0.082
R2273 S.n1217 S.n1214 0.082
R2274 S.n1253 S.n1250 0.082
R2275 S.n1839 S.n1836 0.082
R2276 S.n2879 S.n2877 0.082
R2277 S.n2930 S.n2927 0.082
R2278 S.n3445 S.n3442 0.082
R2279 S.n3951 S.n3948 0.082
R2280 S.n4422 S.n4419 0.082
R2281 S.n5457 S.n5454 0.082
R2282 S.n5278 S.n5274 0.082
R2283 S.n4481 S.n4480 0.08
R2284 S.n3957 S.n3956 0.08
R2285 S.n3483 S.n3482 0.08
R2286 S.n2997 S.n2996 0.08
R2287 S.n2459 S.n2458 0.08
R2288 S.n1967 S.n1966 0.08
R2289 S.n1420 S.n1419 0.08
R2290 S.n911 S.n910 0.08
R2291 S.n883 S.n882 0.08
R2292 S.n5444 S.n5443 0.079
R2293 S.n1236 S.n1235 0.079
R2294 S.n1822 S.n1821 0.079
R2295 S.n2893 S.n2892 0.079
R2296 S.n2913 S.n2912 0.079
R2297 S.n3428 S.n3427 0.079
R2298 S.n3934 S.n3933 0.079
R2299 S.n1102 S.n1101 0.077
R2300 S.n1659 S.n1658 0.077
R2301 S.n2255 S.n2254 0.077
R2302 S.n2751 S.n2750 0.077
R2303 S.n3270 S.n3269 0.077
R2304 S.n3647 S.n3646 0.077
R2305 S.n4236 S.n4235 0.077
R2306 S.n214 S.n213 0.077
R2307 S.n233 S.n232 0.077
R2308 S.n4680 S.n4679 0.076
R2309 S.n1239 S.n1238 0.075
R2310 S.n1825 S.n1824 0.075
R2311 S.n2896 S.n2895 0.075
R2312 S.n2916 S.n2915 0.075
R2313 S.n3431 S.n3430 0.075
R2314 S.n3937 S.n3936 0.075
R2315 S.n5044 S.n5043 0.074
R2316 S.n4225 S.n4224 0.074
R2317 S.n5667 S.n5666 0.074
R2318 S.n3618 S.n3617 0.074
R2319 S.n3223 S.n3222 0.074
R2320 S.n2686 S.n2685 0.074
R2321 S.n2172 S.n2171 0.074
R2322 S.n1558 S.n1557 0.074
R2323 S.n984 S.n983 0.074
R2324 S.n96 S.n95 0.074
R2325 S.n5367 S.n5366 0.073
R2326 S.n5375 S.n5374 0.073
R2327 S.n5383 S.n5382 0.073
R2328 S.n5391 S.n5390 0.073
R2329 S.n5399 S.n5398 0.073
R2330 S.n5407 S.n5406 0.073
R2331 S.n5415 S.n5414 0.073
R2332 S.n5420 S.n5419 0.073
R2333 S.n3964 S.n3963 0.071
R2334 S.n3490 S.n3489 0.071
R2335 S.n3004 S.n3003 0.071
R2336 S.n2466 S.n2465 0.071
R2337 S.n1974 S.n1973 0.071
R2338 S.n1427 S.n1426 0.071
R2339 S.n877 S.n876 0.071
R2340 S.n905 S.n904 0.071
R2341 S.n5707 S.n5706 0.07
R2342 S.t283 S.n5357 0.068
R2343 S.n641 S.n639 0.067
R2344 S.n641 S.n640 0.067
R2345 S.n563 S.n561 0.067
R2346 S.n563 S.n562 0.067
R2347 S.n605 S.n603 0.067
R2348 S.n605 S.n604 0.067
R2349 S.n635 S.n633 0.067
R2350 S.n635 S.n634 0.067
R2351 S.n399 S.n397 0.067
R2352 S.n399 S.n398 0.067
R2353 S.n550 S.n548 0.067
R2354 S.n550 S.n549 0.067
R2355 S.n430 S.n428 0.067
R2356 S.n430 S.n429 0.067
R2357 S.n538 S.n536 0.067
R2358 S.n538 S.n537 0.067
R2359 S.n461 S.n459 0.067
R2360 S.n461 S.n460 0.067
R2361 S.n525 S.n523 0.067
R2362 S.n525 S.n524 0.067
R2363 S.n465 S.n464 0.067
R2364 S.n465 S.n463 0.067
R2365 S.n370 S.n360 0.067
R2366 S.n370 S.n358 0.067
R2367 S.n1253 S.n1244 0.067
R2368 S.n1253 S.n1243 0.067
R2369 S.n1839 S.n1830 0.067
R2370 S.n1839 S.n1829 0.067
R2371 S.n2879 S.n2878 0.067
R2372 S.n2930 S.n2921 0.067
R2373 S.n2930 S.n2920 0.067
R2374 S.n3445 S.n3436 0.067
R2375 S.n3445 S.n3435 0.067
R2376 S.n3951 S.n3942 0.067
R2377 S.n3951 S.n3941 0.067
R2378 S.n4422 S.n4413 0.067
R2379 S.n4422 S.n4412 0.067
R2380 S.n5278 S.n5268 0.067
R2381 S.n5457 S.n5448 0.067
R2382 S.n5457 S.n5447 0.067
R2383 S.n5278 S.n5277 0.067
R2384 S.n2879 S.n2869 0.067
R2385 S.n518 S.n517 0.066
R2386 S.n600 S.n599 0.066
R2387 S.n371 S.n356 0.065
R2388 S.n636 S.n632 0.063
R2389 S.n5458 S.n5457 0.063
R2390 S.n636 S.n635 0.063
R2391 S.n935 S.n934 0.063
R2392 S.n1500 S.n1499 0.063
R2393 S.n1709 S.n1708 0.063
R2394 S.n2044 S.n2043 0.063
R2395 S.n2305 S.n2304 0.063
R2396 S.n2536 S.n2535 0.063
R2397 S.n2801 S.n2800 0.063
R2398 S.n3074 S.n3073 0.063
R2399 S.n3323 S.n3322 0.063
R2400 S.n3560 S.n3559 0.063
R2401 S.n3697 S.n3696 0.063
R2402 S.n4034 S.n4033 0.063
R2403 S.n4286 S.n4285 0.063
R2404 S.n4471 S.n4470 0.063
R2405 S.n4719 S.n4718 0.063
R2406 S.n5484 S.n5483 0.063
R2407 S.n5687 S.n5686 0.063
R2408 S.n348 S.n335 0.063
R2409 S.n254 S.n243 0.063
R2410 S.n851 S.n827 0.063
R2411 S.n1411 S.n1410 0.063
R2412 S.n1649 S.n1648 0.063
R2413 S.n1958 S.n1957 0.063
R2414 S.n2245 S.n2244 0.063
R2415 S.n2450 S.n2449 0.063
R2416 S.n2741 S.n2740 0.063
R2417 S.n2988 S.n2987 0.063
R2418 S.n3260 S.n3259 0.063
R2419 S.n3474 S.n3473 0.063
R2420 S.n3637 S.n3636 0.063
R2421 S.n913 S.n893 0.063
R2422 S.n1466 S.n1453 0.063
R2423 S.n2012 S.n2000 0.063
R2424 S.n2504 S.n2492 0.063
R2425 S.n3042 S.n3030 0.063
R2426 S.n3528 S.n3516 0.063
R2427 S.n4002 S.n3990 0.063
R2428 S.n4439 S.n4427 0.063
R2429 S.n327 S.n313 0.063
R2430 S.n2956 S.n2935 0.063
R2431 S.n2418 S.n2397 0.063
R2432 S.n1926 S.n1905 0.063
R2433 S.n1376 S.n1355 0.063
R2434 S.n817 S.n798 0.063
R2435 S.n394 S.n6 0.063
R2436 S.n789 S.n788 0.063
R2437 S.n1347 S.n1346 0.063
R2438 S.n1613 S.n1612 0.063
R2439 S.n1897 S.n1896 0.063
R2440 S.n2209 S.n2208 0.063
R2441 S.n2389 S.n2388 0.063
R2442 S.n2705 S.n2704 0.063
R2443 S.n1865 S.n1844 0.063
R2444 S.n1313 S.n1292 0.063
R2445 S.n759 S.n739 0.063
R2446 S.n425 S.n407 0.063
R2447 S.n730 S.n729 0.063
R2448 S.n1284 S.n1283 0.063
R2449 S.n1577 S.n1576 0.063
R2450 S.n700 S.n680 0.063
R2451 S.n456 S.n438 0.063
R2452 S.n494 S.n493 0.063
R2453 S.n642 S.n641 0.062
R2454 S.n551 S.n550 0.062
R2455 S.n539 S.n538 0.062
R2456 S.n526 S.n525 0.062
R2457 S.n616 S.n605 0.061
R2458 S.n400 S.n399 0.06
R2459 S.n431 S.n430 0.06
R2460 S.n462 S.n461 0.06
R2461 S.n466 S.n465 0.06
R2462 S.n5232 S.n5231 0.059
R2463 S.n5493 S.n5492 0.059
R2464 S.n1394 S.n1384 0.059
R2465 S.n564 S.n563 0.059
R2466 S.n5279 S.n5278 0.058
R2467 S.n1225 S.n1224 0.058
R2468 S.n1811 S.n1810 0.058
R2469 S.n2882 S.n2881 0.058
R2470 S.n2902 S.n2901 0.058
R2471 S.n3417 S.n3416 0.058
R2472 S.n3923 S.n3922 0.058
R2473 S.n371 S.n370 0.058
R2474 S.n498 S.n497 0.056
R2475 S.n2 S.n1 0.056
R2476 S.n403 S.n402 0.056
R2477 S.n434 S.n433 0.056
R2478 S.n4375 S.n4374 0.055
R2479 S.n521 S.n502 0.055
R2480 S.n5882 S.n5881 0.055
R2481 S.n383 S.n382 0.055
R2482 S.n1206 S.n1205 0.055
R2483 S.n1801 S.n1800 0.055
R2484 S.n2351 S.n2350 0.055
R2485 S.n2866 S.n2865 0.055
R2486 S.n3407 S.n3406 0.055
R2487 S.n3913 S.n3912 0.055
R2488 S.n4394 S.n4393 0.055
R2489 S.n4848 S.n4847 0.055
R2490 S.n5266 S.n4857 0.054
R2491 S.n98 S.n81 0.054
R2492 S.n5046 S.n5029 0.054
R2493 S.n3226 S.n3209 0.054
R2494 S.n3620 S.n3602 0.054
R2495 S.n4228 S.n4211 0.054
R2496 S.n4682 S.n4661 0.054
R2497 S.n5670 S.n5651 0.054
R2498 S.n2175 S.n2158 0.054
R2499 S.n2688 S.n2670 0.054
R2500 S.n987 S.n970 0.054
R2501 S.n1560 S.n1542 0.054
R2502 S.n5289 S.n5288 0.054
R2503 S.n5024 S.n5023 0.054
R2504 S.n5263 S.n5262 0.054
R2505 S.n5714 S.n5713 0.054
R2506 S.n484 S.n483 0.054
R2507 S.n351 S.n350 0.054
R2508 S.n938 S.n937 0.054
R2509 S.n5239 S.n5238 0.054
R2510 S.n5690 S.n5689 0.054
R2511 S.n5487 S.n5486 0.054
R2512 S.n4722 S.n4721 0.054
R2513 S.n4474 S.n4473 0.054
R2514 S.n4289 S.n4288 0.054
R2515 S.n4037 S.n4036 0.054
R2516 S.n3700 S.n3699 0.054
R2517 S.n3563 S.n3562 0.054
R2518 S.n3310 S.n3309 0.054
R2519 S.n3077 S.n3076 0.054
R2520 S.n2804 S.n2803 0.054
R2521 S.n2539 S.n2538 0.054
R2522 S.n2308 S.n2307 0.054
R2523 S.n2047 S.n2046 0.054
R2524 S.n1712 S.n1711 0.054
R2525 S.n1503 S.n1502 0.054
R2526 S.n1153 S.n1152 0.054
R2527 S.n257 S.n256 0.054
R2528 S.n73 S.n72 0.054
R2529 S.n792 S.n791 0.054
R2530 S.n3106 S.n3105 0.054
R2531 S.n2708 S.n2707 0.054
R2532 S.n2392 S.n2391 0.054
R2533 S.n2212 S.n2211 0.054
R2534 S.n1900 S.n1899 0.054
R2535 S.n1616 S.n1615 0.054
R2536 S.n1350 S.n1349 0.054
R2537 S.n1056 S.n1055 0.054
R2538 S.n389 S.n388 0.054
R2539 S.n3597 S.n3596 0.054
R2540 S.n3244 S.n3243 0.054
R2541 S.n2959 S.n2958 0.054
R2542 S.n2725 S.n2724 0.054
R2543 S.n2421 S.n2420 0.054
R2544 S.n2229 S.n2228 0.054
R2545 S.n1929 S.n1928 0.054
R2546 S.n1633 S.n1632 0.054
R2547 S.n1379 S.n1378 0.054
R2548 S.n1075 S.n1074 0.054
R2549 S.n1095 S.n1094 0.054
R2550 S.n854 S.n853 0.054
R2551 S.n285 S.n284 0.054
R2552 S.n308 S.n307 0.054
R2553 S.n1414 S.n1413 0.054
R2554 S.n1961 S.n1960 0.054
R2555 S.n2453 S.n2452 0.054
R2556 S.n2991 S.n2990 0.054
R2557 S.n3477 S.n3476 0.054
R2558 S.n4069 S.n4068 0.054
R2559 S.n3640 S.n3639 0.054
R2560 S.n3263 S.n3262 0.054
R2561 S.n2744 S.n2743 0.054
R2562 S.n2248 S.n2247 0.054
R2563 S.n1652 S.n1651 0.054
R2564 S.n888 S.n887 0.054
R2565 S.n218 S.n217 0.054
R2566 S.n590 S.n589 0.054
R2567 S.n4504 S.n4503 0.054
R2568 S.n4250 S.n4249 0.054
R2569 S.n3985 S.n3984 0.054
R2570 S.n3661 S.n3660 0.054
R2571 S.n3511 S.n3510 0.054
R2572 S.n3284 S.n3283 0.054
R2573 S.n3025 S.n3024 0.054
R2574 S.n2765 S.n2764 0.054
R2575 S.n2487 S.n2486 0.054
R2576 S.n2269 S.n2268 0.054
R2577 S.n1995 S.n1994 0.054
R2578 S.n1673 S.n1672 0.054
R2579 S.n1448 S.n1447 0.054
R2580 S.n1116 S.n1115 0.054
R2581 S.n916 S.n915 0.054
R2582 S.n237 S.n236 0.054
R2583 S.n1136 S.n1135 0.054
R2584 S.n1469 S.n1468 0.054
R2585 S.n1693 S.n1692 0.054
R2586 S.n2015 S.n2014 0.054
R2587 S.n2289 S.n2288 0.054
R2588 S.n2507 S.n2506 0.054
R2589 S.n2785 S.n2784 0.054
R2590 S.n3045 S.n3044 0.054
R2591 S.n3304 S.n3303 0.054
R2592 S.n3531 S.n3530 0.054
R2593 S.n3681 S.n3680 0.054
R2594 S.n4005 S.n4004 0.054
R2595 S.n4270 S.n4269 0.054
R2596 S.n4442 S.n4441 0.054
R2597 S.n4703 S.n4702 0.054
R2598 S.n5515 S.n5514 0.054
R2599 S.n330 S.n329 0.054
R2600 S.n820 S.n819 0.054
R2601 S.n198 S.n197 0.054
R2602 S.n181 S.n180 0.054
R2603 S.n52 S.n51 0.054
R2604 S.n733 S.n732 0.054
R2605 S.n2076 S.n2075 0.054
R2606 S.n1580 S.n1579 0.054
R2607 S.n1287 S.n1286 0.054
R2608 S.n1022 S.n1021 0.054
R2609 S.n420 S.n419 0.054
R2610 S.n2573 S.n2572 0.054
R2611 S.n2193 S.n2192 0.054
R2612 S.n1868 S.n1867 0.054
R2613 S.n1597 S.n1596 0.054
R2614 S.n1316 S.n1315 0.054
R2615 S.n1039 S.n1038 0.054
R2616 S.n762 S.n761 0.054
R2617 S.n165 S.n164 0.054
R2618 S.n148 S.n147 0.054
R2619 S.n31 S.n30 0.054
R2620 S.n965 S.n964 0.054
R2621 S.n451 S.n450 0.054
R2622 S.n1537 S.n1536 0.054
R2623 S.n1005 S.n1004 0.054
R2624 S.n703 S.n702 0.054
R2625 S.n132 S.n131 0.054
R2626 S.n115 S.n114 0.054
R2627 S.n279 S.n278 0.054
R2628 S.n1201 S.n1200 0.054
R2629 S.n1179 S.n1178 0.054
R2630 S.n1769 S.n1768 0.054
R2631 S.n1742 S.n1741 0.054
R2632 S.n2113 S.n2112 0.054
R2633 S.n2086 S.n2085 0.054
R2634 S.n2610 S.n2609 0.054
R2635 S.n2583 S.n2582 0.054
R2636 S.n3143 S.n3142 0.054
R2637 S.n3116 S.n3115 0.054
R2638 S.n3820 S.n3819 0.054
R2639 S.n3793 S.n3792 0.054
R2640 S.n4106 S.n4105 0.054
R2641 S.n4079 S.n4078 0.054
R2642 S.n4541 S.n4540 0.054
R2643 S.n4514 S.n4513 0.054
R2644 S.n5535 S.n5534 0.054
R2645 S.n5735 S.n5734 0.054
R2646 S.n5211 S.n5210 0.054
R2647 S.n5187 S.n5186 0.054
R2648 S.n1173 S.n1172 0.054
R2649 S.n1799 S.n1798 0.054
R2650 S.n4981 S.n4980 0.054
R2651 S.n4993 S.n4992 0.054
R2652 S.n5750 S.n5749 0.054
R2653 S.n5551 S.n5550 0.054
R2654 S.n4557 S.n4556 0.054
R2655 S.n4572 S.n4571 0.054
R2656 S.n4122 S.n4121 0.054
R2657 S.n4137 S.n4136 0.054
R2658 S.n3836 S.n3835 0.054
R2659 S.n3851 S.n3850 0.054
R2660 S.n3159 S.n3158 0.054
R2661 S.n3174 S.n3173 0.054
R2662 S.n2626 S.n2625 0.054
R2663 S.n2641 S.n2640 0.054
R2664 S.n2132 S.n2131 0.054
R2665 S.n2144 S.n2143 0.054
R2666 S.n1785 S.n1784 0.054
R2667 S.n1736 S.n1735 0.054
R2668 S.n2349 S.n2348 0.054
R2669 S.n5062 S.n5061 0.054
R2670 S.n4962 S.n4961 0.054
R2671 S.n5766 S.n5765 0.054
R2672 S.n5566 S.n5565 0.054
R2673 S.n4742 S.n4741 0.054
R2674 S.n4587 S.n4586 0.054
R2675 S.n4309 S.n4308 0.054
R2676 S.n4152 S.n4151 0.054
R2677 S.n3720 S.n3719 0.054
R2678 S.n3866 S.n3865 0.054
R2679 S.n3343 S.n3342 0.054
R2680 S.n3189 S.n3188 0.054
R2681 S.n2824 S.n2823 0.054
R2682 S.n2656 S.n2655 0.054
R2683 S.n2335 S.n2334 0.054
R2684 S.n2332 S.n2331 0.054
R2685 S.n2861 S.n2860 0.054
R2686 S.n5078 S.n5077 0.054
R2687 S.n4947 S.n4946 0.054
R2688 S.n5782 S.n5781 0.054
R2689 S.n5581 S.n5580 0.054
R2690 S.n4758 S.n4757 0.054
R2691 S.n4602 S.n4601 0.054
R2692 S.n4325 S.n4324 0.054
R2693 S.n4167 S.n4166 0.054
R2694 S.n3736 S.n3735 0.054
R2695 S.n3881 S.n3880 0.054
R2696 S.n3359 S.n3358 0.054
R2697 S.n3204 S.n3203 0.054
R2698 S.n2847 S.n2846 0.054
R2699 S.n4617 S.n4616 0.054
R2700 S.n5094 S.n5093 0.054
R2701 S.n4932 S.n4931 0.054
R2702 S.n5798 S.n5797 0.054
R2703 S.n5596 S.n5595 0.054
R2704 S.n4774 S.n4773 0.054
R2705 S.n4182 S.n4181 0.054
R2706 S.n3752 S.n3751 0.054
R2707 S.n3896 S.n3895 0.054
R2708 S.n3385 S.n3384 0.054
R2709 S.n3405 S.n3404 0.054
R2710 S.n2844 S.n2843 0.054
R2711 S.n3379 S.n3378 0.054
R2712 S.n3911 S.n3910 0.054
R2713 S.n5110 S.n5109 0.054
R2714 S.n4917 S.n4916 0.054
R2715 S.n5814 S.n5813 0.054
R2716 S.n5611 S.n5610 0.054
R2717 S.n4790 S.n4789 0.054
R2718 S.n4632 S.n4631 0.054
R2719 S.n4341 S.n4340 0.054
R2720 S.n4197 S.n4196 0.054
R2721 S.n3767 S.n3766 0.054
R2722 S.n3787 S.n3786 0.054
R2723 S.n4392 S.n4391 0.054
R2724 S.n5126 S.n5125 0.054
R2725 S.n4902 S.n4901 0.054
R2726 S.n5830 S.n5829 0.054
R2727 S.n5626 S.n5625 0.054
R2728 S.n4806 S.n4805 0.054
R2729 S.n4647 S.n4646 0.054
R2730 S.n4378 S.n4377 0.054
R2731 S.n4361 S.n4360 0.054
R2732 S.n4846 S.n4845 0.054
R2733 S.n5142 S.n5141 0.054
R2734 S.n4887 S.n4886 0.054
R2735 S.n5846 S.n5845 0.054
R2736 S.n5641 S.n5640 0.054
R2737 S.n4832 S.n4831 0.054
R2738 S.n4829 S.n4828 0.054
R2739 S.n5877 S.n5876 0.054
R2740 S.n5158 S.n5157 0.054
R2741 S.n4872 S.n4871 0.054
R2742 S.n5852 S.n5851 0.054
R2743 S.n5181 S.n5180 0.054
R2744 S.n5442 S.n5290 0.053
R2745 S.n94 S.n93 0.052
R2746 S.n982 S.n981 0.052
R2747 S.n1556 S.n1555 0.052
R2748 S.n2170 S.n2169 0.052
R2749 S.n2684 S.n2683 0.052
R2750 S.n3221 S.n3220 0.052
R2751 S.n3616 S.n3615 0.052
R2752 S.n4223 S.n4222 0.052
R2753 S.n4678 S.n4677 0.052
R2754 S.n5665 S.n5664 0.052
R2755 S.n5042 S.n5041 0.052
R2756 S.n677 S.n676 0.052
R2757 S.n1235 S.n1234 0.052
R2758 S.n1807 S.n1806 0.052
R2759 S.n1821 S.n1820 0.052
R2760 S.n2357 S.n2356 0.052
R2761 S.n2892 S.n2891 0.052
R2762 S.n2912 S.n2911 0.052
R2763 S.n3413 S.n3412 0.052
R2764 S.n3427 S.n3426 0.052
R2765 S.n3919 S.n3918 0.052
R2766 S.n3933 S.n3932 0.052
R2767 S.n4400 S.n4399 0.052
R2768 S.n4854 S.n4853 0.052
R2769 S.n5898 S.n5897 0.052
R2770 S.n5706 S.n5705 0.052
R2771 S.n2363 S.n2362 0.052
R2772 S.n292 S.n291 0.051
R2773 S.n4061 S.n4059 0.051
R2774 S.n3570 S.n3569 0.051
R2775 S.n3098 S.n3096 0.051
R2776 S.n2546 S.n2545 0.051
R2777 S.n2068 S.n2066 0.051
R2778 S.n1510 S.n1509 0.051
R2779 S.n957 S.n955 0.051
R2780 S.n470 S.n469 0.051
R2781 S.n5296 S.n5295 0.051
R2782 S.n5431 S.n5430 0.051
R2783 S.n360 S.n359 0.051
R2784 S.n358 S.n357 0.051
R2785 S.n5236 S.n5235 0.05
R2786 S.n4063 S.n4062 0.05
R2787 S.n5509 S.n5496 0.05
R2788 S.n321 S.n320 0.05
R2789 S.n3586 S.n3585 0.05
R2790 S.n3591 S.n3572 0.05
R2791 S.n3100 S.n3099 0.05
R2792 S.n2562 S.n2561 0.05
R2793 S.n2567 S.n2548 0.05
R2794 S.n2070 S.n2069 0.05
R2795 S.n1526 S.n1525 0.05
R2796 S.n1531 S.n1512 0.05
R2797 S.n959 S.n958 0.05
R2798 S.n494 S.n472 0.05
R2799 S.n338 S.n337 0.05
R2800 S.n1105 S.n1104 0.049
R2801 S.n1662 S.n1661 0.049
R2802 S.n2258 S.n2257 0.049
R2803 S.n2754 S.n2753 0.049
R2804 S.n3273 S.n3272 0.049
R2805 S.n3650 S.n3649 0.049
R2806 S.n4239 S.n4238 0.049
R2807 S.n212 S.n211 0.049
R2808 S.n231 S.n230 0.049
R2809 S.n4405 S.n4403 0.049
R2810 S.n4822 S.n4821 0.048
R2811 S.n1218 S.n1217 0.048
R2812 S.n1254 S.n1253 0.048
R2813 S.n1840 S.n1839 0.048
R2814 S.n2880 S.n2879 0.048
R2815 S.n2931 S.n2930 0.048
R2816 S.n3446 S.n3445 0.048
R2817 S.n3952 S.n3951 0.048
R2818 S.n4423 S.n4422 0.048
R2819 S.n4 S.n3 0.047
R2820 S.n405 S.n404 0.047
R2821 S.n436 S.n435 0.047
R2822 S.n5018 S.n5016 0.047
R2823 S.n5257 S.n5255 0.047
R2824 S.n5711 S.n5702 0.047
R2825 S.n5900 S.n5884 0.047
R2826 S.n494 S.n487 0.047
R2827 S.n348 S.n346 0.047
R2828 S.n935 S.n924 0.047
R2829 S.n5236 S.n5221 0.047
R2830 S.n5687 S.n5679 0.047
R2831 S.n5484 S.n5472 0.047
R2832 S.n4719 S.n4711 0.047
R2833 S.n4471 S.n4459 0.047
R2834 S.n4286 S.n4278 0.047
R2835 S.n4034 S.n4022 0.047
R2836 S.n3697 S.n3689 0.047
R2837 S.n3560 S.n3548 0.047
R2838 S.n3323 S.n3315 0.047
R2839 S.n3074 S.n3062 0.047
R2840 S.n2801 S.n2793 0.047
R2841 S.n2536 S.n2524 0.047
R2842 S.n2305 S.n2297 0.047
R2843 S.n2044 S.n2032 0.047
R2844 S.n1709 S.n1701 0.047
R2845 S.n1500 S.n1486 0.047
R2846 S.n1150 S.n1144 0.047
R2847 S.n254 S.n252 0.047
R2848 S.n70 S.n68 0.047
R2849 S.n789 S.n779 0.047
R2850 S.n3100 S.n3086 0.047
R2851 S.n2705 S.n2697 0.047
R2852 S.n2389 S.n2377 0.047
R2853 S.n2209 S.n2201 0.047
R2854 S.n1897 S.n1885 0.047
R2855 S.n1613 S.n1605 0.047
R2856 S.n1347 S.n1333 0.047
R2857 S.n1053 S.n1047 0.047
R2858 S.n394 S.n392 0.047
R2859 S.n3591 S.n3582 0.047
R2860 S.n3241 S.n3239 0.047
R2861 S.n2956 S.n2945 0.047
R2862 S.n2722 S.n2720 0.047
R2863 S.n2418 S.n2407 0.047
R2864 S.n2226 S.n2224 0.047
R2865 S.n1926 S.n1915 0.047
R2866 S.n1630 S.n1628 0.047
R2867 S.n1376 S.n1365 0.047
R2868 S.n1072 S.n1068 0.047
R2869 S.n1092 S.n1087 0.047
R2870 S.n851 S.n836 0.047
R2871 S.n290 S.n288 0.047
R2872 S.n305 S.n299 0.047
R2873 S.n1411 S.n1397 0.047
R2874 S.n1958 S.n1946 0.047
R2875 S.n2450 S.n2438 0.047
R2876 S.n2988 S.n2976 0.047
R2877 S.n3474 S.n3462 0.047
R2878 S.n4063 S.n4049 0.047
R2879 S.n3637 S.n3629 0.047
R2880 S.n3260 S.n3252 0.047
R2881 S.n2741 S.n2733 0.047
R2882 S.n2245 S.n2237 0.047
R2883 S.n1649 S.n1641 0.047
R2884 S.n885 S.n875 0.047
R2885 S.n215 S.n209 0.047
R2886 S.n600 S.n593 0.047
R2887 S.n4498 S.n4490 0.047
R2888 S.n4247 S.n4242 0.047
R2889 S.n3982 S.n3967 0.047
R2890 S.n3658 S.n3653 0.047
R2891 S.n3508 S.n3493 0.047
R2892 S.n3281 S.n3276 0.047
R2893 S.n3022 S.n3007 0.047
R2894 S.n2762 S.n2757 0.047
R2895 S.n2484 S.n2469 0.047
R2896 S.n2266 S.n2261 0.047
R2897 S.n1992 S.n1977 0.047
R2898 S.n1670 S.n1665 0.047
R2899 S.n1445 S.n1430 0.047
R2900 S.n1113 S.n1108 0.047
R2901 S.n913 S.n903 0.047
R2902 S.n234 S.n229 0.047
R2903 S.n1133 S.n1127 0.047
R2904 S.n1466 S.n1463 0.047
R2905 S.n1690 S.n1685 0.047
R2906 S.n2012 S.n2010 0.047
R2907 S.n2286 S.n2281 0.047
R2908 S.n2504 S.n2502 0.047
R2909 S.n2782 S.n2777 0.047
R2910 S.n3042 S.n3040 0.047
R2911 S.n3301 S.n3296 0.047
R2912 S.n3528 S.n3526 0.047
R2913 S.n3678 S.n3673 0.047
R2914 S.n4002 S.n4000 0.047
R2915 S.n4267 S.n4262 0.047
R2916 S.n4439 S.n4437 0.047
R2917 S.n4700 S.n4695 0.047
R2918 S.n5509 S.n5507 0.047
R2919 S.n327 S.n319 0.047
R2920 S.n817 S.n807 0.047
R2921 S.n195 S.n193 0.047
R2922 S.n178 S.n176 0.047
R2923 S.n49 S.n47 0.047
R2924 S.n730 S.n720 0.047
R2925 S.n2070 S.n2056 0.047
R2926 S.n1577 S.n1569 0.047
R2927 S.n1284 S.n1270 0.047
R2928 S.n1019 S.n1013 0.047
R2929 S.n425 S.n423 0.047
R2930 S.n2567 S.n2558 0.047
R2931 S.n2190 S.n2188 0.047
R2932 S.n1865 S.n1854 0.047
R2933 S.n1594 S.n1592 0.047
R2934 S.n1313 S.n1302 0.047
R2935 S.n1036 S.n1034 0.047
R2936 S.n759 S.n748 0.047
R2937 S.n162 S.n160 0.047
R2938 S.n145 S.n143 0.047
R2939 S.n28 S.n26 0.047
R2940 S.n959 S.n947 0.047
R2941 S.n456 S.n454 0.047
R2942 S.n1531 S.n1522 0.047
R2943 S.n1002 S.n1000 0.047
R2944 S.n700 S.n689 0.047
R2945 S.n129 S.n127 0.047
R2946 S.n112 S.n110 0.047
R2947 S.n378 S.n373 0.047
R2948 S.n273 S.n269 0.047
R2949 S.n1195 S.n1193 0.047
R2950 S.n1186 S.n1182 0.047
R2951 S.n1763 S.n1757 0.047
R2952 S.n1749 S.n1745 0.047
R2953 S.n2107 S.n2101 0.047
R2954 S.n2093 S.n2089 0.047
R2955 S.n2604 S.n2598 0.047
R2956 S.n2590 S.n2586 0.047
R2957 S.n3137 S.n3131 0.047
R2958 S.n3123 S.n3119 0.047
R2959 S.n3814 S.n3808 0.047
R2960 S.n3800 S.n3796 0.047
R2961 S.n4100 S.n4094 0.047
R2962 S.n4086 S.n4082 0.047
R2963 S.n4535 S.n4529 0.047
R2964 S.n4521 S.n4517 0.047
R2965 S.n5529 S.n5523 0.047
R2966 S.n5729 S.n5725 0.047
R2967 S.n5208 S.n5202 0.047
R2968 S.n5194 S.n5190 0.047
R2969 S.n1222 S.n1208 0.047
R2970 S.n1167 S.n1165 0.047
R2971 S.n1793 S.n1774 0.047
R2972 S.n4988 S.n4978 0.047
R2973 S.n4990 S.n4970 0.047
R2974 S.n5744 S.n5740 0.047
R2975 S.n5545 S.n5540 0.047
R2976 S.n4564 S.n4554 0.047
R2977 S.n4566 S.n4546 0.047
R2978 S.n4129 S.n4119 0.047
R2979 S.n4131 S.n4111 0.047
R2980 S.n3843 S.n3833 0.047
R2981 S.n3845 S.n3825 0.047
R2982 S.n3166 S.n3156 0.047
R2983 S.n3168 S.n3148 0.047
R2984 S.n2633 S.n2623 0.047
R2985 S.n2635 S.n2615 0.047
R2986 S.n2139 S.n2129 0.047
R2987 S.n2141 S.n2118 0.047
R2988 S.n1792 S.n1782 0.047
R2989 S.n1809 S.n1256 0.047
R2990 S.n1730 S.n1724 0.047
R2991 S.n2343 S.n2149 0.047
R2992 S.n5056 S.n5051 0.047
R2993 S.n4959 S.n4955 0.047
R2994 S.n5760 S.n5755 0.047
R2995 S.n5560 S.n5556 0.047
R2996 S.n4736 S.n4731 0.047
R2997 S.n4581 S.n4577 0.047
R2998 S.n4303 S.n4298 0.047
R2999 S.n4146 S.n4142 0.047
R3000 S.n3714 S.n3709 0.047
R3001 S.n3860 S.n3856 0.047
R3002 S.n3337 S.n3332 0.047
R3003 S.n3183 S.n3179 0.047
R3004 S.n2818 S.n2813 0.047
R3005 S.n2650 S.n2646 0.047
R3006 S.n2342 S.n2157 0.047
R3007 S.n2359 S.n1842 0.047
R3008 S.n2326 S.n2320 0.047
R3009 S.n2855 S.n2661 0.047
R3010 S.n5072 S.n5067 0.047
R3011 S.n4944 S.n4940 0.047
R3012 S.n5776 S.n5771 0.047
R3013 S.n5575 S.n5571 0.047
R3014 S.n4752 S.n4747 0.047
R3015 S.n4596 S.n4592 0.047
R3016 S.n4319 S.n4314 0.047
R3017 S.n4161 S.n4157 0.047
R3018 S.n3730 S.n3725 0.047
R3019 S.n3875 S.n3871 0.047
R3020 S.n3353 S.n3348 0.047
R3021 S.n3198 S.n3194 0.047
R3022 S.n2854 S.n2669 0.047
R3023 S.n4611 S.n4607 0.047
R3024 S.n5088 S.n5083 0.047
R3025 S.n4929 S.n4925 0.047
R3026 S.n5792 S.n5787 0.047
R3027 S.n5590 S.n5586 0.047
R3028 S.n4768 S.n4763 0.047
R3029 S.n4176 S.n4174 0.047
R3030 S.n3746 S.n3744 0.047
R3031 S.n3890 S.n3888 0.047
R3032 S.n3390 S.n3388 0.047
R3033 S.n3399 S.n3397 0.047
R3034 S.n2838 S.n2832 0.047
R3035 S.n2900 S.n2868 0.047
R3036 S.n3415 S.n2933 0.047
R3037 S.n3373 S.n3367 0.047
R3038 S.n3905 S.n3901 0.047
R3039 S.n5104 S.n5099 0.047
R3040 S.n4914 S.n4910 0.047
R3041 S.n5808 S.n5803 0.047
R3042 S.n5605 S.n5601 0.047
R3043 S.n4784 S.n4779 0.047
R3044 S.n4626 S.n4622 0.047
R3045 S.n4335 S.n4330 0.047
R3046 S.n4191 S.n4187 0.047
R3047 S.n3761 S.n3757 0.047
R3048 S.n3921 S.n3448 0.047
R3049 S.n3781 S.n3775 0.047
R3050 S.n4386 S.n4202 0.047
R3051 S.n5120 S.n5115 0.047
R3052 S.n4899 S.n4895 0.047
R3053 S.n5824 S.n5819 0.047
R3054 S.n5620 S.n5616 0.047
R3055 S.n4800 S.n4795 0.047
R3056 S.n4641 S.n4637 0.047
R3057 S.n4385 S.n4210 0.047
R3058 S.n4402 S.n3954 0.047
R3059 S.n4355 S.n4349 0.047
R3060 S.n4840 S.n4652 0.047
R3061 S.n5136 S.n5131 0.047
R3062 S.n4884 S.n4880 0.047
R3063 S.n5840 S.n5835 0.047
R3064 S.n5635 S.n5631 0.047
R3065 S.n4839 S.n4660 0.047
R3066 S.n4856 S.n4425 0.047
R3067 S.n4823 S.n4812 0.047
R3068 S.n5871 S.n5868 0.047
R3069 S.n5152 S.n5150 0.047
R3070 S.n4869 S.n4867 0.047
R3071 S.n5857 S.n5855 0.047
R3072 S.n5175 S.n5173 0.047
R3073 S.n4372 S.n4371 0.047
R3074 S.n849 S.n844 0.047
R3075 S.n3458 S.n3457 0.047
R3076 S.n2972 S.n2971 0.047
R3077 S.n2434 S.n2433 0.047
R3078 S.n1942 S.n1941 0.047
R3079 S.n1393 S.n1392 0.047
R3080 S.n624 S.n623 0.046
R3081 S.t241 S.n565 0.046
R3082 S.t241 S.n555 0.046
R3083 S.t241 S.n543 0.046
R3084 S.t241 S.n531 0.046
R3085 S.n1195 S.n1186 0.046
R3086 S.n1793 S.n1792 0.046
R3087 S.n2343 S.n2342 0.045
R3088 S.n2855 S.n2854 0.045
R3089 S.n4386 S.n4385 0.045
R3090 S.n4840 S.n4839 0.045
R3091 S.n3399 S.n3390 0.045
R3092 S.n572 S.n570 0.045
R3093 S.n5870 S.n5869 0.045
R3094 S.n5427 S.n5426 0.045
R3095 S.n5429 S.n5428 0.045
R3096 S.n580 S.n579 0.045
R3097 S.n866 S.n858 0.045
R3098 S.n1442 S.n1434 0.045
R3099 S.n1989 S.n1981 0.045
R3100 S.n2481 S.n2473 0.045
R3101 S.n3019 S.n3011 0.045
R3102 S.n3505 S.n3497 0.045
R3103 S.n3979 S.n3971 0.045
R3104 S.n1227 S.n1226 0.045
R3105 S.n1813 S.n1812 0.045
R3106 S.n2884 S.n2883 0.045
R3107 S.n2904 S.n2903 0.045
R3108 S.n3419 S.n3418 0.045
R3109 S.n3925 S.n3924 0.045
R3110 S.n5294 S.n5293 0.045
R3111 S.n5871 S.n5857 0.044
R3112 S.n616 S.n615 0.044
R3113 S.n1763 S.n1750 0.044
R3114 S.n2107 S.n2094 0.044
R3115 S.n2604 S.n2591 0.044
R3116 S.n3137 S.n3124 0.044
R3117 S.n3814 S.n3801 0.044
R3118 S.n4100 S.n4087 0.044
R3119 S.n4535 S.n4522 0.044
R3120 S.n5529 S.n5516 0.044
R3121 S.n5208 S.n5195 0.044
R3122 S.n2141 S.n2140 0.044
R3123 S.n2635 S.n2634 0.044
R3124 S.n3168 S.n3167 0.044
R3125 S.n3845 S.n3844 0.044
R3126 S.n4131 S.n4130 0.044
R3127 S.n4566 S.n4565 0.044
R3128 S.n5545 S.n5544 0.044
R3129 S.n4990 S.n4989 0.044
R3130 S.n5351 S.n5349 0.044
R3131 S.n9 S.n8 0.044
R3132 S.n410 S.n409 0.044
R3133 S.n441 S.n440 0.044
R3134 S.n5235 S.n5234 0.043
R3135 S.n5496 S.n5495 0.043
R3136 S.n628 S.n627 0.043
R3137 S.n800 S.n799 0.042
R3138 S.n1357 S.n1356 0.042
R3139 S.n1907 S.n1906 0.042
R3140 S.n2399 S.n2398 0.042
R3141 S.n2937 S.n2936 0.042
R3142 S.n741 S.n740 0.042
R3143 S.n1294 S.n1293 0.042
R3144 S.n1846 S.n1845 0.042
R3145 S.n682 S.n681 0.042
R3146 S.n5480 S.n5477 0.042
R3147 S.n4467 S.n4464 0.042
R3148 S.n4030 S.n4027 0.042
R3149 S.n3556 S.n3553 0.042
R3150 S.n3070 S.n3067 0.042
R3151 S.n2532 S.n2529 0.042
R3152 S.n2040 S.n2037 0.042
R3153 S.n1496 S.n1491 0.042
R3154 S.n931 S.n929 0.042
R3155 S.n245 S.n244 0.042
R3156 S.n2385 S.n2382 0.042
R3157 S.n1893 S.n1890 0.042
R3158 S.n1343 S.n1338 0.042
R3159 S.n3470 S.n3467 0.042
R3160 S.n2984 S.n2981 0.042
R3161 S.n2446 S.n2443 0.042
R3162 S.n1954 S.n1951 0.042
R3163 S.n1407 S.n1402 0.042
R3164 S.n1280 S.n1275 0.042
R3165 S.n496 S.n495 0.042
R3166 S.n396 S.n395 0.042
R3167 S.n602 S.n601 0.042
R3168 S.n427 S.n426 0.042
R3169 S.n458 S.n457 0.042
R3170 S.n4429 S.n4428 0.042
R3171 S.n3992 S.n3991 0.042
R3172 S.n3518 S.n3517 0.042
R3173 S.n3032 S.n3031 0.042
R3174 S.n2494 S.n2493 0.042
R3175 S.n2002 S.n2001 0.042
R3176 S.n1455 S.n1454 0.042
R3177 S.n895 S.n894 0.042
R3178 S.n5035 S.n5034 0.042
R3179 S.n632 S.n631 0.041
R3180 S.n4046 S.n4045 0.041
R3181 S.n500 S.n499 0.041
R3182 S.n375 S.n374 0.041
R3183 S.n519 S.n508 0.04
R3184 S.n490 S.n489 0.04
R3185 S.n94 S.n85 0.04
R3186 S.n982 S.n973 0.04
R3187 S.n1556 S.n1547 0.04
R3188 S.n2170 S.n2161 0.04
R3189 S.n2684 S.n2675 0.04
R3190 S.n3221 S.n3212 0.04
R3191 S.n3616 S.n3607 0.04
R3192 S.n4223 S.n4214 0.04
R3193 S.n4678 S.n4669 0.04
R3194 S.n5665 S.n5656 0.04
R3195 S.n5318 S.n5317 0.04
R3196 S.n5316 S.n5315 0.04
R3197 S.n5314 S.n5313 0.04
R3198 S.n5312 S.n5311 0.04
R3199 S.n5310 S.n5309 0.04
R3200 S.n5308 S.n5307 0.04
R3201 S.n5306 S.n5305 0.04
R3202 S.n5304 S.n5303 0.04
R3203 S.n5374 S.n5373 0.039
R3204 S.n5382 S.n5381 0.039
R3205 S.n5390 S.n5389 0.039
R3206 S.n5398 S.n5397 0.039
R3207 S.n5406 S.n5405 0.039
R3208 S.n5414 S.n5413 0.039
R3209 S.n5419 S.n5418 0.039
R3210 S.n507 S.n506 0.039
R3211 S.n5889 S.n5888 0.039
R3212 S.n1228 S.n1227 0.039
R3213 S.n1233 S.n1232 0.039
R3214 S.n1814 S.n1813 0.039
R3215 S.n1819 S.n1818 0.039
R3216 S.n2885 S.n2884 0.039
R3217 S.n2890 S.n2889 0.039
R3218 S.n2905 S.n2904 0.039
R3219 S.n2910 S.n2909 0.039
R3220 S.n3420 S.n3419 0.039
R3221 S.n3425 S.n3424 0.039
R3222 S.n3926 S.n3925 0.039
R3223 S.n3931 S.n3930 0.039
R3224 S.n5298 S.n5297 0.039
R3225 S.n5433 S.n5432 0.039
R3226 S.n93 S.n86 0.039
R3227 S.n981 S.n974 0.039
R3228 S.n1555 S.n1548 0.039
R3229 S.n2169 S.n2162 0.039
R3230 S.n2683 S.n2676 0.039
R3231 S.n3220 S.n3213 0.039
R3232 S.n3615 S.n3608 0.039
R3233 S.n4222 S.n4215 0.039
R3234 S.n4677 S.n4670 0.039
R3235 S.n5664 S.n5657 0.039
R3236 S.n5033 S.n5031 0.038
R3237 S.n5654 S.n5652 0.038
R3238 S.n5468 S.n5467 0.038
R3239 S.n4455 S.n4454 0.038
R3240 S.n4018 S.n4017 0.038
R3241 S.n3544 S.n3543 0.038
R3242 S.n3058 S.n3057 0.038
R3243 S.n2520 S.n2519 0.038
R3244 S.n2028 S.n2027 0.038
R3245 S.n1482 S.n1481 0.038
R3246 S.n2373 S.n2372 0.038
R3247 S.n1881 S.n1880 0.038
R3248 S.n1329 S.n1328 0.038
R3249 S.n775 S.n774 0.038
R3250 S.n2954 S.n2949 0.038
R3251 S.n2416 S.n2411 0.038
R3252 S.n1924 S.n1919 0.038
R3253 S.n1374 S.n1369 0.038
R3254 S.n815 S.n811 0.038
R3255 S.n1266 S.n1265 0.038
R3256 S.n716 S.n715 0.038
R3257 S.n1863 S.n1858 0.038
R3258 S.n1311 S.n1306 0.038
R3259 S.n757 S.n752 0.038
R3260 S.n698 S.n693 0.038
R3261 S.n4497 S.n4495 0.037
R3262 S.n5889 S.n5886 0.037
R3263 S.n5888 S.n5887 0.037
R3264 S.n1445 S.n1427 0.037
R3265 S.n1992 S.n1974 0.037
R3266 S.n2484 S.n2466 0.037
R3267 S.n3022 S.n3004 0.037
R3268 S.n3508 S.n3490 0.037
R3269 S.n3982 S.n3964 0.037
R3270 S.n4498 S.n4487 0.037
R3271 S.n913 S.n905 0.037
R3272 S.n885 S.n877 0.037
R3273 S.n1233 S.n1230 0.037
R3274 S.n1232 S.n1231 0.037
R3275 S.n1819 S.n1816 0.037
R3276 S.n1818 S.n1817 0.037
R3277 S.n2890 S.n2887 0.037
R3278 S.n2889 S.n2888 0.037
R3279 S.n2910 S.n2907 0.037
R3280 S.n2909 S.n2908 0.037
R3281 S.n3425 S.n3422 0.037
R3282 S.n3424 S.n3423 0.037
R3283 S.n3931 S.n3928 0.037
R3284 S.n3930 S.n3929 0.037
R3285 S.n4860 S.n4859 0.037
R3286 S.n5861 S.n5860 0.037
R3287 S.n378 S.n375 0.036
R3288 S.n1132 S.n1131 0.036
R3289 S.n1678 S.n1677 0.036
R3290 S.n2274 S.n2273 0.036
R3291 S.n2770 S.n2769 0.036
R3292 S.n3289 S.n3288 0.036
R3293 S.n3666 S.n3665 0.036
R3294 S.n4255 S.n4254 0.036
R3295 S.n4688 S.n4687 0.036
R3296 S.n92 S.n87 0.036
R3297 S.n980 S.n975 0.036
R3298 S.n1554 S.n1549 0.036
R3299 S.n2168 S.n2163 0.036
R3300 S.n2682 S.n2677 0.036
R3301 S.n3219 S.n3214 0.036
R3302 S.n3614 S.n3609 0.036
R3303 S.n4221 S.n4216 0.036
R3304 S.n4676 S.n4671 0.036
R3305 S.n5663 S.n5658 0.036
R3306 S.n5284 S.n5281 0.036
R3307 S.n3232 S.n3231 0.035
R3308 S.n2713 S.n2712 0.035
R3309 S.n2217 S.n2216 0.035
R3310 S.n1621 S.n1620 0.035
R3311 S.n1061 S.n1060 0.035
R3312 S.n2181 S.n2180 0.035
R3313 S.n1585 S.n1584 0.035
R3314 S.n1027 S.n1026 0.035
R3315 S.n993 S.n992 0.035
R3316 S.n5248 S.n5247 0.035
R3317 S.n5216 S.n5215 0.035
R3318 S.n102 S.n101 0.035
R3319 S.n5026 S.n5025 0.035
R3320 S.n3230 S.n3229 0.035
R3321 S.n3624 S.n3623 0.035
R3322 S.n4232 S.n4231 0.035
R3323 S.n4686 S.n4685 0.035
R3324 S.n5674 S.n5673 0.035
R3325 S.n2179 S.n2178 0.035
R3326 S.n2692 S.n2691 0.035
R3327 S.n991 S.n990 0.035
R3328 S.n1564 S.n1563 0.035
R3329 S.n5890 S.n5889 0.035
R3330 S.n5468 S.n5463 0.035
R3331 S.n4455 S.n4450 0.035
R3332 S.n4018 S.n4013 0.035
R3333 S.n3544 S.n3539 0.035
R3334 S.n3058 S.n3053 0.035
R3335 S.n2520 S.n2515 0.035
R3336 S.n2028 S.n2023 0.035
R3337 S.n1482 S.n1477 0.035
R3338 S.n2373 S.n2368 0.035
R3339 S.n1881 S.n1876 0.035
R3340 S.n1329 S.n1324 0.035
R3341 S.n775 S.n770 0.035
R3342 S.n4063 S.n4046 0.035
R3343 S.n815 S.n814 0.035
R3344 S.n1374 S.n1373 0.035
R3345 S.n1924 S.n1923 0.035
R3346 S.n2416 S.n2415 0.035
R3347 S.n2954 S.n2953 0.035
R3348 S.n1266 S.n1261 0.035
R3349 S.n716 S.n711 0.035
R3350 S.n757 S.n756 0.035
R3351 S.n1311 S.n1310 0.035
R3352 S.n1863 S.n1862 0.035
R3353 S.n698 S.n697 0.035
R3354 S.n1226 S.n1225 0.035
R3355 S.n1236 S.n1233 0.035
R3356 S.n1812 S.n1811 0.035
R3357 S.n1822 S.n1819 0.035
R3358 S.n2883 S.n2882 0.035
R3359 S.n2893 S.n2890 0.035
R3360 S.n2903 S.n2902 0.035
R3361 S.n2913 S.n2910 0.035
R3362 S.n3418 S.n3417 0.035
R3363 S.n3428 S.n3425 0.035
R3364 S.n3924 S.n3923 0.035
R3365 S.n3934 S.n3931 0.035
R3366 S.t283 S.n5439 0.035
R3367 S.t241 S.n648 0.035
R3368 S.t241 S.n644 0.035
R3369 S.t241 S.n553 0.035
R3370 S.t241 S.n660 0.035
R3371 S.t241 S.n567 0.035
R3372 S.t241 S.n578 0.035
R3373 S.t241 S.n626 0.035
R3374 S.t241 S.n541 0.035
R3375 S.t241 S.n656 0.035
R3376 S.t241 S.n528 0.035
R3377 S.t241 S.n652 0.035
R3378 S.t283 S.n5353 0.035
R3379 S.t283 S.n5364 0.035
R3380 S.t283 S.n5371 0.035
R3381 S.t283 S.n5379 0.035
R3382 S.t283 S.n5387 0.035
R3383 S.t283 S.n5395 0.035
R3384 S.t283 S.n5403 0.035
R3385 S.t283 S.n5411 0.035
R3386 S.t283 S.n5422 0.035
R3387 S.t283 S.n5345 0.035
R3388 S.n5356 S.n5355 0.035
R3389 S.n4410 S.n4409 0.034
R3390 S.n564 S.n560 0.034
R3391 S.n557 S.n556 0.034
R3392 S.n545 S.n544 0.034
R3393 S.n533 S.n532 0.034
R3394 S.n5194 S.n5191 0.034
R3395 S.n5208 S.n5204 0.034
R3396 S.n5729 S.n5726 0.034
R3397 S.n5529 S.n5525 0.034
R3398 S.n4521 S.n4518 0.034
R3399 S.n4535 S.n4531 0.034
R3400 S.n4086 S.n4083 0.034
R3401 S.n4100 S.n4096 0.034
R3402 S.n3800 S.n3797 0.034
R3403 S.n3814 S.n3810 0.034
R3404 S.n3123 S.n3120 0.034
R3405 S.n3137 S.n3133 0.034
R3406 S.n2590 S.n2587 0.034
R3407 S.n2604 S.n2600 0.034
R3408 S.n2093 S.n2090 0.034
R3409 S.n2107 S.n2103 0.034
R3410 S.n1749 S.n1746 0.034
R3411 S.n1763 S.n1759 0.034
R3412 S.n1186 S.n1183 0.034
R3413 S.n1222 S.n674 0.034
R3414 S.n1809 S.n1808 0.034
R3415 S.n2359 S.n2358 0.034
R3416 S.n3415 S.n3414 0.034
R3417 S.n3921 S.n3920 0.034
R3418 S.n4402 S.n4401 0.034
R3419 S.n4856 S.n4855 0.034
R3420 S.n5900 S.n5899 0.034
R3421 S.n2900 S.n2360 0.034
R3422 S.n4225 S.n4212 0.034
R3423 S.n3618 S.n3605 0.034
R3424 S.n3223 S.n3210 0.034
R3425 S.n2686 S.n2673 0.034
R3426 S.n2172 S.n2159 0.034
R3427 S.n1558 S.n1545 0.034
R3428 S.n984 S.n971 0.034
R3429 S.n96 S.n83 0.034
R3430 S.t283 S.n5438 0.034
R3431 S.t241 S.n651 0.034
R3432 S.t241 S.n643 0.034
R3433 S.t241 S.n552 0.034
R3434 S.t241 S.n663 0.034
R3435 S.t241 S.n566 0.034
R3436 S.t241 S.n577 0.034
R3437 S.t241 S.n625 0.034
R3438 S.t241 S.n540 0.034
R3439 S.t241 S.n659 0.034
R3440 S.t241 S.n527 0.034
R3441 S.t241 S.n655 0.034
R3442 S.t283 S.n5352 0.034
R3443 S.t283 S.n5365 0.034
R3444 S.t283 S.n5372 0.034
R3445 S.t283 S.n5380 0.034
R3446 S.t283 S.n5388 0.034
R3447 S.t283 S.n5396 0.034
R3448 S.t283 S.n5404 0.034
R3449 S.t283 S.n5412 0.034
R3450 S.t283 S.n5421 0.034
R3451 S.t283 S.n5348 0.034
R3452 S.n519 S.n518 0.033
R3453 S.n1091 S.n1090 0.033
R3454 S.n5044 S.n5033 0.032
R3455 S.n5667 S.n5654 0.032
R3456 S.n4663 S.n4662 0.032
R3457 S.n952 S.n951 0.031
R3458 S.t35 S.n5216 0.031
R3459 S.t255 S.n102 0.031
R3460 S.t64 S.n5026 0.031
R3461 S.t12 S.n3230 0.031
R3462 S.t10 S.n3624 0.031
R3463 S.t57 S.n4232 0.031
R3464 S.t8 S.n4686 0.031
R3465 S.t4 S.n5674 0.031
R3466 S.t16 S.n2179 0.031
R3467 S.t0 S.n2692 0.031
R3468 S.t6 S.n991 0.031
R3469 S.t21 S.n1564 0.031
R3470 S.n5463 S.n5462 0.031
R3471 S.n4450 S.n4449 0.031
R3472 S.n4013 S.n4012 0.031
R3473 S.n3539 S.n3538 0.031
R3474 S.n3053 S.n3052 0.031
R3475 S.n2515 S.n2514 0.031
R3476 S.n2023 S.n2022 0.031
R3477 S.n1477 S.n1476 0.031
R3478 S.n2368 S.n2367 0.031
R3479 S.n1876 S.n1875 0.031
R3480 S.n1324 S.n1323 0.031
R3481 S.n770 S.n769 0.031
R3482 S.n814 S.n813 0.031
R3483 S.n1373 S.n1372 0.031
R3484 S.n1923 S.n1922 0.031
R3485 S.n2415 S.n2414 0.031
R3486 S.n2953 S.n2952 0.031
R3487 S.n1261 S.n1260 0.031
R3488 S.n711 S.n710 0.031
R3489 S.n756 S.n755 0.031
R3490 S.n1310 S.n1309 0.031
R3491 S.n1862 S.n1861 0.031
R3492 S.n697 S.n696 0.031
R3493 S.n666 S.n665 0.031
R3494 S.n667 S.n666 0.031
R3495 S.n668 S.n667 0.031
R3496 S.n669 S.n668 0.031
R3497 S.n670 S.n669 0.031
R3498 S.n671 S.n670 0.031
R3499 S.n672 S.n671 0.031
R3500 S.n673 S.n672 0.031
R3501 S.n377 S.n376 0.031
R3502 S.n5910 S.n5909 0.031
R3503 S.n5909 S.n5908 0.031
R3504 S.n5908 S.n5907 0.031
R3505 S.n5907 S.n5906 0.031
R3506 S.n5906 S.n5905 0.031
R3507 S.n5905 S.n5904 0.031
R3508 S.n5904 S.n5903 0.031
R3509 S.n5903 S.n5902 0.031
R3510 S.n5902 S.n5901 0.031
R3511 S.n5901 S.n5446 0.031
R3512 S.n5206 S.n5205 0.031
R3513 S.n5527 S.n5526 0.031
R3514 S.n4533 S.n4532 0.031
R3515 S.n4098 S.n4097 0.031
R3516 S.n3812 S.n3811 0.031
R3517 S.n3135 S.n3134 0.031
R3518 S.n2602 S.n2601 0.031
R3519 S.n2105 S.n2104 0.031
R3520 S.n1761 S.n1760 0.031
R3521 S.n3589 S.n3588 0.031
R3522 S.n2565 S.n2564 0.031
R3523 S.n1529 S.n1528 0.031
R3524 S.n3574 S.n3573 0.03
R3525 S.n2550 S.n2549 0.03
R3526 S.n1514 S.n1513 0.03
R3527 S.n3976 S.n3975 0.03
R3528 S.n3502 S.n3501 0.03
R3529 S.n3016 S.n3015 0.03
R3530 S.n2478 S.n2477 0.03
R3531 S.n1986 S.n1985 0.03
R3532 S.n1439 S.n1438 0.03
R3533 S.n863 S.n862 0.03
R3534 S.n610 S.n609 0.03
R3535 S.n474 S.n473 0.03
R3536 S.n3093 S.n3090 0.029
R3537 S.n4056 S.n4053 0.029
R3538 S.n2063 S.n2060 0.029
R3539 S.n931 S.n930 0.029
R3540 S.n1496 S.n1495 0.029
R3541 S.n2040 S.n2039 0.029
R3542 S.n2532 S.n2531 0.029
R3543 S.n3070 S.n3069 0.029
R3544 S.n3556 S.n3555 0.029
R3545 S.n4030 S.n4029 0.029
R3546 S.n4467 S.n4466 0.029
R3547 S.n5480 S.n5479 0.029
R3548 S.n1407 S.n1406 0.029
R3549 S.n1954 S.n1953 0.029
R3550 S.n2446 S.n2445 0.029
R3551 S.n2984 S.n2983 0.029
R3552 S.n3470 S.n3469 0.029
R3553 S.n1343 S.n1342 0.029
R3554 S.n1893 S.n1892 0.029
R3555 S.n2385 S.n2384 0.029
R3556 S.n1280 S.n1279 0.029
R3557 S.n1943 S.n1942 0.029
R3558 S.n2435 S.n2434 0.029
R3559 S.n2973 S.n2972 0.029
R3560 S.n3459 S.n3458 0.029
R3561 S.n3975 S.n3974 0.029
R3562 S.n3501 S.n3500 0.029
R3563 S.n3015 S.n3014 0.029
R3564 S.n2477 S.n2476 0.029
R3565 S.n1985 S.n1984 0.029
R3566 S.n1438 S.n1437 0.029
R3567 S.n862 S.n861 0.029
R3568 S.n609 S.n608 0.029
R3569 S.n5463 S.n5460 0.028
R3570 S.n4450 S.n4447 0.028
R3571 S.n4013 S.n4010 0.028
R3572 S.n3539 S.n3536 0.028
R3573 S.n3053 S.n3050 0.028
R3574 S.n2515 S.n2512 0.028
R3575 S.n2023 S.n2020 0.028
R3576 S.n1477 S.n1474 0.028
R3577 S.n2368 S.n2365 0.028
R3578 S.n1876 S.n1873 0.028
R3579 S.n1324 S.n1321 0.028
R3580 S.n770 S.n767 0.028
R3581 S.n1373 S.n1370 0.028
R3582 S.n1923 S.n1920 0.028
R3583 S.n2415 S.n2412 0.028
R3584 S.n2953 S.n2950 0.028
R3585 S.n1261 S.n1258 0.028
R3586 S.n711 S.n708 0.028
R3587 S.n756 S.n753 0.028
R3588 S.n1310 S.n1307 0.028
R3589 S.n1862 S.n1859 0.028
R3590 S.n697 S.n694 0.028
R3591 S.n1423 S.n1422 0.028
R3592 S.n1425 S.n1423 0.028
R3593 S.n1970 S.n1969 0.028
R3594 S.n1972 S.n1970 0.028
R3595 S.n2462 S.n2461 0.028
R3596 S.n2464 S.n2462 0.028
R3597 S.n3000 S.n2999 0.028
R3598 S.n3002 S.n3000 0.028
R3599 S.n3486 S.n3485 0.028
R3600 S.n3488 S.n3486 0.028
R3601 S.n3960 S.n3959 0.028
R3602 S.n3962 S.n3960 0.028
R3603 S.n4484 S.n4483 0.028
R3604 S.n4486 S.n4484 0.028
R3605 S.n879 S.n878 0.028
R3606 S.n881 S.n879 0.028
R3607 S.n907 S.n906 0.028
R3608 S.n909 S.n907 0.028
R3609 S.n5229 S.n5228 0.028
R3610 S.n4056 S.n4055 0.028
R3611 S.n3093 S.n3092 0.028
R3612 S.n2063 S.n2062 0.028
R3613 S.n1394 S.n1393 0.028
R3614 S.n367 S.n362 0.028
R3615 S.n1214 S.n1210 0.028
R3616 S.n1250 S.n1246 0.028
R3617 S.n1836 S.n1832 0.028
R3618 S.n2877 S.n2873 0.028
R3619 S.n2927 S.n2923 0.028
R3620 S.n3442 S.n3438 0.028
R3621 S.n3948 S.n3944 0.028
R3622 S.n4419 S.n4415 0.028
R3623 S.n5454 S.n5450 0.028
R3624 S.n5274 S.n5270 0.028
R3625 S.n4860 S.n4858 0.027
R3626 S.n5861 S.n5859 0.027
R3627 S.n600 S.n595 0.027
R3628 S.n323 S.n322 0.027
R3629 S.n3588 S.n3587 0.027
R3630 S.n2564 S.n2563 0.027
R3631 S.n1528 S.n1527 0.027
R3632 S.n1222 S.n1221 0.027
R3633 S.n1759 S.n1758 0.027
R3634 S.n2103 S.n2102 0.027
R3635 S.n2600 S.n2599 0.027
R3636 S.n3133 S.n3132 0.027
R3637 S.n3810 S.n3809 0.027
R3638 S.n4096 S.n4095 0.027
R3639 S.n4531 S.n4530 0.027
R3640 S.n5525 S.n5524 0.027
R3641 S.n5204 S.n5203 0.027
R3642 S.n1070 S.n1069 0.027
R3643 S.n935 S.n932 0.026
R3644 S.n1150 S.n1149 0.026
R3645 S.n1500 S.n1497 0.026
R3646 S.n1709 S.n1706 0.026
R3647 S.n2044 S.n2041 0.026
R3648 S.n2305 S.n2302 0.026
R3649 S.n2536 S.n2533 0.026
R3650 S.n2801 S.n2798 0.026
R3651 S.n3074 S.n3071 0.026
R3652 S.n3323 S.n3320 0.026
R3653 S.n3560 S.n3557 0.026
R3654 S.n3697 S.n3694 0.026
R3655 S.n4034 S.n4031 0.026
R3656 S.n4286 S.n4283 0.026
R3657 S.n4471 S.n4468 0.026
R3658 S.n4719 S.n4716 0.026
R3659 S.n5484 S.n5481 0.026
R3660 S.n5687 S.n5684 0.026
R3661 S.n5236 S.n5230 0.026
R3662 S.n254 S.n246 0.026
R3663 S.n851 S.n829 0.026
R3664 S.n1092 S.n1080 0.026
R3665 S.n1411 S.n1408 0.026
R3666 S.n1649 S.n1646 0.026
R3667 S.n1958 S.n1955 0.026
R3668 S.n2245 S.n2242 0.026
R3669 S.n2450 S.n2447 0.026
R3670 S.n2741 S.n2738 0.026
R3671 S.n2988 S.n2985 0.026
R3672 S.n3260 S.n3257 0.026
R3673 S.n3474 S.n3471 0.026
R3674 S.n3637 S.n3634 0.026
R3675 S.n4063 S.n4057 0.026
R3676 S.n1102 S.n1100 0.026
R3677 S.n1659 S.n1657 0.026
R3678 S.n2255 S.n2253 0.026
R3679 S.n2751 S.n2749 0.026
R3680 S.n3270 S.n3268 0.026
R3681 S.n3647 S.n3645 0.026
R3682 S.n4236 S.n4234 0.026
R3683 S.n4699 S.n4698 0.026
R3684 S.n4266 S.n4265 0.026
R3685 S.n3677 S.n3676 0.026
R3686 S.n3300 S.n3299 0.026
R3687 S.n2781 S.n2780 0.026
R3688 S.n2285 S.n2284 0.026
R3689 S.n1689 S.n1688 0.026
R3690 S.n1122 S.n1121 0.026
R3691 S.n913 S.n896 0.026
R3692 S.n1466 S.n1456 0.026
R3693 S.n2012 S.n2003 0.026
R3694 S.n2504 S.n2495 0.026
R3695 S.n3042 S.n3033 0.026
R3696 S.n3528 S.n3519 0.026
R3697 S.n4002 S.n3993 0.026
R3698 S.n4439 S.n4430 0.026
R3699 S.n5509 S.n5500 0.026
R3700 S.n3591 S.n3575 0.026
R3701 S.n2956 S.n2938 0.026
R3702 S.n2418 S.n2400 0.026
R3703 S.n1926 S.n1908 0.026
R3704 S.n1376 S.n1358 0.026
R3705 S.n817 S.n801 0.026
R3706 S.n789 S.n784 0.026
R3707 S.n1053 S.n1052 0.026
R3708 S.n1347 S.n1344 0.026
R3709 S.n1613 S.n1610 0.026
R3710 S.n1897 S.n1894 0.026
R3711 S.n2209 S.n2206 0.026
R3712 S.n2389 S.n2386 0.026
R3713 S.n2705 S.n2702 0.026
R3714 S.n3100 S.n3094 0.026
R3715 S.n2567 S.n2551 0.026
R3716 S.n1865 S.n1847 0.026
R3717 S.n1313 S.n1295 0.026
R3718 S.n759 S.n742 0.026
R3719 S.n730 S.n725 0.026
R3720 S.n1019 S.n1018 0.026
R3721 S.n1284 S.n1281 0.026
R3722 S.n1577 S.n1574 0.026
R3723 S.n2070 S.n2064 0.026
R3724 S.n1531 S.n1515 0.026
R3725 S.n700 S.n683 0.026
R3726 S.n959 S.n953 0.026
R3727 S.n494 S.n491 0.026
R3728 S.n494 S.n475 0.026
R3729 S.n5711 S.n5695 0.026
R3730 S.n5166 S.n5165 0.026
R3731 S.n305 S.n304 0.026
R3732 S.n5009 S.n5008 0.026
R3733 S.t241 S.n500 0.025
R3734 S.t241 S.n4 0.025
R3735 S.t241 S.n405 0.025
R3736 S.t241 S.n436 0.025
R3737 S.n619 S.n618 0.024
R3738 S.n1216 S.n1215 0.024
R3739 S.n1252 S.n1251 0.024
R3740 S.n1838 S.n1837 0.024
R3741 S.n2871 S.n2870 0.024
R3742 S.n2929 S.n2928 0.024
R3743 S.n3444 S.n3443 0.024
R3744 S.n3950 S.n3949 0.024
R3745 S.n4421 S.n4420 0.024
R3746 S.n5456 S.n5455 0.024
R3747 S.n5276 S.n5275 0.024
R3748 S.n5287 S.n5286 0.024
R3749 S.n3458 S.n3453 0.024
R3750 S.n2972 S.n2967 0.024
R3751 S.n2434 S.n2429 0.024
R3752 S.n1942 S.n1937 0.024
R3753 S.n1393 S.n1388 0.024
R3754 S.n1445 S.n1421 0.024
R3755 S.n1992 S.n1968 0.024
R3756 S.n2484 S.n2460 0.024
R3757 S.n3022 S.n2998 0.024
R3758 S.n3508 S.n3484 0.024
R3759 S.n3982 S.n3958 0.024
R3760 S.n4498 S.n4482 0.024
R3761 S.n913 S.n912 0.024
R3762 S.n885 S.n884 0.024
R3763 S.n849 S.n848 0.024
R3764 S.n1221 S.n1220 0.024
R3765 S.n618 S.n617 0.024
R3766 S.n2363 S.n2361 0.023
R3767 S.n5704 S.n5703 0.023
R3768 S.n5898 S.n5885 0.023
R3769 S.n5437 S.n5429 0.023
R3770 S.n60 S.n59 0.023
R3771 S.n301 S.n300 0.023
R3772 S.n303 S.n301 0.023
R3773 S.n884 S.n883 0.023
R3774 S.t241 S.n619 0.023
R3775 S.n4664 S.n4663 0.023
R3776 S.n4482 S.n4481 0.023
R3777 S.n3958 S.n3957 0.023
R3778 S.n3484 S.n3483 0.023
R3779 S.n2998 S.n2997 0.023
R3780 S.n2460 S.n2459 0.023
R3781 S.n1968 S.n1967 0.023
R3782 S.n1421 S.n1420 0.023
R3783 S.n1445 S.n1425 0.023
R3784 S.n1992 S.n1972 0.023
R3785 S.n2484 S.n2464 0.023
R3786 S.n3022 S.n3002 0.023
R3787 S.n3508 S.n3488 0.023
R3788 S.n3982 S.n3962 0.023
R3789 S.n4498 S.n4486 0.023
R3790 S.n212 S.n210 0.023
R3791 S.n912 S.n911 0.023
R3792 S.n324 S.n323 0.023
R3793 S.n913 S.n909 0.023
R3794 S.n885 S.n881 0.023
R3795 S.n61 S.n57 0.023
R3796 S.n39 S.n38 0.023
R3797 S.n40 S.n36 0.023
R3798 S.n18 S.n17 0.023
R3799 S.n19 S.n15 0.023
R3800 S.n5356 S.n5354 0.023
R3801 S.n677 S.n675 0.023
R3802 S.n1219 S.n1218 0.023
R3803 S.n1807 S.n1805 0.023
R3804 S.n1230 S.n1229 0.023
R3805 S.n2357 S.n2355 0.023
R3806 S.n1816 S.n1815 0.023
R3807 S.n2887 S.n2886 0.023
R3808 S.n3413 S.n3411 0.023
R3809 S.n2907 S.n2906 0.023
R3810 S.n3919 S.n3917 0.023
R3811 S.n3422 S.n3421 0.023
R3812 S.n4400 S.n4398 0.023
R3813 S.n3928 S.n3927 0.023
R3814 S.n4854 S.n4852 0.023
R3815 S.n5302 S.n5294 0.023
R3816 S.n3453 S.n3451 0.023
R3817 S.n2967 S.n2964 0.023
R3818 S.n2429 S.n2427 0.023
R3819 S.n1937 S.n1934 0.023
R3820 S.n1388 S.n1386 0.023
R3821 S.n848 S.n845 0.023
R3822 S.n840 S.n839 0.023
R3823 S.n5234 S.n5233 0.022
R3824 S.n839 S.n838 0.022
R3825 S.n3977 S.n3973 0.022
R3826 S.n3503 S.n3499 0.022
R3827 S.n3017 S.n3013 0.022
R3828 S.n2479 S.n2475 0.022
R3829 S.n1987 S.n1983 0.022
R3830 S.n1440 S.n1436 0.022
R3831 S.n864 S.n860 0.022
R3832 S.n611 S.n607 0.022
R3833 S.n5495 S.n5494 0.022
R3834 S.n1239 S.n1237 0.022
R3835 S.n1825 S.n1823 0.022
R3836 S.n2896 S.n2894 0.022
R3837 S.n2916 S.n2914 0.022
R3838 S.n3431 S.n3429 0.022
R3839 S.n3937 S.n3935 0.022
R3840 S.n4061 S.n4060 0.022
R3841 S.n3570 S.n3568 0.022
R3842 S.n3098 S.n3097 0.022
R3843 S.n2546 S.n2544 0.022
R3844 S.n2068 S.n2067 0.022
R3845 S.n1510 S.n1508 0.022
R3846 S.n957 S.n956 0.022
R3847 S.n470 S.n468 0.022
R3848 S.n5499 S.n5498 0.022
R3849 S.n5229 S.n5226 0.021
R3850 S.n929 S.n928 0.021
R3851 S.n1495 S.n1494 0.021
R3852 S.n1491 S.n1490 0.021
R3853 S.n2039 S.n2038 0.021
R3854 S.n2037 S.n2036 0.021
R3855 S.n2531 S.n2530 0.021
R3856 S.n2529 S.n2528 0.021
R3857 S.n3069 S.n3068 0.021
R3858 S.n3067 S.n3066 0.021
R3859 S.n3555 S.n3554 0.021
R3860 S.n3553 S.n3552 0.021
R3861 S.n4029 S.n4028 0.021
R3862 S.n4027 S.n4026 0.021
R3863 S.n4466 S.n4465 0.021
R3864 S.n4464 S.n4463 0.021
R3865 S.n5479 S.n5478 0.021
R3866 S.n5477 S.n5476 0.021
R3867 S.n5228 S.n5227 0.021
R3868 S.n337 S.n336 0.021
R3869 S.n826 S.n825 0.021
R3870 S.n1406 S.n1405 0.021
R3871 S.n1402 S.n1401 0.021
R3872 S.n1953 S.n1952 0.021
R3873 S.n1951 S.n1950 0.021
R3874 S.n2445 S.n2444 0.021
R3875 S.n2443 S.n2442 0.021
R3876 S.n2983 S.n2982 0.021
R3877 S.n2981 S.n2980 0.021
R3878 S.n3469 S.n3468 0.021
R3879 S.n3467 S.n3466 0.021
R3880 S.n4055 S.n4054 0.021
R3881 S.n787 S.n786 0.021
R3882 S.n1342 S.n1341 0.021
R3883 S.n1338 S.n1337 0.021
R3884 S.n1892 S.n1891 0.021
R3885 S.n1890 S.n1889 0.021
R3886 S.n2384 S.n2383 0.021
R3887 S.n2382 S.n2381 0.021
R3888 S.n3092 S.n3091 0.021
R3889 S.n728 S.n727 0.021
R3890 S.n1279 S.n1278 0.021
R3891 S.n1275 S.n1274 0.021
R3892 S.n2062 S.n2061 0.021
R3893 S.n4667 S.n4666 0.021
R3894 S.n5462 S.n5461 0.021
R3895 S.n4449 S.n4448 0.021
R3896 S.n4012 S.n4011 0.021
R3897 S.n3538 S.n3537 0.021
R3898 S.n3052 S.n3051 0.021
R3899 S.n2514 S.n2513 0.021
R3900 S.n2022 S.n2021 0.021
R3901 S.n1476 S.n1475 0.021
R3902 S.n335 S.n334 0.021
R3903 S.n2367 S.n2366 0.021
R3904 S.n1875 S.n1874 0.021
R3905 S.n1323 S.n1322 0.021
R3906 S.n769 S.n768 0.021
R3907 S.n4062 S.n4061 0.021
R3908 S.n4497 S.n4496 0.021
R3909 S.n813 S.n812 0.021
R3910 S.n1372 S.n1371 0.021
R3911 S.n1922 S.n1921 0.021
R3912 S.n2414 S.n2413 0.021
R3913 S.n2952 S.n2951 0.021
R3914 S.n3572 S.n3570 0.021
R3915 S.n6 S.n5 0.021
R3916 S.n3099 S.n3098 0.021
R3917 S.n1260 S.n1259 0.021
R3918 S.n710 S.n709 0.021
R3919 S.n755 S.n754 0.021
R3920 S.n1309 S.n1308 0.021
R3921 S.n1861 S.n1860 0.021
R3922 S.n2548 S.n2546 0.021
R3923 S.n407 S.n406 0.021
R3924 S.n2069 S.n2068 0.021
R3925 S.n696 S.n695 0.021
R3926 S.n1512 S.n1510 0.021
R3927 S.n438 S.n437 0.021
R3928 S.n958 S.n957 0.021
R3929 S.n472 S.n470 0.021
R3930 S.n5363 S.n5361 0.021
R3931 S.n4406 S.n4405 0.021
R3932 S.n5301 S.n5298 0.02
R3933 S.n5436 S.n5433 0.02
R3934 S.n631 S.n630 0.02
R3935 S.n8 S.n7 0.02
R3936 S.n409 S.n408 0.02
R3937 S.n440 S.n439 0.02
R3938 S.n489 S.n488 0.02
R3939 S.n5247 S.n5246 0.02
R3940 S.n5235 S.n5232 0.02
R3941 S.n3453 S.n3452 0.02
R3942 S.n2967 S.n2966 0.02
R3943 S.n2429 S.n2428 0.02
R3944 S.n1937 S.n1936 0.02
R3945 S.n1388 S.n1387 0.02
R3946 S.n4062 S.n4058 0.02
R3947 S.n5496 S.n5493 0.02
R3948 S.n848 S.n847 0.02
R3949 S.n3572 S.n3571 0.02
R3950 S.n3099 S.n3095 0.02
R3951 S.n2548 S.n2547 0.02
R3952 S.n2069 S.n2065 0.02
R3953 S.n1512 S.n1511 0.02
R3954 S.n958 S.n954 0.02
R3955 S.n472 S.n471 0.02
R3956 S.n623 S.n622 0.02
R3957 S.t241 S.n572 0.019
R3958 S.n1105 S.n1103 0.019
R3959 S.n1662 S.n1660 0.019
R3960 S.n2258 S.n2256 0.019
R3961 S.n2754 S.n2752 0.019
R3962 S.n3273 S.n3271 0.019
R3963 S.n3650 S.n3648 0.019
R3964 S.n4239 S.n4237 0.019
R3965 S.n581 S.n580 0.019
R3966 S.n1124 S.n1123 0.019
R3967 S.n367 S.n366 0.019
R3968 S.n1214 S.n1213 0.019
R3969 S.n1250 S.n1249 0.019
R3970 S.n1836 S.n1835 0.019
R3971 S.n2877 S.n2876 0.019
R3972 S.n2927 S.n2926 0.019
R3973 S.n3442 S.n3441 0.019
R3974 S.n3948 S.n3947 0.019
R3975 S.n4419 S.n4418 0.019
R3976 S.n5454 S.n5453 0.019
R3977 S.n5274 S.n5273 0.019
R3978 S.n3981 S.n3980 0.019
R3979 S.n3507 S.n3506 0.019
R3980 S.n3021 S.n3020 0.019
R3981 S.n2483 S.n2482 0.019
R3982 S.n1991 S.n1990 0.019
R3983 S.n1444 S.n1443 0.019
R3984 S.n868 S.n867 0.019
R3985 S.n5646 S.n5645 0.019
R3986 S.n597 S.n596 0.018
R3987 S.n572 S.n571 0.018
R3988 S.n57 S.n56 0.018
R3989 S.n36 S.n35 0.018
R3990 S.n15 S.n14 0.018
R3991 S S.n673 0.018
R3992 S.n4819 S.n4818 0.018
R3993 S.n576 S.n575 0.018
R3994 S.n847 S.n846 0.018
R3995 S.n2966 S.n2965 0.018
R3996 S.n1936 S.n1935 0.018
R3997 S.n4816 S.n4815 0.017
R3998 S.n5163 S.n5162 0.017
R3999 S.n5006 S.n5005 0.017
R4000 S.n4823 S.n4820 0.017
R4001 S.n5895 S.n5894 0.017
R4002 S.n5894 S.n5893 0.017
R4003 S.n1242 S.n1241 0.017
R4004 S.n1828 S.n1827 0.017
R4005 S.n2899 S.n2898 0.017
R4006 S.n2919 S.n2918 0.017
R4007 S.n3434 S.n3433 0.017
R4008 S.n3940 S.n3939 0.017
R4009 S.n851 S.n840 0.016
R4010 S.n1092 S.n1088 0.016
R4011 S.n3591 S.n3583 0.016
R4012 S.n2567 S.n2559 0.016
R4013 S.n1531 S.n1523 0.016
R4014 S.n1240 S.n1239 0.016
R4015 S.n1826 S.n1825 0.016
R4016 S.n2897 S.n2896 0.016
R4017 S.n2917 S.n2916 0.016
R4018 S.n3432 S.n3431 0.016
R4019 S.n3938 S.n3937 0.016
R4020 S.n3451 S.n3450 0.015
R4021 S.n2427 S.n2426 0.015
R4022 S.n1386 S.n1385 0.015
R4023 S.n5859 S.n5858 0.015
R4024 S.n851 S.n850 0.015
R4025 S.n5226 S.n5225 0.015
R4026 S.n3979 S.n3978 0.015
R4027 S.n3978 S.n3977 0.015
R4028 S.n3977 S.n3976 0.015
R4029 S.n3505 S.n3504 0.015
R4030 S.n3504 S.n3503 0.015
R4031 S.n3503 S.n3502 0.015
R4032 S.n3019 S.n3018 0.015
R4033 S.n3018 S.n3017 0.015
R4034 S.n3017 S.n3016 0.015
R4035 S.n2481 S.n2480 0.015
R4036 S.n2480 S.n2479 0.015
R4037 S.n2479 S.n2478 0.015
R4038 S.n1989 S.n1988 0.015
R4039 S.n1988 S.n1987 0.015
R4040 S.n1987 S.n1986 0.015
R4041 S.n1442 S.n1441 0.015
R4042 S.n1441 S.n1440 0.015
R4043 S.n1440 S.n1439 0.015
R4044 S.n866 S.n865 0.015
R4045 S.n865 S.n864 0.015
R4046 S.n864 S.n863 0.015
R4047 S.n612 S.n611 0.015
R4048 S.n611 S.n610 0.015
R4049 S.n5498 S.n5497 0.015
R4050 S.n326 S.n325 0.015
R4051 S.t283 S.n5356 0.015
R4052 S.n1809 S.n1254 0.015
R4053 S.n2359 S.n1840 0.015
R4054 S.n2900 S.n2880 0.015
R4055 S.n3415 S.n2931 0.015
R4056 S.n3921 S.n3446 0.015
R4057 S.n4402 S.n3952 0.015
R4058 S.n5644 S.n5643 0.015
R4059 S.n5643 S.n5642 0.015
R4060 S.n4818 S.n4817 0.015
R4061 S.n4856 S.n4423 0.015
R4062 S.n5465 S.n5464 0.015
R4063 S.n4452 S.n4451 0.015
R4064 S.n4015 S.n4014 0.015
R4065 S.n3541 S.n3540 0.015
R4066 S.n3055 S.n3054 0.015
R4067 S.n2517 S.n2516 0.015
R4068 S.n2025 S.n2024 0.015
R4069 S.n1479 S.n1478 0.015
R4070 S.n2370 S.n2369 0.015
R4071 S.n1878 S.n1877 0.015
R4072 S.n1326 S.n1325 0.015
R4073 S.n772 S.n771 0.015
R4074 S.n2947 S.n2946 0.015
R4075 S.n2409 S.n2408 0.015
R4076 S.n1917 S.n1916 0.015
R4077 S.n1367 S.n1366 0.015
R4078 S.n809 S.n808 0.015
R4079 S.n1263 S.n1262 0.015
R4080 S.n713 S.n712 0.015
R4081 S.n1856 S.n1855 0.015
R4082 S.n1304 S.n1303 0.015
R4083 S.n750 S.n749 0.015
R4084 S.n691 S.n690 0.015
R4085 S.n615 S.n614 0.014
R4086 S.n4409 S.n4407 0.014
R4087 S.n776 S.n775 0.014
R4088 S.n1375 S.n1374 0.014
R4089 S.n1925 S.n1924 0.014
R4090 S.n2417 S.n2416 0.014
R4091 S.n2955 S.n2954 0.014
R4092 S.n717 S.n716 0.014
R4093 S.n1312 S.n1311 0.014
R4094 S.n1864 S.n1863 0.014
R4095 S.n4869 S.n4860 0.014
R4096 S.n5871 S.n5861 0.014
R4097 S.n850 S.n849 0.014
R4098 S.n1071 S.n1070 0.014
R4099 S.n1729 S.n1728 0.014
R4100 S.n2325 S.n2324 0.014
R4101 S.n3372 S.n3371 0.014
R4102 S.n3780 S.n3779 0.014
R4103 S.n4354 S.n4353 0.014
R4104 S.n5710 S.n5709 0.014
R4105 S.n2837 S.n2836 0.014
R4106 S.n5469 S.n5468 0.013
R4107 S.n4456 S.n4455 0.013
R4108 S.n4019 S.n4018 0.013
R4109 S.n3545 S.n3544 0.013
R4110 S.n3059 S.n3058 0.013
R4111 S.n2521 S.n2520 0.013
R4112 S.n2029 S.n2028 0.013
R4113 S.n1483 S.n1482 0.013
R4114 S.n2374 S.n2373 0.013
R4115 S.n1882 S.n1881 0.013
R4116 S.n1330 S.n1329 0.013
R4117 S.n816 S.n815 0.013
R4118 S.n1267 S.n1266 0.013
R4119 S.n758 S.n757 0.013
R4120 S.n699 S.n698 0.013
R4121 S.n4495 S.n4494 0.013
R4122 S.n1728 S.n1727 0.013
R4123 S.n2324 S.n2323 0.013
R4124 S.n2836 S.n2835 0.013
R4125 S.n3371 S.n3370 0.013
R4126 S.n3779 S.n3778 0.013
R4127 S.n4353 S.n4352 0.013
R4128 S.n5709 S.n5708 0.013
R4129 S.t241 S.n0 0.012
R4130 S.t241 S.n401 0.012
R4131 S.t241 S.n432 0.012
R4132 S.t241 S.n501 0.012
R4133 S.n4423 S.n4411 0.012
R4134 S.n5891 S.n5890 0.012
R4135 S.n5466 S.n5465 0.012
R4136 S.n4453 S.n4452 0.012
R4137 S.n4016 S.n4015 0.012
R4138 S.n3542 S.n3541 0.012
R4139 S.n3056 S.n3055 0.012
R4140 S.n2518 S.n2517 0.012
R4141 S.n2026 S.n2025 0.012
R4142 S.n1480 S.n1479 0.012
R4143 S.n348 S.n339 0.012
R4144 S.n2371 S.n2370 0.012
R4145 S.n1879 S.n1878 0.012
R4146 S.n1327 S.n1326 0.012
R4147 S.n773 S.n772 0.012
R4148 S.n2948 S.n2947 0.012
R4149 S.n2410 S.n2409 0.012
R4150 S.n1918 S.n1917 0.012
R4151 S.n1368 S.n1367 0.012
R4152 S.n843 S.n842 0.012
R4153 S.n3456 S.n3455 0.012
R4154 S.n2970 S.n2969 0.012
R4155 S.n2432 S.n2431 0.012
R4156 S.n1940 S.n1939 0.012
R4157 S.n1391 S.n1390 0.012
R4158 S.n810 S.n809 0.012
R4159 S.n394 S.n10 0.012
R4160 S.n1264 S.n1263 0.012
R4161 S.n714 S.n713 0.012
R4162 S.n1857 S.n1856 0.012
R4163 S.n1305 S.n1304 0.012
R4164 S.n751 S.n750 0.012
R4165 S.n425 S.n411 0.012
R4166 S.n692 S.n691 0.012
R4167 S.n456 S.n442 0.012
R4168 S.n1727 S.n1726 0.012
R4169 S.n1237 S.n1236 0.012
R4170 S.n2323 S.n2322 0.012
R4171 S.n1823 S.n1822 0.012
R4172 S.n2894 S.n2893 0.012
R4173 S.n2835 S.n2834 0.012
R4174 S.n3370 S.n3369 0.012
R4175 S.n2914 S.n2913 0.012
R4176 S.n3778 S.n3777 0.012
R4177 S.n3429 S.n3428 0.012
R4178 S.n4352 S.n4351 0.012
R4179 S.n3935 S.n3934 0.012
R4180 S.n5297 S.n5296 0.012
R4181 S.n5432 S.n5431 0.012
R4182 S.n5708 S.n5707 0.012
R4183 S.n5018 S.n5009 0.011
R4184 S.n5175 S.n5166 0.011
R4185 S.n4823 S.n4816 0.01
R4186 S.n186 S.n185 0.01
R4187 S.n153 S.n152 0.01
R4188 S.n120 S.n119 0.01
R4189 S.n4044 S.n4043 0.01
R4190 S.n305 S.n303 0.01
R4191 S.n1113 S.n1105 0.01
R4192 S.n1670 S.n1662 0.01
R4193 S.n2266 S.n2258 0.01
R4194 S.n2762 S.n2754 0.01
R4195 S.n3281 S.n3273 0.01
R4196 S.n3658 S.n3650 0.01
R4197 S.n4247 S.n4239 0.01
R4198 S.n215 S.n212 0.01
R4199 S.n4700 S.n4696 0.01
R4200 S.n4267 S.n4263 0.01
R4201 S.n3678 S.n3674 0.01
R4202 S.n3301 S.n3297 0.01
R4203 S.n2782 S.n2778 0.01
R4204 S.n2286 S.n2282 0.01
R4205 S.n1690 S.n1686 0.01
R4206 S.n1133 S.n1124 0.01
R4207 S.n234 S.n231 0.01
R4208 S.n61 S.n60 0.01
R4209 S.n40 S.n39 0.01
R4210 S.n19 S.n18 0.01
R4211 S.n273 S.n270 0.01
R4212 S.n1222 S.n1219 0.01
R4213 S.n1222 S.n677 0.01
R4214 S.n1809 S.n1807 0.01
R4215 S.n2359 S.n2357 0.01
R4216 S.n3415 S.n3413 0.01
R4217 S.n3921 S.n3919 0.01
R4218 S.n4402 S.n4400 0.01
R4219 S.n4856 S.n4854 0.01
R4220 S.n5175 S.n5163 0.01
R4221 S.n5018 S.n5006 0.01
R4222 S.n5900 S.n5898 0.01
R4223 S.n2900 S.n2363 0.01
R4224 S.n10 S.n9 0.01
R4225 S.n411 S.n410 0.01
R4226 S.n442 S.n441 0.01
R4227 S.n5893 S.n5891 0.01
R4228 S.n1091 S.n1089 0.01
R4229 S.n59 S.n58 0.01
R4230 S.n38 S.n37 0.01
R4231 S.n17 S.n16 0.01
R4232 S.n4681 S.n4667 0.01
R4233 S.n3619 S.n3604 0.01
R4234 S.n2687 S.n2672 0.01
R4235 S.n1559 S.n1544 0.01
R4236 S.n5280 S.n5267 0.009
R4237 S.n5896 S.n5895 0.009
R4238 S.n4498 S.n4497 0.009
R4239 S.t283 S.n5363 0.009
R4240 S.n5900 S.n5458 0.009
R4241 S.n5162 S.n5161 0.008
R4242 S.n5005 S.n5004 0.008
R4243 S.n5301 S.n5300 0.008
R4244 S.n5436 S.n5435 0.008
R4245 S.n5467 S.n5466 0.008
R4246 S.n4454 S.n4453 0.008
R4247 S.n4017 S.n4016 0.008
R4248 S.n3543 S.n3542 0.008
R4249 S.n3057 S.n3056 0.008
R4250 S.n2519 S.n2518 0.008
R4251 S.n2027 S.n2026 0.008
R4252 S.n1481 S.n1480 0.008
R4253 S.n2372 S.n2371 0.008
R4254 S.n1880 S.n1879 0.008
R4255 S.n1328 S.n1327 0.008
R4256 S.n774 S.n773 0.008
R4257 S.n2949 S.n2948 0.008
R4258 S.n2411 S.n2410 0.008
R4259 S.n1919 S.n1918 0.008
R4260 S.n1369 S.n1368 0.008
R4261 S.n811 S.n810 0.008
R4262 S.n1265 S.n1264 0.008
R4263 S.n715 S.n714 0.008
R4264 S.n1858 S.n1857 0.008
R4265 S.n1306 S.n1305 0.008
R4266 S.n752 S.n751 0.008
R4267 S.n693 S.n692 0.008
R4268 S.n934 S.n933 0.008
R4269 S.n1493 S.n1492 0.008
R4270 S.n1499 S.n1498 0.008
R4271 S.n1708 S.n1707 0.008
R4272 S.n2043 S.n2042 0.008
R4273 S.n2304 S.n2303 0.008
R4274 S.n2535 S.n2534 0.008
R4275 S.n2800 S.n2799 0.008
R4276 S.n3073 S.n3072 0.008
R4277 S.n3322 S.n3321 0.008
R4278 S.n3559 S.n3558 0.008
R4279 S.n3696 S.n3695 0.008
R4280 S.n4033 S.n4032 0.008
R4281 S.n4285 S.n4284 0.008
R4282 S.n4470 S.n4469 0.008
R4283 S.n4718 S.n4717 0.008
R4284 S.n5483 S.n5482 0.008
R4285 S.n5686 S.n5685 0.008
R4286 S.n243 S.n242 0.008
R4287 S.n827 S.n824 0.008
R4288 S.n1404 S.n1403 0.008
R4289 S.n1410 S.n1409 0.008
R4290 S.n1648 S.n1647 0.008
R4291 S.n1957 S.n1956 0.008
R4292 S.n2244 S.n2243 0.008
R4293 S.n2449 S.n2448 0.008
R4294 S.n2740 S.n2739 0.008
R4295 S.n2987 S.n2986 0.008
R4296 S.n3259 S.n3258 0.008
R4297 S.n3473 S.n3472 0.008
R4298 S.n3636 S.n3635 0.008
R4299 S.n1113 S.n1102 0.008
R4300 S.n1670 S.n1659 0.008
R4301 S.n2266 S.n2255 0.008
R4302 S.n2762 S.n2751 0.008
R4303 S.n3281 S.n3270 0.008
R4304 S.n3658 S.n3647 0.008
R4305 S.n4247 S.n4236 0.008
R4306 S.n215 S.n214 0.008
R4307 S.n4700 S.n4699 0.008
R4308 S.n4267 S.n4266 0.008
R4309 S.n3678 S.n3677 0.008
R4310 S.n3301 S.n3300 0.008
R4311 S.n2782 S.n2781 0.008
R4312 S.n2286 S.n2285 0.008
R4313 S.n1690 S.n1689 0.008
R4314 S.n1133 S.n1122 0.008
R4315 S.n893 S.n892 0.008
R4316 S.n1453 S.n1452 0.008
R4317 S.n2000 S.n1999 0.008
R4318 S.n2492 S.n2491 0.008
R4319 S.n3030 S.n3029 0.008
R4320 S.n3516 S.n3515 0.008
R4321 S.n3990 S.n3989 0.008
R4322 S.n4427 S.n4426 0.008
R4323 S.n313 S.n312 0.008
R4324 S.n325 S.n321 0.008
R4325 S.n325 S.n324 0.008
R4326 S.n234 S.n233 0.008
R4327 S.n3590 S.n3586 0.008
R4328 S.n2935 S.n2934 0.008
R4329 S.n2397 S.n2396 0.008
R4330 S.n1905 S.n1904 0.008
R4331 S.n1355 S.n1354 0.008
R4332 S.n798 S.n797 0.008
R4333 S.n788 S.n785 0.008
R4334 S.n1340 S.n1339 0.008
R4335 S.n1346 S.n1345 0.008
R4336 S.n1612 S.n1611 0.008
R4337 S.n1896 S.n1895 0.008
R4338 S.n2208 S.n2207 0.008
R4339 S.n2388 S.n2387 0.008
R4340 S.n2704 S.n2703 0.008
R4341 S.n2566 S.n2562 0.008
R4342 S.n1844 S.n1843 0.008
R4343 S.n1292 S.n1291 0.008
R4344 S.n739 S.n738 0.008
R4345 S.n729 S.n726 0.008
R4346 S.n1277 S.n1276 0.008
R4347 S.n1283 S.n1282 0.008
R4348 S.n1576 S.n1575 0.008
R4349 S.n1530 S.n1526 0.008
R4350 S.n680 S.n679 0.008
R4351 S.n493 S.n492 0.008
R4352 S.n273 S.n272 0.008
R4353 S.n378 S.n377 0.008
R4354 S.n4823 S.n4822 0.008
R4355 S.n5245 S.n5244 0.008
R4356 S.n599 S.n598 0.008
R4357 S.n599 S.n597 0.007
R4358 S.t241 S.n564 0.007
R4359 S.t241 S.n557 0.007
R4360 S.t241 S.n545 0.007
R4361 S.t241 S.n533 0.007
R4362 S.n614 S.n613 0.007
R4363 S.n4815 S.n4814 0.007
R4364 S.t283 S.n5370 0.006
R4365 S.t283 S.n5378 0.006
R4366 S.t283 S.n5386 0.006
R4367 S.t283 S.n5394 0.006
R4368 S.t283 S.n5402 0.006
R4369 S.t283 S.n5410 0.006
R4370 S.t283 S.n5423 0.006
R4371 S.n1494 S.n1493 0.006
R4372 S.n827 S.n826 0.006
R4373 S.n1405 S.n1404 0.006
R4374 S.n788 S.n787 0.006
R4375 S.n1341 S.n1340 0.006
R4376 S.n729 S.n728 0.006
R4377 S.n1278 S.n1277 0.006
R4378 S.n5246 S.n5245 0.006
R4379 S.n5302 S.n5301 0.006
R4380 S.n5437 S.n5436 0.006
R4381 S.n70 S.n61 0.006
R4382 S.n49 S.n40 0.006
R4383 S.n28 S.n19 0.006
R4384 S.n305 S.n292 0.005
R4385 S.n844 S.n843 0.005
R4386 S.n3457 S.n3456 0.005
R4387 S.n2971 S.n2970 0.005
R4388 S.n2433 S.n2432 0.005
R4389 S.n1941 S.n1940 0.005
R4390 S.n1392 S.n1391 0.005
R4391 S.t241 S.n569 0.005
R4392 S.n3585 S.n3584 0.005
R4393 S.n2561 S.n2560 0.005
R4394 S.n1525 S.n1524 0.005
R4395 S.n5300 S.n5299 0.005
R4396 S.n5435 S.n5434 0.005
R4397 S.t241 S.n616 0.005
R4398 S.n5016 S.n5015 0.004
R4399 S.n5255 S.n5254 0.004
R4400 S.n5702 S.n5701 0.004
R4401 S.n5884 S.n5883 0.004
R4402 S.n487 S.n486 0.004
R4403 S.n346 S.n345 0.004
R4404 S.n924 S.n923 0.004
R4405 S.n5221 S.n5220 0.004
R4406 S.n5679 S.n5678 0.004
R4407 S.n5472 S.n5471 0.004
R4408 S.n4711 S.n4710 0.004
R4409 S.n4459 S.n4458 0.004
R4410 S.n4278 S.n4277 0.004
R4411 S.n4022 S.n4021 0.004
R4412 S.n3689 S.n3688 0.004
R4413 S.n3548 S.n3547 0.004
R4414 S.n3315 S.n3314 0.004
R4415 S.n3062 S.n3061 0.004
R4416 S.n2793 S.n2792 0.004
R4417 S.n2524 S.n2523 0.004
R4418 S.n2297 S.n2296 0.004
R4419 S.n2032 S.n2031 0.004
R4420 S.n1701 S.n1700 0.004
R4421 S.n1486 S.n1485 0.004
R4422 S.n1144 S.n1143 0.004
R4423 S.n252 S.n251 0.004
R4424 S.n68 S.n67 0.004
R4425 S.n779 S.n778 0.004
R4426 S.n3086 S.n3085 0.004
R4427 S.n2697 S.n2696 0.004
R4428 S.n2377 S.n2376 0.004
R4429 S.n2201 S.n2200 0.004
R4430 S.n1885 S.n1884 0.004
R4431 S.n1605 S.n1604 0.004
R4432 S.n1333 S.n1332 0.004
R4433 S.n1047 S.n1046 0.004
R4434 S.n392 S.n391 0.004
R4435 S.n3582 S.n3581 0.004
R4436 S.n3239 S.n3238 0.004
R4437 S.n2945 S.n2944 0.004
R4438 S.n2720 S.n2719 0.004
R4439 S.n2407 S.n2406 0.004
R4440 S.n2224 S.n2223 0.004
R4441 S.n1915 S.n1914 0.004
R4442 S.n1628 S.n1627 0.004
R4443 S.n1365 S.n1364 0.004
R4444 S.n1068 S.n1067 0.004
R4445 S.n1087 S.n1086 0.004
R4446 S.n836 S.n835 0.004
R4447 S.n288 S.n287 0.004
R4448 S.n299 S.n298 0.004
R4449 S.n1397 S.n1396 0.004
R4450 S.n1946 S.n1945 0.004
R4451 S.n2438 S.n2437 0.004
R4452 S.n2976 S.n2975 0.004
R4453 S.n3462 S.n3461 0.004
R4454 S.n4049 S.n4048 0.004
R4455 S.n3629 S.n3628 0.004
R4456 S.n3252 S.n3251 0.004
R4457 S.n2733 S.n2732 0.004
R4458 S.n2237 S.n2236 0.004
R4459 S.n1641 S.n1640 0.004
R4460 S.n875 S.n874 0.004
R4461 S.n209 S.n208 0.004
R4462 S.n593 S.n592 0.004
R4463 S.n4490 S.n4489 0.004
R4464 S.n4242 S.n4241 0.004
R4465 S.n3967 S.n3966 0.004
R4466 S.n3653 S.n3652 0.004
R4467 S.n3493 S.n3492 0.004
R4468 S.n3276 S.n3275 0.004
R4469 S.n3007 S.n3006 0.004
R4470 S.n2757 S.n2756 0.004
R4471 S.n2469 S.n2468 0.004
R4472 S.n2261 S.n2260 0.004
R4473 S.n1977 S.n1976 0.004
R4474 S.n1665 S.n1664 0.004
R4475 S.n1430 S.n1429 0.004
R4476 S.n1108 S.n1107 0.004
R4477 S.n903 S.n902 0.004
R4478 S.n229 S.n228 0.004
R4479 S.n1127 S.n1126 0.004
R4480 S.n1463 S.n1462 0.004
R4481 S.n1685 S.n1684 0.004
R4482 S.n2010 S.n2009 0.004
R4483 S.n2281 S.n2280 0.004
R4484 S.n2502 S.n2501 0.004
R4485 S.n2777 S.n2776 0.004
R4486 S.n3040 S.n3039 0.004
R4487 S.n3296 S.n3295 0.004
R4488 S.n3526 S.n3525 0.004
R4489 S.n3673 S.n3672 0.004
R4490 S.n4000 S.n3999 0.004
R4491 S.n4262 S.n4261 0.004
R4492 S.n4437 S.n4436 0.004
R4493 S.n4695 S.n4694 0.004
R4494 S.n5507 S.n5506 0.004
R4495 S.n319 S.n318 0.004
R4496 S.n807 S.n806 0.004
R4497 S.n193 S.n192 0.004
R4498 S.n176 S.n175 0.004
R4499 S.n47 S.n46 0.004
R4500 S.n720 S.n719 0.004
R4501 S.n2056 S.n2055 0.004
R4502 S.n1569 S.n1568 0.004
R4503 S.n1270 S.n1269 0.004
R4504 S.n1013 S.n1012 0.004
R4505 S.n423 S.n422 0.004
R4506 S.n2558 S.n2557 0.004
R4507 S.n2188 S.n2187 0.004
R4508 S.n1854 S.n1853 0.004
R4509 S.n1592 S.n1591 0.004
R4510 S.n1302 S.n1301 0.004
R4511 S.n1034 S.n1033 0.004
R4512 S.n748 S.n747 0.004
R4513 S.n160 S.n159 0.004
R4514 S.n143 S.n142 0.004
R4515 S.n26 S.n25 0.004
R4516 S.n947 S.n946 0.004
R4517 S.n454 S.n453 0.004
R4518 S.n1522 S.n1521 0.004
R4519 S.n1000 S.n999 0.004
R4520 S.n689 S.n688 0.004
R4521 S.n127 S.n126 0.004
R4522 S.n110 S.n109 0.004
R4523 S.n373 S.n372 0.004
R4524 S.n269 S.n268 0.004
R4525 S.n1193 S.n1192 0.004
R4526 S.n1182 S.n1181 0.004
R4527 S.n1757 S.n1756 0.004
R4528 S.n1745 S.n1744 0.004
R4529 S.n2101 S.n2100 0.004
R4530 S.n2089 S.n2088 0.004
R4531 S.n2598 S.n2597 0.004
R4532 S.n2586 S.n2585 0.004
R4533 S.n3131 S.n3130 0.004
R4534 S.n3119 S.n3118 0.004
R4535 S.n3808 S.n3807 0.004
R4536 S.n3796 S.n3795 0.004
R4537 S.n4094 S.n4093 0.004
R4538 S.n4082 S.n4081 0.004
R4539 S.n4529 S.n4528 0.004
R4540 S.n4517 S.n4516 0.004
R4541 S.n5523 S.n5522 0.004
R4542 S.n5725 S.n5724 0.004
R4543 S.n5202 S.n5201 0.004
R4544 S.n5190 S.n5189 0.004
R4545 S.n1208 S.n1207 0.004
R4546 S.n1165 S.n1164 0.004
R4547 S.n1774 S.n1773 0.004
R4548 S.n4978 S.n4977 0.004
R4549 S.n4970 S.n4969 0.004
R4550 S.n5740 S.n5739 0.004
R4551 S.n5540 S.n5539 0.004
R4552 S.n4554 S.n4553 0.004
R4553 S.n4546 S.n4545 0.004
R4554 S.n4119 S.n4118 0.004
R4555 S.n4111 S.n4110 0.004
R4556 S.n3833 S.n3832 0.004
R4557 S.n3825 S.n3824 0.004
R4558 S.n3156 S.n3155 0.004
R4559 S.n3148 S.n3147 0.004
R4560 S.n2623 S.n2622 0.004
R4561 S.n2615 S.n2614 0.004
R4562 S.n2129 S.n2128 0.004
R4563 S.n2118 S.n2117 0.004
R4564 S.n1782 S.n1781 0.004
R4565 S.n1256 S.n1255 0.004
R4566 S.n1724 S.n1723 0.004
R4567 S.n2149 S.n2148 0.004
R4568 S.n5051 S.n5050 0.004
R4569 S.n4955 S.n4954 0.004
R4570 S.n5755 S.n5754 0.004
R4571 S.n5556 S.n5555 0.004
R4572 S.n4731 S.n4730 0.004
R4573 S.n4577 S.n4576 0.004
R4574 S.n4298 S.n4297 0.004
R4575 S.n4142 S.n4141 0.004
R4576 S.n3709 S.n3708 0.004
R4577 S.n3856 S.n3855 0.004
R4578 S.n3332 S.n3331 0.004
R4579 S.n3179 S.n3178 0.004
R4580 S.n2813 S.n2812 0.004
R4581 S.n2646 S.n2645 0.004
R4582 S.n2157 S.n2156 0.004
R4583 S.n1842 S.n1841 0.004
R4584 S.n2320 S.n2319 0.004
R4585 S.n2661 S.n2660 0.004
R4586 S.n5067 S.n5066 0.004
R4587 S.n4940 S.n4939 0.004
R4588 S.n5771 S.n5770 0.004
R4589 S.n5571 S.n5570 0.004
R4590 S.n4747 S.n4746 0.004
R4591 S.n4592 S.n4591 0.004
R4592 S.n4314 S.n4313 0.004
R4593 S.n4157 S.n4156 0.004
R4594 S.n3725 S.n3724 0.004
R4595 S.n3871 S.n3870 0.004
R4596 S.n3348 S.n3347 0.004
R4597 S.n3194 S.n3193 0.004
R4598 S.n2669 S.n2668 0.004
R4599 S.n4607 S.n4606 0.004
R4600 S.n5083 S.n5082 0.004
R4601 S.n4925 S.n4924 0.004
R4602 S.n5787 S.n5786 0.004
R4603 S.n5586 S.n5585 0.004
R4604 S.n4763 S.n4762 0.004
R4605 S.n4174 S.n4173 0.004
R4606 S.n3744 S.n3743 0.004
R4607 S.n3888 S.n3887 0.004
R4608 S.n3388 S.n3387 0.004
R4609 S.n3397 S.n3396 0.004
R4610 S.n2832 S.n2831 0.004
R4611 S.n2868 S.n2867 0.004
R4612 S.n2933 S.n2932 0.004
R4613 S.n3367 S.n3366 0.004
R4614 S.n3901 S.n3900 0.004
R4615 S.n5099 S.n5098 0.004
R4616 S.n4910 S.n4909 0.004
R4617 S.n5803 S.n5802 0.004
R4618 S.n5601 S.n5600 0.004
R4619 S.n4779 S.n4778 0.004
R4620 S.n4622 S.n4621 0.004
R4621 S.n4330 S.n4329 0.004
R4622 S.n4187 S.n4186 0.004
R4623 S.n3757 S.n3756 0.004
R4624 S.n3448 S.n3447 0.004
R4625 S.n3775 S.n3774 0.004
R4626 S.n4202 S.n4201 0.004
R4627 S.n5115 S.n5114 0.004
R4628 S.n4895 S.n4894 0.004
R4629 S.n5819 S.n5818 0.004
R4630 S.n5616 S.n5615 0.004
R4631 S.n4795 S.n4794 0.004
R4632 S.n4637 S.n4636 0.004
R4633 S.n4210 S.n4209 0.004
R4634 S.n3954 S.n3953 0.004
R4635 S.n4349 S.n4348 0.004
R4636 S.n4652 S.n4651 0.004
R4637 S.n5131 S.n5130 0.004
R4638 S.n4880 S.n4879 0.004
R4639 S.n5835 S.n5834 0.004
R4640 S.n5631 S.n5630 0.004
R4641 S.n4660 S.n4659 0.004
R4642 S.n4425 S.n4424 0.004
R4643 S.n4812 S.n4811 0.004
R4644 S.n5868 S.n5867 0.004
R4645 S.n5150 S.n5149 0.004
R4646 S.n4867 S.n4866 0.004
R4647 S.n5855 S.n5854 0.004
R4648 S.n5173 S.n5172 0.004
R4649 S.n4371 S.n4370 0.004
R4650 S.t241 S.n576 0.004
R4651 S.n348 S.n347 0.004
R4652 S.n394 S.n393 0.004
R4653 S.n70 S.n69 0.004
R4654 S.n425 S.n424 0.004
R4655 S.n49 S.n48 0.004
R4656 S.n456 S.n455 0.004
R4657 S.n28 S.n27 0.004
R4658 S.t241 S.n624 0.004
R4659 S.n97 S.n82 0.004
R4660 S.n4227 S.n4226 0.004
R4661 S.n3973 S.n3972 0.004
R4662 S.n3499 S.n3498 0.004
R4663 S.n3013 S.n3012 0.004
R4664 S.n2475 S.n2474 0.004
R4665 S.n1983 S.n1982 0.004
R4666 S.n1436 S.n1435 0.004
R4667 S.n860 S.n859 0.004
R4668 S.n607 S.n606 0.004
R4669 S.n5045 S.n5044 0.004
R4670 S.n4227 S.n4225 0.004
R4671 S.n234 S.n222 0.004
R4672 S.n1133 S.n1132 0.004
R4673 S.n1690 S.n1678 0.004
R4674 S.n2286 S.n2274 0.004
R4675 S.n2782 S.n2770 0.004
R4676 S.n3301 S.n3289 0.004
R4677 S.n3678 S.n3666 0.004
R4678 S.n4267 S.n4255 0.004
R4679 S.n4700 S.n4688 0.004
R4680 S.n5669 S.n5667 0.004
R4681 S.n3619 S.n3618 0.004
R4682 S.n195 S.n186 0.004
R4683 S.n3225 S.n3223 0.004
R4684 S.n2687 S.n2686 0.004
R4685 S.n162 S.n153 0.004
R4686 S.n2174 S.n2172 0.004
R4687 S.n1559 S.n1558 0.004
R4688 S.n129 S.n120 0.004
R4689 S.n986 S.n984 0.004
R4690 S.n97 S.n96 0.004
R4691 S.n842 S.n841 0.004
R4692 S.n3455 S.n3454 0.004
R4693 S.n2969 S.n2968 0.004
R4694 S.n2431 S.n2430 0.004
R4695 S.n1939 S.n1938 0.004
R4696 S.n1390 S.n1389 0.004
R4697 S.n4681 S.n4664 0.004
R4698 S.n3981 S.n3979 0.004
R4699 S.n3507 S.n3505 0.004
R4700 S.n3021 S.n3019 0.004
R4701 S.n2483 S.n2481 0.004
R4702 S.n1991 S.n1989 0.004
R4703 S.n1444 S.n1442 0.004
R4704 S.n868 S.n866 0.004
R4705 S.n1092 S.n1091 0.004
R4706 S.n3591 S.n3590 0.004
R4707 S.n3619 S.n3603 0.004
R4708 S.n2567 S.n2566 0.004
R4709 S.n2687 S.n2671 0.004
R4710 S.n1531 S.n1530 0.004
R4711 S.n1559 S.n1543 0.004
R4712 S.n1242 S.n1228 0.004
R4713 S.n1809 S.n1242 0.004
R4714 S.n1828 S.n1814 0.004
R4715 S.n2359 S.n1828 0.004
R4716 S.n2900 S.n2899 0.004
R4717 S.n2899 S.n2885 0.004
R4718 S.n2919 S.n2905 0.004
R4719 S.n3415 S.n2919 0.004
R4720 S.n3434 S.n3420 0.004
R4721 S.n3921 S.n3434 0.004
R4722 S.n3940 S.n3926 0.004
R4723 S.n4402 S.n3940 0.004
R4724 S.n5646 S.n5644 0.004
R4725 S.n4411 S.n4410 0.004
R4726 S.n4856 S.n4406 0.004
R4727 S.t283 S.n5367 0.004
R4728 S.t283 S.n5375 0.004
R4729 S.t283 S.n5383 0.004
R4730 S.t283 S.n5391 0.004
R4731 S.t283 S.n5399 0.004
R4732 S.t283 S.n5407 0.004
R4733 S.t283 S.n5415 0.004
R4734 S.t283 S.n5420 0.004
R4735 S.t255 S.n100 0.004
R4736 S.t241 S.n650 0.004
R4737 S.t241 S.n647 0.004
R4738 S.t64 S.n5028 0.004
R4739 S.t241 S.n559 0.004
R4740 S.t12 S.n3228 0.004
R4741 S.t241 S.n662 0.004
R4742 S.t10 S.n3622 0.004
R4743 S.t241 S.n574 0.004
R4744 S.t57 S.n4230 0.004
R4745 S.t241 S.n621 0.004
R4746 S.t8 S.n4684 0.004
R4747 S.t4 S.n5672 0.004
R4748 S.t241 S.n638 0.004
R4749 S.t241 S.n547 0.004
R4750 S.t16 S.n2177 0.004
R4751 S.t241 S.n658 0.004
R4752 S.t0 S.n2690 0.004
R4753 S.t241 S.n535 0.004
R4754 S.t6 S.n989 0.004
R4755 S.t241 S.n654 0.004
R4756 S.t21 S.n1562 0.004
R4757 S.t241 S.n522 0.004
R4758 S.t283 S.n5441 0.004
R4759 S.t283 S.n5359 0.004
R4760 S.t283 S.n5369 0.004
R4761 S.t283 S.n5377 0.004
R4762 S.t283 S.n5385 0.004
R4763 S.t283 S.n5393 0.004
R4764 S.t283 S.n5401 0.004
R4765 S.t283 S.n5409 0.004
R4766 S.t283 S.n5417 0.004
R4767 S.t283 S.n5425 0.004
R4768 S.t283 S.n5347 0.004
R4769 S.t241 S.n645 0.004
R4770 S.t283 S.n5351 0.004
R4771 S.t35 S.n5265 0.004
R4772 S.t241 S.n400 0.004
R4773 S.t241 S.n431 0.004
R4774 S.t241 S.n462 0.004
R4775 S.t241 S.n466 0.004
R4776 S.n290 S.n289 0.004
R4777 S.t241 S.n642 0.004
R4778 S.t241 S.n551 0.004
R4779 S.t241 S.n539 0.004
R4780 S.t241 S.n526 0.004
R4781 S.n5669 S.n5668 0.004
R4782 S.n3637 S.n3626 0.004
R4783 S.n3260 S.n3249 0.004
R4784 S.n2741 S.n2730 0.004
R4785 S.n2245 S.n2234 0.004
R4786 S.n1649 S.n1638 0.004
R4787 S.n5021 S.n5020 0.003
R4788 S.n5260 S.n5259 0.003
R4789 S.n5717 S.n5716 0.003
R4790 S.n5880 S.n5879 0.003
R4791 S.n481 S.n480 0.003
R4792 S.n354 S.n353 0.003
R4793 S.n941 S.n940 0.003
R4794 S.n5242 S.n5241 0.003
R4795 S.n5693 S.n5692 0.003
R4796 S.n5490 S.n5489 0.003
R4797 S.n4725 S.n4724 0.003
R4798 S.n4477 S.n4476 0.003
R4799 S.n4292 S.n4291 0.003
R4800 S.n4040 S.n4039 0.003
R4801 S.n3703 S.n3702 0.003
R4802 S.n3566 S.n3565 0.003
R4803 S.n3326 S.n3325 0.003
R4804 S.n3080 S.n3079 0.003
R4805 S.n2807 S.n2806 0.003
R4806 S.n2542 S.n2541 0.003
R4807 S.n2311 S.n2310 0.003
R4808 S.n2050 S.n2049 0.003
R4809 S.n1715 S.n1714 0.003
R4810 S.n1506 S.n1505 0.003
R4811 S.n1156 S.n1155 0.003
R4812 S.n260 S.n259 0.003
R4813 S.n76 S.n75 0.003
R4814 S.n795 S.n794 0.003
R4815 S.n3103 S.n3102 0.003
R4816 S.n2711 S.n2710 0.003
R4817 S.n2395 S.n2394 0.003
R4818 S.n2215 S.n2214 0.003
R4819 S.n1903 S.n1902 0.003
R4820 S.n1619 S.n1618 0.003
R4821 S.n1353 S.n1352 0.003
R4822 S.n1059 S.n1058 0.003
R4823 S.n386 S.n385 0.003
R4824 S.n3594 S.n3593 0.003
R4825 S.n3247 S.n3246 0.003
R4826 S.n2962 S.n2961 0.003
R4827 S.n2728 S.n2727 0.003
R4828 S.n2424 S.n2423 0.003
R4829 S.n2232 S.n2231 0.003
R4830 S.n1932 S.n1931 0.003
R4831 S.n1636 S.n1635 0.003
R4832 S.n1382 S.n1381 0.003
R4833 S.n1078 S.n1077 0.003
R4834 S.n1098 S.n1097 0.003
R4835 S.n857 S.n856 0.003
R4836 S.n282 S.n281 0.003
R4837 S.n311 S.n310 0.003
R4838 S.n1417 S.n1416 0.003
R4839 S.n1964 S.n1963 0.003
R4840 S.n2456 S.n2455 0.003
R4841 S.n2994 S.n2993 0.003
R4842 S.n3480 S.n3479 0.003
R4843 S.n4066 S.n4065 0.003
R4844 S.n3643 S.n3642 0.003
R4845 S.n3266 S.n3265 0.003
R4846 S.n2747 S.n2746 0.003
R4847 S.n2251 S.n2250 0.003
R4848 S.n1655 S.n1654 0.003
R4849 S.n891 S.n890 0.003
R4850 S.n221 S.n220 0.003
R4851 S.n587 S.n586 0.003
R4852 S.n4501 S.n4500 0.003
R4853 S.n4253 S.n4252 0.003
R4854 S.n3988 S.n3987 0.003
R4855 S.n3664 S.n3663 0.003
R4856 S.n3514 S.n3513 0.003
R4857 S.n3287 S.n3286 0.003
R4858 S.n3028 S.n3027 0.003
R4859 S.n2768 S.n2767 0.003
R4860 S.n2490 S.n2489 0.003
R4861 S.n2272 S.n2271 0.003
R4862 S.n1998 S.n1997 0.003
R4863 S.n1676 S.n1675 0.003
R4864 S.n1451 S.n1450 0.003
R4865 S.n1119 S.n1118 0.003
R4866 S.n919 S.n918 0.003
R4867 S.n240 S.n239 0.003
R4868 S.n1139 S.n1138 0.003
R4869 S.n1472 S.n1471 0.003
R4870 S.n1696 S.n1695 0.003
R4871 S.n2018 S.n2017 0.003
R4872 S.n2292 S.n2291 0.003
R4873 S.n2510 S.n2509 0.003
R4874 S.n2788 S.n2787 0.003
R4875 S.n3048 S.n3047 0.003
R4876 S.n3307 S.n3306 0.003
R4877 S.n3534 S.n3533 0.003
R4878 S.n3684 S.n3683 0.003
R4879 S.n4008 S.n4007 0.003
R4880 S.n4273 S.n4272 0.003
R4881 S.n4445 S.n4444 0.003
R4882 S.n4706 S.n4705 0.003
R4883 S.n5512 S.n5511 0.003
R4884 S.n333 S.n332 0.003
R4885 S.n823 S.n822 0.003
R4886 S.n201 S.n200 0.003
R4887 S.n184 S.n183 0.003
R4888 S.n55 S.n54 0.003
R4889 S.n736 S.n735 0.003
R4890 S.n2073 S.n2072 0.003
R4891 S.n1583 S.n1582 0.003
R4892 S.n1290 S.n1289 0.003
R4893 S.n1025 S.n1024 0.003
R4894 S.n417 S.n416 0.003
R4895 S.n2570 S.n2569 0.003
R4896 S.n2196 S.n2195 0.003
R4897 S.n1871 S.n1870 0.003
R4898 S.n1600 S.n1599 0.003
R4899 S.n1319 S.n1318 0.003
R4900 S.n1042 S.n1041 0.003
R4901 S.n765 S.n764 0.003
R4902 S.n168 S.n167 0.003
R4903 S.n151 S.n150 0.003
R4904 S.n34 S.n33 0.003
R4905 S.n962 S.n961 0.003
R4906 S.n448 S.n447 0.003
R4907 S.n1534 S.n1533 0.003
R4908 S.n1008 S.n1007 0.003
R4909 S.n706 S.n705 0.003
R4910 S.n135 S.n134 0.003
R4911 S.n118 S.n117 0.003
R4912 S.n381 S.n380 0.003
R4913 S.n276 S.n275 0.003
R4914 S.n1198 S.n1197 0.003
R4915 S.n1176 S.n1175 0.003
R4916 S.n1766 S.n1765 0.003
R4917 S.n1739 S.n1738 0.003
R4918 S.n2110 S.n2109 0.003
R4919 S.n2083 S.n2082 0.003
R4920 S.n2607 S.n2606 0.003
R4921 S.n2580 S.n2579 0.003
R4922 S.n3140 S.n3139 0.003
R4923 S.n3113 S.n3112 0.003
R4924 S.n3817 S.n3816 0.003
R4925 S.n3790 S.n3789 0.003
R4926 S.n4103 S.n4102 0.003
R4927 S.n4076 S.n4075 0.003
R4928 S.n4538 S.n4537 0.003
R4929 S.n4511 S.n4510 0.003
R4930 S.n5532 S.n5531 0.003
R4931 S.n5732 S.n5731 0.003
R4932 S.n5214 S.n5213 0.003
R4933 S.n5184 S.n5183 0.003
R4934 S.n1204 S.n1203 0.003
R4935 S.n1170 S.n1169 0.003
R4936 S.n1796 S.n1795 0.003
R4937 S.n4984 S.n4983 0.003
R4938 S.n4996 S.n4995 0.003
R4939 S.n5747 S.n5746 0.003
R4940 S.n5548 S.n5547 0.003
R4941 S.n4560 S.n4559 0.003
R4942 S.n4569 S.n4568 0.003
R4943 S.n4125 S.n4124 0.003
R4944 S.n4134 S.n4133 0.003
R4945 S.n3839 S.n3838 0.003
R4946 S.n3848 S.n3847 0.003
R4947 S.n3162 S.n3161 0.003
R4948 S.n3171 S.n3170 0.003
R4949 S.n2629 S.n2628 0.003
R4950 S.n2638 S.n2637 0.003
R4951 S.n2135 S.n2134 0.003
R4952 S.n2121 S.n2120 0.003
R4953 S.n1788 S.n1787 0.003
R4954 S.n1804 S.n1803 0.003
R4955 S.n1733 S.n1732 0.003
R4956 S.n2346 S.n2345 0.003
R4957 S.n5059 S.n5058 0.003
R4958 S.n4965 S.n4964 0.003
R4959 S.n5763 S.n5762 0.003
R4960 S.n5563 S.n5562 0.003
R4961 S.n4739 S.n4738 0.003
R4962 S.n4584 S.n4583 0.003
R4963 S.n4306 S.n4305 0.003
R4964 S.n4149 S.n4148 0.003
R4965 S.n3717 S.n3716 0.003
R4966 S.n3863 S.n3862 0.003
R4967 S.n3340 S.n3339 0.003
R4968 S.n3186 S.n3185 0.003
R4969 S.n2821 S.n2820 0.003
R4970 S.n2653 S.n2652 0.003
R4971 S.n2338 S.n2337 0.003
R4972 S.n2354 S.n2353 0.003
R4973 S.n2329 S.n2328 0.003
R4974 S.n2858 S.n2857 0.003
R4975 S.n5075 S.n5074 0.003
R4976 S.n4950 S.n4949 0.003
R4977 S.n5779 S.n5778 0.003
R4978 S.n5578 S.n5577 0.003
R4979 S.n4755 S.n4754 0.003
R4980 S.n4599 S.n4598 0.003
R4981 S.n4322 S.n4321 0.003
R4982 S.n4164 S.n4163 0.003
R4983 S.n3733 S.n3732 0.003
R4984 S.n3878 S.n3877 0.003
R4985 S.n3356 S.n3355 0.003
R4986 S.n3201 S.n3200 0.003
R4987 S.n2850 S.n2849 0.003
R4988 S.n4614 S.n4613 0.003
R4989 S.n5091 S.n5090 0.003
R4990 S.n4935 S.n4934 0.003
R4991 S.n5795 S.n5794 0.003
R4992 S.n5593 S.n5592 0.003
R4993 S.n4771 S.n4770 0.003
R4994 S.n4179 S.n4178 0.003
R4995 S.n3749 S.n3748 0.003
R4996 S.n3893 S.n3892 0.003
R4997 S.n3382 S.n3381 0.003
R4998 S.n3402 S.n3401 0.003
R4999 S.n2841 S.n2840 0.003
R5000 S.n2864 S.n2863 0.003
R5001 S.n3410 S.n3409 0.003
R5002 S.n3376 S.n3375 0.003
R5003 S.n3908 S.n3907 0.003
R5004 S.n5107 S.n5106 0.003
R5005 S.n4920 S.n4919 0.003
R5006 S.n5811 S.n5810 0.003
R5007 S.n5608 S.n5607 0.003
R5008 S.n4787 S.n4786 0.003
R5009 S.n4629 S.n4628 0.003
R5010 S.n4338 S.n4337 0.003
R5011 S.n4194 S.n4193 0.003
R5012 S.n3764 S.n3763 0.003
R5013 S.n3916 S.n3915 0.003
R5014 S.n3784 S.n3783 0.003
R5015 S.n4389 S.n4388 0.003
R5016 S.n5123 S.n5122 0.003
R5017 S.n4905 S.n4904 0.003
R5018 S.n5827 S.n5826 0.003
R5019 S.n5623 S.n5622 0.003
R5020 S.n4803 S.n4802 0.003
R5021 S.n4644 S.n4643 0.003
R5022 S.n4381 S.n4380 0.003
R5023 S.n4397 S.n4396 0.003
R5024 S.n4358 S.n4357 0.003
R5025 S.n4843 S.n4842 0.003
R5026 S.n5139 S.n5138 0.003
R5027 S.n4890 S.n4889 0.003
R5028 S.n5843 S.n5842 0.003
R5029 S.n5638 S.n5637 0.003
R5030 S.n4835 S.n4834 0.003
R5031 S.n4851 S.n4850 0.003
R5032 S.n4826 S.n4825 0.003
R5033 S.n5874 S.n5873 0.003
R5034 S.n5155 S.n5154 0.003
R5035 S.n4875 S.n4874 0.003
R5036 S.n5849 S.n5848 0.003
R5037 S.n5178 S.n5177 0.003
R5038 S.n1072 S.n1071 0.003
R5039 S.n5018 S.n5013 0.003
R5040 S.n5257 S.n5252 0.003
R5041 S.n5711 S.n5699 0.003
R5042 S.n494 S.n478 0.003
R5043 S.n348 S.n343 0.003
R5044 S.n935 S.n927 0.003
R5045 S.n5236 S.n5224 0.003
R5046 S.n5687 S.n5682 0.003
R5047 S.n5484 S.n5475 0.003
R5048 S.n4719 S.n4714 0.003
R5049 S.n4471 S.n4462 0.003
R5050 S.n4286 S.n4281 0.003
R5051 S.n4034 S.n4025 0.003
R5052 S.n3697 S.n3692 0.003
R5053 S.n3560 S.n3551 0.003
R5054 S.n3323 S.n3318 0.003
R5055 S.n3074 S.n3065 0.003
R5056 S.n2801 S.n2796 0.003
R5057 S.n2536 S.n2527 0.003
R5058 S.n2305 S.n2300 0.003
R5059 S.n2044 S.n2035 0.003
R5060 S.n1709 S.n1704 0.003
R5061 S.n1500 S.n1489 0.003
R5062 S.n1150 S.n1147 0.003
R5063 S.n254 S.n249 0.003
R5064 S.n70 S.n65 0.003
R5065 S.n789 S.n782 0.003
R5066 S.n3100 S.n3089 0.003
R5067 S.n2705 S.n2700 0.003
R5068 S.n2389 S.n2380 0.003
R5069 S.n2209 S.n2204 0.003
R5070 S.n1897 S.n1888 0.003
R5071 S.n1613 S.n1608 0.003
R5072 S.n1347 S.n1336 0.003
R5073 S.n1053 S.n1050 0.003
R5074 S.n394 S.n13 0.003
R5075 S.n3591 S.n3579 0.003
R5076 S.n3241 S.n3236 0.003
R5077 S.n2956 S.n2942 0.003
R5078 S.n2722 S.n2717 0.003
R5079 S.n2418 S.n2404 0.003
R5080 S.n2226 S.n2221 0.003
R5081 S.n1926 S.n1912 0.003
R5082 S.n1630 S.n1625 0.003
R5083 S.n1376 S.n1362 0.003
R5084 S.n1072 S.n1065 0.003
R5085 S.n1092 S.n1084 0.003
R5086 S.n851 S.n833 0.003
R5087 S.n290 S.n80 0.003
R5088 S.n305 S.n296 0.003
R5089 S.n1411 S.n1400 0.003
R5090 S.n1958 S.n1949 0.003
R5091 S.n2450 S.n2441 0.003
R5092 S.n2988 S.n2979 0.003
R5093 S.n3474 S.n3465 0.003
R5094 S.n4063 S.n4052 0.003
R5095 S.n3637 S.n3632 0.003
R5096 S.n3260 S.n3255 0.003
R5097 S.n2741 S.n2736 0.003
R5098 S.n2245 S.n2240 0.003
R5099 S.n1649 S.n1644 0.003
R5100 S.n885 S.n872 0.003
R5101 S.n215 S.n206 0.003
R5102 S.n600 S.n584 0.003
R5103 S.n4498 S.n4493 0.003
R5104 S.n4247 S.n4245 0.003
R5105 S.n3982 S.n3970 0.003
R5106 S.n3658 S.n3656 0.003
R5107 S.n3508 S.n3496 0.003
R5108 S.n3281 S.n3279 0.003
R5109 S.n3022 S.n3010 0.003
R5110 S.n2762 S.n2760 0.003
R5111 S.n2484 S.n2472 0.003
R5112 S.n2266 S.n2264 0.003
R5113 S.n1992 S.n1980 0.003
R5114 S.n1670 S.n1668 0.003
R5115 S.n1445 S.n1433 0.003
R5116 S.n1113 S.n1111 0.003
R5117 S.n913 S.n900 0.003
R5118 S.n234 S.n226 0.003
R5119 S.n1133 S.n1130 0.003
R5120 S.n1466 S.n1460 0.003
R5121 S.n1690 S.n1682 0.003
R5122 S.n2012 S.n2007 0.003
R5123 S.n2286 S.n2278 0.003
R5124 S.n2504 S.n2499 0.003
R5125 S.n2782 S.n2774 0.003
R5126 S.n3042 S.n3037 0.003
R5127 S.n3301 S.n3293 0.003
R5128 S.n3528 S.n3523 0.003
R5129 S.n3678 S.n3670 0.003
R5130 S.n4002 S.n3997 0.003
R5131 S.n4267 S.n4259 0.003
R5132 S.n4439 S.n4434 0.003
R5133 S.n4700 S.n4692 0.003
R5134 S.n5509 S.n5504 0.003
R5135 S.n327 S.n316 0.003
R5136 S.n817 S.n804 0.003
R5137 S.n195 S.n190 0.003
R5138 S.n178 S.n173 0.003
R5139 S.n49 S.n44 0.003
R5140 S.n730 S.n723 0.003
R5141 S.n2070 S.n2059 0.003
R5142 S.n1577 S.n1572 0.003
R5143 S.n1284 S.n1273 0.003
R5144 S.n1019 S.n1016 0.003
R5145 S.n425 S.n414 0.003
R5146 S.n2567 S.n2555 0.003
R5147 S.n2190 S.n2185 0.003
R5148 S.n1865 S.n1851 0.003
R5149 S.n1594 S.n1589 0.003
R5150 S.n1313 S.n1299 0.003
R5151 S.n1036 S.n1031 0.003
R5152 S.n759 S.n745 0.003
R5153 S.n162 S.n157 0.003
R5154 S.n145 S.n140 0.003
R5155 S.n28 S.n23 0.003
R5156 S.n959 S.n950 0.003
R5157 S.n456 S.n445 0.003
R5158 S.n1531 S.n1519 0.003
R5159 S.n1002 S.n997 0.003
R5160 S.n700 S.n686 0.003
R5161 S.n129 S.n124 0.003
R5162 S.n112 S.n107 0.003
R5163 S.n273 S.n266 0.003
R5164 S.n1195 S.n1190 0.003
R5165 S.n1186 S.n969 0.003
R5166 S.n1763 S.n1754 0.003
R5167 S.n1749 S.n1541 0.003
R5168 S.n2107 S.n2098 0.003
R5169 S.n2093 S.n2080 0.003
R5170 S.n2604 S.n2595 0.003
R5171 S.n2590 S.n2577 0.003
R5172 S.n3137 S.n3128 0.003
R5173 S.n3123 S.n3110 0.003
R5174 S.n3814 S.n3805 0.003
R5175 S.n3800 S.n3601 0.003
R5176 S.n4100 S.n4091 0.003
R5177 S.n4086 S.n4073 0.003
R5178 S.n4535 S.n4526 0.003
R5179 S.n4521 S.n4508 0.003
R5180 S.n5529 S.n5520 0.003
R5181 S.n5729 S.n5722 0.003
R5182 S.n5208 S.n5199 0.003
R5183 S.n5194 S.n5000 0.003
R5184 S.n1167 S.n1162 0.003
R5185 S.n1793 S.n1777 0.003
R5186 S.n4988 S.n4987 0.003
R5187 S.n4990 S.n4973 0.003
R5188 S.n5744 S.n5743 0.003
R5189 S.n5545 S.n5543 0.003
R5190 S.n4564 S.n4563 0.003
R5191 S.n4566 S.n4549 0.003
R5192 S.n4129 S.n4128 0.003
R5193 S.n4131 S.n4114 0.003
R5194 S.n3843 S.n3842 0.003
R5195 S.n3845 S.n3828 0.003
R5196 S.n3166 S.n3165 0.003
R5197 S.n3168 S.n3151 0.003
R5198 S.n2633 S.n2632 0.003
R5199 S.n2635 S.n2618 0.003
R5200 S.n2139 S.n2138 0.003
R5201 S.n2141 S.n2124 0.003
R5202 S.n1792 S.n1791 0.003
R5203 S.n1730 S.n1721 0.003
R5204 S.n2343 S.n2152 0.003
R5205 S.n5056 S.n5054 0.003
R5206 S.n4959 S.n4958 0.003
R5207 S.n5760 S.n5758 0.003
R5208 S.n5560 S.n5559 0.003
R5209 S.n4736 S.n4734 0.003
R5210 S.n4581 S.n4580 0.003
R5211 S.n4303 S.n4301 0.003
R5212 S.n4146 S.n4145 0.003
R5213 S.n3714 S.n3712 0.003
R5214 S.n3860 S.n3859 0.003
R5215 S.n3337 S.n3335 0.003
R5216 S.n3183 S.n3182 0.003
R5217 S.n2818 S.n2816 0.003
R5218 S.n2650 S.n2649 0.003
R5219 S.n2342 S.n2341 0.003
R5220 S.n2326 S.n2317 0.003
R5221 S.n2855 S.n2664 0.003
R5222 S.n5072 S.n5070 0.003
R5223 S.n4944 S.n4943 0.003
R5224 S.n5776 S.n5774 0.003
R5225 S.n5575 S.n5574 0.003
R5226 S.n4752 S.n4750 0.003
R5227 S.n4596 S.n4595 0.003
R5228 S.n4319 S.n4317 0.003
R5229 S.n4161 S.n4160 0.003
R5230 S.n3730 S.n3728 0.003
R5231 S.n3875 S.n3874 0.003
R5232 S.n3353 S.n3351 0.003
R5233 S.n3198 S.n3197 0.003
R5234 S.n2854 S.n2853 0.003
R5235 S.n4611 S.n4610 0.003
R5236 S.n5088 S.n5086 0.003
R5237 S.n4929 S.n4928 0.003
R5238 S.n5792 S.n5790 0.003
R5239 S.n5590 S.n5589 0.003
R5240 S.n4768 S.n4766 0.003
R5241 S.n4176 S.n4171 0.003
R5242 S.n3746 S.n3741 0.003
R5243 S.n3890 S.n3885 0.003
R5244 S.n3390 S.n3208 0.003
R5245 S.n3399 S.n3394 0.003
R5246 S.n2838 S.n2829 0.003
R5247 S.n3373 S.n3364 0.003
R5248 S.n3905 S.n3904 0.003
R5249 S.n5104 S.n5102 0.003
R5250 S.n4914 S.n4913 0.003
R5251 S.n5808 S.n5806 0.003
R5252 S.n5605 S.n5604 0.003
R5253 S.n4784 S.n4782 0.003
R5254 S.n4626 S.n4625 0.003
R5255 S.n4335 S.n4333 0.003
R5256 S.n4191 S.n4190 0.003
R5257 S.n3761 S.n3760 0.003
R5258 S.n3781 S.n3772 0.003
R5259 S.n4386 S.n4205 0.003
R5260 S.n5120 S.n5118 0.003
R5261 S.n4899 S.n4898 0.003
R5262 S.n5824 S.n5822 0.003
R5263 S.n5620 S.n5619 0.003
R5264 S.n4800 S.n4798 0.003
R5265 S.n4641 S.n4640 0.003
R5266 S.n4385 S.n4384 0.003
R5267 S.n4355 S.n4346 0.003
R5268 S.n4840 S.n4655 0.003
R5269 S.n5136 S.n5134 0.003
R5270 S.n4884 S.n4883 0.003
R5271 S.n5840 S.n5838 0.003
R5272 S.n5635 S.n5634 0.003
R5273 S.n4839 S.n4838 0.003
R5274 S.n4823 S.n4809 0.003
R5275 S.n5871 S.n5865 0.003
R5276 S.n5152 S.n5147 0.003
R5277 S.n4869 S.n4864 0.003
R5278 S.n5857 S.n5650 0.003
R5279 S.n5175 S.n5170 0.003
R5280 S.n378 S.n371 0.003
R5281 S.n4 S.n2 0.003
R5282 S.n405 S.n403 0.003
R5283 S.n436 S.n434 0.003
R5284 S.n500 S.n498 0.003
R5285 S.n5445 S.n5444 0.003
R5286 S.n5445 S.n5289 0.003
R5287 S.n4681 S.n4680 0.003
R5288 S.n491 S.n490 0.003
R5289 S.n4372 S.n4363 0.003
R5290 S.n4372 S.n4365 0.003
R5291 S.n303 S.n302 0.003
R5292 S.n4666 S.n4665 0.003
R5293 S.n3982 S.n3981 0.003
R5294 S.n3508 S.n3507 0.003
R5295 S.n3022 S.n3021 0.003
R5296 S.n2484 S.n2483 0.003
R5297 S.n1992 S.n1991 0.003
R5298 S.n1445 S.n1444 0.003
R5299 S.n885 S.n868 0.003
R5300 S.n5857 S.n5646 0.003
R5301 S.n5280 S.n5279 0.003
R5302 S.t283 S.n5291 0.003
R5303 S.n5045 S.n5030 0.003
R5304 S.n3225 S.n3224 0.003
R5305 S.n2174 S.n2173 0.003
R5306 S.n986 S.n985 0.003
R5307 S.n5500 S.n5499 0.003
R5308 S.n3241 S.n3232 0.003
R5309 S.n2722 S.n2713 0.003
R5310 S.n2226 S.n2217 0.003
R5311 S.n1630 S.n1621 0.003
R5312 S.n1072 S.n1061 0.003
R5313 S.n2190 S.n2181 0.003
R5314 S.n1594 S.n1585 0.003
R5315 S.n1036 S.n1027 0.003
R5316 S.n1002 S.n993 0.003
R5317 S.n5257 S.n5248 0.003
R5318 S.t283 S.n5344 0.003
R5319 S.t283 S.n5427 0.003
R5320 S.n953 S.n952 0.003
R5321 S.n339 S.n338 0.003
R5322 S.n613 S.n612 0.003
R5323 S.n395 S.n394 0.002
R5324 S.n195 S.n187 0.002
R5325 S.n817 S.n796 0.002
R5326 S.n1072 S.n1062 0.002
R5327 S.n1376 S.n1359 0.002
R5328 S.n1630 S.n1622 0.002
R5329 S.n1926 S.n1909 0.002
R5330 S.n2226 S.n2218 0.002
R5331 S.n2418 S.n2401 0.002
R5332 S.n2722 S.n2714 0.002
R5333 S.n2956 S.n2939 0.002
R5334 S.n3241 S.n3233 0.002
R5335 S.n601 S.n600 0.002
R5336 S.n215 S.n203 0.002
R5337 S.n885 S.n869 0.002
R5338 S.n1113 S.n1099 0.002
R5339 S.n1445 S.n1418 0.002
R5340 S.n1670 S.n1656 0.002
R5341 S.n1992 S.n1965 0.002
R5342 S.n2266 S.n2252 0.002
R5343 S.n2484 S.n2457 0.002
R5344 S.n2762 S.n2748 0.002
R5345 S.n3022 S.n2995 0.002
R5346 S.n3281 S.n3267 0.002
R5347 S.n3508 S.n3481 0.002
R5348 S.n3658 S.n3644 0.002
R5349 S.n3982 S.n3955 0.002
R5350 S.n4247 S.n4233 0.002
R5351 S.n4700 S.n4689 0.002
R5352 S.n4439 S.n4431 0.002
R5353 S.n4267 S.n4256 0.002
R5354 S.n4002 S.n3994 0.002
R5355 S.n3678 S.n3667 0.002
R5356 S.n3528 S.n3520 0.002
R5357 S.n3301 S.n3290 0.002
R5358 S.n3042 S.n3034 0.002
R5359 S.n2782 S.n2771 0.002
R5360 S.n2504 S.n2496 0.002
R5361 S.n2286 S.n2275 0.002
R5362 S.n2012 S.n2004 0.002
R5363 S.n1690 S.n1679 0.002
R5364 S.n1466 S.n1457 0.002
R5365 S.n1133 S.n1120 0.002
R5366 S.n913 S.n897 0.002
R5367 S.n234 S.n223 0.002
R5368 S.n426 S.n425 0.002
R5369 S.n162 S.n154 0.002
R5370 S.n759 S.n737 0.002
R5371 S.n1036 S.n1028 0.002
R5372 S.n1313 S.n1296 0.002
R5373 S.n1594 S.n1586 0.002
R5374 S.n1865 S.n1848 0.002
R5375 S.n2190 S.n2182 0.002
R5376 S.n457 S.n456 0.002
R5377 S.n129 S.n121 0.002
R5378 S.n700 S.n678 0.002
R5379 S.n1002 S.n994 0.002
R5380 S.n5194 S.n4997 0.002
R5381 S.n5208 S.n5196 0.002
R5382 S.n5729 S.n5719 0.002
R5383 S.n5529 S.n5517 0.002
R5384 S.n4521 S.n4505 0.002
R5385 S.n4535 S.n4523 0.002
R5386 S.n4086 S.n4070 0.002
R5387 S.n4100 S.n4088 0.002
R5388 S.n3800 S.n3598 0.002
R5389 S.n3814 S.n3802 0.002
R5390 S.n3123 S.n3107 0.002
R5391 S.n3137 S.n3125 0.002
R5392 S.n2590 S.n2574 0.002
R5393 S.n2604 S.n2592 0.002
R5394 S.n2093 S.n2077 0.002
R5395 S.n2107 S.n2095 0.002
R5396 S.n1749 S.n1538 0.002
R5397 S.n1763 S.n1751 0.002
R5398 S.n1186 S.n966 0.002
R5399 S.n1195 S.n1187 0.002
R5400 S.n4988 S.n4974 0.002
R5401 S.n4990 S.n4966 0.002
R5402 S.n5744 S.n5736 0.002
R5403 S.n5545 S.n5536 0.002
R5404 S.n4564 S.n4550 0.002
R5405 S.n4566 S.n4542 0.002
R5406 S.n4129 S.n4115 0.002
R5407 S.n4131 S.n4107 0.002
R5408 S.n3843 S.n3829 0.002
R5409 S.n3845 S.n3821 0.002
R5410 S.n3166 S.n3152 0.002
R5411 S.n3168 S.n3144 0.002
R5412 S.n2633 S.n2619 0.002
R5413 S.n2635 S.n2611 0.002
R5414 S.n2139 S.n2125 0.002
R5415 S.n2141 S.n2114 0.002
R5416 S.n1792 S.n1778 0.002
R5417 S.n1793 S.n1770 0.002
R5418 S.n1167 S.n1159 0.002
R5419 S.n5056 S.n5047 0.002
R5420 S.n4959 S.n4951 0.002
R5421 S.n5760 S.n5751 0.002
R5422 S.n5560 S.n5552 0.002
R5423 S.n4736 S.n4727 0.002
R5424 S.n4581 S.n4573 0.002
R5425 S.n4303 S.n4294 0.002
R5426 S.n4146 S.n4138 0.002
R5427 S.n3714 S.n3705 0.002
R5428 S.n3860 S.n3852 0.002
R5429 S.n3337 S.n3328 0.002
R5430 S.n3183 S.n3175 0.002
R5431 S.n2818 S.n2809 0.002
R5432 S.n2650 S.n2642 0.002
R5433 S.n2342 S.n2153 0.002
R5434 S.n2343 S.n2145 0.002
R5435 S.n1730 S.n1718 0.002
R5436 S.n5072 S.n5063 0.002
R5437 S.n4944 S.n4936 0.002
R5438 S.n5776 S.n5767 0.002
R5439 S.n5575 S.n5567 0.002
R5440 S.n4752 S.n4743 0.002
R5441 S.n4596 S.n4588 0.002
R5442 S.n4319 S.n4310 0.002
R5443 S.n4161 S.n4153 0.002
R5444 S.n3730 S.n3721 0.002
R5445 S.n3875 S.n3867 0.002
R5446 S.n3353 S.n3344 0.002
R5447 S.n3198 S.n3190 0.002
R5448 S.n2854 S.n2665 0.002
R5449 S.n2855 S.n2657 0.002
R5450 S.n2326 S.n2314 0.002
R5451 S.n5088 S.n5079 0.002
R5452 S.n4929 S.n4921 0.002
R5453 S.n5792 S.n5783 0.002
R5454 S.n5590 S.n5582 0.002
R5455 S.n4768 S.n4759 0.002
R5456 S.n4611 S.n4603 0.002
R5457 S.n4372 S.n4367 0.002
R5458 S.n4176 S.n4168 0.002
R5459 S.n3746 S.n3738 0.002
R5460 S.n3890 S.n3882 0.002
R5461 S.n3390 S.n3205 0.002
R5462 S.n3399 S.n3391 0.002
R5463 S.n2838 S.n2826 0.002
R5464 S.n5104 S.n5095 0.002
R5465 S.n4914 S.n4906 0.002
R5466 S.n5808 S.n5799 0.002
R5467 S.n5605 S.n5597 0.002
R5468 S.n4784 S.n4775 0.002
R5469 S.n4626 S.n4618 0.002
R5470 S.n4335 S.n4326 0.002
R5471 S.n4191 S.n4183 0.002
R5472 S.n3761 S.n3753 0.002
R5473 S.n3905 S.n3897 0.002
R5474 S.n3373 S.n3361 0.002
R5475 S.n5120 S.n5111 0.002
R5476 S.n4899 S.n4891 0.002
R5477 S.n5824 S.n5815 0.002
R5478 S.n5620 S.n5612 0.002
R5479 S.n4800 S.n4791 0.002
R5480 S.n4641 S.n4633 0.002
R5481 S.n4385 S.n4206 0.002
R5482 S.n4386 S.n4198 0.002
R5483 S.n3781 S.n3769 0.002
R5484 S.n5136 S.n5127 0.002
R5485 S.n4884 S.n4876 0.002
R5486 S.n5840 S.n5831 0.002
R5487 S.n5635 S.n5627 0.002
R5488 S.n4839 S.n4656 0.002
R5489 S.n4840 S.n4648 0.002
R5490 S.n4355 S.n4343 0.002
R5491 S.n5857 S.n5647 0.002
R5492 S.n4869 S.n4861 0.002
R5493 S.n5152 S.n5144 0.002
R5494 S.n4823 S.n4813 0.002
R5495 S.n5871 S.n5862 0.002
R5496 S.n5711 S.n5696 0.002
R5497 S.n5257 S.n5249 0.002
R5498 S.n5018 S.n5010 0.002
R5499 S.n495 S.n494 0.002
R5500 S.n3591 S.n3576 0.002
R5501 S.n4498 S.n4479 0.002
R5502 S.n5509 S.n5501 0.002
R5503 S.n2567 S.n2552 0.002
R5504 S.n1531 S.n1516 0.002
R5505 S.n1241 S.n1240 0.002
R5506 S.n1827 S.n1826 0.002
R5507 S.n2898 S.n2897 0.002
R5508 S.n2918 S.n2917 0.002
R5509 S.n3433 S.n3432 0.002
R5510 S.n3939 S.n3938 0.002
R5511 S.n5161 S.n5160 0.002
R5512 S.n5004 S.n5003 0.002
R5513 S.n5320 S.n5319 0.002
R5514 S.n5323 S.n5322 0.002
R5515 S.n5326 S.n5325 0.002
R5516 S.n5329 S.n5328 0.002
R5517 S.n5332 S.n5331 0.002
R5518 S.n5335 S.n5334 0.002
R5519 S.n5338 S.n5337 0.002
R5520 S.n5341 S.n5340 0.002
R5521 S.t241 S.n636 0.002
R5522 S.n1195 S.n1194 0.002
R5523 S.n475 S.n474 0.002
R5524 S.n5230 S.n5229 0.002
R5525 S.n4057 S.n4056 0.002
R5526 S.n3094 S.n3093 0.002
R5527 S.n2064 S.n2063 0.002
R5528 S.n935 S.n921 0.002
R5529 S.n789 S.n776 0.002
R5530 S.n1376 S.n1375 0.002
R5531 S.n1630 S.n1629 0.002
R5532 S.n1926 S.n1925 0.002
R5533 S.n2226 S.n2225 0.002
R5534 S.n2418 S.n2417 0.002
R5535 S.n2722 S.n2721 0.002
R5536 S.n2956 S.n2955 0.002
R5537 S.n3241 S.n3240 0.002
R5538 S.n730 S.n717 0.002
R5539 S.n1036 S.n1035 0.002
R5540 S.n1313 S.n1312 0.002
R5541 S.n1594 S.n1593 0.002
R5542 S.n1865 S.n1864 0.002
R5543 S.n2190 S.n2189 0.002
R5544 S.n1002 S.n1001 0.002
R5545 S.n1793 S.n1771 0.002
R5546 S.n2343 S.n2146 0.002
R5547 S.n2855 S.n2658 0.002
R5548 S.n4611 S.n4604 0.002
R5549 S.n2838 S.n2837 0.002
R5550 S.n3399 S.n3398 0.002
R5551 S.n3390 S.n3389 0.002
R5552 S.n3890 S.n3889 0.002
R5553 S.n3746 S.n3745 0.002
R5554 S.n4176 S.n4175 0.002
R5555 S.n4372 S.n4366 0.002
R5556 S.n3905 S.n3898 0.002
R5557 S.n4386 S.n4199 0.002
R5558 S.n4840 S.n4649 0.002
R5559 S.n5857 S.n5856 0.002
R5560 S.n4869 S.n4868 0.002
R5561 S.n5152 S.n5151 0.002
R5562 S.n5711 S.n5710 0.002
R5563 S.n5257 S.n5256 0.002
R5564 S.n5018 S.n5017 0.002
R5565 S.n3575 S.n3574 0.002
R5566 S.n2551 S.n2550 0.002
R5567 S.n1515 S.n1514 0.002
R5568 S.n5687 S.n5676 0.002
R5569 S.n5484 S.n5469 0.002
R5570 S.n4719 S.n4708 0.002
R5571 S.n4471 S.n4456 0.002
R5572 S.n4286 S.n4275 0.002
R5573 S.n4034 S.n4019 0.002
R5574 S.n3697 S.n3686 0.002
R5575 S.n3560 S.n3545 0.002
R5576 S.n3323 S.n3312 0.002
R5577 S.n3074 S.n3059 0.002
R5578 S.n2801 S.n2790 0.002
R5579 S.n2536 S.n2521 0.002
R5580 S.n2305 S.n2294 0.002
R5581 S.n2044 S.n2029 0.002
R5582 S.n1709 S.n1698 0.002
R5583 S.n1500 S.n1483 0.002
R5584 S.n1150 S.n1141 0.002
R5585 S.n254 S.n253 0.002
R5586 S.n2705 S.n2694 0.002
R5587 S.n2389 S.n2374 0.002
R5588 S.n2209 S.n2198 0.002
R5589 S.n1897 S.n1882 0.002
R5590 S.n1613 S.n1602 0.002
R5591 S.n1347 S.n1330 0.002
R5592 S.n1053 S.n1044 0.002
R5593 S.n817 S.n816 0.002
R5594 S.n195 S.n194 0.002
R5595 S.n178 S.n177 0.002
R5596 S.n1577 S.n1566 0.002
R5597 S.n1284 S.n1267 0.002
R5598 S.n1019 S.n1010 0.002
R5599 S.n759 S.n758 0.002
R5600 S.n162 S.n161 0.002
R5601 S.n145 S.n144 0.002
R5602 S.n700 S.n699 0.002
R5603 S.n129 S.n128 0.002
R5604 S.n112 S.n111 0.002
R5605 S.n4988 S.n4975 0.002
R5606 S.n4990 S.n4967 0.002
R5607 S.n5744 S.n5737 0.002
R5608 S.n5545 S.n5537 0.002
R5609 S.n4564 S.n4551 0.002
R5610 S.n4566 S.n4543 0.002
R5611 S.n4129 S.n4116 0.002
R5612 S.n4131 S.n4108 0.002
R5613 S.n3843 S.n3830 0.002
R5614 S.n3845 S.n3822 0.002
R5615 S.n3166 S.n3153 0.002
R5616 S.n3168 S.n3145 0.002
R5617 S.n2633 S.n2620 0.002
R5618 S.n2635 S.n2612 0.002
R5619 S.n2139 S.n2126 0.002
R5620 S.n2141 S.n2115 0.002
R5621 S.n1792 S.n1779 0.002
R5622 S.n1167 S.n1166 0.002
R5623 S.n5056 S.n5048 0.002
R5624 S.n4959 S.n4952 0.002
R5625 S.n5760 S.n5752 0.002
R5626 S.n5560 S.n5553 0.002
R5627 S.n4736 S.n4728 0.002
R5628 S.n4581 S.n4574 0.002
R5629 S.n4303 S.n4295 0.002
R5630 S.n4146 S.n4139 0.002
R5631 S.n3714 S.n3706 0.002
R5632 S.n3860 S.n3853 0.002
R5633 S.n3337 S.n3329 0.002
R5634 S.n3183 S.n3176 0.002
R5635 S.n2818 S.n2810 0.002
R5636 S.n2650 S.n2643 0.002
R5637 S.n2342 S.n2154 0.002
R5638 S.n1730 S.n1729 0.002
R5639 S.n5072 S.n5064 0.002
R5640 S.n4944 S.n4937 0.002
R5641 S.n5776 S.n5768 0.002
R5642 S.n5575 S.n5568 0.002
R5643 S.n4752 S.n4744 0.002
R5644 S.n4596 S.n4589 0.002
R5645 S.n4319 S.n4311 0.002
R5646 S.n4161 S.n4154 0.002
R5647 S.n3730 S.n3722 0.002
R5648 S.n3875 S.n3868 0.002
R5649 S.n3353 S.n3345 0.002
R5650 S.n3198 S.n3191 0.002
R5651 S.n2854 S.n2666 0.002
R5652 S.n2326 S.n2325 0.002
R5653 S.n5088 S.n5080 0.002
R5654 S.n4929 S.n4922 0.002
R5655 S.n5792 S.n5784 0.002
R5656 S.n5590 S.n5583 0.002
R5657 S.n4768 S.n4760 0.002
R5658 S.n5104 S.n5096 0.002
R5659 S.n4914 S.n4907 0.002
R5660 S.n5808 S.n5800 0.002
R5661 S.n5605 S.n5598 0.002
R5662 S.n4784 S.n4776 0.002
R5663 S.n4626 S.n4619 0.002
R5664 S.n4335 S.n4327 0.002
R5665 S.n4191 S.n4184 0.002
R5666 S.n3761 S.n3754 0.002
R5667 S.n3373 S.n3372 0.002
R5668 S.n5120 S.n5112 0.002
R5669 S.n4899 S.n4892 0.002
R5670 S.n5824 S.n5816 0.002
R5671 S.n5620 S.n5613 0.002
R5672 S.n4800 S.n4792 0.002
R5673 S.n4641 S.n4634 0.002
R5674 S.n4385 S.n4207 0.002
R5675 S.n3781 S.n3780 0.002
R5676 S.n5136 S.n5128 0.002
R5677 S.n4884 S.n4877 0.002
R5678 S.n5840 S.n5832 0.002
R5679 S.n5635 S.n5628 0.002
R5680 S.n4839 S.n4657 0.002
R5681 S.n4355 S.n4354 0.002
R5682 S.n5871 S.n5870 0.002
R5683 S.n5175 S.n5174 0.002
R5684 S.n600 S.n581 0.002
R5685 S.n327 S.n326 0.002
R5686 S.n4823 S.n4819 0.002
R5687 S.n516 S.n513 0.002
R5688 S.t283 S.n5302 0.002
R5689 S.t283 S.n5437 0.002
R5690 S.n1223 S.n1222 0.002
R5691 S.n5236 S.n5218 0.002
R5692 S.n3100 S.n3083 0.002
R5693 S.n2070 S.n2053 0.002
R5694 S.n959 S.n944 0.002
R5695 S.n520 S.n519 0.002
R5696 S.n5509 S.n5508 0.002
R5697 S.n4439 S.n4438 0.002
R5698 S.n4002 S.n4001 0.002
R5699 S.n3528 S.n3527 0.002
R5700 S.n3042 S.n3041 0.002
R5701 S.n2504 S.n2503 0.002
R5702 S.n2012 S.n2011 0.002
R5703 S.n1466 S.n1465 0.002
R5704 S.n1730 S.n1717 0.002
R5705 S.n2818 S.n2817 0.002
R5706 S.n3337 S.n3336 0.002
R5707 S.n3714 S.n3713 0.002
R5708 S.n4303 S.n4302 0.002
R5709 S.n4736 S.n4735 0.002
R5710 S.n5760 S.n5759 0.002
R5711 S.n5056 S.n5055 0.002
R5712 S.n2326 S.n2313 0.002
R5713 S.n3353 S.n3352 0.002
R5714 S.n3730 S.n3729 0.002
R5715 S.n4319 S.n4318 0.002
R5716 S.n4752 S.n4751 0.002
R5717 S.n5776 S.n5775 0.002
R5718 S.n5072 S.n5071 0.002
R5719 S.n4768 S.n4767 0.002
R5720 S.n5792 S.n5791 0.002
R5721 S.n5088 S.n5087 0.002
R5722 S.n3373 S.n3360 0.002
R5723 S.n4335 S.n4334 0.002
R5724 S.n4784 S.n4783 0.002
R5725 S.n5808 S.n5807 0.002
R5726 S.n5104 S.n5103 0.002
R5727 S.n3781 S.n3768 0.002
R5728 S.n4800 S.n4799 0.002
R5729 S.n5824 S.n5823 0.002
R5730 S.n5120 S.n5119 0.002
R5731 S.n4355 S.n4342 0.002
R5732 S.n5840 S.n5839 0.002
R5733 S.n5136 S.n5135 0.002
R5734 S.n5152 S.n5143 0.002
R5735 S.n2838 S.n2825 0.002
R5736 S.n3746 S.n3737 0.002
R5737 S.n4372 S.n4368 0.002
R5738 S.n4247 S.n4246 0.002
R5739 S.n3658 S.n3657 0.002
R5740 S.n3281 S.n3280 0.002
R5741 S.n2762 S.n2761 0.002
R5742 S.n2266 S.n2265 0.002
R5743 S.n1670 S.n1669 0.002
R5744 S.n1113 S.n1112 0.002
R5745 S.n215 S.n202 0.002
R5746 S.n273 S.n262 0.002
R5747 S.n1750 S.n1749 0.002
R5748 S.n2094 S.n2093 0.002
R5749 S.n2591 S.n2590 0.002
R5750 S.n3124 S.n3123 0.002
R5751 S.n3801 S.n3800 0.002
R5752 S.n4087 S.n4086 0.002
R5753 S.n4522 S.n4521 0.002
R5754 S.n5195 S.n5194 0.002
R5755 S.n1167 S.n1158 0.002
R5756 S.n2140 S.n2139 0.002
R5757 S.n2634 S.n2633 0.002
R5758 S.n3167 S.n3166 0.002
R5759 S.n3844 S.n3843 0.002
R5760 S.n4130 S.n4129 0.002
R5761 S.n4565 S.n4564 0.002
R5762 S.n4989 S.n4988 0.002
R5763 S.n5236 S.n5217 0.002
R5764 S.n5687 S.n5675 0.002
R5765 S.n5484 S.n5459 0.002
R5766 S.n4719 S.n4707 0.002
R5767 S.n4471 S.n4446 0.002
R5768 S.n4286 S.n4274 0.002
R5769 S.n4034 S.n4009 0.002
R5770 S.n3697 S.n3685 0.002
R5771 S.n3560 S.n3535 0.002
R5772 S.n3323 S.n3311 0.002
R5773 S.n3074 S.n3049 0.002
R5774 S.n2801 S.n2789 0.002
R5775 S.n2536 S.n2511 0.002
R5776 S.n2305 S.n2293 0.002
R5777 S.n2044 S.n2019 0.002
R5778 S.n1709 S.n1697 0.002
R5779 S.n1500 S.n1473 0.002
R5780 S.n1150 S.n1140 0.002
R5781 S.n935 S.n920 0.002
R5782 S.n254 S.n241 0.002
R5783 S.n348 S.n340 0.002
R5784 S.n4063 S.n4042 0.002
R5785 S.n3637 S.n3625 0.002
R5786 S.n3474 S.n3449 0.002
R5787 S.n3260 S.n3248 0.002
R5788 S.n2988 S.n2963 0.002
R5789 S.n2741 S.n2729 0.002
R5790 S.n2450 S.n2425 0.002
R5791 S.n2245 S.n2233 0.002
R5792 S.n1958 S.n1933 0.002
R5793 S.n1649 S.n1637 0.002
R5794 S.n1411 S.n1383 0.002
R5795 S.n1092 S.n1081 0.002
R5796 S.n851 S.n830 0.002
R5797 S.n305 S.n293 0.002
R5798 S.n290 S.n77 0.002
R5799 S.n3100 S.n3082 0.002
R5800 S.n2705 S.n2693 0.002
R5801 S.n2389 S.n2364 0.002
R5802 S.n2209 S.n2197 0.002
R5803 S.n1897 S.n1872 0.002
R5804 S.n1613 S.n1601 0.002
R5805 S.n1347 S.n1320 0.002
R5806 S.n1053 S.n1043 0.002
R5807 S.n789 S.n766 0.002
R5808 S.n178 S.n169 0.002
R5809 S.n70 S.n62 0.002
R5810 S.n2070 S.n2052 0.002
R5811 S.n1577 S.n1565 0.002
R5812 S.n1284 S.n1257 0.002
R5813 S.n1019 S.n1009 0.002
R5814 S.n730 S.n707 0.002
R5815 S.n145 S.n136 0.002
R5816 S.n49 S.n41 0.002
R5817 S.n959 S.n943 0.002
R5818 S.n112 S.n103 0.002
R5819 S.n28 S.n20 0.002
R5820 S.n5175 S.n5167 0.002
R5821 S.n5445 S.n5442 0.002
R5822 S.n632 S.n629 0.002
R5823 S.n5343 S.n5321 0.001
R5824 S.n5343 S.n5324 0.001
R5825 S.n5343 S.n5327 0.001
R5826 S.n5343 S.n5330 0.001
R5827 S.n5343 S.n5333 0.001
R5828 S.n5343 S.n5336 0.001
R5829 S.n5343 S.n5339 0.001
R5830 S.n5343 S.n5342 0.001
R5831 S.n829 S.n828 0.001
R5832 S.n784 S.n783 0.001
R5833 S.n725 S.n724 0.001
R5834 S.n5283 S.n5282 0.001
R5835 S.n521 S.n520 0.001
R5836 S.t241 S.n521 0.001
R5837 S.n4430 S.n4429 0.001
R5838 S.n3993 S.n3992 0.001
R5839 S.n3519 S.n3518 0.001
R5840 S.n3033 S.n3032 0.001
R5841 S.n2495 S.n2494 0.001
R5842 S.n2003 S.n2002 0.001
R5843 S.n1456 S.n1455 0.001
R5844 S.n896 S.n895 0.001
R5845 S.n5442 S.t283 0.001
R5846 S.n4409 S.n4408 0.001
R5847 S.n1411 S.n1394 0.001
R5848 S.n3590 S.n3589 0.001
R5849 S.n2566 S.n2565 0.001
R5850 S.n1530 S.n1529 0.001
R5851 S.n5897 S.n5896 0.001
R5852 S.n932 S.n931 0.001
R5853 S.n1149 S.n1148 0.001
R5854 S.n1497 S.n1496 0.001
R5855 S.n1706 S.n1705 0.001
R5856 S.n2041 S.n2040 0.001
R5857 S.n2302 S.n2301 0.001
R5858 S.n2533 S.n2532 0.001
R5859 S.n2798 S.n2797 0.001
R5860 S.n3071 S.n3070 0.001
R5861 S.n3320 S.n3319 0.001
R5862 S.n3557 S.n3556 0.001
R5863 S.n3694 S.n3693 0.001
R5864 S.n4031 S.n4030 0.001
R5865 S.n4283 S.n4282 0.001
R5866 S.n4468 S.n4467 0.001
R5867 S.n4716 S.n4715 0.001
R5868 S.n5481 S.n5480 0.001
R5869 S.n5684 S.n5683 0.001
R5870 S.n246 S.n245 0.001
R5871 S.n1080 S.n1079 0.001
R5872 S.n1408 S.n1407 0.001
R5873 S.n1646 S.n1645 0.001
R5874 S.n1955 S.n1954 0.001
R5875 S.n2242 S.n2241 0.001
R5876 S.n2447 S.n2446 0.001
R5877 S.n2738 S.n2737 0.001
R5878 S.n2985 S.n2984 0.001
R5879 S.n3257 S.n3256 0.001
R5880 S.n3471 S.n3470 0.001
R5881 S.n3634 S.n3633 0.001
R5882 S.n1052 S.n1051 0.001
R5883 S.n1344 S.n1343 0.001
R5884 S.n1610 S.n1609 0.001
R5885 S.n1894 S.n1893 0.001
R5886 S.n2206 S.n2205 0.001
R5887 S.n2386 S.n2385 0.001
R5888 S.n2702 S.n2701 0.001
R5889 S.n1018 S.n1017 0.001
R5890 S.n1281 S.n1280 0.001
R5891 S.n1574 S.n1573 0.001
R5892 S.n2938 S.n2937 0.001
R5893 S.n2400 S.n2399 0.001
R5894 S.n1908 S.n1907 0.001
R5895 S.n1358 S.n1357 0.001
R5896 S.n801 S.n800 0.001
R5897 S.n1847 S.n1846 0.001
R5898 S.n1295 S.n1294 0.001
R5899 S.n742 S.n741 0.001
R5900 S.n683 S.n682 0.001
R5901 S.n273 S.n263 0.001
R5902 S.n93 S.n92 0.001
R5903 S.n981 S.n980 0.001
R5904 S.n1555 S.n1554 0.001
R5905 S.n2169 S.n2168 0.001
R5906 S.n2683 S.n2682 0.001
R5907 S.n3220 S.n3219 0.001
R5908 S.n3615 S.n3614 0.001
R5909 S.n4222 S.n4221 0.001
R5910 S.n4677 S.n4676 0.001
R5911 S.n5664 S.n5663 0.001
R5912 S.n5285 S.n5284 0.001
R5913 S.t241 S.n496 0.001
R5914 S.t241 S.n396 0.001
R5915 S.t241 S.n568 0.001
R5916 S.t241 S.n602 0.001
R5917 S.t241 S.n427 0.001
R5918 S.t241 S.n458 0.001
R5919 S.n664 S.t241 0.001
R5920 S.t241 S.n628 0.001
R5921 S.t241 S.n554 0.001
R5922 S.t241 S.n542 0.001
R5923 S.t241 S.n530 0.001
R5924 S.n517 S.n516 0.001
R5925 S.n3474 S.n3459 0.001
R5926 S.n2988 S.n2973 0.001
R5927 S.n2450 S.n2435 0.001
R5928 S.n1958 S.n1943 0.001
R5929 S.n5046 S.n5045 0.001
R5930 S.n3226 S.n3225 0.001
R5931 S.n4228 S.n4227 0.001
R5932 S.n4682 S.n4681 0.001
R5933 S.n5670 S.n5669 0.001
R5934 S.n3620 S.n3619 0.001
R5935 S.n2175 S.n2174 0.001
R5936 S.n2688 S.n2687 0.001
R5937 S.n987 S.n986 0.001
R5938 S.n1560 S.n1559 0.001
R5939 S.n98 S.n97 0.001
R5940 S.n5280 S.n5266 0.001
R5941 S.n516 S.n515 0.001
R5942 S.n4063 S.n4044 0.001
R5943 S.n5194 S.n5193 0.001
R5944 S.n5208 S.n5207 0.001
R5945 S.n5729 S.n5728 0.001
R5946 S.n5529 S.n5528 0.001
R5947 S.n4521 S.n4520 0.001
R5948 S.n4535 S.n4534 0.001
R5949 S.n4086 S.n4085 0.001
R5950 S.n4100 S.n4099 0.001
R5951 S.n3800 S.n3799 0.001
R5952 S.n3814 S.n3813 0.001
R5953 S.n3123 S.n3122 0.001
R5954 S.n3137 S.n3136 0.001
R5955 S.n2590 S.n2589 0.001
R5956 S.n2604 S.n2603 0.001
R5957 S.n2093 S.n2092 0.001
R5958 S.n2107 S.n2106 0.001
R5959 S.n1749 S.n1748 0.001
R5960 S.n1763 S.n1762 0.001
R5961 S.n1186 S.n1185 0.001
R5962 S.n5165 S.n5164 0.001
R5963 S.n5008 S.n5007 0.001
R5964 S.n91 S.n90 0.001
R5965 S.n979 S.n978 0.001
R5966 S.n1553 S.n1552 0.001
R5967 S.n2167 S.n2166 0.001
R5968 S.n2681 S.n2680 0.001
R5969 S.n3218 S.n3217 0.001
R5970 S.n3613 S.n3612 0.001
R5971 S.n4220 S.n4219 0.001
R5972 S.n4675 S.n4674 0.001
R5973 S.n5662 S.n5661 0.001
R5974 S.n5039 S.n5038 0.001
R5975 S.n5266 S.t35 0.001
R5976 S.t255 S.n98 0.001
R5977 S.t64 S.n5046 0.001
R5978 S.t12 S.n3226 0.001
R5979 S.t10 S.n3620 0.001
R5980 S.t57 S.n4228 0.001
R5981 S.t8 S.n4682 0.001
R5982 S.t4 S.n5670 0.001
R5983 S.t16 S.n2175 0.001
R5984 S.t0 S.n2688 0.001
R5985 S.t6 S.n987 0.001
R5986 S.t21 S.n1560 0.001
R5987 S.n5284 S.n5283 0.001
R5988 S.n92 S.n91 0.001
R5989 S.n980 S.n979 0.001
R5990 S.n1554 S.n1553 0.001
R5991 S.n2168 S.n2167 0.001
R5992 S.n2682 S.n2681 0.001
R5993 S.n3219 S.n3218 0.001
R5994 S.n3614 S.n3613 0.001
R5995 S.n4221 S.n4220 0.001
R5996 S.n4676 S.n4675 0.001
R5997 S.n5663 S.n5662 0.001
R5998 S.n5041 S.n5035 0.001
R5999 S.n5343 S.n5318 0.001
R6000 S.n5695 S.n5694 0.001
R6001 S.n291 S.n290 0.001
R6002 S.n178 S.n170 0.001
R6003 S.n145 S.n137 0.001
R6004 S.n112 S.n104 0.001
R6005 S.n366 S.n365 0.001
R6006 S.n1213 S.n1212 0.001
R6007 S.n1249 S.n1248 0.001
R6008 S.n1835 S.n1834 0.001
R6009 S.n2876 S.n2875 0.001
R6010 S.n2926 S.n2925 0.001
R6011 S.n3441 S.n3440 0.001
R6012 S.n3947 S.n3946 0.001
R6013 S.n4418 S.n4417 0.001
R6014 S.n5453 S.n5452 0.001
R6015 S.n5273 S.n5272 0.001
R6016 S.n595 S.n594 0.001
R6017 S.n516 S.n509 0.001
R6018 S.n516 S.n512 0.001
R6019 S.n516 S.n511 0.001
R6020 S.n516 S.n510 0.001
R6021 S.n5013 S.n5012 0.001
R6022 S.n5252 S.n5251 0.001
R6023 S.n5699 S.n5698 0.001
R6024 S.n478 S.n477 0.001
R6025 S.n343 S.n342 0.001
R6026 S.n927 S.n926 0.001
R6027 S.n5224 S.n5223 0.001
R6028 S.n5682 S.n5681 0.001
R6029 S.n5475 S.n5474 0.001
R6030 S.n4714 S.n4713 0.001
R6031 S.n4462 S.n4461 0.001
R6032 S.n4281 S.n4280 0.001
R6033 S.n4025 S.n4024 0.001
R6034 S.n3692 S.n3691 0.001
R6035 S.n3551 S.n3550 0.001
R6036 S.n3318 S.n3317 0.001
R6037 S.n3065 S.n3064 0.001
R6038 S.n2796 S.n2795 0.001
R6039 S.n2527 S.n2526 0.001
R6040 S.n2300 S.n2299 0.001
R6041 S.n2035 S.n2034 0.001
R6042 S.n1704 S.n1703 0.001
R6043 S.n1489 S.n1488 0.001
R6044 S.n1147 S.n1146 0.001
R6045 S.n249 S.n248 0.001
R6046 S.n65 S.n64 0.001
R6047 S.n782 S.n781 0.001
R6048 S.n3089 S.n3088 0.001
R6049 S.n2700 S.n2699 0.001
R6050 S.n2380 S.n2379 0.001
R6051 S.n2204 S.n2203 0.001
R6052 S.n1888 S.n1887 0.001
R6053 S.n1608 S.n1607 0.001
R6054 S.n1336 S.n1335 0.001
R6055 S.n1050 S.n1049 0.001
R6056 S.n13 S.n12 0.001
R6057 S.n3579 S.n3578 0.001
R6058 S.n3236 S.n3235 0.001
R6059 S.n2942 S.n2941 0.001
R6060 S.n2717 S.n2716 0.001
R6061 S.n2404 S.n2403 0.001
R6062 S.n2221 S.n2220 0.001
R6063 S.n1912 S.n1911 0.001
R6064 S.n1625 S.n1624 0.001
R6065 S.n1362 S.n1361 0.001
R6066 S.n1065 S.n1064 0.001
R6067 S.n1084 S.n1083 0.001
R6068 S.n833 S.n832 0.001
R6069 S.n80 S.n79 0.001
R6070 S.n296 S.n295 0.001
R6071 S.n1400 S.n1399 0.001
R6072 S.n1949 S.n1948 0.001
R6073 S.n2441 S.n2440 0.001
R6074 S.n2979 S.n2978 0.001
R6075 S.n3465 S.n3464 0.001
R6076 S.n4052 S.n4051 0.001
R6077 S.n3632 S.n3631 0.001
R6078 S.n3255 S.n3254 0.001
R6079 S.n2736 S.n2735 0.001
R6080 S.n2240 S.n2239 0.001
R6081 S.n1644 S.n1643 0.001
R6082 S.n872 S.n871 0.001
R6083 S.n206 S.n205 0.001
R6084 S.n584 S.n583 0.001
R6085 S.n4493 S.n4492 0.001
R6086 S.n4245 S.n4244 0.001
R6087 S.n3970 S.n3969 0.001
R6088 S.n3656 S.n3655 0.001
R6089 S.n3496 S.n3495 0.001
R6090 S.n3279 S.n3278 0.001
R6091 S.n3010 S.n3009 0.001
R6092 S.n2760 S.n2759 0.001
R6093 S.n2472 S.n2471 0.001
R6094 S.n2264 S.n2263 0.001
R6095 S.n1980 S.n1979 0.001
R6096 S.n1668 S.n1667 0.001
R6097 S.n1433 S.n1432 0.001
R6098 S.n1111 S.n1110 0.001
R6099 S.n900 S.n899 0.001
R6100 S.n226 S.n225 0.001
R6101 S.n1130 S.n1129 0.001
R6102 S.n1460 S.n1459 0.001
R6103 S.n1682 S.n1681 0.001
R6104 S.n2007 S.n2006 0.001
R6105 S.n2278 S.n2277 0.001
R6106 S.n2499 S.n2498 0.001
R6107 S.n2774 S.n2773 0.001
R6108 S.n3037 S.n3036 0.001
R6109 S.n3293 S.n3292 0.001
R6110 S.n3523 S.n3522 0.001
R6111 S.n3670 S.n3669 0.001
R6112 S.n3997 S.n3996 0.001
R6113 S.n4259 S.n4258 0.001
R6114 S.n4434 S.n4433 0.001
R6115 S.n4692 S.n4691 0.001
R6116 S.n5504 S.n5503 0.001
R6117 S.n316 S.n315 0.001
R6118 S.n804 S.n803 0.001
R6119 S.n190 S.n189 0.001
R6120 S.n173 S.n172 0.001
R6121 S.n44 S.n43 0.001
R6122 S.n723 S.n722 0.001
R6123 S.n2059 S.n2058 0.001
R6124 S.n1572 S.n1571 0.001
R6125 S.n1273 S.n1272 0.001
R6126 S.n1016 S.n1015 0.001
R6127 S.n414 S.n413 0.001
R6128 S.n2555 S.n2554 0.001
R6129 S.n2185 S.n2184 0.001
R6130 S.n1851 S.n1850 0.001
R6131 S.n1589 S.n1588 0.001
R6132 S.n1299 S.n1298 0.001
R6133 S.n1031 S.n1030 0.001
R6134 S.n745 S.n744 0.001
R6135 S.n157 S.n156 0.001
R6136 S.n140 S.n139 0.001
R6137 S.n23 S.n22 0.001
R6138 S.n950 S.n949 0.001
R6139 S.n445 S.n444 0.001
R6140 S.n1519 S.n1518 0.001
R6141 S.n997 S.n996 0.001
R6142 S.n686 S.n685 0.001
R6143 S.n124 S.n123 0.001
R6144 S.n107 S.n106 0.001
R6145 S.n266 S.n265 0.001
R6146 S.n1190 S.n1189 0.001
R6147 S.n969 S.n968 0.001
R6148 S.n1754 S.n1753 0.001
R6149 S.n1541 S.n1540 0.001
R6150 S.n2098 S.n2097 0.001
R6151 S.n2080 S.n2079 0.001
R6152 S.n2595 S.n2594 0.001
R6153 S.n2577 S.n2576 0.001
R6154 S.n3128 S.n3127 0.001
R6155 S.n3110 S.n3109 0.001
R6156 S.n3805 S.n3804 0.001
R6157 S.n3601 S.n3600 0.001
R6158 S.n4091 S.n4090 0.001
R6159 S.n4073 S.n4072 0.001
R6160 S.n4526 S.n4525 0.001
R6161 S.n4508 S.n4507 0.001
R6162 S.n5520 S.n5519 0.001
R6163 S.n5722 S.n5721 0.001
R6164 S.n5199 S.n5198 0.001
R6165 S.n5000 S.n4999 0.001
R6166 S.n1162 S.n1161 0.001
R6167 S.n1777 S.n1776 0.001
R6168 S.n4987 S.n4986 0.001
R6169 S.n4973 S.n4972 0.001
R6170 S.n5743 S.n5742 0.001
R6171 S.n5543 S.n5542 0.001
R6172 S.n4563 S.n4562 0.001
R6173 S.n4549 S.n4548 0.001
R6174 S.n4128 S.n4127 0.001
R6175 S.n4114 S.n4113 0.001
R6176 S.n3842 S.n3841 0.001
R6177 S.n3828 S.n3827 0.001
R6178 S.n3165 S.n3164 0.001
R6179 S.n3151 S.n3150 0.001
R6180 S.n2632 S.n2631 0.001
R6181 S.n2618 S.n2617 0.001
R6182 S.n2138 S.n2137 0.001
R6183 S.n2124 S.n2123 0.001
R6184 S.n1791 S.n1790 0.001
R6185 S.n1721 S.n1720 0.001
R6186 S.n2152 S.n2151 0.001
R6187 S.n5054 S.n5053 0.001
R6188 S.n4958 S.n4957 0.001
R6189 S.n5758 S.n5757 0.001
R6190 S.n5559 S.n5558 0.001
R6191 S.n4734 S.n4733 0.001
R6192 S.n4580 S.n4579 0.001
R6193 S.n4301 S.n4300 0.001
R6194 S.n4145 S.n4144 0.001
R6195 S.n3712 S.n3711 0.001
R6196 S.n3859 S.n3858 0.001
R6197 S.n3335 S.n3334 0.001
R6198 S.n3182 S.n3181 0.001
R6199 S.n2816 S.n2815 0.001
R6200 S.n2649 S.n2648 0.001
R6201 S.n2341 S.n2340 0.001
R6202 S.n2317 S.n2316 0.001
R6203 S.n2664 S.n2663 0.001
R6204 S.n5070 S.n5069 0.001
R6205 S.n4943 S.n4942 0.001
R6206 S.n5774 S.n5773 0.001
R6207 S.n5574 S.n5573 0.001
R6208 S.n4750 S.n4749 0.001
R6209 S.n4595 S.n4594 0.001
R6210 S.n4317 S.n4316 0.001
R6211 S.n4160 S.n4159 0.001
R6212 S.n3728 S.n3727 0.001
R6213 S.n3874 S.n3873 0.001
R6214 S.n3351 S.n3350 0.001
R6215 S.n3197 S.n3196 0.001
R6216 S.n2853 S.n2852 0.001
R6217 S.n4610 S.n4609 0.001
R6218 S.n5086 S.n5085 0.001
R6219 S.n4928 S.n4927 0.001
R6220 S.n5790 S.n5789 0.001
R6221 S.n5589 S.n5588 0.001
R6222 S.n4766 S.n4765 0.001
R6223 S.n4171 S.n4170 0.001
R6224 S.n3741 S.n3740 0.001
R6225 S.n3885 S.n3884 0.001
R6226 S.n3208 S.n3207 0.001
R6227 S.n3394 S.n3393 0.001
R6228 S.n2829 S.n2828 0.001
R6229 S.n3364 S.n3363 0.001
R6230 S.n3904 S.n3903 0.001
R6231 S.n5102 S.n5101 0.001
R6232 S.n4913 S.n4912 0.001
R6233 S.n5806 S.n5805 0.001
R6234 S.n5604 S.n5603 0.001
R6235 S.n4782 S.n4781 0.001
R6236 S.n4625 S.n4624 0.001
R6237 S.n4333 S.n4332 0.001
R6238 S.n4190 S.n4189 0.001
R6239 S.n3760 S.n3759 0.001
R6240 S.n3772 S.n3771 0.001
R6241 S.n4205 S.n4204 0.001
R6242 S.n5118 S.n5117 0.001
R6243 S.n4898 S.n4897 0.001
R6244 S.n5822 S.n5821 0.001
R6245 S.n5619 S.n5618 0.001
R6246 S.n4798 S.n4797 0.001
R6247 S.n4640 S.n4639 0.001
R6248 S.n4384 S.n4383 0.001
R6249 S.n4346 S.n4345 0.001
R6250 S.n4655 S.n4654 0.001
R6251 S.n5134 S.n5133 0.001
R6252 S.n4883 S.n4882 0.001
R6253 S.n5838 S.n5837 0.001
R6254 S.n5634 S.n5633 0.001
R6255 S.n4838 S.n4837 0.001
R6256 S.n4809 S.n4808 0.001
R6257 S.n5865 S.n5864 0.001
R6258 S.n5147 S.n5146 0.001
R6259 S.n4864 S.n4863 0.001
R6260 S.n5650 S.n5649 0.001
R6261 S.n5170 S.n5169 0.001
R6262 S.n5321 S.n5320 0.001
R6263 S.n5324 S.n5323 0.001
R6264 S.n5327 S.n5326 0.001
R6265 S.n5330 S.n5329 0.001
R6266 S.n5333 S.n5332 0.001
R6267 S.n5336 S.n5335 0.001
R6268 S.n5339 S.n5338 0.001
R6269 S.n5342 S.n5341 0.001
R6270 S.n516 S.n514 0.001
R6271 S.n5043 S.n5042 0.001
R6272 S.n5666 S.n5665 0.001
R6273 S.n4679 S.n4678 0.001
R6274 S.n4224 S.n4223 0.001
R6275 S.n3617 S.n3616 0.001
R6276 S.n3222 S.n3221 0.001
R6277 S.n2685 S.n2684 0.001
R6278 S.n2171 S.n2170 0.001
R6279 S.n1557 S.n1556 0.001
R6280 S.n983 S.n982 0.001
R6281 S.n95 S.n94 0.001
R6282 S.t64 S.n5021 0.001
R6283 S.t64 S.n5024 0.001
R6284 S.t35 S.n5260 0.001
R6285 S.t35 S.n5263 0.001
R6286 S.t4 S.n5717 0.001
R6287 S.t4 S.n5714 0.001
R6288 S.n5714 S.n5711 0.001
R6289 S.n5880 S.t25 0.001
R6290 S.n5900 S.n5882 0.001
R6291 S.n494 S.n484 0.001
R6292 S.t198 S.n354 0.001
R6293 S.t198 S.n351 0.001
R6294 S.n351 S.n348 0.001
R6295 S.t59 S.n941 0.001
R6296 S.t59 S.n938 0.001
R6297 S.n938 S.n935 0.001
R6298 S.t35 S.n5242 0.001
R6299 S.t35 S.n5239 0.001
R6300 S.n5239 S.n5236 0.001
R6301 S.t4 S.n5693 0.001
R6302 S.t4 S.n5690 0.001
R6303 S.n5690 S.n5687 0.001
R6304 S.t25 S.n5490 0.001
R6305 S.t25 S.n5487 0.001
R6306 S.n5487 S.n5484 0.001
R6307 S.t8 S.n4725 0.001
R6308 S.t8 S.n4722 0.001
R6309 S.n4722 S.n4719 0.001
R6310 S.t71 S.n4477 0.001
R6311 S.t71 S.n4474 0.001
R6312 S.n4474 S.n4471 0.001
R6313 S.t57 S.n4292 0.001
R6314 S.t57 S.n4289 0.001
R6315 S.n4289 S.n4286 0.001
R6316 S.t54 S.n4040 0.001
R6317 S.t54 S.n4037 0.001
R6318 S.n4037 S.n4034 0.001
R6319 S.t10 S.n3703 0.001
R6320 S.t10 S.n3700 0.001
R6321 S.n3700 S.n3697 0.001
R6322 S.t42 S.n3566 0.001
R6323 S.t42 S.n3563 0.001
R6324 S.n3563 S.n3560 0.001
R6325 S.t12 S.n3326 0.001
R6326 S.t12 S.n3310 0.001
R6327 S.t14 S.n3080 0.001
R6328 S.t14 S.n3077 0.001
R6329 S.n3077 S.n3074 0.001
R6330 S.t0 S.n2807 0.001
R6331 S.t0 S.n2804 0.001
R6332 S.n2804 S.n2801 0.001
R6333 S.t66 S.n2542 0.001
R6334 S.t66 S.n2539 0.001
R6335 S.n2539 S.n2536 0.001
R6336 S.t16 S.n2311 0.001
R6337 S.t16 S.n2308 0.001
R6338 S.n2308 S.n2305 0.001
R6339 S.t47 S.n2050 0.001
R6340 S.t47 S.n2047 0.001
R6341 S.n2047 S.n2044 0.001
R6342 S.t21 S.n1715 0.001
R6343 S.t21 S.n1712 0.001
R6344 S.n1712 S.n1709 0.001
R6345 S.t23 S.n1506 0.001
R6346 S.t23 S.n1503 0.001
R6347 S.n1503 S.n1500 0.001
R6348 S.t6 S.n1156 0.001
R6349 S.t6 S.n1153 0.001
R6350 S.n1153 S.n1150 0.001
R6351 S.t255 S.n260 0.001
R6352 S.t255 S.n257 0.001
R6353 S.n257 S.n254 0.001
R6354 S.t198 S.n76 0.001
R6355 S.t198 S.n73 0.001
R6356 S.n73 S.n70 0.001
R6357 S.t59 S.n795 0.001
R6358 S.t59 S.n792 0.001
R6359 S.n792 S.n789 0.001
R6360 S.t14 S.n3103 0.001
R6361 S.t14 S.n3106 0.001
R6362 S.t0 S.n2711 0.001
R6363 S.t0 S.n2708 0.001
R6364 S.n2708 S.n2705 0.001
R6365 S.t66 S.n2395 0.001
R6366 S.t66 S.n2392 0.001
R6367 S.n2392 S.n2389 0.001
R6368 S.t16 S.n2215 0.001
R6369 S.t16 S.n2212 0.001
R6370 S.n2212 S.n2209 0.001
R6371 S.t47 S.n1903 0.001
R6372 S.t47 S.n1900 0.001
R6373 S.n1900 S.n1897 0.001
R6374 S.t21 S.n1619 0.001
R6375 S.t21 S.n1616 0.001
R6376 S.n1616 S.n1613 0.001
R6377 S.t23 S.n1353 0.001
R6378 S.t23 S.n1350 0.001
R6379 S.n1350 S.n1347 0.001
R6380 S.t6 S.n1059 0.001
R6381 S.t6 S.n1056 0.001
R6382 S.n1056 S.n1053 0.001
R6383 S.n386 S.t198 0.001
R6384 S.n394 S.n389 0.001
R6385 S.t42 S.n3594 0.001
R6386 S.t42 S.n3597 0.001
R6387 S.t12 S.n3247 0.001
R6388 S.t12 S.n3244 0.001
R6389 S.n3244 S.n3241 0.001
R6390 S.t14 S.n2962 0.001
R6391 S.t14 S.n2959 0.001
R6392 S.n2959 S.n2956 0.001
R6393 S.t0 S.n2728 0.001
R6394 S.t0 S.n2725 0.001
R6395 S.n2725 S.n2722 0.001
R6396 S.t66 S.n2424 0.001
R6397 S.t66 S.n2421 0.001
R6398 S.n2421 S.n2418 0.001
R6399 S.t16 S.n2232 0.001
R6400 S.t16 S.n2229 0.001
R6401 S.n2229 S.n2226 0.001
R6402 S.t47 S.n1932 0.001
R6403 S.t47 S.n1929 0.001
R6404 S.n1929 S.n1926 0.001
R6405 S.t21 S.n1636 0.001
R6406 S.t21 S.n1633 0.001
R6407 S.n1633 S.n1630 0.001
R6408 S.t23 S.n1382 0.001
R6409 S.t23 S.n1379 0.001
R6410 S.n1379 S.n1376 0.001
R6411 S.t6 S.n1078 0.001
R6412 S.t6 S.n1075 0.001
R6413 S.n1075 S.n1072 0.001
R6414 S.t6 S.n1098 0.001
R6415 S.t6 S.n1095 0.001
R6416 S.n1095 S.n1092 0.001
R6417 S.t59 S.n857 0.001
R6418 S.t59 S.n854 0.001
R6419 S.n854 S.n851 0.001
R6420 S.n282 S.t255 0.001
R6421 S.n290 S.n285 0.001
R6422 S.t198 S.n311 0.001
R6423 S.t198 S.n308 0.001
R6424 S.n308 S.n305 0.001
R6425 S.t23 S.n1417 0.001
R6426 S.t23 S.n1414 0.001
R6427 S.n1414 S.n1411 0.001
R6428 S.t47 S.n1964 0.001
R6429 S.t47 S.n1961 0.001
R6430 S.n1961 S.n1958 0.001
R6431 S.t66 S.n2456 0.001
R6432 S.t66 S.n2453 0.001
R6433 S.n2453 S.n2450 0.001
R6434 S.t14 S.n2994 0.001
R6435 S.t14 S.n2991 0.001
R6436 S.n2991 S.n2988 0.001
R6437 S.t42 S.n3480 0.001
R6438 S.t42 S.n3477 0.001
R6439 S.n3477 S.n3474 0.001
R6440 S.t54 S.n4066 0.001
R6441 S.t54 S.n4069 0.001
R6442 S.t10 S.n3643 0.001
R6443 S.t10 S.n3640 0.001
R6444 S.n3640 S.n3637 0.001
R6445 S.t12 S.n3266 0.001
R6446 S.t12 S.n3263 0.001
R6447 S.n3263 S.n3260 0.001
R6448 S.t0 S.n2747 0.001
R6449 S.t0 S.n2744 0.001
R6450 S.n2744 S.n2741 0.001
R6451 S.t16 S.n2251 0.001
R6452 S.t16 S.n2248 0.001
R6453 S.n2248 S.n2245 0.001
R6454 S.t21 S.n1655 0.001
R6455 S.t21 S.n1652 0.001
R6456 S.n1652 S.n1649 0.001
R6457 S.t59 S.n891 0.001
R6458 S.t59 S.n888 0.001
R6459 S.n888 S.n885 0.001
R6460 S.t255 S.n221 0.001
R6461 S.t255 S.n218 0.001
R6462 S.n218 S.n215 0.001
R6463 S.n600 S.n590 0.001
R6464 S.t71 S.n4501 0.001
R6465 S.t71 S.n4504 0.001
R6466 S.t57 S.n4253 0.001
R6467 S.t57 S.n4250 0.001
R6468 S.n4250 S.n4247 0.001
R6469 S.t54 S.n3988 0.001
R6470 S.t54 S.n3985 0.001
R6471 S.n3985 S.n3982 0.001
R6472 S.t10 S.n3664 0.001
R6473 S.t10 S.n3661 0.001
R6474 S.n3661 S.n3658 0.001
R6475 S.t42 S.n3514 0.001
R6476 S.t42 S.n3511 0.001
R6477 S.n3511 S.n3508 0.001
R6478 S.t12 S.n3287 0.001
R6479 S.t12 S.n3284 0.001
R6480 S.n3284 S.n3281 0.001
R6481 S.t14 S.n3028 0.001
R6482 S.t14 S.n3025 0.001
R6483 S.n3025 S.n3022 0.001
R6484 S.t0 S.n2768 0.001
R6485 S.t0 S.n2765 0.001
R6486 S.n2765 S.n2762 0.001
R6487 S.t66 S.n2490 0.001
R6488 S.t66 S.n2487 0.001
R6489 S.n2487 S.n2484 0.001
R6490 S.t16 S.n2272 0.001
R6491 S.t16 S.n2269 0.001
R6492 S.n2269 S.n2266 0.001
R6493 S.t47 S.n1998 0.001
R6494 S.t47 S.n1995 0.001
R6495 S.n1995 S.n1992 0.001
R6496 S.t21 S.n1676 0.001
R6497 S.t21 S.n1673 0.001
R6498 S.n1673 S.n1670 0.001
R6499 S.t23 S.n1451 0.001
R6500 S.t23 S.n1448 0.001
R6501 S.n1448 S.n1445 0.001
R6502 S.t6 S.n1119 0.001
R6503 S.t6 S.n1116 0.001
R6504 S.n1116 S.n1113 0.001
R6505 S.t59 S.n919 0.001
R6506 S.t59 S.n916 0.001
R6507 S.n916 S.n913 0.001
R6508 S.t255 S.n240 0.001
R6509 S.t255 S.n237 0.001
R6510 S.n237 S.n234 0.001
R6511 S.t6 S.n1139 0.001
R6512 S.t6 S.n1136 0.001
R6513 S.n1136 S.n1133 0.001
R6514 S.t23 S.n1472 0.001
R6515 S.t23 S.n1469 0.001
R6516 S.n1469 S.n1466 0.001
R6517 S.t21 S.n1696 0.001
R6518 S.t21 S.n1693 0.001
R6519 S.n1693 S.n1690 0.001
R6520 S.t47 S.n2018 0.001
R6521 S.t47 S.n2015 0.001
R6522 S.n2015 S.n2012 0.001
R6523 S.t16 S.n2292 0.001
R6524 S.t16 S.n2289 0.001
R6525 S.n2289 S.n2286 0.001
R6526 S.t66 S.n2510 0.001
R6527 S.t66 S.n2507 0.001
R6528 S.n2507 S.n2504 0.001
R6529 S.t0 S.n2788 0.001
R6530 S.t0 S.n2785 0.001
R6531 S.n2785 S.n2782 0.001
R6532 S.t14 S.n3048 0.001
R6533 S.t14 S.n3045 0.001
R6534 S.n3045 S.n3042 0.001
R6535 S.t12 S.n3307 0.001
R6536 S.t12 S.n3304 0.001
R6537 S.n3304 S.n3301 0.001
R6538 S.t42 S.n3534 0.001
R6539 S.t42 S.n3531 0.001
R6540 S.n3531 S.n3528 0.001
R6541 S.t10 S.n3684 0.001
R6542 S.t10 S.n3681 0.001
R6543 S.n3681 S.n3678 0.001
R6544 S.t54 S.n4008 0.001
R6545 S.t54 S.n4005 0.001
R6546 S.n4005 S.n4002 0.001
R6547 S.t57 S.n4273 0.001
R6548 S.t57 S.n4270 0.001
R6549 S.n4270 S.n4267 0.001
R6550 S.t71 S.n4445 0.001
R6551 S.t71 S.n4442 0.001
R6552 S.n4442 S.n4439 0.001
R6553 S.t8 S.n4706 0.001
R6554 S.t8 S.n4703 0.001
R6555 S.n4703 S.n4700 0.001
R6556 S.t25 S.n5512 0.001
R6557 S.t25 S.n5515 0.001
R6558 S.t198 S.n333 0.001
R6559 S.t198 S.n330 0.001
R6560 S.n330 S.n327 0.001
R6561 S.t59 S.n823 0.001
R6562 S.t59 S.n820 0.001
R6563 S.n820 S.n817 0.001
R6564 S.t255 S.n201 0.001
R6565 S.t255 S.n198 0.001
R6566 S.n198 S.n195 0.001
R6567 S.t255 S.n184 0.001
R6568 S.t255 S.n181 0.001
R6569 S.n181 S.n178 0.001
R6570 S.t198 S.n55 0.001
R6571 S.t198 S.n52 0.001
R6572 S.n52 S.n49 0.001
R6573 S.t59 S.n736 0.001
R6574 S.t59 S.n733 0.001
R6575 S.n733 S.n730 0.001
R6576 S.t47 S.n2073 0.001
R6577 S.t47 S.n2076 0.001
R6578 S.t21 S.n1583 0.001
R6579 S.t21 S.n1580 0.001
R6580 S.n1580 S.n1577 0.001
R6581 S.t23 S.n1290 0.001
R6582 S.t23 S.n1287 0.001
R6583 S.n1287 S.n1284 0.001
R6584 S.t6 S.n1025 0.001
R6585 S.t6 S.n1022 0.001
R6586 S.n1022 S.n1019 0.001
R6587 S.n425 S.n420 0.001
R6588 S.t66 S.n2570 0.001
R6589 S.t66 S.n2573 0.001
R6590 S.t16 S.n2196 0.001
R6591 S.t16 S.n2193 0.001
R6592 S.n2193 S.n2190 0.001
R6593 S.t47 S.n1871 0.001
R6594 S.t47 S.n1868 0.001
R6595 S.n1868 S.n1865 0.001
R6596 S.t21 S.n1600 0.001
R6597 S.t21 S.n1597 0.001
R6598 S.n1597 S.n1594 0.001
R6599 S.t23 S.n1319 0.001
R6600 S.t23 S.n1316 0.001
R6601 S.n1316 S.n1313 0.001
R6602 S.t6 S.n1042 0.001
R6603 S.t6 S.n1039 0.001
R6604 S.n1039 S.n1036 0.001
R6605 S.t59 S.n765 0.001
R6606 S.t59 S.n762 0.001
R6607 S.n762 S.n759 0.001
R6608 S.t255 S.n168 0.001
R6609 S.t255 S.n165 0.001
R6610 S.n165 S.n162 0.001
R6611 S.t255 S.n151 0.001
R6612 S.t255 S.n148 0.001
R6613 S.n148 S.n145 0.001
R6614 S.t198 S.n34 0.001
R6615 S.t198 S.n31 0.001
R6616 S.n31 S.n28 0.001
R6617 S.t59 S.n962 0.001
R6618 S.t59 S.n965 0.001
R6619 S.n456 S.n451 0.001
R6620 S.t23 S.n1534 0.001
R6621 S.t23 S.n1537 0.001
R6622 S.t6 S.n1008 0.001
R6623 S.t6 S.n1005 0.001
R6624 S.n1005 S.n1002 0.001
R6625 S.t59 S.n706 0.001
R6626 S.t59 S.n703 0.001
R6627 S.n703 S.n700 0.001
R6628 S.t255 S.n135 0.001
R6629 S.t255 S.n132 0.001
R6630 S.n132 S.n129 0.001
R6631 S.t255 S.n118 0.001
R6632 S.t255 S.n115 0.001
R6633 S.n115 S.n112 0.001
R6634 S.t198 S.n381 0.001
R6635 S.t198 S.n383 0.001
R6636 S.t255 S.n276 0.001
R6637 S.t255 S.n279 0.001
R6638 S.t59 S.n1198 0.001
R6639 S.t59 S.n1201 0.001
R6640 S.n1176 S.t6 0.001
R6641 S.n1186 S.n1179 0.001
R6642 S.t23 S.n1766 0.001
R6643 S.t23 S.n1769 0.001
R6644 S.n1739 S.t21 0.001
R6645 S.n1749 S.n1742 0.001
R6646 S.t47 S.n2110 0.001
R6647 S.t47 S.n2113 0.001
R6648 S.n2093 S.n2086 0.001
R6649 S.t66 S.n2607 0.001
R6650 S.t66 S.n2610 0.001
R6651 S.n2590 S.n2583 0.001
R6652 S.t14 S.n3140 0.001
R6653 S.t14 S.n3143 0.001
R6654 S.n3123 S.n3116 0.001
R6655 S.t42 S.n3817 0.001
R6656 S.t42 S.n3820 0.001
R6657 S.n3790 S.t10 0.001
R6658 S.n3800 S.n3793 0.001
R6659 S.t54 S.n4103 0.001
R6660 S.t54 S.n4106 0.001
R6661 S.n4086 S.n4079 0.001
R6662 S.t71 S.n4538 0.001
R6663 S.t71 S.n4541 0.001
R6664 S.n4521 S.n4514 0.001
R6665 S.t25 S.n5532 0.001
R6666 S.t25 S.n5535 0.001
R6667 S.t4 S.n5732 0.001
R6668 S.t4 S.n5735 0.001
R6669 S.t35 S.n5214 0.001
R6670 S.t35 S.n5211 0.001
R6671 S.n5211 S.n5208 0.001
R6672 S.n5184 S.t64 0.001
R6673 S.n5194 S.n5187 0.001
R6674 S.n5193 S.n5192 0.001
R6675 S.n5207 S.n5206 0.001
R6676 S.n5728 S.n5727 0.001
R6677 S.n5528 S.n5527 0.001
R6678 S.n4520 S.n4519 0.001
R6679 S.n4534 S.n4533 0.001
R6680 S.n4085 S.n4084 0.001
R6681 S.n4099 S.n4098 0.001
R6682 S.n3799 S.n3798 0.001
R6683 S.n3813 S.n3812 0.001
R6684 S.n3122 S.n3121 0.001
R6685 S.n3136 S.n3135 0.001
R6686 S.n2589 S.n2588 0.001
R6687 S.n2603 S.n2602 0.001
R6688 S.n2092 S.n2091 0.001
R6689 S.n2106 S.n2105 0.001
R6690 S.n1748 S.n1747 0.001
R6691 S.n1762 S.n1761 0.001
R6692 S.n1185 S.n1184 0.001
R6693 S.n1204 S.t59 0.001
R6694 S.n1222 S.n1206 0.001
R6695 S.t6 S.n1170 0.001
R6696 S.t6 S.n1173 0.001
R6697 S.t23 S.n1796 0.001
R6698 S.t23 S.n1799 0.001
R6699 S.n4988 S.n4981 0.001
R6700 S.t35 S.n4996 0.001
R6701 S.t35 S.n4993 0.001
R6702 S.n4993 S.n4990 0.001
R6703 S.t4 S.n5747 0.001
R6704 S.t4 S.n5750 0.001
R6705 S.t25 S.n5548 0.001
R6706 S.t25 S.n5551 0.001
R6707 S.n4564 S.n4557 0.001
R6708 S.t71 S.n4569 0.001
R6709 S.t71 S.n4572 0.001
R6710 S.n4129 S.n4122 0.001
R6711 S.t54 S.n4134 0.001
R6712 S.t54 S.n4137 0.001
R6713 S.n3843 S.n3836 0.001
R6714 S.t42 S.n3848 0.001
R6715 S.t42 S.n3851 0.001
R6716 S.n3166 S.n3159 0.001
R6717 S.t14 S.n3171 0.001
R6718 S.t14 S.n3174 0.001
R6719 S.n2633 S.n2626 0.001
R6720 S.t66 S.n2638 0.001
R6721 S.t66 S.n2641 0.001
R6722 S.n2139 S.n2132 0.001
R6723 S.t47 S.n2144 0.001
R6724 S.n2144 S.n2141 0.001
R6725 S.n1792 S.n1785 0.001
R6726 S.n1801 S.t23 0.001
R6727 S.n1809 S.n1801 0.001
R6728 S.t21 S.n1733 0.001
R6729 S.t21 S.n1736 0.001
R6730 S.t47 S.n2346 0.001
R6731 S.t47 S.n2349 0.001
R6732 S.t64 S.n5059 0.001
R6733 S.t64 S.n5062 0.001
R6734 S.t35 S.n4965 0.001
R6735 S.t35 S.n4962 0.001
R6736 S.n4962 S.n4959 0.001
R6737 S.t4 S.n5763 0.001
R6738 S.t4 S.n5766 0.001
R6739 S.t25 S.n5563 0.001
R6740 S.t25 S.n5566 0.001
R6741 S.t8 S.n4739 0.001
R6742 S.t8 S.n4742 0.001
R6743 S.t71 S.n4584 0.001
R6744 S.t71 S.n4587 0.001
R6745 S.t57 S.n4306 0.001
R6746 S.t57 S.n4309 0.001
R6747 S.t54 S.n4149 0.001
R6748 S.t54 S.n4152 0.001
R6749 S.t10 S.n3717 0.001
R6750 S.t10 S.n3720 0.001
R6751 S.t42 S.n3863 0.001
R6752 S.t42 S.n3866 0.001
R6753 S.t12 S.n3340 0.001
R6754 S.t12 S.n3343 0.001
R6755 S.t14 S.n3186 0.001
R6756 S.t14 S.n3189 0.001
R6757 S.t0 S.n2821 0.001
R6758 S.t0 S.n2824 0.001
R6759 S.t66 S.n2653 0.001
R6760 S.t66 S.n2656 0.001
R6761 S.n2335 S.t16 0.001
R6762 S.n2342 S.n2335 0.001
R6763 S.n2351 S.t47 0.001
R6764 S.n2359 S.n2351 0.001
R6765 S.t16 S.n2329 0.001
R6766 S.t16 S.n2332 0.001
R6767 S.t66 S.n2858 0.001
R6768 S.t66 S.n2861 0.001
R6769 S.t64 S.n5075 0.001
R6770 S.t64 S.n5078 0.001
R6771 S.t35 S.n4950 0.001
R6772 S.t35 S.n4947 0.001
R6773 S.n4947 S.n4944 0.001
R6774 S.t4 S.n5779 0.001
R6775 S.t4 S.n5782 0.001
R6776 S.t25 S.n5578 0.001
R6777 S.t25 S.n5581 0.001
R6778 S.t8 S.n4755 0.001
R6779 S.t8 S.n4758 0.001
R6780 S.t71 S.n4599 0.001
R6781 S.t71 S.n4602 0.001
R6782 S.t57 S.n4322 0.001
R6783 S.t57 S.n4325 0.001
R6784 S.t54 S.n4164 0.001
R6785 S.t54 S.n4167 0.001
R6786 S.t10 S.n3733 0.001
R6787 S.t10 S.n3736 0.001
R6788 S.t42 S.n3878 0.001
R6789 S.t42 S.n3881 0.001
R6790 S.t12 S.n3356 0.001
R6791 S.t12 S.n3359 0.001
R6792 S.t14 S.n3201 0.001
R6793 S.t14 S.n3204 0.001
R6794 S.n2847 S.t0 0.001
R6795 S.n2854 S.n2847 0.001
R6796 S.t71 S.n4614 0.001
R6797 S.t71 S.n4617 0.001
R6798 S.t64 S.n5091 0.001
R6799 S.t64 S.n5094 0.001
R6800 S.t35 S.n4935 0.001
R6801 S.t35 S.n4932 0.001
R6802 S.n4932 S.n4929 0.001
R6803 S.t4 S.n5795 0.001
R6804 S.t4 S.n5798 0.001
R6805 S.t25 S.n5593 0.001
R6806 S.t25 S.n5596 0.001
R6807 S.t8 S.n4771 0.001
R6808 S.t8 S.n4774 0.001
R6809 S.t54 S.n4179 0.001
R6810 S.t54 S.n4182 0.001
R6811 S.t10 S.n3749 0.001
R6812 S.t10 S.n3752 0.001
R6813 S.t42 S.n3893 0.001
R6814 S.t42 S.n3896 0.001
R6815 S.n3382 S.t12 0.001
R6816 S.n3390 S.n3385 0.001
R6817 S.t14 S.n3402 0.001
R6818 S.t14 S.n3405 0.001
R6819 S.t0 S.n2841 0.001
R6820 S.t0 S.n2844 0.001
R6821 S.n2864 S.t66 0.001
R6822 S.n2900 S.n2866 0.001
R6823 S.n3407 S.t14 0.001
R6824 S.n3415 S.n3407 0.001
R6825 S.t12 S.n3376 0.001
R6826 S.t12 S.n3379 0.001
R6827 S.t42 S.n3908 0.001
R6828 S.t42 S.n3911 0.001
R6829 S.t64 S.n5107 0.001
R6830 S.t64 S.n5110 0.001
R6831 S.t35 S.n4920 0.001
R6832 S.t35 S.n4917 0.001
R6833 S.n4917 S.n4914 0.001
R6834 S.t4 S.n5811 0.001
R6835 S.t4 S.n5814 0.001
R6836 S.t25 S.n5608 0.001
R6837 S.t25 S.n5611 0.001
R6838 S.t8 S.n4787 0.001
R6839 S.t8 S.n4790 0.001
R6840 S.t71 S.n4629 0.001
R6841 S.t71 S.n4632 0.001
R6842 S.t57 S.n4338 0.001
R6843 S.t57 S.n4341 0.001
R6844 S.t54 S.n4194 0.001
R6845 S.t54 S.n4197 0.001
R6846 S.t10 S.n3764 0.001
R6847 S.t10 S.n3767 0.001
R6848 S.n3913 S.t42 0.001
R6849 S.n3921 S.n3913 0.001
R6850 S.t10 S.n3784 0.001
R6851 S.t10 S.n3787 0.001
R6852 S.t54 S.n4389 0.001
R6853 S.t54 S.n4392 0.001
R6854 S.t64 S.n5123 0.001
R6855 S.t64 S.n5126 0.001
R6856 S.t35 S.n4905 0.001
R6857 S.t35 S.n4902 0.001
R6858 S.n4902 S.n4899 0.001
R6859 S.t4 S.n5827 0.001
R6860 S.t4 S.n5830 0.001
R6861 S.t25 S.n5623 0.001
R6862 S.t25 S.n5626 0.001
R6863 S.t8 S.n4803 0.001
R6864 S.t8 S.n4806 0.001
R6865 S.t71 S.n4644 0.001
R6866 S.t71 S.n4647 0.001
R6867 S.n4378 S.t57 0.001
R6868 S.n4385 S.n4378 0.001
R6869 S.n4394 S.t54 0.001
R6870 S.n4402 S.n4394 0.001
R6871 S.t57 S.n4358 0.001
R6872 S.t57 S.n4361 0.001
R6873 S.t71 S.n4843 0.001
R6874 S.t71 S.n4846 0.001
R6875 S.t64 S.n5139 0.001
R6876 S.t64 S.n5142 0.001
R6877 S.t35 S.n4890 0.001
R6878 S.t35 S.n4887 0.001
R6879 S.n4887 S.n4884 0.001
R6880 S.t4 S.n5843 0.001
R6881 S.t4 S.n5846 0.001
R6882 S.t25 S.n5638 0.001
R6883 S.t25 S.n5641 0.001
R6884 S.n4832 S.t8 0.001
R6885 S.n4839 S.n4832 0.001
R6886 S.n4848 S.t71 0.001
R6887 S.n4856 S.n4848 0.001
R6888 S.t8 S.n4826 0.001
R6889 S.t8 S.n4829 0.001
R6890 S.t25 S.n5874 0.001
R6891 S.t25 S.n5877 0.001
R6892 S.t64 S.n5155 0.001
R6893 S.t64 S.n5158 0.001
R6894 S.t35 S.n4875 0.001
R6895 S.t35 S.n4872 0.001
R6896 S.n4872 S.n4869 0.001
R6897 S.n5849 S.t4 0.001
R6898 S.n5857 S.n5852 0.001
R6899 S.n504 S.n503 0.001
R6900 S.n508 S.n507 0.001
R6901 S.n5278 S.n5276 0.001
R6902 S.n5457 S.n5456 0.001
R6903 S.n370 S.n369 0.001
R6904 S.n1217 S.n1216 0.001
R6905 S.n1253 S.n1252 0.001
R6906 S.n1839 S.n1838 0.001
R6907 S.n2879 S.n2871 0.001
R6908 S.n2930 S.n2929 0.001
R6909 S.n3445 S.n3444 0.001
R6910 S.n3951 S.n3950 0.001
R6911 S.n4422 S.n4421 0.001
R6912 S.n5288 S.n5287 0.001
R6913 S.n5343 S.n5316 0.001
R6914 S.n5343 S.n5314 0.001
R6915 S.n5343 S.n5312 0.001
R6916 S.n5343 S.n5310 0.001
R6917 S.n5343 S.n5308 0.001
R6918 S.n5343 S.n5306 0.001
R6919 S.n5343 S.n5304 0.001
R6920 S.n5040 S.n5039 0.001
R6921 S.n5021 S.n5018 0.001
R6922 S.n5260 S.n5257 0.001
R6923 S.n5900 S.n5880 0.001
R6924 S.n3326 S.n3323 0.001
R6925 S.n5512 S.n5509 0.001
R6926 S.n4501 S.n4498 0.001
R6927 S.n600 S.n587 0.001
R6928 S.n290 S.n282 0.001
R6929 S.n4066 S.n4063 0.001
R6930 S.n3594 S.n3591 0.001
R6931 S.n394 S.n386 0.001
R6932 S.n3103 S.n3100 0.001
R6933 S.n2570 S.n2567 0.001
R6934 S.n425 S.n417 0.001
R6935 S.n2073 S.n2070 0.001
R6936 S.n1534 S.n1531 0.001
R6937 S.n456 S.n448 0.001
R6938 S.n962 S.n959 0.001
R6939 S.n494 S.n481 0.001
R6940 S.n381 S.n378 0.001
R6941 S.n5194 S.n5184 0.001
R6942 S.n5732 S.n5729 0.001
R6943 S.n5532 S.n5529 0.001
R6944 S.n4521 S.n4511 0.001
R6945 S.n4538 S.n4535 0.001
R6946 S.n4086 S.n4076 0.001
R6947 S.n4103 S.n4100 0.001
R6948 S.n3800 S.n3790 0.001
R6949 S.n3817 S.n3814 0.001
R6950 S.n3123 S.n3113 0.001
R6951 S.n3140 S.n3137 0.001
R6952 S.n2590 S.n2580 0.001
R6953 S.n2607 S.n2604 0.001
R6954 S.n2093 S.n2083 0.001
R6955 S.n2110 S.n2107 0.001
R6956 S.n1749 S.n1739 0.001
R6957 S.n1766 S.n1763 0.001
R6958 S.n1186 S.n1176 0.001
R6959 S.n1198 S.n1195 0.001
R6960 S.n276 S.n273 0.001
R6961 S.n1222 S.n1204 0.001
R6962 S.n4988 S.n4984 0.001
R6963 S.n5747 S.n5744 0.001
R6964 S.n5548 S.n5545 0.001
R6965 S.n4564 S.n4560 0.001
R6966 S.n4569 S.n4566 0.001
R6967 S.n4129 S.n4125 0.001
R6968 S.n4134 S.n4131 0.001
R6969 S.n3843 S.n3839 0.001
R6970 S.n3848 S.n3845 0.001
R6971 S.n3166 S.n3162 0.001
R6972 S.n3171 S.n3168 0.001
R6973 S.n2633 S.n2629 0.001
R6974 S.n2638 S.n2635 0.001
R6975 S.n2139 S.n2135 0.001
R6976 S.n2141 S.n2121 0.001
R6977 S.n1792 S.n1788 0.001
R6978 S.n1796 S.n1793 0.001
R6979 S.n1170 S.n1167 0.001
R6980 S.n1809 S.n1804 0.001
R6981 S.n1733 S.n1730 0.001
R6982 S.n2346 S.n2343 0.001
R6983 S.n2342 S.n2338 0.001
R6984 S.n2653 S.n2650 0.001
R6985 S.n2821 S.n2818 0.001
R6986 S.n3186 S.n3183 0.001
R6987 S.n3340 S.n3337 0.001
R6988 S.n3863 S.n3860 0.001
R6989 S.n3717 S.n3714 0.001
R6990 S.n4149 S.n4146 0.001
R6991 S.n4306 S.n4303 0.001
R6992 S.n4584 S.n4581 0.001
R6993 S.n4739 S.n4736 0.001
R6994 S.n5563 S.n5560 0.001
R6995 S.n5763 S.n5760 0.001
R6996 S.n5059 S.n5056 0.001
R6997 S.n2359 S.n2354 0.001
R6998 S.n2329 S.n2326 0.001
R6999 S.n2858 S.n2855 0.001
R7000 S.n2854 S.n2850 0.001
R7001 S.n3201 S.n3198 0.001
R7002 S.n3356 S.n3353 0.001
R7003 S.n3878 S.n3875 0.001
R7004 S.n3733 S.n3730 0.001
R7005 S.n4164 S.n4161 0.001
R7006 S.n4322 S.n4319 0.001
R7007 S.n4599 S.n4596 0.001
R7008 S.n4755 S.n4752 0.001
R7009 S.n5578 S.n5575 0.001
R7010 S.n5779 S.n5776 0.001
R7011 S.n5075 S.n5072 0.001
R7012 S.n2900 S.n2864 0.001
R7013 S.n2841 S.n2838 0.001
R7014 S.n3402 S.n3399 0.001
R7015 S.n3390 S.n3382 0.001
R7016 S.n3893 S.n3890 0.001
R7017 S.n3749 S.n3746 0.001
R7018 S.n4179 S.n4176 0.001
R7019 S.n4614 S.n4611 0.001
R7020 S.n4771 S.n4768 0.001
R7021 S.n5593 S.n5590 0.001
R7022 S.n5795 S.n5792 0.001
R7023 S.n5091 S.n5088 0.001
R7024 S.n3415 S.n3410 0.001
R7025 S.n3376 S.n3373 0.001
R7026 S.n3908 S.n3905 0.001
R7027 S.n3764 S.n3761 0.001
R7028 S.n4194 S.n4191 0.001
R7029 S.n4338 S.n4335 0.001
R7030 S.n4629 S.n4626 0.001
R7031 S.n4787 S.n4784 0.001
R7032 S.n5608 S.n5605 0.001
R7033 S.n5811 S.n5808 0.001
R7034 S.n5107 S.n5104 0.001
R7035 S.n3921 S.n3916 0.001
R7036 S.n3784 S.n3781 0.001
R7037 S.n4389 S.n4386 0.001
R7038 S.n4385 S.n4381 0.001
R7039 S.n4644 S.n4641 0.001
R7040 S.n4803 S.n4800 0.001
R7041 S.n5623 S.n5620 0.001
R7042 S.n5827 S.n5824 0.001
R7043 S.n5123 S.n5120 0.001
R7044 S.n4402 S.n4397 0.001
R7045 S.n4358 S.n4355 0.001
R7046 S.n4843 S.n4840 0.001
R7047 S.n4839 S.n4835 0.001
R7048 S.n5638 S.n5635 0.001
R7049 S.n5843 S.n5840 0.001
R7050 S.n5139 S.n5136 0.001
R7051 S.n4856 S.n4851 0.001
R7052 S.n4826 S.n4823 0.001
R7053 S.n5874 S.n5871 0.001
R7054 S.n5857 S.n5849 0.001
R7055 S.n5155 S.n5152 0.001
R7056 S.n5041 S.n5040 0.001
R7057 S.t64 S.n5178 0.001
R7058 S.t64 S.n5181 0.001
R7059 S.n5178 S.n5175 0.001
R7060 S.t57 S.n4375 0.001
R7061 S.n4375 S.n4372 0.001
C0 DNW S 2936.40fF
C1 DNW G 6.22fF
C2 S G 1404.81fF
C3 DNW D 355.65fF
C4 S D 2210.84fF
C5 G D 1015.86fF
C6 D SUB -46.48fF
C7 G SUB -129.60fF
C8 S SUB 181.73fF $ **FLOATING
C9 DNW SUB 6933.01fF $ **FLOATING
C10 S.n0 SUB 0.95fF $ **FLOATING
C11 S.n1 SUB 0.93fF $ **FLOATING
C12 S.n2 SUB 0.34fF $ **FLOATING
C13 S.n3 SUB 0.46fF $ **FLOATING
C14 S.n4 SUB 0.33fF $ **FLOATING
C15 S.n5 SUB 0.18fF $ **FLOATING
C16 S.n6 SUB 0.09fF $ **FLOATING
C17 S.n7 SUB 0.76fF $ **FLOATING
C18 S.n8 SUB 0.21fF $ **FLOATING
C19 S.n9 SUB 0.35fF $ **FLOATING
C20 S.n10 SUB 0.53fF $ **FLOATING
C21 S.n11 SUB 0.12fF $ **FLOATING
C22 S.t613 SUB 0.02fF
C23 S.n12 SUB 0.14fF $ **FLOATING
C24 S.n14 SUB 0.64fF $ **FLOATING
C25 S.n15 SUB 0.43fF $ **FLOATING
C26 S.n16 SUB 1.60fF $ **FLOATING
C27 S.n17 SUB 0.49fF $ **FLOATING
C28 S.n18 SUB 0.45fF $ **FLOATING
C29 S.n19 SUB 0.45fF $ **FLOATING
C30 S.n20 SUB 1.82fF $ **FLOATING
C31 S.n21 SUB 0.12fF $ **FLOATING
C32 S.t936 SUB 0.02fF
C33 S.n22 SUB 0.14fF $ **FLOATING
C34 S.t18 SUB 0.02fF
C35 S.n24 SUB 0.24fF $ **FLOATING
C36 S.n25 SUB 0.35fF $ **FLOATING
C37 S.n26 SUB 0.60fF $ **FLOATING
C38 S.n27 SUB 2.46fF $ **FLOATING
C39 S.n28 SUB 2.00fF $ **FLOATING
C40 S.t553 SUB 0.02fF
C41 S.n29 SUB 0.24fF $ **FLOATING
C42 S.n30 SUB 0.90fF $ **FLOATING
C43 S.n31 SUB 0.05fF $ **FLOATING
C44 S.t1022 SUB 0.02fF
C45 S.n32 SUB 0.12fF $ **FLOATING
C46 S.n33 SUB 0.14fF $ **FLOATING
C47 S.n35 SUB 0.64fF $ **FLOATING
C48 S.n36 SUB 0.43fF $ **FLOATING
C49 S.n37 SUB 1.60fF $ **FLOATING
C50 S.n38 SUB 0.49fF $ **FLOATING
C51 S.n39 SUB 0.45fF $ **FLOATING
C52 S.n40 SUB 0.45fF $ **FLOATING
C53 S.n41 SUB 1.82fF $ **FLOATING
C54 S.n42 SUB 0.12fF $ **FLOATING
C55 S.t595 SUB 0.02fF
C56 S.n43 SUB 0.14fF $ **FLOATING
C57 S.t811 SUB 0.02fF
C58 S.n45 SUB 0.24fF $ **FLOATING
C59 S.n46 SUB 0.35fF $ **FLOATING
C60 S.n47 SUB 0.60fF $ **FLOATING
C61 S.n48 SUB 2.46fF $ **FLOATING
C62 S.n49 SUB 2.00fF $ **FLOATING
C63 S.t381 SUB 0.02fF
C64 S.n50 SUB 0.24fF $ **FLOATING
C65 S.n51 SUB 0.90fF $ **FLOATING
C66 S.n52 SUB 0.05fF $ **FLOATING
C67 S.t659 SUB 0.02fF
C68 S.n53 SUB 0.12fF $ **FLOATING
C69 S.n54 SUB 0.14fF $ **FLOATING
C70 S.n56 SUB 0.64fF $ **FLOATING
C71 S.n57 SUB 0.43fF $ **FLOATING
C72 S.n58 SUB 1.60fF $ **FLOATING
C73 S.n59 SUB 0.49fF $ **FLOATING
C74 S.n60 SUB 0.45fF $ **FLOATING
C75 S.n61 SUB 0.45fF $ **FLOATING
C76 S.n62 SUB 1.82fF $ **FLOATING
C77 S.n63 SUB 0.12fF $ **FLOATING
C78 S.t921 SUB 0.02fF
C79 S.n64 SUB 0.14fF $ **FLOATING
C80 S.t3 SUB 0.02fF
C81 S.n66 SUB 0.24fF $ **FLOATING
C82 S.n67 SUB 0.35fF $ **FLOATING
C83 S.n68 SUB 0.60fF $ **FLOATING
C84 S.n69 SUB 2.46fF $ **FLOATING
C85 S.n70 SUB 2.00fF $ **FLOATING
C86 S.t713 SUB 0.02fF
C87 S.n71 SUB 0.24fF $ **FLOATING
C88 S.n72 SUB 0.90fF $ **FLOATING
C89 S.n73 SUB 0.05fF $ **FLOATING
C90 S.t1017 SUB 0.02fF
C91 S.n74 SUB 0.12fF $ **FLOATING
C92 S.n75 SUB 0.14fF $ **FLOATING
C93 S.n77 SUB 1.87fF $ **FLOATING
C94 S.n78 SUB 0.12fF $ **FLOATING
C95 S.t292 SUB 0.02fF
C96 S.n79 SUB 0.14fF $ **FLOATING
C97 S.t1074 SUB 0.02fF
C98 S.n81 SUB 1.20fF $ **FLOATING
C99 S.n82 SUB 2.27fF $ **FLOATING
C100 S.n83 SUB 0.60fF $ **FLOATING
C101 S.n84 SUB 0.35fF $ **FLOATING
C102 S.n85 SUB 0.62fF $ **FLOATING
C103 S.n86 SUB 1.14fF $ **FLOATING
C104 S.n87 SUB 2.18fF $ **FLOATING
C105 S.n88 SUB 0.59fF $ **FLOATING
C106 S.n89 SUB 0.02fF $ **FLOATING
C107 S.n90 SUB 0.96fF $ **FLOATING
C108 S.t259 SUB 14.50fF
C109 S.n91 SUB 14.37fF $ **FLOATING
C110 S.n93 SUB 0.37fF $ **FLOATING
C111 S.n94 SUB 0.23fF $ **FLOATING
C112 S.n95 SUB 2.86fF $ **FLOATING
C113 S.n96 SUB 2.43fF $ **FLOATING
C114 S.n97 SUB 4.25fF $ **FLOATING
C115 S.n98 SUB 0.25fF $ **FLOATING
C116 S.n99 SUB 0.01fF $ **FLOATING
C117 S.t991 SUB 0.02fF
C118 S.n100 SUB 0.25fF $ **FLOATING
C119 S.t705 SUB 0.02fF
C120 S.n101 SUB 0.94fF $ **FLOATING
C121 S.n102 SUB 0.70fF $ **FLOATING
C122 S.n103 SUB 1.87fF $ **FLOATING
C123 S.n104 SUB 1.76fF $ **FLOATING
C124 S.n105 SUB 0.12fF $ **FLOATING
C125 S.t655 SUB 0.02fF
C126 S.n106 SUB 0.14fF $ **FLOATING
C127 S.t692 SUB 0.02fF
C128 S.n108 SUB 0.24fF $ **FLOATING
C129 S.n109 SUB 0.35fF $ **FLOATING
C130 S.n110 SUB 0.60fF $ **FLOATING
C131 S.n111 SUB 2.71fF $ **FLOATING
C132 S.n112 SUB 2.03fF $ **FLOATING
C133 S.t327 SUB 0.02fF
C134 S.n113 SUB 0.24fF $ **FLOATING
C135 S.n114 SUB 0.90fF $ **FLOATING
C136 S.n115 SUB 0.05fF $ **FLOATING
C137 S.t961 SUB 0.02fF
C138 S.n116 SUB 0.12fF $ **FLOATING
C139 S.n117 SUB 0.14fF $ **FLOATING
C140 S.n119 SUB 1.23fF $ **FLOATING
C141 S.n120 SUB 1.27fF $ **FLOATING
C142 S.n121 SUB 1.86fF $ **FLOATING
C143 S.n122 SUB 0.12fF $ **FLOATING
C144 S.t1059 SUB 0.02fF
C145 S.n123 SUB 0.14fF $ **FLOATING
C146 S.t742 SUB 0.02fF
C147 S.n125 SUB 0.24fF $ **FLOATING
C148 S.n126 SUB 0.35fF $ **FLOATING
C149 S.n127 SUB 0.60fF $ **FLOATING
C150 S.n128 SUB 2.72fF $ **FLOATING
C151 S.n129 SUB 2.14fF $ **FLOATING
C152 S.t447 SUB 0.02fF
C153 S.n130 SUB 0.24fF $ **FLOATING
C154 S.n131 SUB 0.90fF $ **FLOATING
C155 S.n132 SUB 0.05fF $ **FLOATING
C156 S.t578 SUB 0.02fF
C157 S.n133 SUB 0.12fF $ **FLOATING
C158 S.n134 SUB 0.14fF $ **FLOATING
C159 S.n136 SUB 1.87fF $ **FLOATING
C160 S.n137 SUB 1.77fF $ **FLOATING
C161 S.n138 SUB 0.12fF $ **FLOATING
C162 S.t680 SUB 0.02fF
C163 S.n139 SUB 0.14fF $ **FLOATING
C164 S.t357 SUB 0.02fF
C165 S.n141 SUB 0.24fF $ **FLOATING
C166 S.n142 SUB 0.35fF $ **FLOATING
C167 S.n143 SUB 0.60fF $ **FLOATING
C168 S.n144 SUB 2.70fF $ **FLOATING
C169 S.n145 SUB 2.03fF $ **FLOATING
C170 S.t27 SUB 0.02fF
C171 S.n146 SUB 0.24fF $ **FLOATING
C172 S.n147 SUB 0.90fF $ **FLOATING
C173 S.n148 SUB 0.05fF $ **FLOATING
C174 S.t1011 SUB 0.02fF
C175 S.n149 SUB 0.12fF $ **FLOATING
C176 S.n150 SUB 0.14fF $ **FLOATING
C177 S.n152 SUB 1.23fF $ **FLOATING
C178 S.n153 SUB 1.27fF $ **FLOATING
C179 S.n154 SUB 1.86fF $ **FLOATING
C180 S.n155 SUB 0.12fF $ **FLOATING
C181 S.t309 SUB 0.02fF
C182 S.n156 SUB 0.14fF $ **FLOATING
C183 S.t1084 SUB 0.02fF
C184 S.n158 SUB 0.24fF $ **FLOATING
C185 S.n159 SUB 0.35fF $ **FLOATING
C186 S.n160 SUB 0.60fF $ **FLOATING
C187 S.n161 SUB 2.72fF $ **FLOATING
C188 S.n162 SUB 2.14fF $ **FLOATING
C189 S.t776 SUB 0.02fF
C190 S.n163 SUB 0.24fF $ **FLOATING
C191 S.n164 SUB 0.90fF $ **FLOATING
C192 S.n165 SUB 0.05fF $ **FLOATING
C193 S.t638 SUB 0.02fF
C194 S.n166 SUB 0.12fF $ **FLOATING
C195 S.n167 SUB 0.14fF $ **FLOATING
C196 S.n169 SUB 1.87fF $ **FLOATING
C197 S.n170 SUB 1.77fF $ **FLOATING
C198 S.n171 SUB 0.12fF $ **FLOATING
C199 S.t1039 SUB 0.02fF
C200 S.n172 SUB 0.14fF $ **FLOATING
C201 S.t696 SUB 0.02fF
C202 S.n174 SUB 0.24fF $ **FLOATING
C203 S.n175 SUB 0.35fF $ **FLOATING
C204 S.n176 SUB 0.60fF $ **FLOATING
C205 S.n177 SUB 2.70fF $ **FLOATING
C206 S.n178 SUB 2.03fF $ **FLOATING
C207 S.t389 SUB 0.02fF
C208 S.n179 SUB 0.24fF $ **FLOATING
C209 S.n180 SUB 0.90fF $ **FLOATING
C210 S.n181 SUB 0.05fF $ **FLOATING
C211 S.t256 SUB 0.02fF
C212 S.n182 SUB 0.12fF $ **FLOATING
C213 S.n183 SUB 0.14fF $ **FLOATING
C214 S.n185 SUB 1.23fF $ **FLOATING
C215 S.n186 SUB 1.27fF $ **FLOATING
C216 S.n187 SUB 1.86fF $ **FLOATING
C217 S.n188 SUB 0.12fF $ **FLOATING
C218 S.t662 SUB 0.02fF
C219 S.n189 SUB 0.14fF $ **FLOATING
C220 S.t316 SUB 0.02fF
C221 S.n191 SUB 0.24fF $ **FLOATING
C222 S.n192 SUB 0.35fF $ **FLOATING
C223 S.n193 SUB 0.60fF $ **FLOATING
C224 S.n194 SUB 2.72fF $ **FLOATING
C225 S.n195 SUB 2.14fF $ **FLOATING
C226 S.t1111 SUB 0.02fF
C227 S.n196 SUB 0.24fF $ **FLOATING
C228 S.n197 SUB 0.90fF $ **FLOATING
C229 S.n198 SUB 0.05fF $ **FLOATING
C230 S.t978 SUB 0.02fF
C231 S.n199 SUB 0.12fF $ **FLOATING
C232 S.n200 SUB 0.14fF $ **FLOATING
C233 S.n202 SUB 2.58fF $ **FLOATING
C234 S.n203 SUB 1.86fF $ **FLOATING
C235 S.n204 SUB 0.12fF $ **FLOATING
C236 S.t1020 SUB 0.02fF
C237 S.n205 SUB 0.14fF $ **FLOATING
C238 S.t670 SUB 0.02fF
C239 S.n207 SUB 0.24fF $ **FLOATING
C240 S.n208 SUB 0.35fF $ **FLOATING
C241 S.n209 SUB 0.60fF $ **FLOATING
C242 S.n210 SUB 0.89fF $ **FLOATING
C243 S.n211 SUB 0.76fF $ **FLOATING
C244 S.n212 SUB 0.96fF $ **FLOATING
C245 S.n213 SUB 0.09fF $ **FLOATING
C246 S.n214 SUB 0.32fF $ **FLOATING
C247 S.n215 SUB 2.13fF $ **FLOATING
C248 S.t339 SUB 0.02fF
C249 S.n216 SUB 0.24fF $ **FLOATING
C250 S.n217 SUB 0.90fF $ **FLOATING
C251 S.n218 SUB 0.05fF $ **FLOATING
C252 S.t278 SUB 0.02fF
C253 S.n219 SUB 0.12fF $ **FLOATING
C254 S.n220 SUB 0.14fF $ **FLOATING
C255 S.n222 SUB 2.27fF $ **FLOATING
C256 S.n223 SUB 1.86fF $ **FLOATING
C257 S.n224 SUB 0.12fF $ **FLOATING
C258 S.t646 SUB 0.02fF
C259 S.n225 SUB 0.14fF $ **FLOATING
C260 S.t299 SUB 0.02fF
C261 S.n227 SUB 0.24fF $ **FLOATING
C262 S.n228 SUB 0.35fF $ **FLOATING
C263 S.n229 SUB 0.60fF $ **FLOATING
C264 S.n230 SUB 0.76fF $ **FLOATING
C265 S.n231 SUB 0.48fF $ **FLOATING
C266 S.n232 SUB 0.09fF $ **FLOATING
C267 S.n233 SUB 0.32fF $ **FLOATING
C268 S.n234 SUB 2.00fF $ **FLOATING
C269 S.t1067 SUB 0.02fF
C270 S.n235 SUB 0.24fF $ **FLOATING
C271 S.n236 SUB 0.90fF $ **FLOATING
C272 S.n237 SUB 0.05fF $ **FLOATING
C273 S.t997 SUB 0.02fF
C274 S.n238 SUB 0.12fF $ **FLOATING
C275 S.n239 SUB 0.14fF $ **FLOATING
C276 S.n241 SUB 1.87fF $ **FLOATING
C277 S.n242 SUB 0.25fF $ **FLOATING
C278 S.n243 SUB 0.09fF $ **FLOATING
C279 S.n244 SUB 0.22fF $ **FLOATING
C280 S.n245 SUB 1.14fF $ **FLOATING
C281 S.n246 SUB 0.22fF $ **FLOATING
C282 S.n247 SUB 0.12fF $ **FLOATING
C283 S.t271 SUB 0.02fF
C284 S.n248 SUB 0.14fF $ **FLOATING
C285 S.t1030 SUB 0.02fF
C286 S.n250 SUB 0.24fF $ **FLOATING
C287 S.n251 SUB 0.35fF $ **FLOATING
C288 S.n252 SUB 0.60fF $ **FLOATING
C289 S.n253 SUB 2.70fF $ **FLOATING
C290 S.n254 SUB 1.86fF $ **FLOATING
C291 S.t684 SUB 0.02fF
C292 S.n255 SUB 0.24fF $ **FLOATING
C293 S.n256 SUB 0.90fF $ **FLOATING
C294 S.n257 SUB 0.05fF $ **FLOATING
C295 S.t622 SUB 0.02fF
C296 S.n258 SUB 0.12fF $ **FLOATING
C297 S.n259 SUB 0.14fF $ **FLOATING
C298 S.n261 SUB 14.09fF $ **FLOATING
C299 S.n262 SUB 2.69fF $ **FLOATING
C300 S.n263 SUB 1.93fF $ **FLOATING
C301 S.n264 SUB 0.12fF $ **FLOATING
C302 S.t718 SUB 0.02fF
C303 S.n265 SUB 0.14fF $ **FLOATING
C304 S.t679 SUB 0.02fF
C305 S.n267 SUB 0.24fF $ **FLOATING
C306 S.n268 SUB 0.35fF $ **FLOATING
C307 S.n269 SUB 0.60fF $ **FLOATING
C308 S.n270 SUB 1.55fF $ **FLOATING
C309 S.n271 SUB 0.70fF $ **FLOATING
C310 S.n272 SUB 0.28fF $ **FLOATING
C311 S.n273 SUB 2.08fF $ **FLOATING
C312 S.t1051 SUB 0.02fF
C313 S.n274 SUB 0.12fF $ **FLOATING
C314 S.n275 SUB 0.14fF $ **FLOATING
C315 S.t1117 SUB 0.02fF
C316 S.n277 SUB 0.24fF $ **FLOATING
C317 S.n278 SUB 0.90fF $ **FLOATING
C318 S.n279 SUB 0.05fF $ **FLOATING
C319 S.t255 SUB 32.35fF
C320 S.t652 SUB 0.02fF
C321 S.n280 SUB 0.12fF $ **FLOATING
C322 S.n281 SUB 0.14fF $ **FLOATING
C323 S.t721 SUB 0.02fF
C324 S.n283 SUB 0.24fF $ **FLOATING
C325 S.n284 SUB 0.90fF $ **FLOATING
C326 S.n285 SUB 0.05fF $ **FLOATING
C327 S.t1047 SUB 0.02fF
C328 S.n286 SUB 0.24fF $ **FLOATING
C329 S.n287 SUB 0.35fF $ **FLOATING
C330 S.n288 SUB 0.60fF $ **FLOATING
C331 S.n289 SUB 2.21fF $ **FLOATING
C332 S.n290 SUB 2.67fF $ **FLOATING
C333 S.n291 SUB 2.62fF $ **FLOATING
C334 S.n292 SUB 2.34fF $ **FLOATING
C335 S.n293 SUB 1.82fF $ **FLOATING
C336 S.n294 SUB 0.12fF $ **FLOATING
C337 S.t225 SUB 0.02fF
C338 S.n295 SUB 0.14fF $ **FLOATING
C339 S.t457 SUB 0.02fF
C340 S.n297 SUB 0.24fF $ **FLOATING
C341 S.n298 SUB 0.35fF $ **FLOATING
C342 S.n299 SUB 0.60fF $ **FLOATING
C343 S.n300 SUB 0.66fF $ **FLOATING
C344 S.n301 SUB 0.40fF $ **FLOATING
C345 S.n302 SUB 0.54fF $ **FLOATING
C346 S.n303 SUB 0.32fF $ **FLOATING
C347 S.n304 SUB 1.06fF $ **FLOATING
C348 S.n305 SUB 2.11fF $ **FLOATING
C349 S.t1128 SUB 0.02fF
C350 S.n306 SUB 0.24fF $ **FLOATING
C351 S.n307 SUB 0.90fF $ **FLOATING
C352 S.n308 SUB 0.05fF $ **FLOATING
C353 S.t263 SUB 0.02fF
C354 S.n309 SUB 0.12fF $ **FLOATING
C355 S.n310 SUB 0.14fF $ **FLOATING
C356 S.n312 SUB 0.25fF $ **FLOATING
C357 S.n313 SUB 0.09fF $ **FLOATING
C358 S.n314 SUB 0.12fF $ **FLOATING
C359 S.t569 SUB 0.02fF
C360 S.n315 SUB 0.14fF $ **FLOATING
C361 S.t793 SUB 0.02fF
C362 S.n317 SUB 0.24fF $ **FLOATING
C363 S.n318 SUB 0.35fF $ **FLOATING
C364 S.n319 SUB 0.60fF $ **FLOATING
C365 S.n320 SUB 0.82fF $ **FLOATING
C366 S.n321 SUB 0.31fF $ **FLOATING
C367 S.n322 SUB 0.29fF $ **FLOATING
C368 S.n323 SUB 0.25fF $ **FLOATING
C369 S.n324 SUB 0.22fF $ **FLOATING
C370 S.n325 SUB 0.60fF $ **FLOATING
C371 S.n326 SUB 0.27fF $ **FLOATING
C372 S.n327 SUB 1.92fF $ **FLOATING
C373 S.t358 SUB 0.02fF
C374 S.n328 SUB 0.24fF $ **FLOATING
C375 S.n329 SUB 0.90fF $ **FLOATING
C376 S.n330 SUB 0.05fF $ **FLOATING
C377 S.t606 SUB 0.02fF
C378 S.n331 SUB 0.12fF $ **FLOATING
C379 S.n332 SUB 0.14fF $ **FLOATING
C380 S.n334 SUB 0.19fF $ **FLOATING
C381 S.n335 SUB 0.09fF $ **FLOATING
C382 S.n336 SUB 0.67fF $ **FLOATING
C383 S.n337 SUB 0.28fF $ **FLOATING
C384 S.n338 SUB 1.72fF $ **FLOATING
C385 S.n339 SUB 0.21fF $ **FLOATING
C386 S.n340 SUB 1.82fF $ **FLOATING
C387 S.n341 SUB 0.12fF $ **FLOATING
C388 S.t540 SUB 0.02fF
C389 S.n342 SUB 0.14fF $ **FLOATING
C390 S.t1073 SUB 0.02fF
C391 S.n344 SUB 0.24fF $ **FLOATING
C392 S.n345 SUB 0.35fF $ **FLOATING
C393 S.n346 SUB 0.60fF $ **FLOATING
C394 S.n347 SUB 2.46fF $ **FLOATING
C395 S.n348 SUB 1.84fF $ **FLOATING
C396 S.t839 SUB 0.02fF
C397 S.n349 SUB 0.24fF $ **FLOATING
C398 S.n350 SUB 0.90fF $ **FLOATING
C399 S.n351 SUB 0.05fF $ **FLOATING
C400 S.t215 SUB 0.02fF
C401 S.n352 SUB 0.12fF $ **FLOATING
C402 S.n353 SUB 0.14fF $ **FLOATING
C403 S.n355 SUB 14.09fF $ **FLOATING
C404 S.n356 SUB 1.12fF $ **FLOATING
C405 S.n357 SUB 8.87fF $ **FLOATING
C406 S.n358 SUB 20.14fF $ **FLOATING
C407 S.n359 SUB 8.87fF $ **FLOATING
C408 S.n360 SUB 20.14fF $ **FLOATING
C409 S.n361 SUB 0.59fF $ **FLOATING
C410 S.n362 SUB 0.21fF $ **FLOATING
C411 S.n363 SUB 0.87fF $ **FLOATING
C412 S.n364 SUB 0.87fF $ **FLOATING
C413 S.n365 SUB 2.57fF $ **FLOATING
C414 S.n366 SUB 0.29fF $ **FLOATING
C415 S.t2 SUB 14.50fF
C416 S.n367 SUB 15.77fF $ **FLOATING
C417 S.n368 SUB 0.21fF $ **FLOATING
C418 S.n369 SUB 1.40fF $ **FLOATING
C419 S.n370 SUB 4.20fF $ **FLOATING
C420 S.n371 SUB 1.78fF $ **FLOATING
C421 S.t822 SUB 0.02fF
C422 S.n372 SUB 0.63fF $ **FLOATING
C423 S.n373 SUB 0.60fF $ **FLOATING
C424 S.n374 SUB 1.19fF $ **FLOATING
C425 S.n375 SUB 0.36fF $ **FLOATING
C426 S.n376 SUB 1.17fF $ **FLOATING
C427 S.n377 SUB 0.38fF $ **FLOATING
C428 S.n378 SUB 4.17fF $ **FLOATING
C429 S.t219 SUB 0.02fF
C430 S.n379 SUB 0.01fF $ **FLOATING
C431 S.n380 SUB 0.25fF $ **FLOATING
C432 S.t397 SUB 0.02fF
C433 S.n382 SUB 1.18fF $ **FLOATING
C434 S.n383 SUB 0.05fF $ **FLOATING
C435 S.t198 SUB 31.97fF
C436 S.t643 SUB 0.02fF
C437 S.n384 SUB 0.12fF $ **FLOATING
C438 S.n385 SUB 0.14fF $ **FLOATING
C439 S.t409 SUB 0.02fF
C440 S.n387 SUB 0.24fF $ **FLOATING
C441 S.n388 SUB 0.90fF $ **FLOATING
C442 S.n389 SUB 0.05fF $ **FLOATING
C443 S.t831 SUB 0.02fF
C444 S.n390 SUB 0.24fF $ **FLOATING
C445 S.n391 SUB 0.35fF $ **FLOATING
C446 S.n392 SUB 0.60fF $ **FLOATING
C447 S.n393 SUB 2.45fF $ **FLOATING
C448 S.n394 SUB 1.94fF $ **FLOATING
C449 S.n395 SUB 1.48fF $ **FLOATING
C450 S.n396 SUB 2.60fF $ **FLOATING
C451 S.n397 SUB 8.87fF $ **FLOATING
C452 S.n398 SUB 8.87fF $ **FLOATING
C453 S.n399 SUB 5.32fF $ **FLOATING
C454 S.n400 SUB 2.15fF $ **FLOATING
C455 S.n401 SUB 0.95fF $ **FLOATING
C456 S.n402 SUB 0.93fF $ **FLOATING
C457 S.n403 SUB 0.34fF $ **FLOATING
C458 S.n404 SUB 0.46fF $ **FLOATING
C459 S.n405 SUB 0.33fF $ **FLOATING
C460 S.n406 SUB 0.18fF $ **FLOATING
C461 S.n407 SUB 0.09fF $ **FLOATING
C462 S.n408 SUB 0.76fF $ **FLOATING
C463 S.n409 SUB 0.21fF $ **FLOATING
C464 S.n410 SUB 0.35fF $ **FLOATING
C465 S.n411 SUB 0.53fF $ **FLOATING
C466 S.n412 SUB 0.12fF $ **FLOATING
C467 S.t199 SUB 0.02fF
C468 S.n413 SUB 0.14fF $ **FLOATING
C469 S.t290 SUB 0.02fF
C470 S.n415 SUB 0.12fF $ **FLOATING
C471 S.n416 SUB 0.14fF $ **FLOATING
C472 S.t1102 SUB 0.02fF
C473 S.n418 SUB 0.24fF $ **FLOATING
C474 S.n419 SUB 0.90fF $ **FLOATING
C475 S.n420 SUB 0.05fF $ **FLOATING
C476 S.t436 SUB 0.02fF
C477 S.n421 SUB 0.24fF $ **FLOATING
C478 S.n422 SUB 0.35fF $ **FLOATING
C479 S.n423 SUB 0.60fF $ **FLOATING
C480 S.n424 SUB 2.45fF $ **FLOATING
C481 S.n425 SUB 1.94fF $ **FLOATING
C482 S.n426 SUB 1.48fF $ **FLOATING
C483 S.n427 SUB 2.60fF $ **FLOATING
C484 S.n428 SUB 8.87fF $ **FLOATING
C485 S.n429 SUB 8.87fF $ **FLOATING
C486 S.n430 SUB 5.32fF $ **FLOATING
C487 S.n431 SUB 2.15fF $ **FLOATING
C488 S.n432 SUB 0.95fF $ **FLOATING
C489 S.n433 SUB 0.93fF $ **FLOATING
C490 S.n434 SUB 0.34fF $ **FLOATING
C491 S.n435 SUB 0.46fF $ **FLOATING
C492 S.n436 SUB 0.33fF $ **FLOATING
C493 S.n437 SUB 0.18fF $ **FLOATING
C494 S.n438 SUB 0.09fF $ **FLOATING
C495 S.n439 SUB 0.76fF $ **FLOATING
C496 S.n440 SUB 0.21fF $ **FLOATING
C497 S.n441 SUB 0.35fF $ **FLOATING
C498 S.n442 SUB 0.53fF $ **FLOATING
C499 S.n443 SUB 0.12fF $ **FLOATING
C500 S.t973 SUB 0.02fF
C501 S.n444 SUB 0.14fF $ **FLOATING
C502 S.t1035 SUB 0.02fF
C503 S.n446 SUB 0.12fF $ **FLOATING
C504 S.n447 SUB 0.14fF $ **FLOATING
C505 S.t766 SUB 0.02fF
C506 S.n449 SUB 0.24fF $ **FLOATING
C507 S.n450 SUB 0.90fF $ **FLOATING
C508 S.n451 SUB 0.05fF $ **FLOATING
C509 S.t77 SUB 0.02fF
C510 S.n452 SUB 0.24fF $ **FLOATING
C511 S.n453 SUB 0.35fF $ **FLOATING
C512 S.n454 SUB 0.60fF $ **FLOATING
C513 S.n455 SUB 2.45fF $ **FLOATING
C514 S.n456 SUB 1.94fF $ **FLOATING
C515 S.n457 SUB 1.48fF $ **FLOATING
C516 S.n458 SUB 2.60fF $ **FLOATING
C517 S.n459 SUB 8.87fF $ **FLOATING
C518 S.n460 SUB 8.87fF $ **FLOATING
C519 S.n461 SUB 5.32fF $ **FLOATING
C520 S.n462 SUB 2.15fF $ **FLOATING
C521 S.n463 SUB 13.46fF $ **FLOATING
C522 S.n464 SUB 13.46fF $ **FLOATING
C523 S.n465 SUB 5.27fF $ **FLOATING
C524 S.n466 SUB 2.02fF $ **FLOATING
C525 S.n467 SUB 16.29fF $ **FLOATING
C526 S.n468 SUB 0.06fF $ **FLOATING
C527 S.n469 SUB 0.20fF $ **FLOATING
C528 S.n470 SUB 0.09fF $ **FLOATING
C529 S.n471 SUB 0.20fF $ **FLOATING
C530 S.n472 SUB 0.09fF $ **FLOATING
C531 S.n473 SUB 0.30fF $ **FLOATING
C532 S.n474 SUB 0.99fF $ **FLOATING
C533 S.n475 SUB 0.44fF $ **FLOATING
C534 S.n476 SUB 0.12fF $ **FLOATING
C535 S.t211 SUB 0.02fF
C536 S.n477 SUB 0.14fF $ **FLOATING
C537 S.t252 SUB 0.02fF
C538 S.n479 SUB 0.12fF $ **FLOATING
C539 S.n480 SUB 0.14fF $ **FLOATING
C540 S.t931 SUB 0.02fF
C541 S.n482 SUB 0.24fF $ **FLOATING
C542 S.n483 SUB 0.90fF $ **FLOATING
C543 S.n484 SUB 0.05fF $ **FLOATING
C544 S.t442 SUB 0.02fF
C545 S.n485 SUB 0.24fF $ **FLOATING
C546 S.n486 SUB 0.35fF $ **FLOATING
C547 S.n487 SUB 0.60fF $ **FLOATING
C548 S.n488 SUB 0.78fF $ **FLOATING
C549 S.n489 SUB 0.18fF $ **FLOATING
C550 S.n490 SUB 0.39fF $ **FLOATING
C551 S.n491 SUB 0.44fF $ **FLOATING
C552 S.n492 SUB 0.25fF $ **FLOATING
C553 S.n493 SUB 0.09fF $ **FLOATING
C554 S.n494 SUB 1.79fF $ **FLOATING
C555 S.n495 SUB 1.93fF $ **FLOATING
C556 S.n496 SUB 2.60fF $ **FLOATING
C557 S.n497 SUB 0.95fF $ **FLOATING
C558 S.n498 SUB 0.34fF $ **FLOATING
C559 S.n499 SUB 0.43fF $ **FLOATING
C560 S.n500 SUB 0.30fF $ **FLOATING
C561 S.n501 SUB 0.95fF $ **FLOATING
C562 S.t112 SUB 0.02fF
C563 S.n502 SUB 1.29fF $ **FLOATING
C564 S.n503 SUB 38.81fF $ **FLOATING
C565 S.n504 SUB 2.20fF $ **FLOATING
C566 S.n505 SUB 0.35fF $ **FLOATING
C567 S.n506 SUB 0.62fF $ **FLOATING
C568 S.n507 SUB 0.52fF $ **FLOATING
C569 S.n508 SUB 3.62fF $ **FLOATING
C570 S.n509 SUB 4.21fF $ **FLOATING
C571 S.n510 SUB 4.17fF $ **FLOATING
C572 S.n511 SUB 4.17fF $ **FLOATING
C573 S.n512 SUB 4.17fF $ **FLOATING
C574 S.n513 SUB 4.65fF $ **FLOATING
C575 S.n514 SUB 4.25fF $ **FLOATING
C576 S.n515 SUB 4.23fF $ **FLOATING
C577 S.n516 SUB 85.92fF $ **FLOATING
C578 S.n517 SUB 2.17fF $ **FLOATING
C579 S.n518 SUB 12.76fF $ **FLOATING
C580 S.n519 SUB 1.87fF $ **FLOATING
C581 S.n520 SUB 9.30fF $ **FLOATING
C582 S.n521 SUB 0.25fF $ **FLOATING
C583 S.t1078 SUB 0.02fF
C584 S.n522 SUB 0.43fF $ **FLOATING
C585 S.n523 SUB 8.87fF $ **FLOATING
C586 S.n524 SUB 8.87fF $ **FLOATING
C587 S.n525 SUB 5.40fF $ **FLOATING
C588 S.n526 SUB 1.94fF $ **FLOATING
C589 S.t324 SUB 0.02fF
C590 S.n527 SUB 0.88fF $ **FLOATING
C591 S.t672 SUB 0.02fF
C592 S.n528 SUB 0.88fF $ **FLOATING
C593 S.n529 SUB 9.33fF $ **FLOATING
C594 S.n530 SUB 3.23fF $ **FLOATING
C595 S.n531 SUB 0.38fF $ **FLOATING
C596 S.n532 SUB 0.30fF $ **FLOATING
C597 S.n533 SUB 0.99fF $ **FLOATING
C598 S.n534 SUB 0.02fF $ **FLOATING
C599 S.t1112 SUB 0.02fF
C600 S.n535 SUB 0.36fF $ **FLOATING
C601 S.n536 SUB 8.87fF $ **FLOATING
C602 S.n537 SUB 8.87fF $ **FLOATING
C603 S.n538 SUB 5.40fF $ **FLOATING
C604 S.n539 SUB 1.94fF $ **FLOATING
C605 S.t675 SUB 0.02fF
C606 S.n540 SUB 0.88fF $ **FLOATING
C607 S.t1003 SUB 0.02fF
C608 S.n541 SUB 0.88fF $ **FLOATING
C609 S.n542 SUB 3.23fF $ **FLOATING
C610 S.n543 SUB 0.38fF $ **FLOATING
C611 S.n544 SUB 0.30fF $ **FLOATING
C612 S.n545 SUB 0.99fF $ **FLOATING
C613 S.n546 SUB 0.02fF $ **FLOATING
C614 S.t343 SUB 0.02fF
C615 S.n547 SUB 0.36fF $ **FLOATING
C616 S.n548 SUB 8.87fF $ **FLOATING
C617 S.n549 SUB 8.87fF $ **FLOATING
C618 S.n550 SUB 5.40fF $ **FLOATING
C619 S.n551 SUB 1.94fF $ **FLOATING
C620 S.t1032 SUB 0.02fF
C621 S.n552 SUB 0.88fF $ **FLOATING
C622 S.t242 SUB 0.02fF
C623 S.n553 SUB 0.88fF $ **FLOATING
C624 S.n554 SUB 3.23fF $ **FLOATING
C625 S.n555 SUB 0.38fF $ **FLOATING
C626 S.n556 SUB 0.30fF $ **FLOATING
C627 S.n557 SUB 0.99fF $ **FLOATING
C628 S.n558 SUB 0.02fF $ **FLOATING
C629 S.t685 SUB 0.02fF
C630 S.n559 SUB 0.36fF $ **FLOATING
C631 S.n560 SUB 0.30fF $ **FLOATING
C632 S.n561 SUB 8.87fF $ **FLOATING
C633 S.n562 SUB 8.87fF $ **FLOATING
C634 S.n563 SUB 5.16fF $ **FLOATING
C635 S.n564 SUB 0.99fF $ **FLOATING
C636 S.n565 SUB 0.35fF $ **FLOATING
C637 S.t286 SUB 0.02fF
C638 S.n566 SUB 0.88fF $ **FLOATING
C639 S.t644 SUB 0.02fF
C640 S.n567 SUB 0.88fF $ **FLOATING
C641 S.n568 SUB 3.23fF $ **FLOATING
C642 S.n569 SUB 0.27fF $ **FLOATING
C643 S.n570 SUB 1.04fF $ **FLOATING
C644 S.n571 SUB 1.13fF $ **FLOATING
C645 S.n572 SUB 0.42fF $ **FLOATING
C646 S.n573 SUB 0.02fF $ **FLOATING
C647 S.t1044 SUB 0.02fF
C648 S.n574 SUB 0.36fF $ **FLOATING
C649 S.n575 SUB 0.37fF $ **FLOATING
C650 S.n576 SUB 0.82fF $ **FLOATING
C651 S.t1014 SUB 0.02fF
C652 S.n577 SUB 0.88fF $ **FLOATING
C653 S.t265 SUB 0.02fF
C654 S.n578 SUB 0.88fF $ **FLOATING
C655 S.n579 SUB 0.04fF $ **FLOATING
C656 S.n580 SUB 0.48fF $ **FLOATING
C657 S.n581 SUB 0.37fF $ **FLOATING
C658 S.n582 SUB 0.12fF $ **FLOATING
C659 S.t947 SUB 0.02fF
C660 S.n583 SUB 0.14fF $ **FLOATING
C661 S.t983 SUB 0.02fF
C662 S.n585 SUB 0.12fF $ **FLOATING
C663 S.n586 SUB 0.14fF $ **FLOATING
C664 S.t744 SUB 0.02fF
C665 S.n588 SUB 0.24fF $ **FLOATING
C666 S.n589 SUB 0.90fF $ **FLOATING
C667 S.n590 SUB 0.05fF $ **FLOATING
C668 S.t50 SUB 0.02fF
C669 S.n591 SUB 0.24fF $ **FLOATING
C670 S.n592 SUB 0.35fF $ **FLOATING
C671 S.n593 SUB 0.60fF $ **FLOATING
C672 S.n594 SUB 0.35fF $ **FLOATING
C673 S.n595 SUB 0.53fF $ **FLOATING
C674 S.n596 SUB 0.38fF $ **FLOATING
C675 S.n597 SUB 0.18fF $ **FLOATING
C676 S.n598 SUB 0.25fF $ **FLOATING
C677 S.n599 SUB 0.09fF $ **FLOATING
C678 S.n600 SUB 1.94fF $ **FLOATING
C679 S.n601 SUB 1.48fF $ **FLOATING
C680 S.n602 SUB 2.60fF $ **FLOATING
C681 S.n603 SUB 8.87fF $ **FLOATING
C682 S.n604 SUB 8.87fF $ **FLOATING
C683 S.n605 SUB 5.69fF $ **FLOATING
C684 S.n606 SUB 0.03fF $ **FLOATING
C685 S.n607 SUB 0.03fF $ **FLOATING
C686 S.n608 SUB 0.10fF $ **FLOATING
C687 S.n609 SUB 0.36fF $ **FLOATING
C688 S.n610 SUB 0.37fF $ **FLOATING
C689 S.n611 SUB 0.10fF $ **FLOATING
C690 S.n612 SUB 0.12fF $ **FLOATING
C691 S.n613 SUB 0.03fF $ **FLOATING
C692 S.n614 SUB 0.07fF $ **FLOATING
C693 S.n615 SUB 1.39fF $ **FLOATING
C694 S.n616 SUB 1.75fF $ **FLOATING
C695 S.n617 SUB 1.12fF $ **FLOATING
C696 S.n618 SUB 0.00fF $ **FLOATING
C697 S.n619 SUB 0.39fF $ **FLOATING
C698 S.n620 SUB 0.02fF $ **FLOATING
C699 S.t667 SUB 0.02fF
C700 S.n621 SUB 0.36fF $ **FLOATING
C701 S.n622 SUB 0.14fF $ **FLOATING
C702 S.n623 SUB 1.72fF $ **FLOATING
C703 S.n624 SUB 1.60fF $ **FLOATING
C704 S.t640 SUB 0.02fF
C705 S.n625 SUB 0.88fF $ **FLOATING
C706 S.t985 SUB 0.02fF
C707 S.n626 SUB 0.88fF $ **FLOATING
C708 S.n627 SUB 1.48fF $ **FLOATING
C709 S.n628 SUB 2.60fF $ **FLOATING
C710 S.n629 SUB 0.44fF $ **FLOATING
C711 S.n630 SUB 0.77fF $ **FLOATING
C712 S.n631 SUB 0.21fF $ **FLOATING
C713 S.n632 SUB 1.71fF $ **FLOATING
C714 S.n633 SUB 8.87fF $ **FLOATING
C715 S.n634 SUB 8.87fF $ **FLOATING
C716 S.n635 SUB 5.46fF $ **FLOATING
C717 S.n636 SUB 1.49fF $ **FLOATING
C718 S.n637 SUB 0.02fF $ **FLOATING
C719 S.t295 SUB 0.02fF
C720 S.n638 SUB 0.36fF $ **FLOATING
C721 S.n639 SUB 20.57fF $ **FLOATING
C722 S.n640 SUB 20.57fF $ **FLOATING
C723 S.n641 SUB 5.72fF $ **FLOATING
C724 S.n642 SUB 1.94fF $ **FLOATING
C725 S.t254 SUB 0.02fF
C726 S.n643 SUB 0.88fF $ **FLOATING
C727 S.t581 SUB 0.02fF
C728 S.n644 SUB 0.88fF $ **FLOATING
C729 S.n645 SUB 1.61fF $ **FLOATING
C730 S.n646 SUB 0.02fF $ **FLOATING
C731 S.t220 SUB 0.02fF
C732 S.n647 SUB 0.36fF $ **FLOATING
C733 S.t111 SUB 16.30fF
C734 S.t1049 SUB 0.02fF
C735 S.n648 SUB 0.88fF $ **FLOATING
C736 S.n649 SUB 0.02fF $ **FLOATING
C737 S.t845 SUB 0.02fF
C738 S.n650 SUB 0.36fF $ **FLOATING
C739 S.t761 SUB 0.02fF
C740 S.n651 SUB 0.88fF $ **FLOATING
C741 S.t279 SUB 0.02fF
C742 S.n652 SUB 0.88fF $ **FLOATING
C743 S.n653 SUB 0.02fF $ **FLOATING
C744 S.t722 SUB 0.02fF
C745 S.n654 SUB 0.36fF $ **FLOATING
C746 S.t1050 SUB 0.02fF
C747 S.n655 SUB 0.88fF $ **FLOATING
C748 S.t628 SUB 0.02fF
C749 S.n656 SUB 0.88fF $ **FLOATING
C750 S.n657 SUB 0.02fF $ **FLOATING
C751 S.t1065 SUB 0.02fF
C752 S.n658 SUB 0.36fF $ **FLOATING
C753 S.t303 SUB 0.02fF
C754 S.n659 SUB 0.88fF $ **FLOATING
C755 S.t1018 SUB 0.02fF
C756 S.n660 SUB 0.88fF $ **FLOATING
C757 S.n661 SUB 0.02fF $ **FLOATING
C758 S.t312 SUB 0.02fF
C759 S.n662 SUB 0.36fF $ **FLOATING
C760 S.t657 SUB 0.02fF
C761 S.n663 SUB 0.88fF $ **FLOATING
C762 S.t241 SUB 84.23fF
C763 S.n664 SUB 3.23fF $ **FLOATING
C764 S.n665 SUB 9.33fF $ **FLOATING
C765 S.n666 SUB 9.33fF $ **FLOATING
C766 S.n667 SUB 9.33fF $ **FLOATING
C767 S.n668 SUB 9.33fF $ **FLOATING
C768 S.n669 SUB 9.33fF $ **FLOATING
C769 S.n670 SUB 9.33fF $ **FLOATING
C770 S.n671 SUB 9.33fF $ **FLOATING
C771 S.n672 SUB 9.33fF $ **FLOATING
C772 S.n673 SUB 7.65fF $ **FLOATING
C773 S.n674 SUB 0.24fF $ **FLOATING
C774 S.n675 SUB 1.48fF $ **FLOATING
C775 S.n676 SUB 1.29fF $ **FLOATING
C776 S.n677 SUB 0.27fF $ **FLOATING
C777 S.n678 SUB 1.86fF $ **FLOATING
C778 S.n679 SUB 0.25fF $ **FLOATING
C779 S.n680 SUB 0.09fF $ **FLOATING
C780 S.n681 SUB 0.21fF $ **FLOATING
C781 S.n682 SUB 0.79fF $ **FLOATING
C782 S.n683 SUB 0.44fF $ **FLOATING
C783 S.n684 SUB 0.12fF $ **FLOATING
C784 S.t802 SUB 0.02fF
C785 S.n685 SUB 0.14fF $ **FLOATING
C786 S.t1033 SUB 0.02fF
C787 S.n687 SUB 0.24fF $ **FLOATING
C788 S.n688 SUB 0.35fF $ **FLOATING
C789 S.n689 SUB 0.60fF $ **FLOATING
C790 S.n690 SUB 0.02fF $ **FLOATING
C791 S.n691 SUB 0.01fF $ **FLOATING
C792 S.n692 SUB 0.02fF $ **FLOATING
C793 S.n693 SUB 0.08fF $ **FLOATING
C794 S.n694 SUB 0.06fF $ **FLOATING
C795 S.n695 SUB 0.03fF $ **FLOATING
C796 S.n696 SUB 0.03fF $ **FLOATING
C797 S.n697 SUB 0.99fF $ **FLOATING
C798 S.n698 SUB 0.36fF $ **FLOATING
C799 S.n699 SUB 1.83fF $ **FLOATING
C800 S.n700 SUB 1.97fF $ **FLOATING
C801 S.t419 SUB 0.02fF
C802 S.n701 SUB 0.24fF $ **FLOATING
C803 S.n702 SUB 0.90fF $ **FLOATING
C804 S.n703 SUB 0.05fF $ **FLOATING
C805 S.t887 SUB 0.02fF
C806 S.n704 SUB 0.12fF $ **FLOATING
C807 S.n705 SUB 0.14fF $ **FLOATING
C808 S.n707 SUB 1.87fF $ **FLOATING
C809 S.n708 SUB 0.06fF $ **FLOATING
C810 S.n709 SUB 0.03fF $ **FLOATING
C811 S.n710 SUB 0.03fF $ **FLOATING
C812 S.n711 SUB 0.98fF $ **FLOATING
C813 S.n712 SUB 0.02fF $ **FLOATING
C814 S.n713 SUB 0.01fF $ **FLOATING
C815 S.n714 SUB 0.02fF $ **FLOATING
C816 S.n715 SUB 0.08fF $ **FLOATING
C817 S.n716 SUB 0.35fF $ **FLOATING
C818 S.n717 SUB 1.84fF $ **FLOATING
C819 S.t824 SUB 0.02fF
C820 S.n718 SUB 0.24fF $ **FLOATING
C821 S.n719 SUB 0.35fF $ **FLOATING
C822 S.n720 SUB 0.60fF $ **FLOATING
C823 S.n721 SUB 0.12fF $ **FLOATING
C824 S.t605 SUB 0.02fF
C825 S.n722 SUB 0.14fF $ **FLOATING
C826 S.n724 SUB 0.94fF $ **FLOATING
C827 S.n725 SUB 0.58fF $ **FLOATING
C828 S.n726 SUB 0.25fF $ **FLOATING
C829 S.n727 SUB 0.69fF $ **FLOATING
C830 S.n728 SUB 0.22fF $ **FLOATING
C831 S.n729 SUB 0.09fF $ **FLOATING
C832 S.n730 SUB 1.87fF $ **FLOATING
C833 S.t399 SUB 0.02fF
C834 S.n731 SUB 0.24fF $ **FLOATING
C835 S.n732 SUB 0.90fF $ **FLOATING
C836 S.n733 SUB 0.05fF $ **FLOATING
C837 S.t665 SUB 0.02fF
C838 S.n734 SUB 0.12fF $ **FLOATING
C839 S.n735 SUB 0.14fF $ **FLOATING
C840 S.n737 SUB 1.86fF $ **FLOATING
C841 S.n738 SUB 0.25fF $ **FLOATING
C842 S.n739 SUB 0.09fF $ **FLOATING
C843 S.n740 SUB 0.21fF $ **FLOATING
C844 S.n741 SUB 0.79fF $ **FLOATING
C845 S.n742 SUB 0.44fF $ **FLOATING
C846 S.n743 SUB 0.12fF $ **FLOATING
C847 S.t214 SUB 0.02fF
C848 S.n744 SUB 0.14fF $ **FLOATING
C849 S.t450 SUB 0.02fF
C850 S.n746 SUB 0.24fF $ **FLOATING
C851 S.n747 SUB 0.35fF $ **FLOATING
C852 S.n748 SUB 0.60fF $ **FLOATING
C853 S.n749 SUB 0.02fF $ **FLOATING
C854 S.n750 SUB 0.01fF $ **FLOATING
C855 S.n751 SUB 0.02fF $ **FLOATING
C856 S.n752 SUB 0.08fF $ **FLOATING
C857 S.n753 SUB 0.06fF $ **FLOATING
C858 S.n754 SUB 0.03fF $ **FLOATING
C859 S.n755 SUB 0.03fF $ **FLOATING
C860 S.n756 SUB 0.99fF $ **FLOATING
C861 S.n757 SUB 0.36fF $ **FLOATING
C862 S.n758 SUB 1.83fF $ **FLOATING
C863 S.n759 SUB 1.97fF $ **FLOATING
C864 S.t1118 SUB 0.02fF
C865 S.n760 SUB 0.24fF $ **FLOATING
C866 S.n761 SUB 0.90fF $ **FLOATING
C867 S.n762 SUB 0.05fF $ **FLOATING
C868 S.t294 SUB 0.02fF
C869 S.n763 SUB 0.12fF $ **FLOATING
C870 S.n764 SUB 0.14fF $ **FLOATING
C871 S.n766 SUB 1.87fF $ **FLOATING
C872 S.n767 SUB 0.06fF $ **FLOATING
C873 S.n768 SUB 0.03fF $ **FLOATING
C874 S.n769 SUB 0.03fF $ **FLOATING
C875 S.n770 SUB 0.98fF $ **FLOATING
C876 S.n771 SUB 0.02fF $ **FLOATING
C877 S.n772 SUB 0.01fF $ **FLOATING
C878 S.n773 SUB 0.02fF $ **FLOATING
C879 S.n774 SUB 0.08fF $ **FLOATING
C880 S.n775 SUB 0.35fF $ **FLOATING
C881 S.n776 SUB 1.84fF $ **FLOATING
C882 S.t34 SUB 0.02fF
C883 S.n777 SUB 0.24fF $ **FLOATING
C884 S.n778 SUB 0.35fF $ **FLOATING
C885 S.n779 SUB 0.60fF $ **FLOATING
C886 S.n780 SUB 0.12fF $ **FLOATING
C887 S.t940 SUB 0.02fF
C888 S.n781 SUB 0.14fF $ **FLOATING
C889 S.n783 SUB 0.94fF $ **FLOATING
C890 S.n784 SUB 0.58fF $ **FLOATING
C891 S.n785 SUB 0.25fF $ **FLOATING
C892 S.n786 SUB 0.69fF $ **FLOATING
C893 S.n787 SUB 0.22fF $ **FLOATING
C894 S.n788 SUB 0.09fF $ **FLOATING
C895 S.n789 SUB 1.87fF $ **FLOATING
C896 S.t727 SUB 0.02fF
C897 S.n790 SUB 0.24fF $ **FLOATING
C898 S.n791 SUB 0.90fF $ **FLOATING
C899 S.n792 SUB 0.05fF $ **FLOATING
C900 S.t1025 SUB 0.02fF
C901 S.n793 SUB 0.12fF $ **FLOATING
C902 S.n794 SUB 0.14fF $ **FLOATING
C903 S.n796 SUB 1.86fF $ **FLOATING
C904 S.n797 SUB 0.25fF $ **FLOATING
C905 S.n798 SUB 0.09fF $ **FLOATING
C906 S.n799 SUB 0.21fF $ **FLOATING
C907 S.n800 SUB 0.79fF $ **FLOATING
C908 S.n801 SUB 0.44fF $ **FLOATING
C909 S.n802 SUB 0.12fF $ **FLOATING
C910 S.t559 SUB 0.02fF
C911 S.n803 SUB 0.14fF $ **FLOATING
C912 S.t781 SUB 0.02fF
C913 S.n805 SUB 0.24fF $ **FLOATING
C914 S.n806 SUB 0.35fF $ **FLOATING
C915 S.n807 SUB 0.60fF $ **FLOATING
C916 S.n808 SUB 0.02fF $ **FLOATING
C917 S.n809 SUB 0.01fF $ **FLOATING
C918 S.n810 SUB 0.02fF $ **FLOATING
C919 S.n811 SUB 0.08fF $ **FLOATING
C920 S.n812 SUB 0.03fF $ **FLOATING
C921 S.n813 SUB 0.03fF $ **FLOATING
C922 S.n814 SUB 1.01fF $ **FLOATING
C923 S.n815 SUB 0.36fF $ **FLOATING
C924 S.n816 SUB 1.83fF $ **FLOATING
C925 S.n817 SUB 1.97fF $ **FLOATING
C926 S.t346 SUB 0.02fF
C927 S.n818 SUB 0.24fF $ **FLOATING
C928 S.n819 SUB 0.90fF $ **FLOATING
C929 S.n820 SUB 0.05fF $ **FLOATING
C930 S.t651 SUB 0.02fF
C931 S.n821 SUB 0.12fF $ **FLOATING
C932 S.n822 SUB 0.14fF $ **FLOATING
C933 S.n824 SUB 0.25fF $ **FLOATING
C934 S.n825 SUB 0.69fF $ **FLOATING
C935 S.n826 SUB 0.22fF $ **FLOATING
C936 S.n827 SUB 0.09fF $ **FLOATING
C937 S.n828 SUB 0.94fF $ **FLOATING
C938 S.n829 SUB 0.58fF $ **FLOATING
C939 S.n830 SUB 1.87fF $ **FLOATING
C940 S.n831 SUB 0.12fF $ **FLOATING
C941 S.t236 SUB 0.02fF
C942 S.n832 SUB 0.14fF $ **FLOATING
C943 S.t468 SUB 0.02fF
C944 S.n834 SUB 0.24fF $ **FLOATING
C945 S.n835 SUB 0.35fF $ **FLOATING
C946 S.n836 SUB 0.60fF $ **FLOATING
C947 S.n837 SUB 0.18fF $ **FLOATING
C948 S.n838 SUB 0.21fF $ **FLOATING
C949 S.n839 SUB 0.47fF $ **FLOATING
C950 S.n840 SUB 0.33fF $ **FLOATING
C951 S.n841 SUB 0.01fF $ **FLOATING
C952 S.n842 SUB 0.01fF $ **FLOATING
C953 S.n843 SUB 0.01fF $ **FLOATING
C954 S.n844 SUB 0.07fF $ **FLOATING
C955 S.n845 SUB 0.07fF $ **FLOATING
C956 S.n846 SUB 0.04fF $ **FLOATING
C957 S.n847 SUB 0.05fF $ **FLOATING
C958 S.n848 SUB 0.41fF $ **FLOATING
C959 S.n849 SUB 0.57fF $ **FLOATING
C960 S.n850 SUB 0.19fF $ **FLOATING
C961 S.n851 SUB 1.95fF $ **FLOATING
C962 S.t1144 SUB 0.02fF
C963 S.n852 SUB 0.24fF $ **FLOATING
C964 S.n853 SUB 0.90fF $ **FLOATING
C965 S.n854 SUB 0.05fF $ **FLOATING
C966 S.t277 SUB 0.02fF
C967 S.n855 SUB 0.12fF $ **FLOATING
C968 S.n856 SUB 0.14fF $ **FLOATING
C969 S.n858 SUB 0.04fF $ **FLOATING
C970 S.n859 SUB 0.03fF $ **FLOATING
C971 S.n860 SUB 0.03fF $ **FLOATING
C972 S.n861 SUB 0.10fF $ **FLOATING
C973 S.n862 SUB 0.36fF $ **FLOATING
C974 S.n863 SUB 0.37fF $ **FLOATING
C975 S.n864 SUB 0.10fF $ **FLOATING
C976 S.n865 SUB 0.12fF $ **FLOATING
C977 S.n866 SUB 0.07fF $ **FLOATING
C978 S.n867 SUB 0.12fF $ **FLOATING
C979 S.n868 SUB 0.18fF $ **FLOATING
C980 S.n869 SUB 1.86fF $ **FLOATING
C981 S.n870 SUB 0.12fF $ **FLOATING
C982 S.t965 SUB 0.02fF
C983 S.n871 SUB 0.14fF $ **FLOATING
C984 S.t68 SUB 0.02fF
C985 S.n873 SUB 0.24fF $ **FLOATING
C986 S.n874 SUB 0.35fF $ **FLOATING
C987 S.n875 SUB 0.60fF $ **FLOATING
C988 S.n876 SUB 0.41fF $ **FLOATING
C989 S.n877 SUB 0.20fF $ **FLOATING
C990 S.n878 SUB 0.16fF $ **FLOATING
C991 S.n879 SUB 0.28fF $ **FLOATING
C992 S.n880 SUB 0.21fF $ **FLOATING
C993 S.n881 SUB 0.78fF $ **FLOATING
C994 S.n882 SUB 0.31fF $ **FLOATING
C995 S.n883 SUB 0.22fF $ **FLOATING
C996 S.n884 SUB 0.38fF $ **FLOATING
C997 S.n885 SUB 3.57fF $ **FLOATING
C998 S.t756 SUB 0.02fF
C999 S.n886 SUB 0.24fF $ **FLOATING
C1000 S.n887 SUB 0.90fF $ **FLOATING
C1001 S.n888 SUB 0.05fF $ **FLOATING
C1002 S.t995 SUB 0.02fF
C1003 S.n889 SUB 0.12fF $ **FLOATING
C1004 S.n890 SUB 0.14fF $ **FLOATING
C1005 S.n892 SUB 0.25fF $ **FLOATING
C1006 S.n893 SUB 0.09fF $ **FLOATING
C1007 S.n894 SUB 0.21fF $ **FLOATING
C1008 S.n895 SUB 1.27fF $ **FLOATING
C1009 S.n896 SUB 0.52fF $ **FLOATING
C1010 S.n897 SUB 1.86fF $ **FLOATING
C1011 S.n898 SUB 0.12fF $ **FLOATING
C1012 S.t587 SUB 0.02fF
C1013 S.n899 SUB 0.14fF $ **FLOATING
C1014 S.t809 SUB 0.02fF
C1015 S.n901 SUB 0.24fF $ **FLOATING
C1016 S.n902 SUB 0.35fF $ **FLOATING
C1017 S.n903 SUB 0.60fF $ **FLOATING
C1018 S.n904 SUB 0.41fF $ **FLOATING
C1019 S.n905 SUB 0.20fF $ **FLOATING
C1020 S.n906 SUB 0.16fF $ **FLOATING
C1021 S.n907 SUB 0.28fF $ **FLOATING
C1022 S.n908 SUB 0.21fF $ **FLOATING
C1023 S.n909 SUB 0.30fF $ **FLOATING
C1024 S.n910 SUB 0.36fF $ **FLOATING
C1025 S.n911 SUB 0.22fF $ **FLOATING
C1026 S.n912 SUB 0.38fF $ **FLOATING
C1027 S.n913 SUB 2.39fF $ **FLOATING
C1028 S.t372 SUB 0.02fF
C1029 S.n914 SUB 0.24fF $ **FLOATING
C1030 S.n915 SUB 0.90fF $ **FLOATING
C1031 S.n916 SUB 0.05fF $ **FLOATING
C1032 S.t620 SUB 0.02fF
C1033 S.n917 SUB 0.12fF $ **FLOATING
C1034 S.n918 SUB 0.14fF $ **FLOATING
C1035 S.n920 SUB 1.87fF $ **FLOATING
C1036 S.n921 SUB 2.64fF $ **FLOATING
C1037 S.t429 SUB 0.02fF
C1038 S.n922 SUB 0.24fF $ **FLOATING
C1039 S.n923 SUB 0.35fF $ **FLOATING
C1040 S.n924 SUB 0.60fF $ **FLOATING
C1041 S.n925 SUB 0.12fF $ **FLOATING
C1042 S.t192 SUB 0.02fF
C1043 S.n926 SUB 0.14fF $ **FLOATING
C1044 S.n928 SUB 0.69fF $ **FLOATING
C1045 S.n929 SUB 0.22fF $ **FLOATING
C1046 S.n930 SUB 0.69fF $ **FLOATING
C1047 S.n931 SUB 1.14fF $ **FLOATING
C1048 S.n932 SUB 0.22fF $ **FLOATING
C1049 S.n933 SUB 0.25fF $ **FLOATING
C1050 S.n934 SUB 0.09fF $ **FLOATING
C1051 S.n935 SUB 1.87fF $ **FLOATING
C1052 S.t1094 SUB 0.02fF
C1053 S.n936 SUB 0.24fF $ **FLOATING
C1054 S.n937 SUB 0.90fF $ **FLOATING
C1055 S.n938 SUB 0.05fF $ **FLOATING
C1056 S.t232 SUB 0.02fF
C1057 S.n939 SUB 0.12fF $ **FLOATING
C1058 S.n940 SUB 0.14fF $ **FLOATING
C1059 S.n942 SUB 14.09fF $ **FLOATING
C1060 S.n943 SUB 1.70fF $ **FLOATING
C1061 S.n944 SUB 3.02fF $ **FLOATING
C1062 S.t304 SUB 0.02fF
C1063 S.n945 SUB 0.24fF $ **FLOATING
C1064 S.n946 SUB 0.35fF $ **FLOATING
C1065 S.n947 SUB 0.60fF $ **FLOATING
C1066 S.n948 SUB 0.12fF $ **FLOATING
C1067 S.t60 SUB 0.02fF
C1068 S.n949 SUB 0.14fF $ **FLOATING
C1069 S.n951 SUB 0.28fF $ **FLOATING
C1070 S.n952 SUB 0.74fF $ **FLOATING
C1071 S.n953 SUB 0.59fF $ **FLOATING
C1072 S.n954 SUB 0.20fF $ **FLOATING
C1073 S.n955 SUB 0.20fF $ **FLOATING
C1074 S.n956 SUB 0.06fF $ **FLOATING
C1075 S.n957 SUB 0.09fF $ **FLOATING
C1076 S.n958 SUB 0.09fF $ **FLOATING
C1077 S.n959 SUB 1.97fF $ **FLOATING
C1078 S.t99 SUB 0.02fF
C1079 S.n960 SUB 0.12fF $ **FLOATING
C1080 S.n961 SUB 0.14fF $ **FLOATING
C1081 S.t799 SUB 0.02fF
C1082 S.n963 SUB 0.24fF $ **FLOATING
C1083 S.n964 SUB 0.90fF $ **FLOATING
C1084 S.n965 SUB 0.05fF $ **FLOATING
C1085 S.n966 SUB 1.86fF $ **FLOATING
C1086 S.n967 SUB 0.12fF $ **FLOATING
C1087 S.t1148 SUB 0.02fF
C1088 S.n968 SUB 0.14fF $ **FLOATING
C1089 S.t1046 SUB 0.02fF
C1090 S.n970 SUB 1.20fF $ **FLOATING
C1091 S.n971 SUB 0.60fF $ **FLOATING
C1092 S.n972 SUB 0.35fF $ **FLOATING
C1093 S.n973 SUB 0.62fF $ **FLOATING
C1094 S.n974 SUB 1.14fF $ **FLOATING
C1095 S.n975 SUB 2.18fF $ **FLOATING
C1096 S.n976 SUB 0.59fF $ **FLOATING
C1097 S.n977 SUB 0.02fF $ **FLOATING
C1098 S.n978 SUB 0.96fF $ **FLOATING
C1099 S.t91 SUB 14.50fF
C1100 S.n979 SUB 14.37fF $ **FLOATING
C1101 S.n981 SUB 0.37fF $ **FLOATING
C1102 S.n982 SUB 0.23fF $ **FLOATING
C1103 S.n983 SUB 2.87fF $ **FLOATING
C1104 S.n984 SUB 2.43fF $ **FLOATING
C1105 S.n985 SUB 1.94fF $ **FLOATING
C1106 S.n986 SUB 3.89fF $ **FLOATING
C1107 S.n987 SUB 0.25fF $ **FLOATING
C1108 S.n988 SUB 0.01fF $ **FLOATING
C1109 S.t951 SUB 0.02fF
C1110 S.n989 SUB 0.25fF $ **FLOATING
C1111 S.t629 SUB 0.02fF
C1112 S.n990 SUB 0.94fF $ **FLOATING
C1113 S.n991 SUB 0.70fF $ **FLOATING
C1114 S.n992 SUB 0.77fF $ **FLOATING
C1115 S.n993 SUB 1.91fF $ **FLOATING
C1116 S.n994 SUB 1.86fF $ **FLOATING
C1117 S.n995 SUB 0.12fF $ **FLOATING
C1118 S.t637 SUB 0.02fF
C1119 S.n996 SUB 0.14fF $ **FLOATING
C1120 S.t669 SUB 0.02fF
C1121 S.n998 SUB 0.24fF $ **FLOATING
C1122 S.n999 SUB 0.35fF $ **FLOATING
C1123 S.n1000 SUB 0.60fF $ **FLOATING
C1124 S.n1001 SUB 1.50fF $ **FLOATING
C1125 S.n1002 SUB 2.96fF $ **FLOATING
C1126 S.t244 SUB 0.02fF
C1127 S.n1003 SUB 0.24fF $ **FLOATING
C1128 S.n1004 SUB 0.90fF $ **FLOATING
C1129 S.n1005 SUB 0.05fF $ **FLOATING
C1130 S.t907 SUB 0.02fF
C1131 S.n1006 SUB 0.12fF $ **FLOATING
C1132 S.n1007 SUB 0.14fF $ **FLOATING
C1133 S.n1009 SUB 1.87fF $ **FLOATING
C1134 S.n1010 SUB 1.86fF $ **FLOATING
C1135 S.t566 SUB 0.02fF
C1136 S.n1011 SUB 0.24fF $ **FLOATING
C1137 S.n1012 SUB 0.35fF $ **FLOATING
C1138 S.n1013 SUB 0.60fF $ **FLOATING
C1139 S.n1014 SUB 0.12fF $ **FLOATING
C1140 S.t878 SUB 0.02fF
C1141 S.n1015 SUB 0.14fF $ **FLOATING
C1142 S.n1017 SUB 1.14fF $ **FLOATING
C1143 S.n1018 SUB 0.22fF $ **FLOATING
C1144 S.n1019 SUB 1.86fF $ **FLOATING
C1145 S.t49 SUB 0.02fF
C1146 S.n1020 SUB 0.24fF $ **FLOATING
C1147 S.n1021 SUB 0.90fF $ **FLOATING
C1148 S.n1022 SUB 0.05fF $ **FLOATING
C1149 S.t533 SUB 0.02fF
C1150 S.n1023 SUB 0.12fF $ **FLOATING
C1151 S.n1024 SUB 0.14fF $ **FLOATING
C1152 S.n1026 SUB 0.77fF $ **FLOATING
C1153 S.n1027 SUB 1.92fF $ **FLOATING
C1154 S.n1028 SUB 1.86fF $ **FLOATING
C1155 S.n1029 SUB 0.12fF $ **FLOATING
C1156 S.t501 SUB 0.02fF
C1157 S.n1030 SUB 0.14fF $ **FLOATING
C1158 S.t173 SUB 0.02fF
C1159 S.n1032 SUB 0.24fF $ **FLOATING
C1160 S.n1033 SUB 0.35fF $ **FLOATING
C1161 S.n1034 SUB 0.60fF $ **FLOATING
C1162 S.n1035 SUB 1.82fF $ **FLOATING
C1163 S.n1036 SUB 2.96fF $ **FLOATING
C1164 S.t791 SUB 0.02fF
C1165 S.n1037 SUB 0.24fF $ **FLOATING
C1166 S.n1038 SUB 0.90fF $ **FLOATING
C1167 S.n1039 SUB 0.05fF $ **FLOATING
C1168 S.t792 SUB 0.02fF
C1169 S.n1040 SUB 0.12fF $ **FLOATING
C1170 S.n1041 SUB 0.14fF $ **FLOATING
C1171 S.n1043 SUB 1.87fF $ **FLOATING
C1172 S.n1044 SUB 1.86fF $ **FLOATING
C1173 S.t895 SUB 0.02fF
C1174 S.n1045 SUB 0.24fF $ **FLOATING
C1175 S.n1046 SUB 0.35fF $ **FLOATING
C1176 S.n1047 SUB 0.60fF $ **FLOATING
C1177 S.n1048 SUB 0.12fF $ **FLOATING
C1178 S.t113 SUB 0.02fF
C1179 S.n1049 SUB 0.14fF $ **FLOATING
C1180 S.n1051 SUB 1.14fF $ **FLOATING
C1181 S.n1052 SUB 0.22fF $ **FLOATING
C1182 S.n1053 SUB 1.86fF $ **FLOATING
C1183 S.t411 SUB 0.02fF
C1184 S.n1054 SUB 0.24fF $ **FLOATING
C1185 S.n1055 SUB 0.90fF $ **FLOATING
C1186 S.n1056 SUB 0.05fF $ **FLOATING
C1187 S.t412 SUB 0.02fF
C1188 S.n1057 SUB 0.12fF $ **FLOATING
C1189 S.n1058 SUB 0.14fF $ **FLOATING
C1190 S.n1060 SUB 0.77fF $ **FLOATING
C1191 S.n1061 SUB 1.92fF $ **FLOATING
C1192 S.n1062 SUB 1.86fF $ **FLOATING
C1193 S.n1063 SUB 0.12fF $ **FLOATING
C1194 S.t846 SUB 0.02fF
C1195 S.n1064 SUB 0.14fF $ **FLOATING
C1196 S.t522 SUB 0.02fF
C1197 S.n1066 SUB 0.24fF $ **FLOATING
C1198 S.n1067 SUB 0.35fF $ **FLOATING
C1199 S.n1068 SUB 0.60fF $ **FLOATING
C1200 S.n1069 SUB 0.06fF $ **FLOATING
C1201 S.n1070 SUB 0.89fF $ **FLOATING
C1202 S.n1071 SUB 1.09fF $ **FLOATING
C1203 S.n1072 SUB 2.95fF $ **FLOATING
C1204 S.t1125 SUB 0.02fF
C1205 S.n1073 SUB 0.24fF $ **FLOATING
C1206 S.n1074 SUB 0.90fF $ **FLOATING
C1207 S.n1075 SUB 0.05fF $ **FLOATING
C1208 S.t1131 SUB 0.02fF
C1209 S.n1076 SUB 0.12fF $ **FLOATING
C1210 S.n1077 SUB 0.14fF $ **FLOATING
C1211 S.n1079 SUB 1.14fF $ **FLOATING
C1212 S.n1080 SUB 0.22fF $ **FLOATING
C1213 S.n1081 SUB 1.87fF $ **FLOATING
C1214 S.n1082 SUB 0.12fF $ **FLOATING
C1215 S.t471 SUB 0.02fF
C1216 S.n1083 SUB 0.14fF $ **FLOATING
C1217 S.t132 SUB 0.02fF
C1218 S.n1085 SUB 0.24fF $ **FLOATING
C1219 S.n1086 SUB 0.35fF $ **FLOATING
C1220 S.n1087 SUB 0.60fF $ **FLOATING
C1221 S.n1088 SUB 1.09fF $ **FLOATING
C1222 S.n1089 SUB 0.67fF $ **FLOATING
C1223 S.n1090 SUB 0.54fF $ **FLOATING
C1224 S.n1091 SUB 0.31fF $ **FLOATING
C1225 S.n1092 SUB 1.81fF $ **FLOATING
C1226 S.t740 SUB 0.02fF
C1227 S.n1093 SUB 0.24fF $ **FLOATING
C1228 S.n1094 SUB 0.90fF $ **FLOATING
C1229 S.n1095 SUB 0.05fF $ **FLOATING
C1230 S.t741 SUB 0.02fF
C1231 S.n1096 SUB 0.12fF $ **FLOATING
C1232 S.n1097 SUB 0.14fF $ **FLOATING
C1233 S.n1099 SUB 1.86fF $ **FLOATING
C1234 S.n1100 SUB 0.47fF $ **FLOATING
C1235 S.n1101 SUB 0.09fF $ **FLOATING
C1236 S.n1102 SUB 0.32fF $ **FLOATING
C1237 S.n1103 SUB 0.30fF $ **FLOATING
C1238 S.n1104 SUB 0.76fF $ **FLOATING
C1239 S.n1105 SUB 0.58fF $ **FLOATING
C1240 S.t861 SUB 0.02fF
C1241 S.n1106 SUB 0.24fF $ **FLOATING
C1242 S.n1107 SUB 0.35fF $ **FLOATING
C1243 S.n1108 SUB 0.60fF $ **FLOATING
C1244 S.n1109 SUB 0.12fF $ **FLOATING
C1245 S.t69 SUB 0.02fF
C1246 S.n1110 SUB 0.14fF $ **FLOATING
C1247 S.n1112 SUB 2.58fF $ **FLOATING
C1248 S.n1113 SUB 2.13fF $ **FLOATING
C1249 S.t356 SUB 0.02fF
C1250 S.n1114 SUB 0.24fF $ **FLOATING
C1251 S.n1115 SUB 0.90fF $ **FLOATING
C1252 S.n1116 SUB 0.05fF $ **FLOATING
C1253 S.t439 SUB 0.02fF
C1254 S.n1117 SUB 0.12fF $ **FLOATING
C1255 S.n1118 SUB 0.14fF $ **FLOATING
C1256 S.n1120 SUB 1.86fF $ **FLOATING
C1257 S.n1121 SUB 0.47fF $ **FLOATING
C1258 S.n1122 SUB 0.35fF $ **FLOATING
C1259 S.n1123 SUB 0.30fF $ **FLOATING
C1260 S.n1124 SUB 1.26fF $ **FLOATING
C1261 S.t485 SUB 0.02fF
C1262 S.n1125 SUB 0.24fF $ **FLOATING
C1263 S.n1126 SUB 0.35fF $ **FLOATING
C1264 S.n1127 SUB 0.60fF $ **FLOATING
C1265 S.n1128 SUB 0.12fF $ **FLOATING
C1266 S.t808 SUB 0.02fF
C1267 S.n1129 SUB 0.14fF $ **FLOATING
C1268 S.n1131 SUB 0.77fF $ **FLOATING
C1269 S.n1132 SUB 2.27fF $ **FLOATING
C1270 S.n1133 SUB 2.00fF $ **FLOATING
C1271 S.t1081 SUB 0.02fF
C1272 S.n1134 SUB 0.24fF $ **FLOATING
C1273 S.n1135 SUB 0.90fF $ **FLOATING
C1274 S.n1136 SUB 0.05fF $ **FLOATING
C1275 S.t7 SUB 0.02fF
C1276 S.n1137 SUB 0.12fF $ **FLOATING
C1277 S.n1138 SUB 0.14fF $ **FLOATING
C1278 S.n1140 SUB 1.87fF $ **FLOATING
C1279 S.n1141 SUB 2.65fF $ **FLOATING
C1280 S.t92 SUB 0.02fF
C1281 S.n1142 SUB 0.24fF $ **FLOATING
C1282 S.n1143 SUB 0.35fF $ **FLOATING
C1283 S.n1144 SUB 0.60fF $ **FLOATING
C1284 S.n1145 SUB 0.12fF $ **FLOATING
C1285 S.t428 SUB 0.02fF
C1286 S.n1146 SUB 0.14fF $ **FLOATING
C1287 S.n1148 SUB 1.14fF $ **FLOATING
C1288 S.n1149 SUB 0.22fF $ **FLOATING
C1289 S.n1150 SUB 1.86fF $ **FLOATING
C1290 S.t698 SUB 0.02fF
C1291 S.n1151 SUB 0.24fF $ **FLOATING
C1292 S.n1152 SUB 0.90fF $ **FLOATING
C1293 S.n1153 SUB 0.05fF $ **FLOATING
C1294 S.t764 SUB 0.02fF
C1295 S.n1154 SUB 0.12fF $ **FLOATING
C1296 S.n1155 SUB 0.14fF $ **FLOATING
C1297 S.n1157 SUB 14.09fF $ **FLOATING
C1298 S.n1158 SUB 2.69fF $ **FLOATING
C1299 S.n1159 SUB 1.79fF $ **FLOATING
C1300 S.n1160 SUB 0.12fF $ **FLOATING
C1301 S.t956 SUB 0.02fF
C1302 S.n1161 SUB 0.14fF $ **FLOATING
C1303 S.t475 SUB 0.02fF
C1304 S.n1163 SUB 0.24fF $ **FLOATING
C1305 S.n1164 SUB 0.35fF $ **FLOATING
C1306 S.n1165 SUB 0.60fF $ **FLOATING
C1307 S.n1166 SUB 2.34fF $ **FLOATING
C1308 S.n1167 SUB 2.28fF $ **FLOATING
C1309 S.t160 SUB 0.02fF
C1310 S.n1168 SUB 0.12fF $ **FLOATING
C1311 S.n1169 SUB 0.14fF $ **FLOATING
C1312 S.t520 SUB 0.02fF
C1313 S.n1171 SUB 0.24fF $ **FLOATING
C1314 S.n1172 SUB 0.90fF $ **FLOATING
C1315 S.n1173 SUB 0.05fF $ **FLOATING
C1316 S.t6 SUB 32.35fF
C1317 S.t382 SUB 0.02fF
C1318 S.n1174 SUB 0.12fF $ **FLOATING
C1319 S.n1175 SUB 0.14fF $ **FLOATING
C1320 S.t315 SUB 0.02fF
C1321 S.n1177 SUB 0.24fF $ **FLOATING
C1322 S.n1178 SUB 0.90fF $ **FLOATING
C1323 S.n1179 SUB 0.05fF $ **FLOATING
C1324 S.t825 SUB 0.02fF
C1325 S.n1180 SUB 0.24fF $ **FLOATING
C1326 S.n1181 SUB 0.35fF $ **FLOATING
C1327 S.n1182 SUB 0.60fF $ **FLOATING
C1328 S.n1183 SUB 0.31fF $ **FLOATING
C1329 S.n1184 SUB 1.53fF $ **FLOATING
C1330 S.n1185 SUB 0.15fF $ **FLOATING
C1331 S.n1186 SUB 4.92fF $ **FLOATING
C1332 S.n1187 SUB 1.86fF $ **FLOATING
C1333 S.n1188 SUB 0.12fF $ **FLOATING
C1334 S.t1036 SUB 0.02fF
C1335 S.n1189 SUB 0.14fF $ **FLOATING
C1336 S.t498 SUB 0.02fF
C1337 S.n1191 SUB 0.24fF $ **FLOATING
C1338 S.n1192 SUB 0.35fF $ **FLOATING
C1339 S.n1193 SUB 0.60fF $ **FLOATING
C1340 S.n1194 SUB 1.26fF $ **FLOATING
C1341 S.n1195 SUB 5.90fF $ **FLOATING
C1342 S.t954 SUB 0.02fF
C1343 S.n1196 SUB 0.12fF $ **FLOATING
C1344 S.n1197 SUB 0.14fF $ **FLOATING
C1345 S.t260 SUB 0.02fF
C1346 S.n1199 SUB 0.24fF $ **FLOATING
C1347 S.n1200 SUB 0.90fF $ **FLOATING
C1348 S.n1201 SUB 0.05fF $ **FLOATING
C1349 S.t59 SUB 31.97fF
C1350 S.t688 SUB 0.02fF
C1351 S.n1202 SUB 0.01fF $ **FLOATING
C1352 S.n1203 SUB 0.25fF $ **FLOATING
C1353 S.t1133 SUB 0.02fF
C1354 S.n1205 SUB 1.18fF $ **FLOATING
C1355 S.n1206 SUB 0.05fF $ **FLOATING
C1356 S.t459 SUB 0.02fF
C1357 S.n1207 SUB 0.63fF $ **FLOATING
C1358 S.n1208 SUB 0.60fF $ **FLOATING
C1359 S.n1209 SUB 0.59fF $ **FLOATING
C1360 S.n1210 SUB 0.21fF $ **FLOATING
C1361 S.n1211 SUB 0.59fF $ **FLOATING
C1362 S.n1212 SUB 2.57fF $ **FLOATING
C1363 S.n1213 SUB 0.29fF $ **FLOATING
C1364 S.t33 SUB 14.50fF
C1365 S.n1214 SUB 15.77fF $ **FLOATING
C1366 S.n1215 SUB 0.76fF $ **FLOATING
C1367 S.n1216 SUB 0.27fF $ **FLOATING
C1368 S.n1217 SUB 3.96fF $ **FLOATING
C1369 S.n1218 SUB 1.49fF $ **FLOATING
C1370 S.n1219 SUB 0.35fF $ **FLOATING
C1371 S.n1220 SUB 1.28fF $ **FLOATING
C1372 S.n1221 SUB 0.15fF $ **FLOATING
C1373 S.n1222 SUB 1.73fF $ **FLOATING
C1374 S.n1223 SUB 2.26fF $ **FLOATING
C1375 S.n1224 SUB 0.01fF $ **FLOATING
C1376 S.n1225 SUB 0.02fF $ **FLOATING
C1377 S.n1226 SUB 0.03fF $ **FLOATING
C1378 S.n1227 SUB 0.04fF $ **FLOATING
C1379 S.n1228 SUB 0.17fF $ **FLOATING
C1380 S.n1229 SUB 0.01fF $ **FLOATING
C1381 S.n1230 SUB 0.02fF $ **FLOATING
C1382 S.n1231 SUB 0.01fF $ **FLOATING
C1383 S.n1232 SUB 0.01fF $ **FLOATING
C1384 S.n1233 SUB 0.01fF $ **FLOATING
C1385 S.n1234 SUB 0.01fF $ **FLOATING
C1386 S.n1235 SUB 0.01fF $ **FLOATING
C1387 S.n1236 SUB 0.01fF $ **FLOATING
C1388 S.n1237 SUB 0.02fF $ **FLOATING
C1389 S.n1238 SUB 0.05fF $ **FLOATING
C1390 S.n1239 SUB 0.04fF $ **FLOATING
C1391 S.n1240 SUB 0.11fF $ **FLOATING
C1392 S.n1241 SUB 0.37fF $ **FLOATING
C1393 S.n1242 SUB 0.20fF $ **FLOATING
C1394 S.n1243 SUB 8.87fF $ **FLOATING
C1395 S.n1244 SUB 8.87fF $ **FLOATING
C1396 S.n1245 SUB 0.59fF $ **FLOATING
C1397 S.n1246 SUB 0.21fF $ **FLOATING
C1398 S.n1247 SUB 0.59fF $ **FLOATING
C1399 S.n1248 SUB 2.57fF $ **FLOATING
C1400 S.n1249 SUB 0.29fF $ **FLOATING
C1401 S.t141 SUB 14.50fF
C1402 S.n1250 SUB 15.77fF $ **FLOATING
C1403 S.n1251 SUB 0.76fF $ **FLOATING
C1404 S.n1252 SUB 0.27fF $ **FLOATING
C1405 S.n1253 SUB 3.96fF $ **FLOATING
C1406 S.n1254 SUB 1.34fF $ **FLOATING
C1407 S.t998 SUB 0.02fF
C1408 S.n1255 SUB 0.63fF $ **FLOATING
C1409 S.n1256 SUB 0.60fF $ **FLOATING
C1410 S.n1257 SUB 1.87fF $ **FLOATING
C1411 S.n1258 SUB 0.06fF $ **FLOATING
C1412 S.n1259 SUB 0.03fF $ **FLOATING
C1413 S.n1260 SUB 0.03fF $ **FLOATING
C1414 S.n1261 SUB 0.98fF $ **FLOATING
C1415 S.n1262 SUB 0.02fF $ **FLOATING
C1416 S.n1263 SUB 0.01fF $ **FLOATING
C1417 S.n1264 SUB 0.02fF $ **FLOATING
C1418 S.n1265 SUB 0.08fF $ **FLOATING
C1419 S.n1266 SUB 0.36fF $ **FLOATING
C1420 S.n1267 SUB 1.83fF $ **FLOATING
C1421 S.t1113 SUB 0.02fF
C1422 S.n1268 SUB 0.24fF $ **FLOATING
C1423 S.n1269 SUB 0.35fF $ **FLOATING
C1424 S.n1270 SUB 0.60fF $ **FLOATING
C1425 S.n1271 SUB 0.12fF $ **FLOATING
C1426 S.t891 SUB 0.02fF
C1427 S.n1272 SUB 0.14fF $ **FLOATING
C1428 S.n1274 SUB 0.69fF $ **FLOATING
C1429 S.n1275 SUB 0.22fF $ **FLOATING
C1430 S.n1276 SUB 0.25fF $ **FLOATING
C1431 S.n1277 SUB 0.09fF $ **FLOATING
C1432 S.n1278 SUB 0.22fF $ **FLOATING
C1433 S.n1279 SUB 0.69fF $ **FLOATING
C1434 S.n1280 SUB 1.14fF $ **FLOATING
C1435 S.n1281 SUB 0.22fF $ **FLOATING
C1436 S.n1282 SUB 0.25fF $ **FLOATING
C1437 S.n1283 SUB 0.09fF $ **FLOATING
C1438 S.n1284 SUB 1.86fF $ **FLOATING
C1439 S.t371 SUB 0.02fF
C1440 S.n1285 SUB 0.24fF $ **FLOATING
C1441 S.n1286 SUB 0.90fF $ **FLOATING
C1442 S.n1287 SUB 0.05fF $ **FLOATING
C1443 S.t996 SUB 0.02fF
C1444 S.n1288 SUB 0.12fF $ **FLOATING
C1445 S.n1289 SUB 0.14fF $ **FLOATING
C1446 S.n1291 SUB 0.25fF $ **FLOATING
C1447 S.n1292 SUB 0.09fF $ **FLOATING
C1448 S.n1293 SUB 0.21fF $ **FLOATING
C1449 S.n1294 SUB 0.91fF $ **FLOATING
C1450 S.n1295 SUB 0.44fF $ **FLOATING
C1451 S.n1296 SUB 1.86fF $ **FLOATING
C1452 S.n1297 SUB 0.12fF $ **FLOATING
C1453 S.t1093 SUB 0.02fF
C1454 S.n1298 SUB 0.14fF $ **FLOATING
C1455 S.t267 SUB 0.02fF
C1456 S.n1300 SUB 0.24fF $ **FLOATING
C1457 S.n1301 SUB 0.35fF $ **FLOATING
C1458 S.n1302 SUB 0.60fF $ **FLOATING
C1459 S.n1303 SUB 0.02fF $ **FLOATING
C1460 S.n1304 SUB 0.01fF $ **FLOATING
C1461 S.n1305 SUB 0.02fF $ **FLOATING
C1462 S.n1306 SUB 0.08fF $ **FLOATING
C1463 S.n1307 SUB 0.06fF $ **FLOATING
C1464 S.n1308 SUB 0.03fF $ **FLOATING
C1465 S.n1309 SUB 0.03fF $ **FLOATING
C1466 S.n1310 SUB 0.99fF $ **FLOATING
C1467 S.n1311 SUB 0.35fF $ **FLOATING
C1468 S.n1312 SUB 1.85fF $ **FLOATING
C1469 S.n1313 SUB 1.97fF $ **FLOATING
C1470 S.t210 SUB 0.02fF
C1471 S.n1314 SUB 0.24fF $ **FLOATING
C1472 S.n1315 SUB 0.90fF $ **FLOATING
C1473 S.n1316 SUB 0.05fF $ **FLOATING
C1474 S.t81 SUB 0.02fF
C1475 S.n1317 SUB 0.12fF $ **FLOATING
C1476 S.n1318 SUB 0.14fF $ **FLOATING
C1477 S.n1320 SUB 1.87fF $ **FLOATING
C1478 S.n1321 SUB 0.06fF $ **FLOATING
C1479 S.n1322 SUB 0.03fF $ **FLOATING
C1480 S.n1323 SUB 0.03fF $ **FLOATING
C1481 S.n1324 SUB 0.98fF $ **FLOATING
C1482 S.n1325 SUB 0.02fF $ **FLOATING
C1483 S.n1326 SUB 0.01fF $ **FLOATING
C1484 S.n1327 SUB 0.02fF $ **FLOATING
C1485 S.n1328 SUB 0.08fF $ **FLOATING
C1486 S.n1329 SUB 0.36fF $ **FLOATING
C1487 S.n1330 SUB 1.83fF $ **FLOATING
C1488 S.t987 SUB 0.02fF
C1489 S.n1331 SUB 0.24fF $ **FLOATING
C1490 S.n1332 SUB 0.35fF $ **FLOATING
C1491 S.n1333 SUB 0.60fF $ **FLOATING
C1492 S.n1334 SUB 0.12fF $ **FLOATING
C1493 S.t707 SUB 0.02fF
C1494 S.n1335 SUB 0.14fF $ **FLOATING
C1495 S.n1337 SUB 0.69fF $ **FLOATING
C1496 S.n1338 SUB 0.22fF $ **FLOATING
C1497 S.n1339 SUB 0.25fF $ **FLOATING
C1498 S.n1340 SUB 0.09fF $ **FLOATING
C1499 S.n1341 SUB 0.22fF $ **FLOATING
C1500 S.n1342 SUB 0.69fF $ **FLOATING
C1501 S.n1343 SUB 1.14fF $ **FLOATING
C1502 S.n1344 SUB 0.22fF $ **FLOATING
C1503 S.n1345 SUB 0.25fF $ **FLOATING
C1504 S.n1346 SUB 0.09fF $ **FLOATING
C1505 S.n1347 SUB 1.86fF $ **FLOATING
C1506 S.t934 SUB 0.02fF
C1507 S.n1348 SUB 0.24fF $ **FLOATING
C1508 S.n1349 SUB 0.90fF $ **FLOATING
C1509 S.n1350 SUB 0.05fF $ **FLOATING
C1510 S.t819 SUB 0.02fF
C1511 S.n1351 SUB 0.12fF $ **FLOATING
C1512 S.n1352 SUB 0.14fF $ **FLOATING
C1513 S.n1354 SUB 0.25fF $ **FLOATING
C1514 S.n1355 SUB 0.09fF $ **FLOATING
C1515 S.n1356 SUB 0.21fF $ **FLOATING
C1516 S.n1357 SUB 0.91fF $ **FLOATING
C1517 S.n1358 SUB 0.44fF $ **FLOATING
C1518 S.n1359 SUB 1.86fF $ **FLOATING
C1519 S.n1360 SUB 0.12fF $ **FLOATING
C1520 S.t329 SUB 0.02fF
C1521 S.n1361 SUB 0.14fF $ **FLOATING
C1522 S.t608 SUB 0.02fF
C1523 S.n1363 SUB 0.24fF $ **FLOATING
C1524 S.n1364 SUB 0.35fF $ **FLOATING
C1525 S.n1365 SUB 0.60fF $ **FLOATING
C1526 S.n1366 SUB 0.02fF $ **FLOATING
C1527 S.n1367 SUB 0.01fF $ **FLOATING
C1528 S.n1368 SUB 0.02fF $ **FLOATING
C1529 S.n1369 SUB 0.08fF $ **FLOATING
C1530 S.n1370 SUB 0.06fF $ **FLOATING
C1531 S.n1371 SUB 0.03fF $ **FLOATING
C1532 S.n1372 SUB 0.03fF $ **FLOATING
C1533 S.n1373 SUB 0.99fF $ **FLOATING
C1534 S.n1374 SUB 0.35fF $ **FLOATING
C1535 S.n1375 SUB 1.81fF $ **FLOATING
C1536 S.n1376 SUB 1.97fF $ **FLOATING
C1537 S.t555 SUB 0.02fF
C1538 S.n1377 SUB 0.24fF $ **FLOATING
C1539 S.n1378 SUB 0.90fF $ **FLOATING
C1540 S.n1379 SUB 0.05fF $ **FLOATING
C1541 S.t446 SUB 0.02fF
C1542 S.n1380 SUB 0.12fF $ **FLOATING
C1543 S.n1381 SUB 0.14fF $ **FLOATING
C1544 S.n1383 SUB 1.87fF $ **FLOATING
C1545 S.n1384 SUB 0.63fF $ **FLOATING
C1546 S.n1385 SUB 0.04fF $ **FLOATING
C1547 S.n1386 SUB 0.07fF $ **FLOATING
C1548 S.n1387 SUB 0.05fF $ **FLOATING
C1549 S.n1388 SUB 0.86fF $ **FLOATING
C1550 S.n1389 SUB 0.01fF $ **FLOATING
C1551 S.n1390 SUB 0.01fF $ **FLOATING
C1552 S.n1391 SUB 0.01fF $ **FLOATING
C1553 S.n1392 SUB 0.07fF $ **FLOATING
C1554 S.n1393 SUB 0.68fF $ **FLOATING
C1555 S.n1394 SUB 0.13fF $ **FLOATING
C1556 S.t222 SUB 0.02fF
C1557 S.n1395 SUB 0.24fF $ **FLOATING
C1558 S.n1396 SUB 0.35fF $ **FLOATING
C1559 S.n1397 SUB 0.60fF $ **FLOATING
C1560 S.n1398 SUB 0.12fF $ **FLOATING
C1561 S.t1053 SUB 0.02fF
C1562 S.n1399 SUB 0.14fF $ **FLOATING
C1563 S.n1401 SUB 0.69fF $ **FLOATING
C1564 S.n1402 SUB 0.22fF $ **FLOATING
C1565 S.n1403 SUB 0.25fF $ **FLOATING
C1566 S.n1404 SUB 0.09fF $ **FLOATING
C1567 S.n1405 SUB 0.22fF $ **FLOATING
C1568 S.n1406 SUB 0.69fF $ **FLOATING
C1569 S.n1407 SUB 1.14fF $ **FLOATING
C1570 S.n1408 SUB 0.22fF $ **FLOATING
C1571 S.n1409 SUB 0.25fF $ **FLOATING
C1572 S.n1410 SUB 0.09fF $ **FLOATING
C1573 S.n1411 SUB 2.29fF $ **FLOATING
C1574 S.t163 SUB 0.02fF
C1575 S.n1412 SUB 0.24fF $ **FLOATING
C1576 S.n1413 SUB 0.90fF $ **FLOATING
C1577 S.n1414 SUB 0.05fF $ **FLOATING
C1578 S.t24 SUB 0.02fF
C1579 S.n1415 SUB 0.12fF $ **FLOATING
C1580 S.n1416 SUB 0.14fF $ **FLOATING
C1581 S.n1418 SUB 1.86fF $ **FLOATING
C1582 S.n1419 SUB 0.45fF $ **FLOATING
C1583 S.n1420 SUB 0.22fF $ **FLOATING
C1584 S.n1421 SUB 0.38fF $ **FLOATING
C1585 S.n1422 SUB 0.16fF $ **FLOATING
C1586 S.n1423 SUB 0.28fF $ **FLOATING
C1587 S.n1424 SUB 0.21fF $ **FLOATING
C1588 S.n1425 SUB 0.30fF $ **FLOATING
C1589 S.n1426 SUB 0.41fF $ **FLOATING
C1590 S.n1427 SUB 0.20fF $ **FLOATING
C1591 S.t1007 SUB 0.02fF
C1592 S.n1428 SUB 0.24fF $ **FLOATING
C1593 S.n1429 SUB 0.35fF $ **FLOATING
C1594 S.n1430 SUB 0.60fF $ **FLOATING
C1595 S.n1431 SUB 0.12fF $ **FLOATING
C1596 S.t729 SUB 0.02fF
C1597 S.n1432 SUB 0.14fF $ **FLOATING
C1598 S.n1434 SUB 0.04fF $ **FLOATING
C1599 S.n1435 SUB 0.03fF $ **FLOATING
C1600 S.n1436 SUB 0.03fF $ **FLOATING
C1601 S.n1437 SUB 0.10fF $ **FLOATING
C1602 S.n1438 SUB 0.36fF $ **FLOATING
C1603 S.n1439 SUB 0.37fF $ **FLOATING
C1604 S.n1440 SUB 0.10fF $ **FLOATING
C1605 S.n1441 SUB 0.12fF $ **FLOATING
C1606 S.n1442 SUB 0.07fF $ **FLOATING
C1607 S.n1443 SUB 0.12fF $ **FLOATING
C1608 S.n1444 SUB 0.18fF $ **FLOATING
C1609 S.n1445 SUB 3.95fF $ **FLOATING
C1610 S.t964 SUB 0.02fF
C1611 S.n1446 SUB 0.24fF $ **FLOATING
C1612 S.n1447 SUB 0.90fF $ **FLOATING
C1613 S.n1448 SUB 0.05fF $ **FLOATING
C1614 S.t774 SUB 0.02fF
C1615 S.n1449 SUB 0.12fF $ **FLOATING
C1616 S.n1450 SUB 0.14fF $ **FLOATING
C1617 S.n1452 SUB 0.25fF $ **FLOATING
C1618 S.n1453 SUB 0.09fF $ **FLOATING
C1619 S.n1454 SUB 0.21fF $ **FLOATING
C1620 S.n1455 SUB 1.27fF $ **FLOATING
C1621 S.n1456 SUB 0.52fF $ **FLOATING
C1622 S.n1457 SUB 1.86fF $ **FLOATING
C1623 S.n1458 SUB 0.12fF $ **FLOATING
C1624 S.t348 SUB 0.02fF
C1625 S.n1459 SUB 0.14fF $ **FLOATING
C1626 S.t630 SUB 0.02fF
C1627 S.n1461 SUB 0.24fF $ **FLOATING
C1628 S.n1462 SUB 0.35fF $ **FLOATING
C1629 S.n1463 SUB 0.60fF $ **FLOATING
C1630 S.n1464 SUB 0.70fF $ **FLOATING
C1631 S.n1465 SUB 1.56fF $ **FLOATING
C1632 S.n1466 SUB 2.42fF $ **FLOATING
C1633 S.t583 SUB 0.02fF
C1634 S.n1467 SUB 0.24fF $ **FLOATING
C1635 S.n1468 SUB 0.90fF $ **FLOATING
C1636 S.n1469 SUB 0.05fF $ **FLOATING
C1637 S.t388 SUB 0.02fF
C1638 S.n1470 SUB 0.12fF $ **FLOATING
C1639 S.n1471 SUB 0.14fF $ **FLOATING
C1640 S.n1473 SUB 1.87fF $ **FLOATING
C1641 S.n1474 SUB 0.06fF $ **FLOATING
C1642 S.n1475 SUB 0.03fF $ **FLOATING
C1643 S.n1476 SUB 0.03fF $ **FLOATING
C1644 S.n1477 SUB 0.98fF $ **FLOATING
C1645 S.n1478 SUB 0.02fF $ **FLOATING
C1646 S.n1479 SUB 0.01fF $ **FLOATING
C1647 S.n1480 SUB 0.02fF $ **FLOATING
C1648 S.n1481 SUB 0.08fF $ **FLOATING
C1649 S.n1482 SUB 0.36fF $ **FLOATING
C1650 S.n1483 SUB 1.83fF $ **FLOATING
C1651 S.t245 SUB 0.02fF
C1652 S.n1484 SUB 0.24fF $ **FLOATING
C1653 S.n1485 SUB 0.35fF $ **FLOATING
C1654 S.n1486 SUB 0.60fF $ **FLOATING
C1655 S.n1487 SUB 0.12fF $ **FLOATING
C1656 S.t1071 SUB 0.02fF
C1657 S.n1488 SUB 0.14fF $ **FLOATING
C1658 S.n1490 SUB 0.69fF $ **FLOATING
C1659 S.n1491 SUB 0.22fF $ **FLOATING
C1660 S.n1492 SUB 0.25fF $ **FLOATING
C1661 S.n1493 SUB 0.09fF $ **FLOATING
C1662 S.n1494 SUB 0.22fF $ **FLOATING
C1663 S.n1495 SUB 0.69fF $ **FLOATING
C1664 S.n1496 SUB 1.14fF $ **FLOATING
C1665 S.n1497 SUB 0.22fF $ **FLOATING
C1666 S.n1498 SUB 0.25fF $ **FLOATING
C1667 S.n1499 SUB 0.09fF $ **FLOATING
C1668 S.n1500 SUB 1.86fF $ **FLOATING
C1669 S.t189 SUB 0.02fF
C1670 S.n1501 SUB 0.24fF $ **FLOATING
C1671 S.n1502 SUB 0.90fF $ **FLOATING
C1672 S.n1503 SUB 0.05fF $ **FLOATING
C1673 S.t1110 SUB 0.02fF
C1674 S.n1504 SUB 0.12fF $ **FLOATING
C1675 S.n1505 SUB 0.14fF $ **FLOATING
C1676 S.n1507 SUB 14.09fF $ **FLOATING
C1677 S.n1508 SUB 0.06fF $ **FLOATING
C1678 S.n1509 SUB 0.20fF $ **FLOATING
C1679 S.n1510 SUB 0.09fF $ **FLOATING
C1680 S.n1511 SUB 0.20fF $ **FLOATING
C1681 S.n1512 SUB 0.09fF $ **FLOATING
C1682 S.n1513 SUB 0.30fF $ **FLOATING
C1683 S.n1514 SUB 0.69fF $ **FLOATING
C1684 S.n1515 SUB 0.44fF $ **FLOATING
C1685 S.n1516 SUB 2.31fF $ **FLOATING
C1686 S.n1517 SUB 0.12fF $ **FLOATING
C1687 S.t165 SUB 0.02fF
C1688 S.n1518 SUB 0.14fF $ **FLOATING
C1689 S.t392 SUB 0.02fF
C1690 S.n1520 SUB 0.24fF $ **FLOATING
C1691 S.n1521 SUB 0.35fF $ **FLOATING
C1692 S.n1522 SUB 0.60fF $ **FLOATING
C1693 S.n1523 SUB 1.88fF $ **FLOATING
C1694 S.n1524 SUB 0.17fF $ **FLOATING
C1695 S.n1525 SUB 0.76fF $ **FLOATING
C1696 S.n1526 SUB 0.31fF $ **FLOATING
C1697 S.n1527 SUB 0.25fF $ **FLOATING
C1698 S.n1528 SUB 0.29fF $ **FLOATING
C1699 S.n1529 SUB 0.46fF $ **FLOATING
C1700 S.n1530 SUB 0.16fF $ **FLOATING
C1701 S.n1531 SUB 1.91fF $ **FLOATING
C1702 S.t206 SUB 0.02fF
C1703 S.n1532 SUB 0.12fF $ **FLOATING
C1704 S.n1533 SUB 0.14fF $ **FLOATING
C1705 S.t755 SUB 0.02fF
C1706 S.n1535 SUB 0.24fF $ **FLOATING
C1707 S.n1536 SUB 0.90fF $ **FLOATING
C1708 S.n1537 SUB 0.05fF $ **FLOATING
C1709 S.n1538 SUB 1.86fF $ **FLOATING
C1710 S.n1539 SUB 0.12fF $ **FLOATING
C1711 S.t22 SUB 0.02fF
C1712 S.n1540 SUB 0.14fF $ **FLOATING
C1713 S.t952 SUB 0.02fF
C1714 S.n1542 SUB 1.20fF $ **FLOATING
C1715 S.n1543 SUB 0.36fF $ **FLOATING
C1716 S.n1544 SUB 1.21fF $ **FLOATING
C1717 S.n1545 SUB 0.60fF $ **FLOATING
C1718 S.n1546 SUB 0.35fF $ **FLOATING
C1719 S.n1547 SUB 0.62fF $ **FLOATING
C1720 S.n1548 SUB 1.14fF $ **FLOATING
C1721 S.n1549 SUB 2.18fF $ **FLOATING
C1722 S.n1550 SUB 0.59fF $ **FLOATING
C1723 S.n1551 SUB 0.02fF $ **FLOATING
C1724 S.n1552 SUB 0.96fF $ **FLOATING
C1725 S.t106 SUB 14.50fF
C1726 S.n1553 SUB 14.37fF $ **FLOATING
C1727 S.n1555 SUB 0.37fF $ **FLOATING
C1728 S.n1556 SUB 0.23fF $ **FLOATING
C1729 S.n1557 SUB 2.76fF $ **FLOATING
C1730 S.n1558 SUB 2.43fF $ **FLOATING
C1731 S.n1559 SUB 3.95fF $ **FLOATING
C1732 S.n1560 SUB 0.25fF $ **FLOATING
C1733 S.n1561 SUB 0.01fF $ **FLOATING
C1734 S.t814 SUB 0.02fF
C1735 S.n1562 SUB 0.25fF $ **FLOATING
C1736 S.t677 SUB 0.02fF
C1737 S.n1563 SUB 0.94fF $ **FLOATING
C1738 S.n1564 SUB 0.70fF $ **FLOATING
C1739 S.n1565 SUB 1.87fF $ **FLOATING
C1740 S.n1566 SUB 1.86fF $ **FLOATING
C1741 S.t568 SUB 0.02fF
C1742 S.n1567 SUB 0.24fF $ **FLOATING
C1743 S.n1568 SUB 0.35fF $ **FLOATING
C1744 S.n1569 SUB 0.60fF $ **FLOATING
C1745 S.n1570 SUB 0.12fF $ **FLOATING
C1746 S.t494 SUB 0.02fF
C1747 S.n1571 SUB 0.14fF $ **FLOATING
C1748 S.n1573 SUB 1.14fF $ **FLOATING
C1749 S.n1574 SUB 0.22fF $ **FLOATING
C1750 S.n1575 SUB 0.25fF $ **FLOATING
C1751 S.n1576 SUB 0.09fF $ **FLOATING
C1752 S.n1577 SUB 1.86fF $ **FLOATING
C1753 S.t307 SUB 0.02fF
C1754 S.n1578 SUB 0.24fF $ **FLOATING
C1755 S.n1579 SUB 0.90fF $ **FLOATING
C1756 S.n1580 SUB 0.05fF $ **FLOATING
C1757 S.t777 SUB 0.02fF
C1758 S.n1581 SUB 0.12fF $ **FLOATING
C1759 S.n1582 SUB 0.14fF $ **FLOATING
C1760 S.n1584 SUB 0.77fF $ **FLOATING
C1761 S.n1585 SUB 1.92fF $ **FLOATING
C1762 S.n1586 SUB 1.86fF $ **FLOATING
C1763 S.n1587 SUB 0.12fF $ **FLOATING
C1764 S.t515 SUB 0.02fF
C1765 S.n1588 SUB 0.14fF $ **FLOATING
C1766 S.t187 SUB 0.02fF
C1767 S.n1590 SUB 0.24fF $ **FLOATING
C1768 S.n1591 SUB 0.35fF $ **FLOATING
C1769 S.n1592 SUB 0.60fF $ **FLOATING
C1770 S.n1593 SUB 1.82fF $ **FLOATING
C1771 S.n1594 SUB 2.96fF $ **FLOATING
C1772 S.t618 SUB 0.02fF
C1773 S.n1595 SUB 0.24fF $ **FLOATING
C1774 S.n1596 SUB 0.90fF $ **FLOATING
C1775 S.n1597 SUB 0.05fF $ **FLOATING
C1776 S.t395 SUB 0.02fF
C1777 S.n1598 SUB 0.12fF $ **FLOATING
C1778 S.n1599 SUB 0.14fF $ **FLOATING
C1779 S.n1601 SUB 1.87fF $ **FLOATING
C1780 S.n1602 SUB 1.86fF $ **FLOATING
C1781 S.t910 SUB 0.02fF
C1782 S.n1603 SUB 0.24fF $ **FLOATING
C1783 S.n1604 SUB 0.35fF $ **FLOATING
C1784 S.n1605 SUB 0.60fF $ **FLOATING
C1785 S.n1606 SUB 0.12fF $ **FLOATING
C1786 S.t123 SUB 0.02fF
C1787 S.n1607 SUB 0.14fF $ **FLOATING
C1788 S.n1609 SUB 1.14fF $ **FLOATING
C1789 S.n1610 SUB 0.22fF $ **FLOATING
C1790 S.n1611 SUB 0.25fF $ **FLOATING
C1791 S.n1612 SUB 0.09fF $ **FLOATING
C1792 S.n1613 SUB 1.86fF $ **FLOATING
C1793 S.t229 SUB 0.02fF
C1794 S.n1614 SUB 0.24fF $ **FLOATING
C1795 S.n1615 SUB 0.90fF $ **FLOATING
C1796 S.n1616 SUB 0.05fF $ **FLOATING
C1797 S.t427 SUB 0.02fF
C1798 S.n1617 SUB 0.12fF $ **FLOATING
C1799 S.n1618 SUB 0.14fF $ **FLOATING
C1800 S.n1620 SUB 0.77fF $ **FLOATING
C1801 S.n1621 SUB 1.92fF $ **FLOATING
C1802 S.n1622 SUB 1.86fF $ **FLOATING
C1803 S.n1623 SUB 0.12fF $ **FLOATING
C1804 S.t855 SUB 0.02fF
C1805 S.n1624 SUB 0.14fF $ **FLOATING
C1806 S.t532 SUB 0.02fF
C1807 S.n1626 SUB 0.24fF $ **FLOATING
C1808 S.n1627 SUB 0.35fF $ **FLOATING
C1809 S.n1628 SUB 0.60fF $ **FLOATING
C1810 S.n1629 SUB 1.82fF $ **FLOATING
C1811 S.n1630 SUB 2.96fF $ **FLOATING
C1812 S.t953 SUB 0.02fF
C1813 S.n1631 SUB 0.24fF $ **FLOATING
C1814 S.n1632 SUB 0.90fF $ **FLOATING
C1815 S.n1633 SUB 0.05fF $ **FLOATING
C1816 S.t1146 SUB 0.02fF
C1817 S.n1634 SUB 0.12fF $ **FLOATING
C1818 S.n1635 SUB 0.14fF $ **FLOATING
C1819 S.n1637 SUB 1.87fF $ **FLOATING
C1820 S.n1638 SUB 1.73fF $ **FLOATING
C1821 S.t146 SUB 0.02fF
C1822 S.n1639 SUB 0.24fF $ **FLOATING
C1823 S.n1640 SUB 0.35fF $ **FLOATING
C1824 S.n1641 SUB 0.60fF $ **FLOATING
C1825 S.n1642 SUB 0.12fF $ **FLOATING
C1826 S.t479 SUB 0.02fF
C1827 S.n1643 SUB 0.14fF $ **FLOATING
C1828 S.n1645 SUB 1.14fF $ **FLOATING
C1829 S.n1646 SUB 0.22fF $ **FLOATING
C1830 S.n1647 SUB 0.25fF $ **FLOATING
C1831 S.n1648 SUB 0.09fF $ **FLOATING
C1832 S.n1649 SUB 2.41fF $ **FLOATING
C1833 S.t573 SUB 0.02fF
C1834 S.n1650 SUB 0.24fF $ **FLOATING
C1835 S.n1651 SUB 0.90fF $ **FLOATING
C1836 S.n1652 SUB 0.05fF $ **FLOATING
C1837 S.t757 SUB 0.02fF
C1838 S.n1653 SUB 0.12fF $ **FLOATING
C1839 S.n1654 SUB 0.14fF $ **FLOATING
C1840 S.n1656 SUB 1.86fF $ **FLOATING
C1841 S.n1657 SUB 0.47fF $ **FLOATING
C1842 S.n1658 SUB 0.09fF $ **FLOATING
C1843 S.n1659 SUB 0.32fF $ **FLOATING
C1844 S.n1660 SUB 0.30fF $ **FLOATING
C1845 S.n1661 SUB 0.76fF $ **FLOATING
C1846 S.n1662 SUB 0.58fF $ **FLOATING
C1847 S.t874 SUB 0.02fF
C1848 S.n1663 SUB 0.24fF $ **FLOATING
C1849 S.n1664 SUB 0.35fF $ **FLOATING
C1850 S.n1665 SUB 0.60fF $ **FLOATING
C1851 S.n1666 SUB 0.12fF $ **FLOATING
C1852 S.t83 SUB 0.02fF
C1853 S.n1667 SUB 0.14fF $ **FLOATING
C1854 S.n1669 SUB 2.58fF $ **FLOATING
C1855 S.n1670 SUB 2.13fF $ **FLOATING
C1856 S.t176 SUB 0.02fF
C1857 S.n1671 SUB 0.24fF $ **FLOATING
C1858 S.n1672 SUB 0.90fF $ **FLOATING
C1859 S.n1673 SUB 0.05fF $ **FLOATING
C1860 S.t370 SUB 0.02fF
C1861 S.n1674 SUB 0.12fF $ **FLOATING
C1862 S.n1675 SUB 0.14fF $ **FLOATING
C1863 S.n1677 SUB 0.77fF $ **FLOATING
C1864 S.n1678 SUB 2.27fF $ **FLOATING
C1865 S.n1679 SUB 1.86fF $ **FLOATING
C1866 S.n1680 SUB 0.12fF $ **FLOATING
C1867 S.t818 SUB 0.02fF
C1868 S.n1681 SUB 0.14fF $ **FLOATING
C1869 S.t496 SUB 0.02fF
C1870 S.n1683 SUB 0.24fF $ **FLOATING
C1871 S.n1684 SUB 0.35fF $ **FLOATING
C1872 S.n1685 SUB 0.60fF $ **FLOATING
C1873 S.n1686 SUB 1.37fF $ **FLOATING
C1874 S.n1687 SUB 0.70fF $ **FLOATING
C1875 S.n1688 SUB 1.13fF $ **FLOATING
C1876 S.n1689 SUB 0.35fF $ **FLOATING
C1877 S.n1690 SUB 2.00fF $ **FLOATING
C1878 S.t900 SUB 0.02fF
C1879 S.n1691 SUB 0.24fF $ **FLOATING
C1880 S.n1692 SUB 0.90fF $ **FLOATING
C1881 S.n1693 SUB 0.05fF $ **FLOATING
C1882 S.t40 SUB 0.02fF
C1883 S.n1694 SUB 0.12fF $ **FLOATING
C1884 S.n1695 SUB 0.14fF $ **FLOATING
C1885 S.n1697 SUB 1.87fF $ **FLOATING
C1886 S.n1698 SUB 1.86fF $ **FLOATING
C1887 S.t107 SUB 0.02fF
C1888 S.n1699 SUB 0.24fF $ **FLOATING
C1889 S.n1700 SUB 0.35fF $ **FLOATING
C1890 S.n1701 SUB 0.60fF $ **FLOATING
C1891 S.n1702 SUB 0.12fF $ **FLOATING
C1892 S.t444 SUB 0.02fF
C1893 S.n1703 SUB 0.14fF $ **FLOATING
C1894 S.n1705 SUB 1.14fF $ **FLOATING
C1895 S.n1706 SUB 0.22fF $ **FLOATING
C1896 S.n1707 SUB 0.25fF $ **FLOATING
C1897 S.n1708 SUB 0.09fF $ **FLOATING
C1898 S.n1709 SUB 1.86fF $ **FLOATING
C1899 S.t527 SUB 0.02fF
C1900 S.n1710 SUB 0.24fF $ **FLOATING
C1901 S.n1711 SUB 0.90fF $ **FLOATING
C1902 S.n1712 SUB 0.05fF $ **FLOATING
C1903 S.t783 SUB 0.02fF
C1904 S.n1713 SUB 0.12fF $ **FLOATING
C1905 S.n1714 SUB 0.14fF $ **FLOATING
C1906 S.n1716 SUB 14.09fF $ **FLOATING
C1907 S.n1717 SUB 2.70fF $ **FLOATING
C1908 S.n1718 SUB 1.58fF $ **FLOATING
C1909 S.n1719 SUB 0.12fF $ **FLOATING
C1910 S.t318 SUB 0.02fF
C1911 S.n1720 SUB 0.14fF $ **FLOATING
C1912 S.t975 SUB 0.02fF
C1913 S.n1722 SUB 0.24fF $ **FLOATING
C1914 S.n1723 SUB 0.35fF $ **FLOATING
C1915 S.n1724 SUB 0.60fF $ **FLOATING
C1916 S.n1725 SUB 0.07fF $ **FLOATING
C1917 S.n1726 SUB 0.01fF $ **FLOATING
C1918 S.n1727 SUB 0.23fF $ **FLOATING
C1919 S.n1728 SUB 1.15fF $ **FLOATING
C1920 S.n1729 SUB 1.33fF $ **FLOATING
C1921 S.n1730 SUB 2.28fF $ **FLOATING
C1922 S.t664 SUB 0.02fF
C1923 S.n1731 SUB 0.12fF $ **FLOATING
C1924 S.n1732 SUB 0.14fF $ **FLOATING
C1925 S.t1083 SUB 0.02fF
C1926 S.n1734 SUB 0.24fF $ **FLOATING
C1927 S.n1735 SUB 0.90fF $ **FLOATING
C1928 S.n1736 SUB 0.05fF $ **FLOATING
C1929 S.t21 SUB 32.35fF
C1930 S.t398 SUB 0.02fF
C1931 S.n1737 SUB 0.12fF $ **FLOATING
C1932 S.n1738 SUB 0.14fF $ **FLOATING
C1933 S.t142 SUB 0.02fF
C1934 S.n1740 SUB 0.24fF $ **FLOATING
C1935 S.n1741 SUB 0.90fF $ **FLOATING
C1936 S.n1742 SUB 0.05fF $ **FLOATING
C1937 S.t837 SUB 0.02fF
C1938 S.n1743 SUB 0.24fF $ **FLOATING
C1939 S.n1744 SUB 0.35fF $ **FLOATING
C1940 S.n1745 SUB 0.60fF $ **FLOATING
C1941 S.n1746 SUB 0.31fF $ **FLOATING
C1942 S.n1747 SUB 1.08fF $ **FLOATING
C1943 S.n1748 SUB 0.15fF $ **FLOATING
C1944 S.n1749 SUB 2.08fF $ **FLOATING
C1945 S.n1750 SUB 2.91fF $ **FLOATING
C1946 S.n1751 SUB 1.86fF $ **FLOATING
C1947 S.n1752 SUB 0.12fF $ **FLOATING
C1948 S.t689 SUB 0.02fF
C1949 S.n1753 SUB 0.14fF $ **FLOATING
C1950 S.t969 SUB 0.02fF
C1951 S.n1755 SUB 0.24fF $ **FLOATING
C1952 S.n1756 SUB 0.35fF $ **FLOATING
C1953 S.n1757 SUB 0.60fF $ **FLOATING
C1954 S.n1758 SUB 0.91fF $ **FLOATING
C1955 S.n1759 SUB 0.31fF $ **FLOATING
C1956 S.n1760 SUB 0.91fF $ **FLOATING
C1957 S.n1761 SUB 1.08fF $ **FLOATING
C1958 S.n1762 SUB 0.15fF $ **FLOATING
C1959 S.n1763 SUB 4.63fF $ **FLOATING
C1960 S.t720 SUB 0.02fF
C1961 S.n1764 SUB 0.12fF $ **FLOATING
C1962 S.n1765 SUB 0.14fF $ **FLOATING
C1963 S.t912 SUB 0.02fF
C1964 S.n1767 SUB 0.24fF $ **FLOATING
C1965 S.n1768 SUB 0.90fF $ **FLOATING
C1966 S.n1769 SUB 0.05fF $ **FLOATING
C1967 S.n1770 SUB 1.86fF $ **FLOATING
C1968 S.n1771 SUB 2.64fF $ **FLOATING
C1969 S.t989 SUB 0.02fF
C1970 S.n1772 SUB 0.24fF $ **FLOATING
C1971 S.n1773 SUB 0.35fF $ **FLOATING
C1972 S.n1774 SUB 0.60fF $ **FLOATING
C1973 S.n1775 SUB 0.12fF $ **FLOATING
C1974 S.t408 SUB 0.02fF
C1975 S.n1776 SUB 0.14fF $ **FLOATING
C1976 S.n1778 SUB 1.86fF $ **FLOATING
C1977 S.n1779 SUB 2.65fF $ **FLOATING
C1978 S.t463 SUB 0.02fF
C1979 S.n1780 SUB 0.24fF $ **FLOATING
C1980 S.n1781 SUB 0.35fF $ **FLOATING
C1981 S.n1782 SUB 0.60fF $ **FLOATING
C1982 S.t867 SUB 0.02fF
C1983 S.n1783 SUB 0.24fF $ **FLOATING
C1984 S.n1784 SUB 0.90fF $ **FLOATING
C1985 S.n1785 SUB 0.05fF $ **FLOATING
C1986 S.t1120 SUB 0.02fF
C1987 S.n1786 SUB 0.12fF $ **FLOATING
C1988 S.n1787 SUB 0.14fF $ **FLOATING
C1989 S.n1789 SUB 0.12fF $ **FLOATING
C1990 S.t773 SUB 0.02fF
C1991 S.n1790 SUB 0.14fF $ **FLOATING
C1992 S.n1792 SUB 5.12fF $ **FLOATING
C1993 S.n1793 SUB 5.40fF $ **FLOATING
C1994 S.t341 SUB 0.02fF
C1995 S.n1794 SUB 0.12fF $ **FLOATING
C1996 S.n1795 SUB 0.14fF $ **FLOATING
C1997 S.t445 SUB 0.02fF
C1998 S.n1797 SUB 0.24fF $ **FLOATING
C1999 S.n1798 SUB 0.90fF $ **FLOATING
C2000 S.n1799 SUB 0.05fF $ **FLOATING
C2001 S.t23 SUB 31.97fF
C2002 S.t948 SUB 0.02fF
C2003 S.n1800 SUB 1.18fF $ **FLOATING
C2004 S.n1801 SUB 0.05fF $ **FLOATING
C2005 S.t74 SUB 0.02fF
C2006 S.n1802 SUB 0.01fF $ **FLOATING
C2007 S.n1803 SUB 0.25fF $ **FLOATING
C2008 S.n1805 SUB 1.48fF $ **FLOATING
C2009 S.n1806 SUB 1.29fF $ **FLOATING
C2010 S.n1807 SUB 0.27fF $ **FLOATING
C2011 S.n1808 SUB 0.24fF $ **FLOATING
C2012 S.n1809 SUB 4.34fF $ **FLOATING
C2013 S.n1810 SUB 0.01fF $ **FLOATING
C2014 S.n1811 SUB 0.02fF $ **FLOATING
C2015 S.n1812 SUB 0.03fF $ **FLOATING
C2016 S.n1813 SUB 0.04fF $ **FLOATING
C2017 S.n1814 SUB 0.17fF $ **FLOATING
C2018 S.n1815 SUB 0.01fF $ **FLOATING
C2019 S.n1816 SUB 0.02fF $ **FLOATING
C2020 S.n1817 SUB 0.01fF $ **FLOATING
C2021 S.n1818 SUB 0.01fF $ **FLOATING
C2022 S.n1819 SUB 0.01fF $ **FLOATING
C2023 S.n1820 SUB 0.01fF $ **FLOATING
C2024 S.n1821 SUB 0.01fF $ **FLOATING
C2025 S.n1822 SUB 0.01fF $ **FLOATING
C2026 S.n1823 SUB 0.02fF $ **FLOATING
C2027 S.n1824 SUB 0.05fF $ **FLOATING
C2028 S.n1825 SUB 0.04fF $ **FLOATING
C2029 S.n1826 SUB 0.11fF $ **FLOATING
C2030 S.n1827 SUB 0.37fF $ **FLOATING
C2031 S.n1828 SUB 0.20fF $ **FLOATING
C2032 S.n1829 SUB 8.87fF $ **FLOATING
C2033 S.n1830 SUB 8.87fF $ **FLOATING
C2034 S.n1831 SUB 0.59fF $ **FLOATING
C2035 S.n1832 SUB 0.21fF $ **FLOATING
C2036 S.n1833 SUB 0.59fF $ **FLOATING
C2037 S.n1834 SUB 2.57fF $ **FLOATING
C2038 S.n1835 SUB 0.29fF $ **FLOATING
C2039 S.t149 SUB 14.50fF
C2040 S.n1836 SUB 15.77fF $ **FLOATING
C2041 S.n1837 SUB 0.76fF $ **FLOATING
C2042 S.n1838 SUB 0.27fF $ **FLOATING
C2043 S.n1839 SUB 3.96fF $ **FLOATING
C2044 S.n1840 SUB 1.34fF $ **FLOATING
C2045 S.t632 SUB 0.02fF
C2046 S.n1841 SUB 0.63fF $ **FLOATING
C2047 S.n1842 SUB 0.60fF $ **FLOATING
C2048 S.n1843 SUB 0.25fF $ **FLOATING
C2049 S.n1844 SUB 0.09fF $ **FLOATING
C2050 S.n1845 SUB 0.21fF $ **FLOATING
C2051 S.n1846 SUB 0.91fF $ **FLOATING
C2052 S.n1847 SUB 0.44fF $ **FLOATING
C2053 S.n1848 SUB 1.86fF $ **FLOATING
C2054 S.n1849 SUB 0.12fF $ **FLOATING
C2055 S.t754 SUB 0.02fF
C2056 S.n1850 SUB 0.14fF $ **FLOATING
C2057 S.t1015 SUB 0.02fF
C2058 S.n1852 SUB 0.24fF $ **FLOATING
C2059 S.n1853 SUB 0.35fF $ **FLOATING
C2060 S.n1854 SUB 0.60fF $ **FLOATING
C2061 S.n1855 SUB 0.02fF $ **FLOATING
C2062 S.n1856 SUB 0.01fF $ **FLOATING
C2063 S.n1857 SUB 0.02fF $ **FLOATING
C2064 S.n1858 SUB 0.08fF $ **FLOATING
C2065 S.n1859 SUB 0.06fF $ **FLOATING
C2066 S.n1860 SUB 0.03fF $ **FLOATING
C2067 S.n1861 SUB 0.03fF $ **FLOATING
C2068 S.n1862 SUB 0.99fF $ **FLOATING
C2069 S.n1863 SUB 0.35fF $ **FLOATING
C2070 S.n1864 SUB 1.85fF $ **FLOATING
C2071 S.n1865 SUB 1.97fF $ **FLOATING
C2072 S.t280 SUB 0.02fF
C2073 S.n1866 SUB 0.24fF $ **FLOATING
C2074 S.n1867 SUB 0.90fF $ **FLOATING
C2075 S.n1868 SUB 0.05fF $ **FLOATING
C2076 S.t856 SUB 0.02fF
C2077 S.n1869 SUB 0.12fF $ **FLOATING
C2078 S.n1870 SUB 0.14fF $ **FLOATING
C2079 S.n1872 SUB 1.87fF $ **FLOATING
C2080 S.n1873 SUB 0.06fF $ **FLOATING
C2081 S.n1874 SUB 0.03fF $ **FLOATING
C2082 S.n1875 SUB 0.03fF $ **FLOATING
C2083 S.n1876 SUB 0.98fF $ **FLOATING
C2084 S.n1877 SUB 0.02fF $ **FLOATING
C2085 S.n1878 SUB 0.01fF $ **FLOATING
C2086 S.n1879 SUB 0.02fF $ **FLOATING
C2087 S.n1880 SUB 0.08fF $ **FLOATING
C2088 S.n1881 SUB 0.36fF $ **FLOATING
C2089 S.n1882 SUB 1.83fF $ **FLOATING
C2090 S.t1001 SUB 0.02fF
C2091 S.n1883 SUB 0.24fF $ **FLOATING
C2092 S.n1884 SUB 0.35fF $ **FLOATING
C2093 S.n1885 SUB 0.60fF $ **FLOATING
C2094 S.n1886 SUB 0.12fF $ **FLOATING
C2095 S.t719 SUB 0.02fF
C2096 S.n1887 SUB 0.14fF $ **FLOATING
C2097 S.n1889 SUB 0.69fF $ **FLOATING
C2098 S.n1890 SUB 0.22fF $ **FLOATING
C2099 S.n1891 SUB 0.22fF $ **FLOATING
C2100 S.n1892 SUB 0.69fF $ **FLOATING
C2101 S.n1893 SUB 1.14fF $ **FLOATING
C2102 S.n1894 SUB 0.22fF $ **FLOATING
C2103 S.n1895 SUB 0.25fF $ **FLOATING
C2104 S.n1896 SUB 0.09fF $ **FLOATING
C2105 S.n1897 SUB 1.86fF $ **FLOATING
C2106 S.t950 SUB 0.02fF
C2107 S.n1898 SUB 0.24fF $ **FLOATING
C2108 S.n1899 SUB 0.90fF $ **FLOATING
C2109 S.n1900 SUB 0.05fF $ **FLOATING
C2110 S.t830 SUB 0.02fF
C2111 S.n1901 SUB 0.12fF $ **FLOATING
C2112 S.n1902 SUB 0.14fF $ **FLOATING
C2113 S.n1904 SUB 0.25fF $ **FLOATING
C2114 S.n1905 SUB 0.09fF $ **FLOATING
C2115 S.n1906 SUB 0.21fF $ **FLOATING
C2116 S.n1907 SUB 0.91fF $ **FLOATING
C2117 S.n1908 SUB 0.44fF $ **FLOATING
C2118 S.n1909 SUB 1.86fF $ **FLOATING
C2119 S.n1910 SUB 0.12fF $ **FLOATING
C2120 S.t338 SUB 0.02fF
C2121 S.n1911 SUB 0.14fF $ **FLOATING
C2122 S.t624 SUB 0.02fF
C2123 S.n1913 SUB 0.24fF $ **FLOATING
C2124 S.n1914 SUB 0.35fF $ **FLOATING
C2125 S.n1915 SUB 0.60fF $ **FLOATING
C2126 S.n1916 SUB 0.02fF $ **FLOATING
C2127 S.n1917 SUB 0.01fF $ **FLOATING
C2128 S.n1918 SUB 0.02fF $ **FLOATING
C2129 S.n1919 SUB 0.08fF $ **FLOATING
C2130 S.n1920 SUB 0.06fF $ **FLOATING
C2131 S.n1921 SUB 0.03fF $ **FLOATING
C2132 S.n1922 SUB 0.03fF $ **FLOATING
C2133 S.n1923 SUB 0.99fF $ **FLOATING
C2134 S.n1924 SUB 0.35fF $ **FLOATING
C2135 S.n1925 SUB 1.85fF $ **FLOATING
C2136 S.n1926 SUB 1.97fF $ **FLOATING
C2137 S.t571 SUB 0.02fF
C2138 S.n1927 SUB 0.24fF $ **FLOATING
C2139 S.n1928 SUB 0.90fF $ **FLOATING
C2140 S.n1929 SUB 0.05fF $ **FLOATING
C2141 S.t456 SUB 0.02fF
C2142 S.n1930 SUB 0.12fF $ **FLOATING
C2143 S.n1931 SUB 0.14fF $ **FLOATING
C2144 S.n1933 SUB 1.87fF $ **FLOATING
C2145 S.n1934 SUB 0.07fF $ **FLOATING
C2146 S.n1935 SUB 0.04fF $ **FLOATING
C2147 S.n1936 SUB 0.05fF $ **FLOATING
C2148 S.n1937 SUB 0.86fF $ **FLOATING
C2149 S.n1938 SUB 0.01fF $ **FLOATING
C2150 S.n1939 SUB 0.01fF $ **FLOATING
C2151 S.n1940 SUB 0.01fF $ **FLOATING
C2152 S.n1941 SUB 0.07fF $ **FLOATING
C2153 S.n1942 SUB 0.68fF $ **FLOATING
C2154 S.n1943 SUB 0.71fF $ **FLOATING
C2155 S.t234 SUB 0.02fF
C2156 S.n1944 SUB 0.24fF $ **FLOATING
C2157 S.n1945 SUB 0.35fF $ **FLOATING
C2158 S.n1946 SUB 0.60fF $ **FLOATING
C2159 S.n1947 SUB 0.12fF $ **FLOATING
C2160 S.t1066 SUB 0.02fF
C2161 S.n1948 SUB 0.14fF $ **FLOATING
C2162 S.n1950 SUB 0.69fF $ **FLOATING
C2163 S.n1951 SUB 0.22fF $ **FLOATING
C2164 S.n1952 SUB 0.22fF $ **FLOATING
C2165 S.n1953 SUB 0.69fF $ **FLOATING
C2166 S.n1954 SUB 1.14fF $ **FLOATING
C2167 S.n1955 SUB 0.22fF $ **FLOATING
C2168 S.n1956 SUB 0.25fF $ **FLOATING
C2169 S.n1957 SUB 0.09fF $ **FLOATING
C2170 S.n1958 SUB 2.29fF $ **FLOATING
C2171 S.t177 SUB 0.02fF
C2172 S.n1959 SUB 0.24fF $ **FLOATING
C2173 S.n1960 SUB 0.90fF $ **FLOATING
C2174 S.n1961 SUB 0.05fF $ **FLOATING
C2175 S.t48 SUB 0.02fF
C2176 S.n1962 SUB 0.12fF $ **FLOATING
C2177 S.n1963 SUB 0.14fF $ **FLOATING
C2178 S.n1965 SUB 1.86fF $ **FLOATING
C2179 S.n1966 SUB 0.45fF $ **FLOATING
C2180 S.n1967 SUB 0.22fF $ **FLOATING
C2181 S.n1968 SUB 0.38fF $ **FLOATING
C2182 S.n1969 SUB 0.16fF $ **FLOATING
C2183 S.n1970 SUB 0.28fF $ **FLOATING
C2184 S.n1971 SUB 0.21fF $ **FLOATING
C2185 S.n1972 SUB 0.30fF $ **FLOATING
C2186 S.n1973 SUB 0.41fF $ **FLOATING
C2187 S.n1974 SUB 0.20fF $ **FLOATING
C2188 S.t963 SUB 0.02fF
C2189 S.n1975 SUB 0.24fF $ **FLOATING
C2190 S.n1976 SUB 0.35fF $ **FLOATING
C2191 S.n1977 SUB 0.60fF $ **FLOATING
C2192 S.n1978 SUB 0.12fF $ **FLOATING
C2193 S.t683 SUB 0.02fF
C2194 S.n1979 SUB 0.14fF $ **FLOATING
C2195 S.n1981 SUB 0.04fF $ **FLOATING
C2196 S.n1982 SUB 0.03fF $ **FLOATING
C2197 S.n1983 SUB 0.03fF $ **FLOATING
C2198 S.n1984 SUB 0.10fF $ **FLOATING
C2199 S.n1985 SUB 0.36fF $ **FLOATING
C2200 S.n1986 SUB 0.37fF $ **FLOATING
C2201 S.n1987 SUB 0.10fF $ **FLOATING
C2202 S.n1988 SUB 0.12fF $ **FLOATING
C2203 S.n1989 SUB 0.07fF $ **FLOATING
C2204 S.n1990 SUB 0.12fF $ **FLOATING
C2205 S.n1991 SUB 0.18fF $ **FLOATING
C2206 S.n1992 SUB 3.95fF $ **FLOATING
C2207 S.t901 SUB 0.02fF
C2208 S.n1993 SUB 0.24fF $ **FLOATING
C2209 S.n1994 SUB 0.90fF $ **FLOATING
C2210 S.n1995 SUB 0.05fF $ **FLOATING
C2211 S.t790 SUB 0.02fF
C2212 S.n1996 SUB 0.12fF $ **FLOATING
C2213 S.n1997 SUB 0.14fF $ **FLOATING
C2214 S.n1999 SUB 0.25fF $ **FLOATING
C2215 S.n2000 SUB 0.09fF $ **FLOATING
C2216 S.n2001 SUB 0.21fF $ **FLOATING
C2217 S.n2002 SUB 1.27fF $ **FLOATING
C2218 S.n2003 SUB 0.52fF $ **FLOATING
C2219 S.n2004 SUB 1.86fF $ **FLOATING
C2220 S.n2005 SUB 0.12fF $ **FLOATING
C2221 S.t362 SUB 0.02fF
C2222 S.n2006 SUB 0.14fF $ **FLOATING
C2223 S.t641 SUB 0.02fF
C2224 S.n2008 SUB 0.24fF $ **FLOATING
C2225 S.n2009 SUB 0.35fF $ **FLOATING
C2226 S.n2010 SUB 0.60fF $ **FLOATING
C2227 S.n2011 SUB 1.56fF $ **FLOATING
C2228 S.n2012 SUB 2.42fF $ **FLOATING
C2229 S.t599 SUB 0.02fF
C2230 S.n2013 SUB 0.24fF $ **FLOATING
C2231 S.n2014 SUB 0.90fF $ **FLOATING
C2232 S.n2015 SUB 0.05fF $ **FLOATING
C2233 S.t410 SUB 0.02fF
C2234 S.n2016 SUB 0.12fF $ **FLOATING
C2235 S.n2017 SUB 0.14fF $ **FLOATING
C2236 S.n2019 SUB 1.87fF $ **FLOATING
C2237 S.n2020 SUB 0.06fF $ **FLOATING
C2238 S.n2021 SUB 0.03fF $ **FLOATING
C2239 S.n2022 SUB 0.03fF $ **FLOATING
C2240 S.n2023 SUB 0.98fF $ **FLOATING
C2241 S.n2024 SUB 0.02fF $ **FLOATING
C2242 S.n2025 SUB 0.01fF $ **FLOATING
C2243 S.n2026 SUB 0.02fF $ **FLOATING
C2244 S.n2027 SUB 0.08fF $ **FLOATING
C2245 S.n2028 SUB 0.36fF $ **FLOATING
C2246 S.n2029 SUB 1.83fF $ **FLOATING
C2247 S.t258 SUB 0.02fF
C2248 S.n2030 SUB 0.24fF $ **FLOATING
C2249 S.n2031 SUB 0.35fF $ **FLOATING
C2250 S.n2032 SUB 0.60fF $ **FLOATING
C2251 S.n2033 SUB 0.12fF $ **FLOATING
C2252 S.t1088 SUB 0.02fF
C2253 S.n2034 SUB 0.14fF $ **FLOATING
C2254 S.n2036 SUB 0.69fF $ **FLOATING
C2255 S.n2037 SUB 0.22fF $ **FLOATING
C2256 S.n2038 SUB 0.22fF $ **FLOATING
C2257 S.n2039 SUB 0.69fF $ **FLOATING
C2258 S.n2040 SUB 1.14fF $ **FLOATING
C2259 S.n2041 SUB 0.22fF $ **FLOATING
C2260 S.n2042 SUB 0.25fF $ **FLOATING
C2261 S.n2043 SUB 0.09fF $ **FLOATING
C2262 S.n2044 SUB 1.86fF $ **FLOATING
C2263 S.t202 SUB 0.02fF
C2264 S.n2045 SUB 0.24fF $ **FLOATING
C2265 S.n2046 SUB 0.90fF $ **FLOATING
C2266 S.n2047 SUB 0.05fF $ **FLOATING
C2267 S.t1124 SUB 0.02fF
C2268 S.n2048 SUB 0.12fF $ **FLOATING
C2269 S.n2049 SUB 0.14fF $ **FLOATING
C2270 S.n2051 SUB 14.09fF $ **FLOATING
C2271 S.n2052 SUB 1.70fF $ **FLOATING
C2272 S.n2053 SUB 3.01fF $ **FLOATING
C2273 S.t287 SUB 0.02fF
C2274 S.n2054 SUB 0.24fF $ **FLOATING
C2275 S.n2055 SUB 0.35fF $ **FLOATING
C2276 S.n2056 SUB 0.60fF $ **FLOATING
C2277 S.n2057 SUB 0.12fF $ **FLOATING
C2278 S.t1142 SUB 0.02fF
C2279 S.n2058 SUB 0.14fF $ **FLOATING
C2280 S.n2060 SUB 0.31fF $ **FLOATING
C2281 S.n2061 SUB 0.22fF $ **FLOATING
C2282 S.n2062 SUB 0.65fF $ **FLOATING
C2283 S.n2063 SUB 0.94fF $ **FLOATING
C2284 S.n2064 SUB 0.22fF $ **FLOATING
C2285 S.n2065 SUB 0.20fF $ **FLOATING
C2286 S.n2066 SUB 0.20fF $ **FLOATING
C2287 S.n2067 SUB 0.06fF $ **FLOATING
C2288 S.n2068 SUB 0.09fF $ **FLOATING
C2289 S.n2069 SUB 0.09fF $ **FLOATING
C2290 S.n2070 SUB 1.97fF $ **FLOATING
C2291 S.t56 SUB 0.02fF
C2292 S.n2071 SUB 0.12fF $ **FLOATING
C2293 S.n2072 SUB 0.14fF $ **FLOATING
C2294 S.t654 SUB 0.02fF
C2295 S.n2074 SUB 0.24fF $ **FLOATING
C2296 S.n2075 SUB 0.90fF $ **FLOATING
C2297 S.n2076 SUB 0.05fF $ **FLOATING
C2298 S.n2077 SUB 1.86fF $ **FLOATING
C2299 S.n2078 SUB 0.12fF $ **FLOATING
C2300 S.t46 SUB 0.02fF
C2301 S.n2079 SUB 0.14fF $ **FLOATING
C2302 S.t417 SUB 0.02fF
C2303 S.n2081 SUB 0.12fF $ **FLOATING
C2304 S.n2082 SUB 0.14fF $ **FLOATING
C2305 S.t150 SUB 0.02fF
C2306 S.n2084 SUB 0.24fF $ **FLOATING
C2307 S.n2085 SUB 0.90fF $ **FLOATING
C2308 S.n2086 SUB 0.05fF $ **FLOATING
C2309 S.t850 SUB 0.02fF
C2310 S.n2087 SUB 0.24fF $ **FLOATING
C2311 S.n2088 SUB 0.35fF $ **FLOATING
C2312 S.n2089 SUB 0.60fF $ **FLOATING
C2313 S.n2090 SUB 0.31fF $ **FLOATING
C2314 S.n2091 SUB 1.08fF $ **FLOATING
C2315 S.n2092 SUB 0.15fF $ **FLOATING
C2316 S.n2093 SUB 2.08fF $ **FLOATING
C2317 S.n2094 SUB 2.91fF $ **FLOATING
C2318 S.n2095 SUB 1.86fF $ **FLOATING
C2319 S.n2096 SUB 0.12fF $ **FLOATING
C2320 S.t701 SUB 0.02fF
C2321 S.n2097 SUB 0.14fF $ **FLOATING
C2322 S.t980 SUB 0.02fF
C2323 S.n2099 SUB 0.24fF $ **FLOATING
C2324 S.n2100 SUB 0.35fF $ **FLOATING
C2325 S.n2101 SUB 0.60fF $ **FLOATING
C2326 S.n2102 SUB 0.91fF $ **FLOATING
C2327 S.n2103 SUB 0.31fF $ **FLOATING
C2328 S.n2104 SUB 0.91fF $ **FLOATING
C2329 S.n2105 SUB 1.08fF $ **FLOATING
C2330 S.n2106 SUB 0.15fF $ **FLOATING
C2331 S.n2107 SUB 4.90fF $ **FLOATING
C2332 S.t738 SUB 0.02fF
C2333 S.n2108 SUB 0.12fF $ **FLOATING
C2334 S.n2109 SUB 0.14fF $ **FLOATING
C2335 S.t926 SUB 0.02fF
C2336 S.n2111 SUB 0.24fF $ **FLOATING
C2337 S.n2112 SUB 0.90fF $ **FLOATING
C2338 S.n2113 SUB 0.05fF $ **FLOATING
C2339 S.n2114 SUB 1.86fF $ **FLOATING
C2340 S.n2115 SUB 2.64fF $ **FLOATING
C2341 S.t603 SUB 0.02fF
C2342 S.n2116 SUB 0.24fF $ **FLOATING
C2343 S.n2117 SUB 0.35fF $ **FLOATING
C2344 S.n2118 SUB 0.60fF $ **FLOATING
C2345 S.t355 SUB 0.02fF
C2346 S.n2119 SUB 0.12fF $ **FLOATING
C2347 S.n2120 SUB 0.14fF $ **FLOATING
C2348 S.n2122 SUB 0.12fF $ **FLOATING
C2349 S.t322 SUB 0.02fF
C2350 S.n2123 SUB 0.14fF $ **FLOATING
C2351 S.n2125 SUB 1.86fF $ **FLOATING
C2352 S.n2126 SUB 2.64fF $ **FLOATING
C2353 S.t474 SUB 0.02fF
C2354 S.n2127 SUB 0.24fF $ **FLOATING
C2355 S.n2128 SUB 0.35fF $ **FLOATING
C2356 S.n2129 SUB 0.60fF $ **FLOATING
C2357 S.t879 SUB 0.02fF
C2358 S.n2130 SUB 0.24fF $ **FLOATING
C2359 S.n2131 SUB 0.90fF $ **FLOATING
C2360 S.n2132 SUB 0.05fF $ **FLOATING
C2361 S.t1135 SUB 0.02fF
C2362 S.n2133 SUB 0.12fF $ **FLOATING
C2363 S.n2134 SUB 0.14fF $ **FLOATING
C2364 S.n2136 SUB 0.12fF $ **FLOATING
C2365 S.t789 SUB 0.02fF
C2366 S.n2137 SUB 0.14fF $ **FLOATING
C2367 S.n2139 SUB 2.28fF $ **FLOATING
C2368 S.n2140 SUB 2.91fF $ **FLOATING
C2369 S.n2141 SUB 4.83fF $ **FLOATING
C2370 S.t548 SUB 0.02fF
C2371 S.n2142 SUB 0.24fF $ **FLOATING
C2372 S.n2143 SUB 0.90fF $ **FLOATING
C2373 S.n2144 SUB 0.05fF $ **FLOATING
C2374 S.n2145 SUB 1.86fF $ **FLOATING
C2375 S.n2146 SUB 2.64fF $ **FLOATING
C2376 S.t349 SUB 0.02fF
C2377 S.n2147 SUB 0.24fF $ **FLOATING
C2378 S.n2148 SUB 0.35fF $ **FLOATING
C2379 S.n2149 SUB 0.60fF $ **FLOATING
C2380 S.n2150 SUB 0.12fF $ **FLOATING
C2381 S.t919 SUB 0.02fF
C2382 S.n2151 SUB 0.14fF $ **FLOATING
C2383 S.n2153 SUB 1.86fF $ **FLOATING
C2384 S.n2154 SUB 2.65fF $ **FLOATING
C2385 S.t76 SUB 0.02fF
C2386 S.n2155 SUB 0.24fF $ **FLOATING
C2387 S.n2156 SUB 0.35fF $ **FLOATING
C2388 S.n2157 SUB 0.60fF $ **FLOATING
C2389 S.t815 SUB 0.02fF
C2390 S.n2158 SUB 1.20fF $ **FLOATING
C2391 S.n2159 SUB 0.60fF $ **FLOATING
C2392 S.n2160 SUB 0.35fF $ **FLOATING
C2393 S.n2161 SUB 0.62fF $ **FLOATING
C2394 S.n2162 SUB 1.14fF $ **FLOATING
C2395 S.n2163 SUB 2.18fF $ **FLOATING
C2396 S.n2164 SUB 0.59fF $ **FLOATING
C2397 S.n2165 SUB 0.02fF $ **FLOATING
C2398 S.n2166 SUB 0.96fF $ **FLOATING
C2399 S.t75 SUB 14.50fF
C2400 S.n2167 SUB 14.37fF $ **FLOATING
C2401 S.n2169 SUB 0.37fF $ **FLOATING
C2402 S.n2170 SUB 0.23fF $ **FLOATING
C2403 S.n2171 SUB 2.87fF $ **FLOATING
C2404 S.n2172 SUB 2.43fF $ **FLOATING
C2405 S.n2173 SUB 1.94fF $ **FLOATING
C2406 S.n2174 SUB 3.89fF $ **FLOATING
C2407 S.n2175 SUB 0.25fF $ **FLOATING
C2408 S.n2176 SUB 0.01fF $ **FLOATING
C2409 S.t673 SUB 0.02fF
C2410 S.n2177 SUB 0.25fF $ **FLOATING
C2411 S.t592 SUB 0.02fF
C2412 S.n2178 SUB 0.94fF $ **FLOATING
C2413 S.n2179 SUB 0.70fF $ **FLOATING
C2414 S.n2180 SUB 0.77fF $ **FLOATING
C2415 S.n2181 SUB 1.91fF $ **FLOATING
C2416 S.n2182 SUB 1.86fF $ **FLOATING
C2417 S.n2183 SUB 0.12fF $ **FLOATING
C2418 S.t336 SUB 0.02fF
C2419 S.n2184 SUB 0.14fF $ **FLOATING
C2420 S.t437 SUB 0.02fF
C2421 S.n2186 SUB 0.24fF $ **FLOATING
C2422 S.n2187 SUB 0.35fF $ **FLOATING
C2423 S.n2188 SUB 0.60fF $ **FLOATING
C2424 S.n2189 SUB 1.50fF $ **FLOATING
C2425 S.n2190 SUB 2.96fF $ **FLOATING
C2426 S.t195 SUB 0.02fF
C2427 S.n2191 SUB 0.24fF $ **FLOATING
C2428 S.n2192 SUB 0.90fF $ **FLOATING
C2429 S.n2193 SUB 0.05fF $ **FLOATING
C2430 S.t658 SUB 0.02fF
C2431 S.n2194 SUB 0.12fF $ **FLOATING
C2432 S.n2195 SUB 0.14fF $ **FLOATING
C2433 S.n2197 SUB 1.87fF $ **FLOATING
C2434 S.n2198 SUB 1.86fF $ **FLOATING
C2435 S.t925 SUB 0.02fF
C2436 S.n2199 SUB 0.24fF $ **FLOATING
C2437 S.n2200 SUB 0.35fF $ **FLOATING
C2438 S.n2201 SUB 0.60fF $ **FLOATING
C2439 S.n2202 SUB 0.12fF $ **FLOATING
C2440 S.t135 SUB 0.02fF
C2441 S.n2203 SUB 0.14fF $ **FLOATING
C2442 S.n2205 SUB 1.14fF $ **FLOATING
C2443 S.n2206 SUB 0.22fF $ **FLOATING
C2444 S.n2207 SUB 0.25fF $ **FLOATING
C2445 S.n2208 SUB 0.09fF $ **FLOATING
C2446 S.n2209 SUB 1.86fF $ **FLOATING
C2447 S.t243 SUB 0.02fF
C2448 S.n2210 SUB 0.24fF $ **FLOATING
C2449 S.n2211 SUB 0.90fF $ **FLOATING
C2450 S.n2212 SUB 0.05fF $ **FLOATING
C2451 S.t288 SUB 0.02fF
C2452 S.n2213 SUB 0.12fF $ **FLOATING
C2453 S.n2214 SUB 0.14fF $ **FLOATING
C2454 S.n2216 SUB 0.77fF $ **FLOATING
C2455 S.n2217 SUB 1.92fF $ **FLOATING
C2456 S.n2218 SUB 1.86fF $ **FLOATING
C2457 S.n2219 SUB 0.12fF $ **FLOATING
C2458 S.t863 SUB 0.02fF
C2459 S.n2220 SUB 0.14fF $ **FLOATING
C2460 S.t547 SUB 0.02fF
C2461 S.n2222 SUB 0.24fF $ **FLOATING
C2462 S.n2223 SUB 0.35fF $ **FLOATING
C2463 S.n2224 SUB 0.60fF $ **FLOATING
C2464 S.n2225 SUB 1.82fF $ **FLOATING
C2465 S.n2226 SUB 2.96fF $ **FLOATING
C2466 S.t968 SUB 0.02fF
C2467 S.n2227 SUB 0.24fF $ **FLOATING
C2468 S.n2228 SUB 0.90fF $ **FLOATING
C2469 S.n2229 SUB 0.05fF $ **FLOATING
C2470 S.t17 SUB 0.02fF
C2471 S.n2230 SUB 0.12fF $ **FLOATING
C2472 S.n2231 SUB 0.14fF $ **FLOATING
C2473 S.n2233 SUB 1.87fF $ **FLOATING
C2474 S.n2234 SUB 1.73fF $ **FLOATING
C2475 S.t158 SUB 0.02fF
C2476 S.n2235 SUB 0.24fF $ **FLOATING
C2477 S.n2236 SUB 0.35fF $ **FLOATING
C2478 S.n2237 SUB 0.60fF $ **FLOATING
C2479 S.n2238 SUB 0.12fF $ **FLOATING
C2480 S.t488 SUB 0.02fF
C2481 S.n2239 SUB 0.14fF $ **FLOATING
C2482 S.n2241 SUB 1.14fF $ **FLOATING
C2483 S.n2242 SUB 0.22fF $ **FLOATING
C2484 S.n2243 SUB 0.25fF $ **FLOATING
C2485 S.n2244 SUB 0.09fF $ **FLOATING
C2486 S.n2245 SUB 2.41fF $ **FLOATING
C2487 S.t591 SUB 0.02fF
C2488 S.n2246 SUB 0.24fF $ **FLOATING
C2489 S.n2247 SUB 0.90fF $ **FLOATING
C2490 S.n2248 SUB 0.05fF $ **FLOATING
C2491 S.t771 SUB 0.02fF
C2492 S.n2249 SUB 0.12fF $ **FLOATING
C2493 S.n2250 SUB 0.14fF $ **FLOATING
C2494 S.n2252 SUB 1.86fF $ **FLOATING
C2495 S.n2253 SUB 0.47fF $ **FLOATING
C2496 S.n2254 SUB 0.09fF $ **FLOATING
C2497 S.n2255 SUB 0.32fF $ **FLOATING
C2498 S.n2256 SUB 0.30fF $ **FLOATING
C2499 S.n2257 SUB 0.76fF $ **FLOATING
C2500 S.n2258 SUB 0.58fF $ **FLOATING
C2501 S.t886 SUB 0.02fF
C2502 S.n2259 SUB 0.24fF $ **FLOATING
C2503 S.n2260 SUB 0.35fF $ **FLOATING
C2504 S.n2261 SUB 0.60fF $ **FLOATING
C2505 S.n2262 SUB 0.12fF $ **FLOATING
C2506 S.t98 SUB 0.02fF
C2507 S.n2263 SUB 0.14fF $ **FLOATING
C2508 S.n2265 SUB 2.58fF $ **FLOATING
C2509 S.n2266 SUB 2.13fF $ **FLOATING
C2510 S.t194 SUB 0.02fF
C2511 S.n2267 SUB 0.24fF $ **FLOATING
C2512 S.n2268 SUB 0.90fF $ **FLOATING
C2513 S.n2269 SUB 0.05fF $ **FLOATING
C2514 S.t390 SUB 0.02fF
C2515 S.n2270 SUB 0.12fF $ **FLOATING
C2516 S.n2271 SUB 0.14fF $ **FLOATING
C2517 S.n2273 SUB 0.77fF $ **FLOATING
C2518 S.n2274 SUB 2.27fF $ **FLOATING
C2519 S.n2275 SUB 1.86fF $ **FLOATING
C2520 S.n2276 SUB 0.12fF $ **FLOATING
C2521 S.t832 SUB 0.02fF
C2522 S.n2277 SUB 0.14fF $ **FLOATING
C2523 S.t509 SUB 0.02fF
C2524 S.n2279 SUB 0.24fF $ **FLOATING
C2525 S.n2280 SUB 0.35fF $ **FLOATING
C2526 S.n2281 SUB 0.60fF $ **FLOATING
C2527 S.n2282 SUB 1.37fF $ **FLOATING
C2528 S.n2283 SUB 0.70fF $ **FLOATING
C2529 S.n2284 SUB 1.13fF $ **FLOATING
C2530 S.n2285 SUB 0.35fF $ **FLOATING
C2531 S.n2286 SUB 2.00fF $ **FLOATING
C2532 S.t915 SUB 0.02fF
C2533 S.n2287 SUB 0.24fF $ **FLOATING
C2534 S.n2288 SUB 0.90fF $ **FLOATING
C2535 S.n2289 SUB 0.05fF $ **FLOATING
C2536 S.t1109 SUB 0.02fF
C2537 S.n2290 SUB 0.12fF $ **FLOATING
C2538 S.n2291 SUB 0.14fF $ **FLOATING
C2539 S.n2293 SUB 1.87fF $ **FLOATING
C2540 S.n2294 SUB 1.86fF $ **FLOATING
C2541 S.t116 SUB 0.02fF
C2542 S.n2295 SUB 0.24fF $ **FLOATING
C2543 S.n2296 SUB 0.35fF $ **FLOATING
C2544 S.n2297 SUB 0.60fF $ **FLOATING
C2545 S.n2298 SUB 0.12fF $ **FLOATING
C2546 S.t455 SUB 0.02fF
C2547 S.n2299 SUB 0.14fF $ **FLOATING
C2548 S.n2301 SUB 1.14fF $ **FLOATING
C2549 S.n2302 SUB 0.22fF $ **FLOATING
C2550 S.n2303 SUB 0.25fF $ **FLOATING
C2551 S.n2304 SUB 0.09fF $ **FLOATING
C2552 S.n2305 SUB 1.86fF $ **FLOATING
C2553 S.t538 SUB 0.02fF
C2554 S.n2306 SUB 0.24fF $ **FLOATING
C2555 S.n2307 SUB 0.90fF $ **FLOATING
C2556 S.n2308 SUB 0.05fF $ **FLOATING
C2557 S.t798 SUB 0.02fF
C2558 S.n2309 SUB 0.12fF $ **FLOATING
C2559 S.n2310 SUB 0.14fF $ **FLOATING
C2560 S.n2312 SUB 14.09fF $ **FLOATING
C2561 S.n2313 SUB 2.70fF $ **FLOATING
C2562 S.n2314 SUB 1.58fF $ **FLOATING
C2563 S.n2315 SUB 0.12fF $ **FLOATING
C2564 S.t849 SUB 0.02fF
C2565 S.n2316 SUB 0.14fF $ **FLOATING
C2566 S.t323 SUB 0.02fF
C2567 S.n2318 SUB 0.24fF $ **FLOATING
C2568 S.n2319 SUB 0.35fF $ **FLOATING
C2569 S.n2320 SUB 0.60fF $ **FLOATING
C2570 S.n2321 SUB 0.07fF $ **FLOATING
C2571 S.n2322 SUB 0.01fF $ **FLOATING
C2572 S.n2323 SUB 0.23fF $ **FLOATING
C2573 S.n2324 SUB 1.15fF $ **FLOATING
C2574 S.n2325 SUB 1.33fF $ **FLOATING
C2575 S.n2326 SUB 2.28fF $ **FLOATING
C2576 S.t51 SUB 0.02fF
C2577 S.n2327 SUB 0.12fF $ **FLOATING
C2578 S.n2328 SUB 0.14fF $ **FLOATING
C2579 S.t490 SUB 0.02fF
C2580 S.n2330 SUB 0.24fF $ **FLOATING
C2581 S.n2331 SUB 0.90fF $ **FLOATING
C2582 S.n2332 SUB 0.05fF $ **FLOATING
C2583 S.t16 SUB 32.35fF
C2584 S.t502 SUB 0.02fF
C2585 S.n2333 SUB 0.24fF $ **FLOATING
C2586 S.n2334 SUB 0.90fF $ **FLOATING
C2587 S.n2335 SUB 0.05fF $ **FLOATING
C2588 S.t748 SUB 0.02fF
C2589 S.n2336 SUB 0.12fF $ **FLOATING
C2590 S.n2337 SUB 0.14fF $ **FLOATING
C2591 S.n2339 SUB 0.12fF $ **FLOATING
C2592 S.t407 SUB 0.02fF
C2593 S.n2340 SUB 0.14fF $ **FLOATING
C2594 S.n2342 SUB 5.11fF $ **FLOATING
C2595 S.n2343 SUB 5.38fF $ **FLOATING
C2596 S.t1082 SUB 0.02fF
C2597 S.n2344 SUB 0.12fF $ **FLOATING
C2598 S.n2345 SUB 0.14fF $ **FLOATING
C2599 S.t955 SUB 0.02fF
C2600 S.n2347 SUB 0.24fF $ **FLOATING
C2601 S.n2348 SUB 0.90fF $ **FLOATING
C2602 S.n2349 SUB 0.05fF $ **FLOATING
C2603 S.t47 SUB 31.97fF
C2604 S.t588 SUB 0.02fF
C2605 S.n2350 SUB 1.18fF $ **FLOATING
C2606 S.n2351 SUB 0.05fF $ **FLOATING
C2607 S.t610 SUB 0.02fF
C2608 S.n2352 SUB 0.01fF $ **FLOATING
C2609 S.n2353 SUB 0.25fF $ **FLOATING
C2610 S.n2355 SUB 1.48fF $ **FLOATING
C2611 S.n2356 SUB 1.29fF $ **FLOATING
C2612 S.n2357 SUB 0.27fF $ **FLOATING
C2613 S.n2358 SUB 0.24fF $ **FLOATING
C2614 S.n2359 SUB 4.34fF $ **FLOATING
C2615 S.n2360 SUB 0.24fF $ **FLOATING
C2616 S.n2361 SUB 1.48fF $ **FLOATING
C2617 S.n2362 SUB 1.28fF $ **FLOATING
C2618 S.n2363 SUB 0.27fF $ **FLOATING
C2619 S.n2364 SUB 1.87fF $ **FLOATING
C2620 S.n2365 SUB 0.06fF $ **FLOATING
C2621 S.n2366 SUB 0.03fF $ **FLOATING
C2622 S.n2367 SUB 0.03fF $ **FLOATING
C2623 S.n2368 SUB 0.98fF $ **FLOATING
C2624 S.n2369 SUB 0.02fF $ **FLOATING
C2625 S.n2370 SUB 0.01fF $ **FLOATING
C2626 S.n2371 SUB 0.02fF $ **FLOATING
C2627 S.n2372 SUB 0.08fF $ **FLOATING
C2628 S.n2373 SUB 0.36fF $ **FLOATING
C2629 S.n2374 SUB 1.83fF $ **FLOATING
C2630 S.t877 SUB 0.02fF
C2631 S.n2375 SUB 0.24fF $ **FLOATING
C2632 S.n2376 SUB 0.35fF $ **FLOATING
C2633 S.n2377 SUB 0.60fF $ **FLOATING
C2634 S.n2378 SUB 0.12fF $ **FLOATING
C2635 S.t653 SUB 0.02fF
C2636 S.n2379 SUB 0.14fF $ **FLOATING
C2637 S.n2381 SUB 0.69fF $ **FLOATING
C2638 S.n2382 SUB 0.22fF $ **FLOATING
C2639 S.n2383 SUB 0.22fF $ **FLOATING
C2640 S.n2384 SUB 0.69fF $ **FLOATING
C2641 S.n2385 SUB 1.14fF $ **FLOATING
C2642 S.n2386 SUB 0.22fF $ **FLOATING
C2643 S.n2387 SUB 0.25fF $ **FLOATING
C2644 S.n2388 SUB 0.09fF $ **FLOATING
C2645 S.n2389 SUB 1.86fF $ **FLOATING
C2646 S.t134 SUB 0.02fF
C2647 S.n2390 SUB 0.24fF $ **FLOATING
C2648 S.n2391 SUB 0.90fF $ **FLOATING
C2649 S.n2392 SUB 0.05fF $ **FLOATING
C2650 S.t702 SUB 0.02fF
C2651 S.n2393 SUB 0.12fF $ **FLOATING
C2652 S.n2394 SUB 0.14fF $ **FLOATING
C2653 S.n2396 SUB 0.25fF $ **FLOATING
C2654 S.n2397 SUB 0.09fF $ **FLOATING
C2655 S.n2398 SUB 0.21fF $ **FLOATING
C2656 S.n2399 SUB 0.91fF $ **FLOATING
C2657 S.n2400 SUB 0.44fF $ **FLOATING
C2658 S.n2401 SUB 1.86fF $ **FLOATING
C2659 S.n2402 SUB 0.12fF $ **FLOATING
C2660 S.t353 SUB 0.02fF
C2661 S.n2403 SUB 0.14fF $ **FLOATING
C2662 S.t634 SUB 0.02fF
C2663 S.n2405 SUB 0.24fF $ **FLOATING
C2664 S.n2406 SUB 0.35fF $ **FLOATING
C2665 S.n2407 SUB 0.60fF $ **FLOATING
C2666 S.n2408 SUB 0.02fF $ **FLOATING
C2667 S.n2409 SUB 0.01fF $ **FLOATING
C2668 S.n2410 SUB 0.02fF $ **FLOATING
C2669 S.n2411 SUB 0.08fF $ **FLOATING
C2670 S.n2412 SUB 0.06fF $ **FLOATING
C2671 S.n2413 SUB 0.03fF $ **FLOATING
C2672 S.n2414 SUB 0.03fF $ **FLOATING
C2673 S.n2415 SUB 0.99fF $ **FLOATING
C2674 S.n2416 SUB 0.35fF $ **FLOATING
C2675 S.n2417 SUB 1.85fF $ **FLOATING
C2676 S.n2418 SUB 1.97fF $ **FLOATING
C2677 S.t590 SUB 0.02fF
C2678 S.n2419 SUB 0.24fF $ **FLOATING
C2679 S.n2420 SUB 0.90fF $ **FLOATING
C2680 S.n2421 SUB 0.05fF $ **FLOATING
C2681 S.t467 SUB 0.02fF
C2682 S.n2422 SUB 0.12fF $ **FLOATING
C2683 S.n2423 SUB 0.14fF $ **FLOATING
C2684 S.n2425 SUB 1.87fF $ **FLOATING
C2685 S.n2426 SUB 0.04fF $ **FLOATING
C2686 S.n2427 SUB 0.07fF $ **FLOATING
C2687 S.n2428 SUB 0.05fF $ **FLOATING
C2688 S.n2429 SUB 0.86fF $ **FLOATING
C2689 S.n2430 SUB 0.01fF $ **FLOATING
C2690 S.n2431 SUB 0.01fF $ **FLOATING
C2691 S.n2432 SUB 0.01fF $ **FLOATING
C2692 S.n2433 SUB 0.07fF $ **FLOATING
C2693 S.n2434 SUB 0.68fF $ **FLOATING
C2694 S.n2435 SUB 0.71fF $ **FLOATING
C2695 S.t251 SUB 0.02fF
C2696 S.n2436 SUB 0.24fF $ **FLOATING
C2697 S.n2437 SUB 0.35fF $ **FLOATING
C2698 S.n2438 SUB 0.60fF $ **FLOATING
C2699 S.n2439 SUB 0.12fF $ **FLOATING
C2700 S.t1080 SUB 0.02fF
C2701 S.n2440 SUB 0.14fF $ **FLOATING
C2702 S.n2442 SUB 0.69fF $ **FLOATING
C2703 S.n2443 SUB 0.22fF $ **FLOATING
C2704 S.n2444 SUB 0.22fF $ **FLOATING
C2705 S.n2445 SUB 0.69fF $ **FLOATING
C2706 S.n2446 SUB 1.14fF $ **FLOATING
C2707 S.n2447 SUB 0.22fF $ **FLOATING
C2708 S.n2448 SUB 0.25fF $ **FLOATING
C2709 S.n2449 SUB 0.09fF $ **FLOATING
C2710 S.n2450 SUB 2.29fF $ **FLOATING
C2711 S.t193 SUB 0.02fF
C2712 S.n2451 SUB 0.24fF $ **FLOATING
C2713 S.n2452 SUB 0.90fF $ **FLOATING
C2714 S.n2453 SUB 0.05fF $ **FLOATING
C2715 S.t67 SUB 0.02fF
C2716 S.n2454 SUB 0.12fF $ **FLOATING
C2717 S.n2455 SUB 0.14fF $ **FLOATING
C2718 S.n2457 SUB 1.86fF $ **FLOATING
C2719 S.n2458 SUB 0.45fF $ **FLOATING
C2720 S.n2459 SUB 0.22fF $ **FLOATING
C2721 S.n2460 SUB 0.38fF $ **FLOATING
C2722 S.n2461 SUB 0.16fF $ **FLOATING
C2723 S.n2462 SUB 0.28fF $ **FLOATING
C2724 S.n2463 SUB 0.21fF $ **FLOATING
C2725 S.n2464 SUB 0.30fF $ **FLOATING
C2726 S.n2465 SUB 0.41fF $ **FLOATING
C2727 S.n2466 SUB 0.20fF $ **FLOATING
C2728 S.t971 SUB 0.02fF
C2729 S.n2467 SUB 0.24fF $ **FLOATING
C2730 S.n2468 SUB 0.35fF $ **FLOATING
C2731 S.n2469 SUB 0.60fF $ **FLOATING
C2732 S.n2470 SUB 0.12fF $ **FLOATING
C2733 S.t697 SUB 0.02fF
C2734 S.n2471 SUB 0.14fF $ **FLOATING
C2735 S.n2473 SUB 0.04fF $ **FLOATING
C2736 S.n2474 SUB 0.03fF $ **FLOATING
C2737 S.n2475 SUB 0.03fF $ **FLOATING
C2738 S.n2476 SUB 0.10fF $ **FLOATING
C2739 S.n2477 SUB 0.36fF $ **FLOATING
C2740 S.n2478 SUB 0.37fF $ **FLOATING
C2741 S.n2479 SUB 0.10fF $ **FLOATING
C2742 S.n2480 SUB 0.12fF $ **FLOATING
C2743 S.n2481 SUB 0.07fF $ **FLOATING
C2744 S.n2482 SUB 0.12fF $ **FLOATING
C2745 S.n2483 SUB 0.18fF $ **FLOATING
C2746 S.n2484 SUB 3.95fF $ **FLOATING
C2747 S.t916 SUB 0.02fF
C2748 S.n2485 SUB 0.24fF $ **FLOATING
C2749 S.n2486 SUB 0.90fF $ **FLOATING
C2750 S.n2487 SUB 0.05fF $ **FLOATING
C2751 S.t807 SUB 0.02fF
C2752 S.n2488 SUB 0.12fF $ **FLOATING
C2753 S.n2489 SUB 0.14fF $ **FLOATING
C2754 S.n2491 SUB 0.25fF $ **FLOATING
C2755 S.n2492 SUB 0.09fF $ **FLOATING
C2756 S.n2493 SUB 0.21fF $ **FLOATING
C2757 S.n2494 SUB 1.27fF $ **FLOATING
C2758 S.n2495 SUB 0.52fF $ **FLOATING
C2759 S.n2496 SUB 1.86fF $ **FLOATING
C2760 S.n2497 SUB 0.12fF $ **FLOATING
C2761 S.t314 SUB 0.02fF
C2762 S.n2498 SUB 0.14fF $ **FLOATING
C2763 S.t597 SUB 0.02fF
C2764 S.n2500 SUB 0.24fF $ **FLOATING
C2765 S.n2501 SUB 0.35fF $ **FLOATING
C2766 S.n2502 SUB 0.60fF $ **FLOATING
C2767 S.n2503 SUB 1.56fF $ **FLOATING
C2768 S.n2504 SUB 2.42fF $ **FLOATING
C2769 S.t539 SUB 0.02fF
C2770 S.n2505 SUB 0.24fF $ **FLOATING
C2771 S.n2506 SUB 0.90fF $ **FLOATING
C2772 S.n2507 SUB 0.05fF $ **FLOATING
C2773 S.t426 SUB 0.02fF
C2774 S.n2508 SUB 0.12fF $ **FLOATING
C2775 S.n2509 SUB 0.14fF $ **FLOATING
C2776 S.n2511 SUB 1.87fF $ **FLOATING
C2777 S.n2512 SUB 0.06fF $ **FLOATING
C2778 S.n2513 SUB 0.03fF $ **FLOATING
C2779 S.n2514 SUB 0.03fF $ **FLOATING
C2780 S.n2515 SUB 0.98fF $ **FLOATING
C2781 S.n2516 SUB 0.02fF $ **FLOATING
C2782 S.n2517 SUB 0.01fF $ **FLOATING
C2783 S.n2518 SUB 0.02fF $ **FLOATING
C2784 S.n2519 SUB 0.08fF $ **FLOATING
C2785 S.n2520 SUB 0.36fF $ **FLOATING
C2786 S.n2521 SUB 1.83fF $ **FLOATING
C2787 S.t275 SUB 0.02fF
C2788 S.n2522 SUB 0.24fF $ **FLOATING
C2789 S.n2523 SUB 0.35fF $ **FLOATING
C2790 S.n2524 SUB 0.60fF $ **FLOATING
C2791 S.n2525 SUB 0.12fF $ **FLOATING
C2792 S.t1100 SUB 0.02fF
C2793 S.n2526 SUB 0.14fF $ **FLOATING
C2794 S.n2528 SUB 0.69fF $ **FLOATING
C2795 S.n2529 SUB 0.22fF $ **FLOATING
C2796 S.n2530 SUB 0.22fF $ **FLOATING
C2797 S.n2531 SUB 0.69fF $ **FLOATING
C2798 S.n2532 SUB 1.14fF $ **FLOATING
C2799 S.n2533 SUB 0.22fF $ **FLOATING
C2800 S.n2534 SUB 0.25fF $ **FLOATING
C2801 S.n2535 SUB 0.09fF $ **FLOATING
C2802 S.n2536 SUB 1.86fF $ **FLOATING
C2803 S.t221 SUB 0.02fF
C2804 S.n2537 SUB 0.24fF $ **FLOATING
C2805 S.n2538 SUB 0.90fF $ **FLOATING
C2806 S.n2539 SUB 0.05fF $ **FLOATING
C2807 S.t1145 SUB 0.02fF
C2808 S.n2540 SUB 0.12fF $ **FLOATING
C2809 S.n2541 SUB 0.14fF $ **FLOATING
C2810 S.n2543 SUB 14.09fF $ **FLOATING
C2811 S.n2544 SUB 0.06fF $ **FLOATING
C2812 S.n2545 SUB 0.20fF $ **FLOATING
C2813 S.n2546 SUB 0.09fF $ **FLOATING
C2814 S.n2547 SUB 0.20fF $ **FLOATING
C2815 S.n2548 SUB 0.09fF $ **FLOATING
C2816 S.n2549 SUB 0.30fF $ **FLOATING
C2817 S.n2550 SUB 0.69fF $ **FLOATING
C2818 S.n2551 SUB 0.44fF $ **FLOATING
C2819 S.n2552 SUB 2.31fF $ **FLOATING
C2820 S.n2553 SUB 0.12fF $ **FLOATING
C2821 S.t1027 SUB 0.02fF
C2822 S.n2554 SUB 0.14fF $ **FLOATING
C2823 S.t147 SUB 0.02fF
C2824 S.n2556 SUB 0.24fF $ **FLOATING
C2825 S.n2557 SUB 0.35fF $ **FLOATING
C2826 S.n2558 SUB 0.60fF $ **FLOATING
C2827 S.n2559 SUB 1.88fF $ **FLOATING
C2828 S.n2560 SUB 0.17fF $ **FLOATING
C2829 S.n2561 SUB 0.76fF $ **FLOATING
C2830 S.n2562 SUB 0.31fF $ **FLOATING
C2831 S.n2563 SUB 0.25fF $ **FLOATING
C2832 S.n2564 SUB 0.29fF $ **FLOATING
C2833 S.n2565 SUB 0.46fF $ **FLOATING
C2834 S.n2566 SUB 0.16fF $ **FLOATING
C2835 S.n2567 SUB 1.91fF $ **FLOATING
C2836 S.t1043 SUB 0.02fF
C2837 S.n2568 SUB 0.12fF $ **FLOATING
C2838 S.n2569 SUB 0.14fF $ **FLOATING
C2839 S.t524 SUB 0.02fF
C2840 S.n2571 SUB 0.24fF $ **FLOATING
C2841 S.n2572 SUB 0.90fF $ **FLOATING
C2842 S.n2573 SUB 0.05fF $ **FLOATING
C2843 S.n2574 SUB 1.86fF $ **FLOATING
C2844 S.n2575 SUB 0.12fF $ **FLOATING
C2845 S.t61 SUB 0.02fF
C2846 S.n2576 SUB 0.14fF $ **FLOATING
C2847 S.t435 SUB 0.02fF
C2848 S.n2578 SUB 0.12fF $ **FLOATING
C2849 S.n2579 SUB 0.14fF $ **FLOATING
C2850 S.t161 SUB 0.02fF
C2851 S.n2581 SUB 0.24fF $ **FLOATING
C2852 S.n2582 SUB 0.90fF $ **FLOATING
C2853 S.n2583 SUB 0.05fF $ **FLOATING
C2854 S.t859 SUB 0.02fF
C2855 S.n2584 SUB 0.24fF $ **FLOATING
C2856 S.n2585 SUB 0.35fF $ **FLOATING
C2857 S.n2586 SUB 0.60fF $ **FLOATING
C2858 S.n2587 SUB 0.31fF $ **FLOATING
C2859 S.n2588 SUB 1.08fF $ **FLOATING
C2860 S.n2589 SUB 0.15fF $ **FLOATING
C2861 S.n2590 SUB 2.08fF $ **FLOATING
C2862 S.n2591 SUB 2.91fF $ **FLOATING
C2863 S.n2592 SUB 1.86fF $ **FLOATING
C2864 S.n2593 SUB 0.12fF $ **FLOATING
C2865 S.t712 SUB 0.02fF
C2866 S.n2594 SUB 0.14fF $ **FLOATING
C2867 S.t992 SUB 0.02fF
C2868 S.n2596 SUB 0.24fF $ **FLOATING
C2869 S.n2597 SUB 0.35fF $ **FLOATING
C2870 S.n2598 SUB 0.60fF $ **FLOATING
C2871 S.n2599 SUB 0.91fF $ **FLOATING
C2872 S.n2600 SUB 0.31fF $ **FLOATING
C2873 S.n2601 SUB 0.91fF $ **FLOATING
C2874 S.n2602 SUB 1.08fF $ **FLOATING
C2875 S.n2603 SUB 0.15fF $ **FLOATING
C2876 S.n2604 SUB 4.90fF $ **FLOATING
C2877 S.t752 SUB 0.02fF
C2878 S.n2605 SUB 0.12fF $ **FLOATING
C2879 S.n2606 SUB 0.14fF $ **FLOATING
C2880 S.t943 SUB 0.02fF
C2881 S.n2608 SUB 0.24fF $ **FLOATING
C2882 S.n2609 SUB 0.90fF $ **FLOATING
C2883 S.n2610 SUB 0.05fF $ **FLOATING
C2884 S.n2611 SUB 1.86fF $ **FLOATING
C2885 S.n2612 SUB 2.64fF $ **FLOATING
C2886 S.t616 SUB 0.02fF
C2887 S.n2613 SUB 0.24fF $ **FLOATING
C2888 S.n2614 SUB 0.35fF $ **FLOATING
C2889 S.n2615 SUB 0.60fF $ **FLOATING
C2890 S.n2616 SUB 0.12fF $ **FLOATING
C2891 S.t331 SUB 0.02fF
C2892 S.n2617 SUB 0.14fF $ **FLOATING
C2893 S.n2619 SUB 1.86fF $ **FLOATING
C2894 S.n2620 SUB 2.64fF $ **FLOATING
C2895 S.t483 SUB 0.02fF
C2896 S.n2621 SUB 0.24fF $ **FLOATING
C2897 S.n2622 SUB 0.35fF $ **FLOATING
C2898 S.n2623 SUB 0.60fF $ **FLOATING
C2899 S.t888 SUB 0.02fF
C2900 S.n2624 SUB 0.24fF $ **FLOATING
C2901 S.n2625 SUB 0.90fF $ **FLOATING
C2902 S.n2626 SUB 0.05fF $ **FLOATING
C2903 S.t1 SUB 0.02fF
C2904 S.n2627 SUB 0.12fF $ **FLOATING
C2905 S.n2628 SUB 0.14fF $ **FLOATING
C2906 S.n2630 SUB 0.12fF $ **FLOATING
C2907 S.t804 SUB 0.02fF
C2908 S.n2631 SUB 0.14fF $ **FLOATING
C2909 S.n2633 SUB 2.28fF $ **FLOATING
C2910 S.n2634 SUB 2.91fF $ **FLOATING
C2911 S.n2635 SUB 5.10fF $ **FLOATING
C2912 S.t367 SUB 0.02fF
C2913 S.n2636 SUB 0.12fF $ **FLOATING
C2914 S.n2637 SUB 0.14fF $ **FLOATING
C2915 S.t564 SUB 0.02fF
C2916 S.n2639 SUB 0.24fF $ **FLOATING
C2917 S.n2640 SUB 0.90fF $ **FLOATING
C2918 S.n2641 SUB 0.05fF $ **FLOATING
C2919 S.n2642 SUB 1.86fF $ **FLOATING
C2920 S.n2643 SUB 2.64fF $ **FLOATING
C2921 S.t228 SUB 0.02fF
C2922 S.n2644 SUB 0.24fF $ **FLOATING
C2923 S.n2645 SUB 0.35fF $ **FLOATING
C2924 S.n2646 SUB 0.60fF $ **FLOATING
C2925 S.n2647 SUB 0.12fF $ **FLOATING
C2926 S.t1057 SUB 0.02fF
C2927 S.n2648 SUB 0.14fF $ **FLOATING
C2928 S.n2650 SUB 4.84fF $ **FLOATING
C2929 S.t1091 SUB 0.02fF
C2930 S.n2651 SUB 0.12fF $ **FLOATING
C2931 S.n2652 SUB 0.14fF $ **FLOATING
C2932 S.t171 SUB 0.02fF
C2933 S.n2654 SUB 0.24fF $ **FLOATING
C2934 S.n2655 SUB 0.90fF $ **FLOATING
C2935 S.n2656 SUB 0.05fF $ **FLOATING
C2936 S.n2657 SUB 1.86fF $ **FLOATING
C2937 S.n2658 SUB 2.64fF $ **FLOATING
C2938 S.t880 SUB 0.02fF
C2939 S.n2659 SUB 0.24fF $ **FLOATING
C2940 S.n2660 SUB 0.35fF $ **FLOATING
C2941 S.n2661 SUB 0.60fF $ **FLOATING
C2942 S.n2662 SUB 0.12fF $ **FLOATING
C2943 S.t308 SUB 0.02fF
C2944 S.n2663 SUB 0.14fF $ **FLOATING
C2945 S.n2665 SUB 1.86fF $ **FLOATING
C2946 S.n2666 SUB 2.65fF $ **FLOATING
C2947 S.t823 SUB 0.02fF
C2948 S.n2667 SUB 0.24fF $ **FLOATING
C2949 S.n2668 SUB 0.35fF $ **FLOATING
C2950 S.n2669 SUB 0.60fF $ **FLOATING
C2951 S.t674 SUB 0.02fF
C2952 S.n2670 SUB 1.20fF $ **FLOATING
C2953 S.n2671 SUB 0.36fF $ **FLOATING
C2954 S.n2672 SUB 1.21fF $ **FLOATING
C2955 S.n2673 SUB 0.60fF $ **FLOATING
C2956 S.n2674 SUB 0.35fF $ **FLOATING
C2957 S.n2675 SUB 0.62fF $ **FLOATING
C2958 S.n2676 SUB 1.14fF $ **FLOATING
C2959 S.n2677 SUB 2.18fF $ **FLOATING
C2960 S.n2678 SUB 0.59fF $ **FLOATING
C2961 S.n2679 SUB 0.02fF $ **FLOATING
C2962 S.n2680 SUB 0.96fF $ **FLOATING
C2963 S.t89 SUB 14.50fF
C2964 S.n2681 SUB 14.37fF $ **FLOATING
C2965 S.n2683 SUB 0.37fF $ **FLOATING
C2966 S.n2684 SUB 0.23fF $ **FLOATING
C2967 S.n2685 SUB 2.76fF $ **FLOATING
C2968 S.n2686 SUB 2.43fF $ **FLOATING
C2969 S.n2687 SUB 3.95fF $ **FLOATING
C2970 S.n2688 SUB 0.25fF $ **FLOATING
C2971 S.n2689 SUB 0.01fF $ **FLOATING
C2972 S.t579 SUB 0.02fF
C2973 S.n2690 SUB 0.25fF $ **FLOATING
C2974 S.t454 SUB 0.02fF
C2975 S.n2691 SUB 0.94fF $ **FLOATING
C2976 S.n2692 SUB 0.70fF $ **FLOATING
C2977 S.n2693 SUB 1.87fF $ **FLOATING
C2978 S.n2694 SUB 1.86fF $ **FLOATING
C2979 S.t302 SUB 0.02fF
C2980 S.n2695 SUB 0.24fF $ **FLOATING
C2981 S.n2696 SUB 0.35fF $ **FLOATING
C2982 S.n2697 SUB 0.60fF $ **FLOATING
C2983 S.n2698 SUB 0.12fF $ **FLOATING
C2984 S.t257 SUB 0.02fF
C2985 S.n2699 SUB 0.14fF $ **FLOATING
C2986 S.n2701 SUB 1.14fF $ **FLOATING
C2987 S.n2702 SUB 0.22fF $ **FLOATING
C2988 S.n2703 SUB 0.25fF $ **FLOATING
C2989 S.n2704 SUB 0.09fF $ **FLOATING
C2990 S.n2705 SUB 1.86fF $ **FLOATING
C2991 S.t45 SUB 0.02fF
C2992 S.n2706 SUB 0.24fF $ **FLOATING
C2993 S.n2707 SUB 0.90fF $ **FLOATING
C2994 S.n2708 SUB 0.05fF $ **FLOATING
C2995 S.t537 SUB 0.02fF
C2996 S.n2709 SUB 0.12fF $ **FLOATING
C2997 S.n2710 SUB 0.14fF $ **FLOATING
C2998 S.n2712 SUB 0.77fF $ **FLOATING
C2999 S.n2713 SUB 1.92fF $ **FLOATING
C3000 S.n2714 SUB 1.86fF $ **FLOATING
C3001 S.n2715 SUB 0.12fF $ **FLOATING
C3002 S.t876 SUB 0.02fF
C3003 S.n2716 SUB 0.14fF $ **FLOATING
C3004 S.t562 SUB 0.02fF
C3005 S.n2718 SUB 0.24fF $ **FLOATING
C3006 S.n2719 SUB 0.35fF $ **FLOATING
C3007 S.n2720 SUB 0.60fF $ **FLOATING
C3008 S.n2721 SUB 1.82fF $ **FLOATING
C3009 S.n2722 SUB 2.96fF $ **FLOATING
C3010 S.t979 SUB 0.02fF
C3011 S.n2723 SUB 0.24fF $ **FLOATING
C3012 S.n2724 SUB 0.90fF $ **FLOATING
C3013 S.n2725 SUB 0.05fF $ **FLOATING
C3014 S.t148 SUB 0.02fF
C3015 S.n2726 SUB 0.12fF $ **FLOATING
C3016 S.n2727 SUB 0.14fF $ **FLOATING
C3017 S.n2729 SUB 1.87fF $ **FLOATING
C3018 S.n2730 SUB 1.73fF $ **FLOATING
C3019 S.t170 SUB 0.02fF
C3020 S.n2731 SUB 0.24fF $ **FLOATING
C3021 S.n2732 SUB 0.35fF $ **FLOATING
C3022 S.n2733 SUB 0.60fF $ **FLOATING
C3023 S.n2734 SUB 0.12fF $ **FLOATING
C3024 S.t499 SUB 0.02fF
C3025 S.n2735 SUB 0.14fF $ **FLOATING
C3026 S.n2737 SUB 1.14fF $ **FLOATING
C3027 S.n2738 SUB 0.22fF $ **FLOATING
C3028 S.n2739 SUB 0.25fF $ **FLOATING
C3029 S.n2740 SUB 0.09fF $ **FLOATING
C3030 S.n2741 SUB 2.41fF $ **FLOATING
C3031 S.t602 SUB 0.02fF
C3032 S.n2742 SUB 0.24fF $ **FLOATING
C3033 S.n2743 SUB 0.90fF $ **FLOATING
C3034 S.n2744 SUB 0.05fF $ **FLOATING
C3035 S.t788 SUB 0.02fF
C3036 S.n2745 SUB 0.12fF $ **FLOATING
C3037 S.n2746 SUB 0.14fF $ **FLOATING
C3038 S.n2748 SUB 1.86fF $ **FLOATING
C3039 S.n2749 SUB 0.47fF $ **FLOATING
C3040 S.n2750 SUB 0.09fF $ **FLOATING
C3041 S.n2751 SUB 0.32fF $ **FLOATING
C3042 S.n2752 SUB 0.30fF $ **FLOATING
C3043 S.n2753 SUB 0.76fF $ **FLOATING
C3044 S.n2754 SUB 0.58fF $ **FLOATING
C3045 S.t893 SUB 0.02fF
C3046 S.n2755 SUB 0.24fF $ **FLOATING
C3047 S.n2756 SUB 0.35fF $ **FLOATING
C3048 S.n2757 SUB 0.60fF $ **FLOATING
C3049 S.n2758 SUB 0.12fF $ **FLOATING
C3050 S.t110 SUB 0.02fF
C3051 S.n2759 SUB 0.14fF $ **FLOATING
C3052 S.n2761 SUB 2.58fF $ **FLOATING
C3053 S.n2762 SUB 2.13fF $ **FLOATING
C3054 S.t209 SUB 0.02fF
C3055 S.n2763 SUB 0.24fF $ **FLOATING
C3056 S.n2764 SUB 0.90fF $ **FLOATING
C3057 S.n2765 SUB 0.05fF $ **FLOATING
C3058 S.t406 SUB 0.02fF
C3059 S.n2766 SUB 0.12fF $ **FLOATING
C3060 S.n2767 SUB 0.14fF $ **FLOATING
C3061 S.n2769 SUB 0.77fF $ **FLOATING
C3062 S.n2770 SUB 2.27fF $ **FLOATING
C3063 S.n2771 SUB 1.86fF $ **FLOATING
C3064 S.n2772 SUB 0.12fF $ **FLOATING
C3065 S.t843 SUB 0.02fF
C3066 S.n2773 SUB 0.14fF $ **FLOATING
C3067 S.t521 SUB 0.02fF
C3068 S.n2775 SUB 0.24fF $ **FLOATING
C3069 S.n2776 SUB 0.35fF $ **FLOATING
C3070 S.n2777 SUB 0.60fF $ **FLOATING
C3071 S.n2778 SUB 1.37fF $ **FLOATING
C3072 S.n2779 SUB 0.70fF $ **FLOATING
C3073 S.n2780 SUB 1.13fF $ **FLOATING
C3074 S.n2781 SUB 0.35fF $ **FLOATING
C3075 S.n2782 SUB 2.00fF $ **FLOATING
C3076 S.t933 SUB 0.02fF
C3077 S.n2783 SUB 0.24fF $ **FLOATING
C3078 S.n2784 SUB 0.90fF $ **FLOATING
C3079 S.n2785 SUB 0.05fF $ **FLOATING
C3080 S.t1126 SUB 0.02fF
C3081 S.n2786 SUB 0.12fF $ **FLOATING
C3082 S.n2787 SUB 0.14fF $ **FLOATING
C3083 S.n2789 SUB 1.87fF $ **FLOATING
C3084 S.n2790 SUB 1.86fF $ **FLOATING
C3085 S.t130 SUB 0.02fF
C3086 S.n2791 SUB 0.24fF $ **FLOATING
C3087 S.n2792 SUB 0.35fF $ **FLOATING
C3088 S.n2793 SUB 0.60fF $ **FLOATING
C3089 S.n2794 SUB 0.12fF $ **FLOATING
C3090 S.t469 SUB 0.02fF
C3091 S.n2795 SUB 0.14fF $ **FLOATING
C3092 S.n2797 SUB 1.14fF $ **FLOATING
C3093 S.n2798 SUB 0.22fF $ **FLOATING
C3094 S.n2799 SUB 0.25fF $ **FLOATING
C3095 S.n2800 SUB 0.09fF $ **FLOATING
C3096 S.n2801 SUB 1.86fF $ **FLOATING
C3097 S.t551 SUB 0.02fF
C3098 S.n2802 SUB 0.24fF $ **FLOATING
C3099 S.n2803 SUB 0.90fF $ **FLOATING
C3100 S.n2804 SUB 0.05fF $ **FLOATING
C3101 S.t735 SUB 0.02fF
C3102 S.n2805 SUB 0.12fF $ **FLOATING
C3103 S.n2806 SUB 0.14fF $ **FLOATING
C3104 S.n2808 SUB 14.09fF $ **FLOATING
C3105 S.n2809 SUB 1.86fF $ **FLOATING
C3106 S.n2810 SUB 2.64fF $ **FLOATING
C3107 S.t90 SUB 0.02fF
C3108 S.n2811 SUB 0.24fF $ **FLOATING
C3109 S.n2812 SUB 0.35fF $ **FLOATING
C3110 S.n2813 SUB 0.60fF $ **FLOATING
C3111 S.n2814 SUB 0.12fF $ **FLOATING
C3112 S.t425 SUB 0.02fF
C3113 S.n2815 SUB 0.14fF $ **FLOATING
C3114 S.n2817 SUB 2.77fF $ **FLOATING
C3115 S.n2818 SUB 2.28fF $ **FLOATING
C3116 S.t763 SUB 0.02fF
C3117 S.n2819 SUB 0.12fF $ **FLOATING
C3118 S.n2820 SUB 0.14fF $ **FLOATING
C3119 S.t516 SUB 0.02fF
C3120 S.n2822 SUB 0.24fF $ **FLOATING
C3121 S.n2823 SUB 0.90fF $ **FLOATING
C3122 S.n2824 SUB 0.05fF $ **FLOATING
C3123 S.n2825 SUB 2.71fF $ **FLOATING
C3124 S.n2826 SUB 1.56fF $ **FLOATING
C3125 S.n2827 SUB 0.12fF $ **FLOATING
C3126 S.t272 SUB 0.02fF
C3127 S.n2828 SUB 0.14fF $ **FLOATING
C3128 S.t838 SUB 0.02fF
C3129 S.n2830 SUB 0.24fF $ **FLOATING
C3130 S.n2831 SUB 0.35fF $ **FLOATING
C3131 S.n2832 SUB 0.60fF $ **FLOATING
C3132 S.n2833 SUB 0.07fF $ **FLOATING
C3133 S.n2834 SUB 0.01fF $ **FLOATING
C3134 S.n2835 SUB 0.23fF $ **FLOATING
C3135 S.n2836 SUB 1.15fF $ **FLOATING
C3136 S.n2837 SUB 1.33fF $ **FLOATING
C3137 S.n2838 SUB 2.28fF $ **FLOATING
C3138 S.t598 SUB 0.02fF
C3139 S.n2839 SUB 0.12fF $ **FLOATING
C3140 S.n2840 SUB 0.14fF $ **FLOATING
C3141 S.t1000 SUB 0.02fF
C3142 S.n2842 SUB 0.24fF $ **FLOATING
C3143 S.n2843 SUB 0.90fF $ **FLOATING
C3144 S.n2844 SUB 0.05fF $ **FLOATING
C3145 S.t0 SUB 32.35fF
C3146 S.t124 SUB 0.02fF
C3147 S.n2845 SUB 0.24fF $ **FLOATING
C3148 S.n2846 SUB 0.90fF $ **FLOATING
C3149 S.n2847 SUB 0.05fF $ **FLOATING
C3150 S.t379 SUB 0.02fF
C3151 S.n2848 SUB 0.12fF $ **FLOATING
C3152 S.n2849 SUB 0.14fF $ **FLOATING
C3153 S.n2851 SUB 0.12fF $ **FLOATING
C3154 S.t1143 SUB 0.02fF
C3155 S.n2852 SUB 0.14fF $ **FLOATING
C3156 S.n2854 SUB 5.11fF $ **FLOATING
C3157 S.n2855 SUB 5.38fF $ **FLOATING
C3158 S.t706 SUB 0.02fF
C3159 S.n2856 SUB 0.12fF $ **FLOATING
C3160 S.n2857 SUB 0.14fF $ **FLOATING
C3161 S.t321 SUB 0.02fF
C3162 S.n2859 SUB 0.24fF $ **FLOATING
C3163 S.n2860 SUB 0.90fF $ **FLOATING
C3164 S.n2861 SUB 0.05fF $ **FLOATING
C3165 S.t66 SUB 31.97fF
C3166 S.t1072 SUB 0.02fF
C3167 S.n2862 SUB 0.01fF $ **FLOATING
C3168 S.n2863 SUB 0.25fF $ **FLOATING
C3169 S.t207 SUB 0.02fF
C3170 S.n2865 SUB 1.18fF $ **FLOATING
C3171 S.n2866 SUB 0.05fF $ **FLOATING
C3172 S.t261 SUB 0.02fF
C3173 S.n2867 SUB 0.63fF $ **FLOATING
C3174 S.n2868 SUB 0.60fF $ **FLOATING
C3175 S.n2869 SUB 8.87fF $ **FLOATING
C3176 S.n2870 SUB 0.76fF $ **FLOATING
C3177 S.n2871 SUB 0.27fF $ **FLOATING
C3178 S.n2872 SUB 0.59fF $ **FLOATING
C3179 S.n2873 SUB 0.21fF $ **FLOATING
C3180 S.n2874 SUB 0.59fF $ **FLOATING
C3181 S.n2875 SUB 2.57fF $ **FLOATING
C3182 S.n2876 SUB 0.29fF $ **FLOATING
C3183 S.t44 SUB 14.50fF
C3184 S.n2877 SUB 15.77fF $ **FLOATING
C3185 S.n2878 SUB 8.87fF $ **FLOATING
C3186 S.n2879 SUB 3.96fF $ **FLOATING
C3187 S.n2880 SUB 1.34fF $ **FLOATING
C3188 S.n2881 SUB 0.01fF $ **FLOATING
C3189 S.n2882 SUB 0.02fF $ **FLOATING
C3190 S.n2883 SUB 0.03fF $ **FLOATING
C3191 S.n2884 SUB 0.04fF $ **FLOATING
C3192 S.n2885 SUB 0.17fF $ **FLOATING
C3193 S.n2886 SUB 0.01fF $ **FLOATING
C3194 S.n2887 SUB 0.02fF $ **FLOATING
C3195 S.n2888 SUB 0.01fF $ **FLOATING
C3196 S.n2889 SUB 0.01fF $ **FLOATING
C3197 S.n2890 SUB 0.01fF $ **FLOATING
C3198 S.n2891 SUB 0.01fF $ **FLOATING
C3199 S.n2892 SUB 0.01fF $ **FLOATING
C3200 S.n2893 SUB 0.01fF $ **FLOATING
C3201 S.n2894 SUB 0.02fF $ **FLOATING
C3202 S.n2895 SUB 0.05fF $ **FLOATING
C3203 S.n2896 SUB 0.04fF $ **FLOATING
C3204 S.n2897 SUB 0.11fF $ **FLOATING
C3205 S.n2898 SUB 0.37fF $ **FLOATING
C3206 S.n2899 SUB 0.20fF $ **FLOATING
C3207 S.n2900 SUB 4.37fF $ **FLOATING
C3208 S.n2901 SUB 0.01fF $ **FLOATING
C3209 S.n2902 SUB 0.02fF $ **FLOATING
C3210 S.n2903 SUB 0.03fF $ **FLOATING
C3211 S.n2904 SUB 0.04fF $ **FLOATING
C3212 S.n2905 SUB 0.17fF $ **FLOATING
C3213 S.n2906 SUB 0.01fF $ **FLOATING
C3214 S.n2907 SUB 0.02fF $ **FLOATING
C3215 S.n2908 SUB 0.01fF $ **FLOATING
C3216 S.n2909 SUB 0.01fF $ **FLOATING
C3217 S.n2910 SUB 0.01fF $ **FLOATING
C3218 S.n2911 SUB 0.01fF $ **FLOATING
C3219 S.n2912 SUB 0.01fF $ **FLOATING
C3220 S.n2913 SUB 0.01fF $ **FLOATING
C3221 S.n2914 SUB 0.02fF $ **FLOATING
C3222 S.n2915 SUB 0.05fF $ **FLOATING
C3223 S.n2916 SUB 0.04fF $ **FLOATING
C3224 S.n2917 SUB 0.11fF $ **FLOATING
C3225 S.n2918 SUB 0.37fF $ **FLOATING
C3226 S.n2919 SUB 0.20fF $ **FLOATING
C3227 S.n2920 SUB 8.87fF $ **FLOATING
C3228 S.n2921 SUB 8.87fF $ **FLOATING
C3229 S.n2922 SUB 0.59fF $ **FLOATING
C3230 S.n2923 SUB 0.21fF $ **FLOATING
C3231 S.n2924 SUB 0.59fF $ **FLOATING
C3232 S.n2925 SUB 2.57fF $ **FLOATING
C3233 S.n2926 SUB 0.29fF $ **FLOATING
C3234 S.t136 SUB 14.50fF
C3235 S.n2927 SUB 15.77fF $ **FLOATING
C3236 S.n2928 SUB 0.76fF $ **FLOATING
C3237 S.n2929 SUB 0.27fF $ **FLOATING
C3238 S.n2930 SUB 3.96fF $ **FLOATING
C3239 S.n2931 SUB 1.34fF $ **FLOATING
C3240 S.t993 SUB 0.02fF
C3241 S.n2932 SUB 0.63fF $ **FLOATING
C3242 S.n2933 SUB 0.60fF $ **FLOATING
C3243 S.n2934 SUB 0.25fF $ **FLOATING
C3244 S.n2935 SUB 0.09fF $ **FLOATING
C3245 S.n2936 SUB 0.21fF $ **FLOATING
C3246 S.n2937 SUB 0.91fF $ **FLOATING
C3247 S.n2938 SUB 0.44fF $ **FLOATING
C3248 S.n2939 SUB 1.86fF $ **FLOATING
C3249 S.n2940 SUB 0.12fF $ **FLOATING
C3250 S.t523 SUB 0.02fF
C3251 S.n2941 SUB 0.14fF $ **FLOATING
C3252 S.t728 SUB 0.02fF
C3253 S.n2943 SUB 0.24fF $ **FLOATING
C3254 S.n2944 SUB 0.35fF $ **FLOATING
C3255 S.n2945 SUB 0.60fF $ **FLOATING
C3256 S.n2946 SUB 0.02fF $ **FLOATING
C3257 S.n2947 SUB 0.01fF $ **FLOATING
C3258 S.n2948 SUB 0.02fF $ **FLOATING
C3259 S.n2949 SUB 0.08fF $ **FLOATING
C3260 S.n2950 SUB 0.06fF $ **FLOATING
C3261 S.n2951 SUB 0.03fF $ **FLOATING
C3262 S.n2952 SUB 0.03fF $ **FLOATING
C3263 S.n2953 SUB 0.99fF $ **FLOATING
C3264 S.n2954 SUB 0.35fF $ **FLOATING
C3265 S.n2955 SUB 1.85fF $ **FLOATING
C3266 S.n2956 SUB 1.97fF $ **FLOATING
C3267 S.t1099 SUB 0.02fF
C3268 S.n2957 SUB 0.24fF $ **FLOATING
C3269 S.n2958 SUB 0.90fF $ **FLOATING
C3270 S.n2959 SUB 0.05fF $ **FLOATING
C3271 S.t626 SUB 0.02fF
C3272 S.n2960 SUB 0.12fF $ **FLOATING
C3273 S.n2961 SUB 0.14fF $ **FLOATING
C3274 S.n2963 SUB 1.87fF $ **FLOATING
C3275 S.n2964 SUB 0.07fF $ **FLOATING
C3276 S.n2965 SUB 0.04fF $ **FLOATING
C3277 S.n2966 SUB 0.05fF $ **FLOATING
C3278 S.n2967 SUB 0.86fF $ **FLOATING
C3279 S.n2968 SUB 0.01fF $ **FLOATING
C3280 S.n2969 SUB 0.01fF $ **FLOATING
C3281 S.n2970 SUB 0.01fF $ **FLOATING
C3282 S.n2971 SUB 0.07fF $ **FLOATING
C3283 S.n2972 SUB 0.68fF $ **FLOATING
C3284 S.n2973 SUB 0.71fF $ **FLOATING
C3285 S.t264 SUB 0.02fF
C3286 S.n2974 SUB 0.24fF $ **FLOATING
C3287 S.n2975 SUB 0.35fF $ **FLOATING
C3288 S.n2976 SUB 0.60fF $ **FLOATING
C3289 S.n2977 SUB 0.12fF $ **FLOATING
C3290 S.t1090 SUB 0.02fF
C3291 S.n2978 SUB 0.14fF $ **FLOATING
C3292 S.n2980 SUB 0.69fF $ **FLOATING
C3293 S.n2981 SUB 0.22fF $ **FLOATING
C3294 S.n2982 SUB 0.22fF $ **FLOATING
C3295 S.n2983 SUB 0.69fF $ **FLOATING
C3296 S.n2984 SUB 1.14fF $ **FLOATING
C3297 S.n2985 SUB 0.22fF $ **FLOATING
C3298 S.n2986 SUB 0.25fF $ **FLOATING
C3299 S.n2987 SUB 0.09fF $ **FLOATING
C3300 S.n2988 SUB 2.29fF $ **FLOATING
C3301 S.t208 SUB 0.02fF
C3302 S.n2989 SUB 0.24fF $ **FLOATING
C3303 S.n2990 SUB 0.90fF $ **FLOATING
C3304 S.n2991 SUB 0.05fF $ **FLOATING
C3305 S.t79 SUB 0.02fF
C3306 S.n2992 SUB 0.12fF $ **FLOATING
C3307 S.n2993 SUB 0.14fF $ **FLOATING
C3308 S.n2995 SUB 1.86fF $ **FLOATING
C3309 S.n2996 SUB 0.45fF $ **FLOATING
C3310 S.n2997 SUB 0.22fF $ **FLOATING
C3311 S.n2998 SUB 0.38fF $ **FLOATING
C3312 S.n2999 SUB 0.16fF $ **FLOATING
C3313 S.n3000 SUB 0.28fF $ **FLOATING
C3314 S.n3001 SUB 0.21fF $ **FLOATING
C3315 S.n3002 SUB 0.30fF $ **FLOATING
C3316 S.n3003 SUB 0.41fF $ **FLOATING
C3317 S.n3004 SUB 0.20fF $ **FLOATING
C3318 S.t986 SUB 0.02fF
C3319 S.n3005 SUB 0.24fF $ **FLOATING
C3320 S.n3006 SUB 0.35fF $ **FLOATING
C3321 S.n3007 SUB 0.60fF $ **FLOATING
C3322 S.n3008 SUB 0.12fF $ **FLOATING
C3323 S.t704 SUB 0.02fF
C3324 S.n3009 SUB 0.14fF $ **FLOATING
C3325 S.n3011 SUB 0.04fF $ **FLOATING
C3326 S.n3012 SUB 0.03fF $ **FLOATING
C3327 S.n3013 SUB 0.03fF $ **FLOATING
C3328 S.n3014 SUB 0.10fF $ **FLOATING
C3329 S.n3015 SUB 0.36fF $ **FLOATING
C3330 S.n3016 SUB 0.37fF $ **FLOATING
C3331 S.n3017 SUB 0.10fF $ **FLOATING
C3332 S.n3018 SUB 0.12fF $ **FLOATING
C3333 S.n3019 SUB 0.07fF $ **FLOATING
C3334 S.n3020 SUB 0.12fF $ **FLOATING
C3335 S.n3021 SUB 0.18fF $ **FLOATING
C3336 S.n3022 SUB 3.95fF $ **FLOATING
C3337 S.t930 SUB 0.02fF
C3338 S.n3023 SUB 0.24fF $ **FLOATING
C3339 S.n3024 SUB 0.90fF $ **FLOATING
C3340 S.n3025 SUB 0.05fF $ **FLOATING
C3341 S.t817 SUB 0.02fF
C3342 S.n3026 SUB 0.12fF $ **FLOATING
C3343 S.n3027 SUB 0.14fF $ **FLOATING
C3344 S.n3029 SUB 0.25fF $ **FLOATING
C3345 S.n3030 SUB 0.09fF $ **FLOATING
C3346 S.n3031 SUB 0.21fF $ **FLOATING
C3347 S.n3032 SUB 1.27fF $ **FLOATING
C3348 S.n3033 SUB 0.52fF $ **FLOATING
C3349 S.n3034 SUB 1.86fF $ **FLOATING
C3350 S.n3035 SUB 0.12fF $ **FLOATING
C3351 S.t326 SUB 0.02fF
C3352 S.n3036 SUB 0.14fF $ **FLOATING
C3353 S.t609 SUB 0.02fF
C3354 S.n3038 SUB 0.24fF $ **FLOATING
C3355 S.n3039 SUB 0.35fF $ **FLOATING
C3356 S.n3040 SUB 0.60fF $ **FLOATING
C3357 S.n3041 SUB 1.56fF $ **FLOATING
C3358 S.n3042 SUB 2.42fF $ **FLOATING
C3359 S.t552 SUB 0.02fF
C3360 S.n3043 SUB 0.24fF $ **FLOATING
C3361 S.n3044 SUB 0.90fF $ **FLOATING
C3362 S.n3045 SUB 0.05fF $ **FLOATING
C3363 S.t441 SUB 0.02fF
C3364 S.n3046 SUB 0.12fF $ **FLOATING
C3365 S.n3047 SUB 0.14fF $ **FLOATING
C3366 S.n3049 SUB 1.87fF $ **FLOATING
C3367 S.n3050 SUB 0.06fF $ **FLOATING
C3368 S.n3051 SUB 0.03fF $ **FLOATING
C3369 S.n3052 SUB 0.03fF $ **FLOATING
C3370 S.n3053 SUB 0.98fF $ **FLOATING
C3371 S.n3054 SUB 0.02fF $ **FLOATING
C3372 S.n3055 SUB 0.01fF $ **FLOATING
C3373 S.n3056 SUB 0.02fF $ **FLOATING
C3374 S.n3057 SUB 0.08fF $ **FLOATING
C3375 S.n3058 SUB 0.36fF $ **FLOATING
C3376 S.n3059 SUB 1.83fF $ **FLOATING
C3377 S.t217 SUB 0.02fF
C3378 S.n3060 SUB 0.24fF $ **FLOATING
C3379 S.n3061 SUB 0.35fF $ **FLOATING
C3380 S.n3062 SUB 0.60fF $ **FLOATING
C3381 S.n3063 SUB 0.12fF $ **FLOATING
C3382 S.t1052 SUB 0.02fF
C3383 S.n3064 SUB 0.14fF $ **FLOATING
C3384 S.n3066 SUB 0.69fF $ **FLOATING
C3385 S.n3067 SUB 0.22fF $ **FLOATING
C3386 S.n3068 SUB 0.22fF $ **FLOATING
C3387 S.n3069 SUB 0.69fF $ **FLOATING
C3388 S.n3070 SUB 1.14fF $ **FLOATING
C3389 S.n3071 SUB 0.22fF $ **FLOATING
C3390 S.n3072 SUB 0.25fF $ **FLOATING
C3391 S.n3073 SUB 0.09fF $ **FLOATING
C3392 S.n3074 SUB 1.86fF $ **FLOATING
C3393 S.t162 SUB 0.02fF
C3394 S.n3075 SUB 0.24fF $ **FLOATING
C3395 S.n3076 SUB 0.90fF $ **FLOATING
C3396 S.n3077 SUB 0.05fF $ **FLOATING
C3397 S.t15 SUB 0.02fF
C3398 S.n3078 SUB 0.12fF $ **FLOATING
C3399 S.n3079 SUB 0.14fF $ **FLOATING
C3400 S.n3081 SUB 14.09fF $ **FLOATING
C3401 S.n3082 SUB 1.70fF $ **FLOATING
C3402 S.n3083 SUB 3.01fF $ **FLOATING
C3403 S.t1119 SUB 0.02fF
C3404 S.n3084 SUB 0.24fF $ **FLOATING
C3405 S.n3085 SUB 0.35fF $ **FLOATING
C3406 S.n3086 SUB 0.60fF $ **FLOATING
C3407 S.n3087 SUB 0.12fF $ **FLOATING
C3408 S.t896 SUB 0.02fF
C3409 S.n3088 SUB 0.14fF $ **FLOATING
C3410 S.n3090 SUB 0.31fF $ **FLOATING
C3411 S.n3091 SUB 0.22fF $ **FLOATING
C3412 S.n3092 SUB 0.65fF $ **FLOATING
C3413 S.n3093 SUB 0.94fF $ **FLOATING
C3414 S.n3094 SUB 0.22fF $ **FLOATING
C3415 S.n3095 SUB 0.20fF $ **FLOATING
C3416 S.n3096 SUB 0.20fF $ **FLOATING
C3417 S.n3097 SUB 0.06fF $ **FLOATING
C3418 S.n3098 SUB 0.09fF $ **FLOATING
C3419 S.n3099 SUB 0.09fF $ **FLOATING
C3420 S.n3100 SUB 1.97fF $ **FLOATING
C3421 S.t937 SUB 0.02fF
C3422 S.n3101 SUB 0.12fF $ **FLOATING
C3423 S.n3102 SUB 0.14fF $ **FLOATING
C3424 S.t378 SUB 0.02fF
C3425 S.n3104 SUB 0.24fF $ **FLOATING
C3426 S.n3105 SUB 0.90fF $ **FLOATING
C3427 S.n3106 SUB 0.05fF $ **FLOATING
C3428 S.n3107 SUB 1.86fF $ **FLOATING
C3429 S.n3108 SUB 0.12fF $ **FLOATING
C3430 S.t80 SUB 0.02fF
C3431 S.n3109 SUB 0.14fF $ **FLOATING
C3432 S.t366 SUB 0.02fF
C3433 S.n3111 SUB 0.12fF $ **FLOATING
C3434 S.n3112 SUB 0.14fF $ **FLOATING
C3435 S.t174 SUB 0.02fF
C3436 S.n3114 SUB 0.24fF $ **FLOATING
C3437 S.n3115 SUB 0.90fF $ **FLOATING
C3438 S.n3116 SUB 0.05fF $ **FLOATING
C3439 S.t872 SUB 0.02fF
C3440 S.n3117 SUB 0.24fF $ **FLOATING
C3441 S.n3118 SUB 0.35fF $ **FLOATING
C3442 S.n3119 SUB 0.60fF $ **FLOATING
C3443 S.n3120 SUB 0.31fF $ **FLOATING
C3444 S.n3121 SUB 1.08fF $ **FLOATING
C3445 S.n3122 SUB 0.15fF $ **FLOATING
C3446 S.n3123 SUB 2.08fF $ **FLOATING
C3447 S.n3124 SUB 2.91fF $ **FLOATING
C3448 S.n3125 SUB 1.86fF $ **FLOATING
C3449 S.n3126 SUB 0.12fF $ **FLOATING
C3450 S.t726 SUB 0.02fF
C3451 S.n3127 SUB 0.14fF $ **FLOATING
C3452 S.t1005 SUB 0.02fF
C3453 S.n3129 SUB 0.24fF $ **FLOATING
C3454 S.n3130 SUB 0.35fF $ **FLOATING
C3455 S.n3131 SUB 0.60fF $ **FLOATING
C3456 S.n3132 SUB 0.91fF $ **FLOATING
C3457 S.n3133 SUB 0.31fF $ **FLOATING
C3458 S.n3134 SUB 0.91fF $ **FLOATING
C3459 S.n3135 SUB 1.08fF $ **FLOATING
C3460 S.n3136 SUB 0.15fF $ **FLOATING
C3461 S.n3137 SUB 4.90fF $ **FLOATING
C3462 S.t770 SUB 0.02fF
C3463 S.n3138 SUB 0.12fF $ **FLOATING
C3464 S.n3139 SUB 0.14fF $ **FLOATING
C3465 S.t962 SUB 0.02fF
C3466 S.n3141 SUB 0.24fF $ **FLOATING
C3467 S.n3142 SUB 0.90fF $ **FLOATING
C3468 S.n3143 SUB 0.05fF $ **FLOATING
C3469 S.n3144 SUB 1.86fF $ **FLOATING
C3470 S.n3145 SUB 2.64fF $ **FLOATING
C3471 S.t627 SUB 0.02fF
C3472 S.n3146 SUB 0.24fF $ **FLOATING
C3473 S.n3147 SUB 0.35fF $ **FLOATING
C3474 S.n3148 SUB 0.60fF $ **FLOATING
C3475 S.n3149 SUB 0.12fF $ **FLOATING
C3476 S.t345 SUB 0.02fF
C3477 S.n3150 SUB 0.14fF $ **FLOATING
C3478 S.n3152 SUB 1.86fF $ **FLOATING
C3479 S.n3153 SUB 2.64fF $ **FLOATING
C3480 S.t495 SUB 0.02fF
C3481 S.n3154 SUB 0.24fF $ **FLOATING
C3482 S.n3155 SUB 0.35fF $ **FLOATING
C3483 S.n3156 SUB 0.60fF $ **FLOATING
C3484 S.t898 SUB 0.02fF
C3485 S.n3157 SUB 0.24fF $ **FLOATING
C3486 S.n3158 SUB 0.90fF $ **FLOATING
C3487 S.n3159 SUB 0.05fF $ **FLOATING
C3488 S.t32 SUB 0.02fF
C3489 S.n3160 SUB 0.12fF $ **FLOATING
C3490 S.n3161 SUB 0.14fF $ **FLOATING
C3491 S.n3163 SUB 0.12fF $ **FLOATING
C3492 S.t816 SUB 0.02fF
C3493 S.n3164 SUB 0.14fF $ **FLOATING
C3494 S.n3166 SUB 2.28fF $ **FLOATING
C3495 S.n3167 SUB 2.91fF $ **FLOATING
C3496 S.n3168 SUB 5.10fF $ **FLOATING
C3497 S.t386 SUB 0.02fF
C3498 S.n3169 SUB 0.12fF $ **FLOATING
C3499 S.n3170 SUB 0.14fF $ **FLOATING
C3500 S.t582 SUB 0.02fF
C3501 S.n3172 SUB 0.24fF $ **FLOATING
C3502 S.n3173 SUB 0.90fF $ **FLOATING
C3503 S.n3174 SUB 0.05fF $ **FLOATING
C3504 S.n3175 SUB 1.86fF $ **FLOATING
C3505 S.n3176 SUB 2.64fF $ **FLOATING
C3506 S.t238 SUB 0.02fF
C3507 S.n3177 SUB 0.24fF $ **FLOATING
C3508 S.n3178 SUB 0.35fF $ **FLOATING
C3509 S.n3179 SUB 0.60fF $ **FLOATING
C3510 S.n3180 SUB 0.12fF $ **FLOATING
C3511 S.t1070 SUB 0.02fF
C3512 S.n3181 SUB 0.14fF $ **FLOATING
C3513 S.n3183 SUB 5.11fF $ **FLOATING
C3514 S.t1108 SUB 0.02fF
C3515 S.n3184 SUB 0.12fF $ **FLOATING
C3516 S.n3185 SUB 0.14fF $ **FLOATING
C3517 S.t185 SUB 0.02fF
C3518 S.n3187 SUB 0.24fF $ **FLOATING
C3519 S.n3188 SUB 0.90fF $ **FLOATING
C3520 S.n3189 SUB 0.05fF $ **FLOATING
C3521 S.n3190 SUB 1.86fF $ **FLOATING
C3522 S.n3191 SUB 2.64fF $ **FLOATING
C3523 S.t967 SUB 0.02fF
C3524 S.n3192 SUB 0.24fF $ **FLOATING
C3525 S.n3193 SUB 0.35fF $ **FLOATING
C3526 S.n3194 SUB 0.60fF $ **FLOATING
C3527 S.n3195 SUB 0.12fF $ **FLOATING
C3528 S.t687 SUB 0.02fF
C3529 S.n3196 SUB 0.14fF $ **FLOATING
C3530 S.n3198 SUB 4.84fF $ **FLOATING
C3531 S.t717 SUB 0.02fF
C3532 S.n3199 SUB 0.12fF $ **FLOATING
C3533 S.n3200 SUB 0.14fF $ **FLOATING
C3534 S.t908 SUB 0.02fF
C3535 S.n3202 SUB 0.24fF $ **FLOATING
C3536 S.n3203 SUB 0.90fF $ **FLOATING
C3537 S.n3204 SUB 0.05fF $ **FLOATING
C3538 S.n3205 SUB 1.86fF $ **FLOATING
C3539 S.n3206 SUB 0.12fF $ **FLOATING
C3540 S.t769 SUB 0.02fF
C3541 S.n3207 SUB 0.14fF $ **FLOATING
C3542 S.t575 SUB 0.02fF
C3543 S.n3209 SUB 1.20fF $ **FLOATING
C3544 S.n3210 SUB 0.60fF $ **FLOATING
C3545 S.n3211 SUB 0.35fF $ **FLOATING
C3546 S.n3212 SUB 0.62fF $ **FLOATING
C3547 S.n3213 SUB 1.14fF $ **FLOATING
C3548 S.n3214 SUB 2.18fF $ **FLOATING
C3549 S.n3215 SUB 0.59fF $ **FLOATING
C3550 S.n3216 SUB 0.02fF $ **FLOATING
C3551 S.n3217 SUB 0.96fF $ **FLOATING
C3552 S.t103 SUB 14.50fF
C3553 S.n3218 SUB 14.37fF $ **FLOATING
C3554 S.n3220 SUB 0.37fF $ **FLOATING
C3555 S.n3221 SUB 0.23fF $ **FLOATING
C3556 S.n3222 SUB 2.87fF $ **FLOATING
C3557 S.n3223 SUB 2.43fF $ **FLOATING
C3558 S.n3224 SUB 1.94fF $ **FLOATING
C3559 S.n3225 SUB 3.89fF $ **FLOATING
C3560 S.n3226 SUB 0.25fF $ **FLOATING
C3561 S.n3227 SUB 0.01fF $ **FLOATING
C3562 S.t448 SUB 0.02fF
C3563 S.n3228 SUB 0.25fF $ **FLOATING
C3564 S.t310 SUB 0.02fF
C3565 S.n3229 SUB 0.94fF $ **FLOATING
C3566 S.n3230 SUB 0.70fF $ **FLOATING
C3567 S.n3231 SUB 0.77fF $ **FLOATING
C3568 S.n3232 SUB 1.91fF $ **FLOATING
C3569 S.n3233 SUB 1.86fF $ **FLOATING
C3570 S.n3234 SUB 0.12fF $ **FLOATING
C3571 S.t105 SUB 0.02fF
C3572 S.n3235 SUB 0.14fF $ **FLOATING
C3573 S.t181 SUB 0.02fF
C3574 S.n3237 SUB 0.24fF $ **FLOATING
C3575 S.n3238 SUB 0.35fF $ **FLOATING
C3576 S.n3239 SUB 0.60fF $ **FLOATING
C3577 S.n3240 SUB 1.50fF $ **FLOATING
C3578 S.n3241 SUB 2.96fF $ **FLOATING
C3579 S.t1040 SUB 0.02fF
C3580 S.n3242 SUB 0.24fF $ **FLOATING
C3581 S.n3243 SUB 0.90fF $ **FLOATING
C3582 S.n3244 SUB 0.05fF $ **FLOATING
C3583 S.t400 SUB 0.02fF
C3584 S.n3245 SUB 0.12fF $ **FLOATING
C3585 S.n3246 SUB 0.14fF $ **FLOATING
C3586 S.n3248 SUB 1.87fF $ **FLOATING
C3587 S.n3249 SUB 1.73fF $ **FLOATING
C3588 S.t184 SUB 0.02fF
C3589 S.n3250 SUB 0.24fF $ **FLOATING
C3590 S.n3251 SUB 0.35fF $ **FLOATING
C3591 S.n3252 SUB 0.60fF $ **FLOATING
C3592 S.n3253 SUB 0.12fF $ **FLOATING
C3593 S.t512 SUB 0.02fF
C3594 S.n3254 SUB 0.14fF $ **FLOATING
C3595 S.n3256 SUB 1.14fF $ **FLOATING
C3596 S.n3257 SUB 0.22fF $ **FLOATING
C3597 S.n3258 SUB 0.25fF $ **FLOATING
C3598 S.n3259 SUB 0.09fF $ **FLOATING
C3599 S.n3260 SUB 2.41fF $ **FLOATING
C3600 S.t615 SUB 0.02fF
C3601 S.n3261 SUB 0.24fF $ **FLOATING
C3602 S.n3262 SUB 0.90fF $ **FLOATING
C3603 S.n3263 SUB 0.05fF $ **FLOATING
C3604 S.t1121 SUB 0.02fF
C3605 S.n3264 SUB 0.12fF $ **FLOATING
C3606 S.n3265 SUB 0.14fF $ **FLOATING
C3607 S.n3267 SUB 1.86fF $ **FLOATING
C3608 S.n3268 SUB 0.47fF $ **FLOATING
C3609 S.n3269 SUB 0.09fF $ **FLOATING
C3610 S.n3270 SUB 0.32fF $ **FLOATING
C3611 S.n3271 SUB 0.30fF $ **FLOATING
C3612 S.n3272 SUB 0.76fF $ **FLOATING
C3613 S.n3273 SUB 0.58fF $ **FLOATING
C3614 S.t906 SUB 0.02fF
C3615 S.n3274 SUB 0.24fF $ **FLOATING
C3616 S.n3275 SUB 0.35fF $ **FLOATING
C3617 S.n3276 SUB 0.60fF $ **FLOATING
C3618 S.n3277 SUB 0.12fF $ **FLOATING
C3619 S.t121 SUB 0.02fF
C3620 S.n3278 SUB 0.14fF $ **FLOATING
C3621 S.n3280 SUB 2.58fF $ **FLOATING
C3622 S.n3281 SUB 2.13fF $ **FLOATING
C3623 S.t227 SUB 0.02fF
C3624 S.n3282 SUB 0.24fF $ **FLOATING
C3625 S.n3283 SUB 0.90fF $ **FLOATING
C3626 S.n3284 SUB 0.05fF $ **FLOATING
C3627 S.t424 SUB 0.02fF
C3628 S.n3285 SUB 0.12fF $ **FLOATING
C3629 S.n3286 SUB 0.14fF $ **FLOATING
C3630 S.n3288 SUB 0.77fF $ **FLOATING
C3631 S.n3289 SUB 2.27fF $ **FLOATING
C3632 S.n3290 SUB 1.86fF $ **FLOATING
C3633 S.n3291 SUB 0.12fF $ **FLOATING
C3634 S.t854 SUB 0.02fF
C3635 S.n3292 SUB 0.14fF $ **FLOATING
C3636 S.t530 SUB 0.02fF
C3637 S.n3294 SUB 0.24fF $ **FLOATING
C3638 S.n3295 SUB 0.35fF $ **FLOATING
C3639 S.n3296 SUB 0.60fF $ **FLOATING
C3640 S.n3297 SUB 1.37fF $ **FLOATING
C3641 S.n3298 SUB 0.70fF $ **FLOATING
C3642 S.n3299 SUB 1.13fF $ **FLOATING
C3643 S.n3300 SUB 0.35fF $ **FLOATING
C3644 S.n3301 SUB 2.00fF $ **FLOATING
C3645 S.t949 SUB 0.02fF
C3646 S.n3302 SUB 0.24fF $ **FLOATING
C3647 S.n3303 SUB 0.90fF $ **FLOATING
C3648 S.n3304 SUB 0.05fF $ **FLOATING
C3649 S.t1141 SUB 0.02fF
C3650 S.n3305 SUB 0.12fF $ **FLOATING
C3651 S.n3306 SUB 0.14fF $ **FLOATING
C3652 S.t570 SUB 0.02fF
C3653 S.n3308 SUB 0.24fF $ **FLOATING
C3654 S.n3309 SUB 0.90fF $ **FLOATING
C3655 S.n3310 SUB 0.05fF $ **FLOATING
C3656 S.n3311 SUB 1.87fF $ **FLOATING
C3657 S.n3312 SUB 1.86fF $ **FLOATING
C3658 S.t145 SUB 0.02fF
C3659 S.n3313 SUB 0.24fF $ **FLOATING
C3660 S.n3314 SUB 0.35fF $ **FLOATING
C3661 S.n3315 SUB 0.60fF $ **FLOATING
C3662 S.n3316 SUB 0.12fF $ **FLOATING
C3663 S.t478 SUB 0.02fF
C3664 S.n3317 SUB 0.14fF $ **FLOATING
C3665 S.n3319 SUB 1.14fF $ **FLOATING
C3666 S.n3320 SUB 0.22fF $ **FLOATING
C3667 S.n3321 SUB 0.25fF $ **FLOATING
C3668 S.n3322 SUB 0.09fF $ **FLOATING
C3669 S.n3323 SUB 1.86fF $ **FLOATING
C3670 S.t753 SUB 0.02fF
C3671 S.n3324 SUB 0.12fF $ **FLOATING
C3672 S.n3325 SUB 0.14fF $ **FLOATING
C3673 S.n3327 SUB 14.09fF $ **FLOATING
C3674 S.n3328 SUB 1.86fF $ **FLOATING
C3675 S.n3329 SUB 2.64fF $ **FLOATING
C3676 S.t104 SUB 0.02fF
C3677 S.n3330 SUB 0.24fF $ **FLOATING
C3678 S.n3331 SUB 0.35fF $ **FLOATING
C3679 S.n3332 SUB 0.60fF $ **FLOATING
C3680 S.n3333 SUB 0.12fF $ **FLOATING
C3681 S.t440 SUB 0.02fF
C3682 S.n3334 SUB 0.14fF $ **FLOATING
C3683 S.n3336 SUB 2.77fF $ **FLOATING
C3684 S.n3337 SUB 2.28fF $ **FLOATING
C3685 S.t780 SUB 0.02fF
C3686 S.n3338 SUB 0.12fF $ **FLOATING
C3687 S.n3339 SUB 0.14fF $ **FLOATING
C3688 S.t525 SUB 0.02fF
C3689 S.n3341 SUB 0.24fF $ **FLOATING
C3690 S.n3342 SUB 0.90fF $ **FLOATING
C3691 S.n3343 SUB 0.05fF $ **FLOATING
C3692 S.n3344 SUB 1.86fF $ **FLOATING
C3693 S.n3345 SUB 2.64fF $ **FLOATING
C3694 S.t836 SUB 0.02fF
C3695 S.n3346 SUB 0.24fF $ **FLOATING
C3696 S.n3347 SUB 0.35fF $ **FLOATING
C3697 S.n3348 SUB 0.60fF $ **FLOATING
C3698 S.n3349 SUB 0.12fF $ **FLOATING
C3699 S.t13 SUB 0.02fF
C3700 S.n3350 SUB 0.14fF $ **FLOATING
C3701 S.n3352 SUB 2.77fF $ **FLOATING
C3702 S.n3353 SUB 2.28fF $ **FLOATING
C3703 S.t396 SUB 0.02fF
C3704 S.n3354 SUB 0.12fF $ **FLOATING
C3705 S.n3355 SUB 0.14fF $ **FLOATING
C3706 S.t137 SUB 0.02fF
C3707 S.n3357 SUB 0.24fF $ **FLOATING
C3708 S.n3358 SUB 0.90fF $ **FLOATING
C3709 S.n3359 SUB 0.05fF $ **FLOATING
C3710 S.n3360 SUB 2.70fF $ **FLOATING
C3711 S.n3361 SUB 1.58fF $ **FLOATING
C3712 S.n3362 SUB 0.12fF $ **FLOATING
C3713 S.t734 SUB 0.02fF
C3714 S.n3363 SUB 0.14fF $ **FLOATING
C3715 S.t239 SUB 0.02fF
C3716 S.n3365 SUB 0.24fF $ **FLOATING
C3717 S.n3366 SUB 0.35fF $ **FLOATING
C3718 S.n3367 SUB 0.60fF $ **FLOATING
C3719 S.n3368 SUB 0.07fF $ **FLOATING
C3720 S.n3369 SUB 0.01fF $ **FLOATING
C3721 S.n3370 SUB 0.23fF $ **FLOATING
C3722 S.n3371 SUB 1.15fF $ **FLOATING
C3723 S.n3372 SUB 1.33fF $ **FLOATING
C3724 S.n3373 SUB 2.28fF $ **FLOATING
C3725 S.t1058 SUB 0.02fF
C3726 S.n3374 SUB 0.12fF $ **FLOATING
C3727 S.n3375 SUB 0.14fF $ **FLOATING
C3728 S.t342 SUB 0.02fF
C3729 S.n3377 SUB 0.24fF $ **FLOATING
C3730 S.n3378 SUB 0.90fF $ **FLOATING
C3731 S.n3379 SUB 0.05fF $ **FLOATING
C3732 S.t12 SUB 32.35fF
C3733 S.t1116 SUB 0.02fF
C3734 S.n3380 SUB 0.12fF $ **FLOATING
C3735 S.n3381 SUB 0.14fF $ **FLOATING
C3736 S.t865 SUB 0.02fF
C3737 S.n3383 SUB 0.24fF $ **FLOATING
C3738 S.n3384 SUB 0.90fF $ **FLOATING
C3739 S.n3385 SUB 0.05fF $ **FLOATING
C3740 S.t461 SUB 0.02fF
C3741 S.n3386 SUB 0.24fF $ **FLOATING
C3742 S.n3387 SUB 0.35fF $ **FLOATING
C3743 S.n3388 SUB 0.60fF $ **FLOATING
C3744 S.n3389 SUB 2.64fF $ **FLOATING
C3745 S.n3390 SUB 5.11fF $ **FLOATING
C3746 S.n3391 SUB 1.86fF $ **FLOATING
C3747 S.n3392 SUB 0.12fF $ **FLOATING
C3748 S.t826 SUB 0.02fF
C3749 S.n3393 SUB 0.14fF $ **FLOATING
C3750 S.t289 SUB 0.02fF
C3751 S.n3395 SUB 0.24fF $ **FLOATING
C3752 S.n3396 SUB 0.35fF $ **FLOATING
C3753 S.n3397 SUB 0.60fF $ **FLOATING
C3754 S.n3398 SUB 2.64fF $ **FLOATING
C3755 S.n3399 SUB 5.38fF $ **FLOATING
C3756 S.t337 SUB 0.02fF
C3757 S.n3400 SUB 0.12fF $ **FLOATING
C3758 S.n3401 SUB 0.14fF $ **FLOATING
C3759 S.t851 SUB 0.02fF
C3760 S.n3403 SUB 0.24fF $ **FLOATING
C3761 S.n3404 SUB 0.90fF $ **FLOATING
C3762 S.n3405 SUB 0.05fF $ **FLOATING
C3763 S.t14 SUB 31.97fF
C3764 S.t944 SUB 0.02fF
C3765 S.n3406 SUB 1.18fF $ **FLOATING
C3766 S.n3407 SUB 0.05fF $ **FLOATING
C3767 S.t500 SUB 0.02fF
C3768 S.n3408 SUB 0.01fF $ **FLOATING
C3769 S.n3409 SUB 0.25fF $ **FLOATING
C3770 S.n3411 SUB 1.48fF $ **FLOATING
C3771 S.n3412 SUB 1.29fF $ **FLOATING
C3772 S.n3413 SUB 0.27fF $ **FLOATING
C3773 S.n3414 SUB 0.24fF $ **FLOATING
C3774 S.n3415 SUB 4.34fF $ **FLOATING
C3775 S.n3416 SUB 0.01fF $ **FLOATING
C3776 S.n3417 SUB 0.02fF $ **FLOATING
C3777 S.n3418 SUB 0.03fF $ **FLOATING
C3778 S.n3419 SUB 0.04fF $ **FLOATING
C3779 S.n3420 SUB 0.17fF $ **FLOATING
C3780 S.n3421 SUB 0.01fF $ **FLOATING
C3781 S.n3422 SUB 0.02fF $ **FLOATING
C3782 S.n3423 SUB 0.01fF $ **FLOATING
C3783 S.n3424 SUB 0.01fF $ **FLOATING
C3784 S.n3425 SUB 0.01fF $ **FLOATING
C3785 S.n3426 SUB 0.01fF $ **FLOATING
C3786 S.n3427 SUB 0.01fF $ **FLOATING
C3787 S.n3428 SUB 0.01fF $ **FLOATING
C3788 S.n3429 SUB 0.02fF $ **FLOATING
C3789 S.n3430 SUB 0.05fF $ **FLOATING
C3790 S.n3431 SUB 0.04fF $ **FLOATING
C3791 S.n3432 SUB 0.11fF $ **FLOATING
C3792 S.n3433 SUB 0.37fF $ **FLOATING
C3793 S.n3434 SUB 0.20fF $ **FLOATING
C3794 S.n3435 SUB 8.87fF $ **FLOATING
C3795 S.n3436 SUB 8.87fF $ **FLOATING
C3796 S.n3437 SUB 0.59fF $ **FLOATING
C3797 S.n3438 SUB 0.21fF $ **FLOATING
C3798 S.n3439 SUB 0.59fF $ **FLOATING
C3799 S.n3440 SUB 2.57fF $ **FLOATING
C3800 S.n3441 SUB 0.29fF $ **FLOATING
C3801 S.t52 SUB 14.50fF
C3802 S.n3442 SUB 15.77fF $ **FLOATING
C3803 S.n3443 SUB 0.76fF $ **FLOATING
C3804 S.n3444 SUB 0.27fF $ **FLOATING
C3805 S.n3445 SUB 3.96fF $ **FLOATING
C3806 S.n3446 SUB 1.34fF $ **FLOATING
C3807 S.t1002 SUB 0.02fF
C3808 S.n3447 SUB 0.63fF $ **FLOATING
C3809 S.n3448 SUB 0.60fF $ **FLOATING
C3810 S.n3449 SUB 1.87fF $ **FLOATING
C3811 S.n3450 SUB 0.04fF $ **FLOATING
C3812 S.n3451 SUB 0.07fF $ **FLOATING
C3813 S.n3452 SUB 0.05fF $ **FLOATING
C3814 S.n3453 SUB 0.86fF $ **FLOATING
C3815 S.n3454 SUB 0.01fF $ **FLOATING
C3816 S.n3455 SUB 0.01fF $ **FLOATING
C3817 S.n3456 SUB 0.01fF $ **FLOATING
C3818 S.n3457 SUB 0.07fF $ **FLOATING
C3819 S.n3458 SUB 0.68fF $ **FLOATING
C3820 S.n3459 SUB 0.71fF $ **FLOATING
C3821 S.t505 SUB 0.02fF
C3822 S.n3460 SUB 0.24fF $ **FLOATING
C3823 S.n3461 SUB 0.35fF $ **FLOATING
C3824 S.n3462 SUB 0.60fF $ **FLOATING
C3825 S.n3463 SUB 0.12fF $ **FLOATING
C3826 S.t377 SUB 0.02fF
C3827 S.n3464 SUB 0.14fF $ **FLOATING
C3828 S.n3466 SUB 0.69fF $ **FLOATING
C3829 S.n3467 SUB 0.22fF $ **FLOATING
C3830 S.n3468 SUB 0.22fF $ **FLOATING
C3831 S.n3469 SUB 0.69fF $ **FLOATING
C3832 S.n3470 SUB 1.14fF $ **FLOATING
C3833 S.n3471 SUB 0.22fF $ **FLOATING
C3834 S.n3472 SUB 0.25fF $ **FLOATING
C3835 S.n3473 SUB 0.09fF $ **FLOATING
C3836 S.n3474 SUB 2.29fF $ **FLOATING
C3837 S.t1009 SUB 0.02fF
C3838 S.n3475 SUB 0.24fF $ **FLOATING
C3839 S.n3476 SUB 0.90fF $ **FLOATING
C3840 S.n3477 SUB 0.05fF $ **FLOATING
C3841 S.t481 SUB 0.02fF
C3842 S.n3478 SUB 0.12fF $ **FLOATING
C3843 S.n3479 SUB 0.14fF $ **FLOATING
C3844 S.n3481 SUB 1.86fF $ **FLOATING
C3845 S.n3482 SUB 0.45fF $ **FLOATING
C3846 S.n3483 SUB 0.22fF $ **FLOATING
C3847 S.n3484 SUB 0.38fF $ **FLOATING
C3848 S.n3485 SUB 0.16fF $ **FLOATING
C3849 S.n3486 SUB 0.28fF $ **FLOATING
C3850 S.n3487 SUB 0.21fF $ **FLOATING
C3851 S.n3488 SUB 0.30fF $ **FLOATING
C3852 S.n3489 SUB 0.41fF $ **FLOATING
C3853 S.n3490 SUB 0.20fF $ **FLOATING
C3854 S.t268 SUB 0.02fF
C3855 S.n3491 SUB 0.24fF $ **FLOATING
C3856 S.n3492 SUB 0.35fF $ **FLOATING
C3857 S.n3493 SUB 0.60fF $ **FLOATING
C3858 S.n3494 SUB 0.12fF $ **FLOATING
C3859 S.t716 SUB 0.02fF
C3860 S.n3495 SUB 0.14fF $ **FLOATING
C3861 S.n3497 SUB 0.04fF $ **FLOATING
C3862 S.n3498 SUB 0.03fF $ **FLOATING
C3863 S.n3499 SUB 0.03fF $ **FLOATING
C3864 S.n3500 SUB 0.10fF $ **FLOATING
C3865 S.n3501 SUB 0.36fF $ **FLOATING
C3866 S.n3502 SUB 0.37fF $ **FLOATING
C3867 S.n3503 SUB 0.10fF $ **FLOATING
C3868 S.n3504 SUB 0.12fF $ **FLOATING
C3869 S.n3505 SUB 0.07fF $ **FLOATING
C3870 S.n3506 SUB 0.12fF $ **FLOATING
C3871 S.n3507 SUB 0.18fF $ **FLOATING
C3872 S.n3508 SUB 3.95fF $ **FLOATING
C3873 S.t945 SUB 0.02fF
C3874 S.n3509 SUB 0.24fF $ **FLOATING
C3875 S.n3510 SUB 0.90fF $ **FLOATING
C3876 S.n3511 SUB 0.05fF $ **FLOATING
C3877 S.t828 SUB 0.02fF
C3878 S.n3512 SUB 0.12fF $ **FLOATING
C3879 S.n3513 SUB 0.14fF $ **FLOATING
C3880 S.n3515 SUB 0.25fF $ **FLOATING
C3881 S.n3516 SUB 0.09fF $ **FLOATING
C3882 S.n3517 SUB 0.21fF $ **FLOATING
C3883 S.n3518 SUB 1.27fF $ **FLOATING
C3884 S.n3519 SUB 0.52fF $ **FLOATING
C3885 S.n3520 SUB 1.86fF $ **FLOATING
C3886 S.n3521 SUB 0.12fF $ **FLOATING
C3887 S.t335 SUB 0.02fF
C3888 S.n3522 SUB 0.14fF $ **FLOATING
C3889 S.t990 SUB 0.02fF
C3890 S.n3524 SUB 0.24fF $ **FLOATING
C3891 S.n3525 SUB 0.35fF $ **FLOATING
C3892 S.n3526 SUB 0.60fF $ **FLOATING
C3893 S.n3527 SUB 1.56fF $ **FLOATING
C3894 S.n3528 SUB 2.42fF $ **FLOATING
C3895 S.t567 SUB 0.02fF
C3896 S.n3529 SUB 0.24fF $ **FLOATING
C3897 S.n3530 SUB 0.90fF $ **FLOATING
C3898 S.n3531 SUB 0.05fF $ **FLOATING
C3899 S.t453 SUB 0.02fF
C3900 S.n3532 SUB 0.12fF $ **FLOATING
C3901 S.n3533 SUB 0.14fF $ **FLOATING
C3902 S.n3535 SUB 1.87fF $ **FLOATING
C3903 S.n3536 SUB 0.06fF $ **FLOATING
C3904 S.n3537 SUB 0.03fF $ **FLOATING
C3905 S.n3538 SUB 0.03fF $ **FLOATING
C3906 S.n3539 SUB 0.98fF $ **FLOATING
C3907 S.n3540 SUB 0.02fF $ **FLOATING
C3908 S.n3541 SUB 0.01fF $ **FLOATING
C3909 S.n3542 SUB 0.02fF $ **FLOATING
C3910 S.n3543 SUB 0.08fF $ **FLOATING
C3911 S.n3544 SUB 0.36fF $ **FLOATING
C3912 S.n3545 SUB 1.83fF $ **FLOATING
C3913 S.t614 SUB 0.02fF
C3914 S.n3546 SUB 0.24fF $ **FLOATING
C3915 S.n3547 SUB 0.35fF $ **FLOATING
C3916 S.n3548 SUB 0.60fF $ **FLOATING
C3917 S.n3549 SUB 0.12fF $ **FLOATING
C3918 S.t1064 SUB 0.02fF
C3919 S.n3550 SUB 0.14fF $ **FLOATING
C3920 S.n3552 SUB 0.69fF $ **FLOATING
C3921 S.n3553 SUB 0.22fF $ **FLOATING
C3922 S.n3554 SUB 0.22fF $ **FLOATING
C3923 S.n3555 SUB 0.69fF $ **FLOATING
C3924 S.n3556 SUB 1.14fF $ **FLOATING
C3925 S.n3557 SUB 0.22fF $ **FLOATING
C3926 S.n3558 SUB 0.25fF $ **FLOATING
C3927 S.n3559 SUB 0.09fF $ **FLOATING
C3928 S.n3560 SUB 1.86fF $ **FLOATING
C3929 S.t175 SUB 0.02fF
C3930 S.n3561 SUB 0.24fF $ **FLOATING
C3931 S.n3562 SUB 0.90fF $ **FLOATING
C3932 S.n3563 SUB 0.05fF $ **FLOATING
C3933 S.t43 SUB 0.02fF
C3934 S.n3564 SUB 0.12fF $ **FLOATING
C3935 S.n3565 SUB 0.14fF $ **FLOATING
C3936 S.n3567 SUB 14.09fF $ **FLOATING
C3937 S.n3568 SUB 0.06fF $ **FLOATING
C3938 S.n3569 SUB 0.20fF $ **FLOATING
C3939 S.n3570 SUB 0.09fF $ **FLOATING
C3940 S.n3571 SUB 0.20fF $ **FLOATING
C3941 S.n3572 SUB 0.09fF $ **FLOATING
C3942 S.n3573 SUB 0.30fF $ **FLOATING
C3943 S.n3574 SUB 0.69fF $ **FLOATING
C3944 S.n3575 SUB 0.44fF $ **FLOATING
C3945 S.n3576 SUB 2.31fF $ **FLOATING
C3946 S.n3577 SUB 0.12fF $ **FLOATING
C3947 S.t762 SUB 0.02fF
C3948 S.n3578 SUB 0.14fF $ **FLOATING
C3949 S.t885 SUB 0.02fF
C3950 S.n3580 SUB 0.24fF $ **FLOATING
C3951 S.n3581 SUB 0.35fF $ **FLOATING
C3952 S.n3582 SUB 0.60fF $ **FLOATING
C3953 S.n3583 SUB 1.88fF $ **FLOATING
C3954 S.n3584 SUB 0.17fF $ **FLOATING
C3955 S.n3585 SUB 0.76fF $ **FLOATING
C3956 S.n3586 SUB 0.31fF $ **FLOATING
C3957 S.n3587 SUB 0.25fF $ **FLOATING
C3958 S.n3588 SUB 0.29fF $ **FLOATING
C3959 S.n3589 SUB 0.46fF $ **FLOATING
C3960 S.n3590 SUB 0.16fF $ **FLOATING
C3961 S.n3591 SUB 1.91fF $ **FLOATING
C3962 S.t803 SUB 0.02fF
C3963 S.n3592 SUB 0.12fF $ **FLOATING
C3964 S.n3593 SUB 0.14fF $ **FLOATING
C3965 S.t281 SUB 0.02fF
C3966 S.n3595 SUB 0.24fF $ **FLOATING
C3967 S.n3596 SUB 0.90fF $ **FLOATING
C3968 S.n3597 SUB 0.05fF $ **FLOATING
C3969 S.n3598 SUB 1.86fF $ **FLOATING
C3970 S.n3599 SUB 0.12fF $ **FLOATING
C3971 S.t95 SUB 0.02fF
C3972 S.n3600 SUB 0.14fF $ **FLOATING
C3973 S.t443 SUB 0.02fF
C3974 S.n3602 SUB 1.20fF $ **FLOATING
C3975 S.n3603 SUB 0.36fF $ **FLOATING
C3976 S.n3604 SUB 1.21fF $ **FLOATING
C3977 S.n3605 SUB 0.60fF $ **FLOATING
C3978 S.n3606 SUB 0.35fF $ **FLOATING
C3979 S.n3607 SUB 0.62fF $ **FLOATING
C3980 S.n3608 SUB 1.14fF $ **FLOATING
C3981 S.n3609 SUB 2.18fF $ **FLOATING
C3982 S.n3610 SUB 0.59fF $ **FLOATING
C3983 S.n3611 SUB 0.02fF $ **FLOATING
C3984 S.n3612 SUB 0.96fF $ **FLOATING
C3985 S.t19 SUB 14.50fF
C3986 S.n3613 SUB 14.37fF $ **FLOATING
C3987 S.n3615 SUB 0.37fF $ **FLOATING
C3988 S.n3616 SUB 0.23fF $ **FLOATING
C3989 S.n3617 SUB 2.76fF $ **FLOATING
C3990 S.n3618 SUB 2.43fF $ **FLOATING
C3991 S.n3619 SUB 3.95fF $ **FLOATING
C3992 S.n3620 SUB 0.25fF $ **FLOATING
C3993 S.n3621 SUB 0.01fF $ **FLOATING
C3994 S.t306 SUB 0.02fF
C3995 S.n3622 SUB 0.25fF $ **FLOATING
C3996 S.t53 SUB 0.02fF
C3997 S.n3623 SUB 0.94fF $ **FLOATING
C3998 S.n3624 SUB 0.70fF $ **FLOATING
C3999 S.n3625 SUB 1.87fF $ **FLOATING
C4000 S.n3626 SUB 1.71fF $ **FLOATING
C4001 S.t20 SUB 0.02fF
C4002 S.n3627 SUB 0.24fF $ **FLOATING
C4003 S.n3628 SUB 0.35fF $ **FLOATING
C4004 S.n3629 SUB 0.60fF $ **FLOATING
C4005 S.n3630 SUB 0.12fF $ **FLOATING
C4006 S.t1069 SUB 0.02fF
C4007 S.n3631 SUB 0.14fF $ **FLOATING
C4008 S.n3633 SUB 1.14fF $ **FLOATING
C4009 S.n3634 SUB 0.22fF $ **FLOATING
C4010 S.n3635 SUB 0.25fF $ **FLOATING
C4011 S.n3636 SUB 0.09fF $ **FLOATING
C4012 S.n3637 SUB 2.41fF $ **FLOATING
C4013 S.t796 SUB 0.02fF
C4014 S.n3638 SUB 0.24fF $ **FLOATING
C4015 S.n3639 SUB 0.90fF $ **FLOATING
C4016 S.n3640 SUB 0.05fF $ **FLOATING
C4017 S.t291 SUB 0.02fF
C4018 S.n3641 SUB 0.12fF $ **FLOATING
C4019 S.n3642 SUB 0.14fF $ **FLOATING
C4020 S.n3644 SUB 1.86fF $ **FLOATING
C4021 S.n3645 SUB 0.47fF $ **FLOATING
C4022 S.n3646 SUB 0.09fF $ **FLOATING
C4023 S.n3647 SUB 0.32fF $ **FLOATING
C4024 S.n3648 SUB 0.30fF $ **FLOATING
C4025 S.n3649 SUB 0.76fF $ **FLOATING
C4026 S.n3650 SUB 0.58fF $ **FLOATING
C4027 S.t922 SUB 0.02fF
C4028 S.n3651 SUB 0.24fF $ **FLOATING
C4029 S.n3652 SUB 0.35fF $ **FLOATING
C4030 S.n3653 SUB 0.60fF $ **FLOATING
C4031 S.n3654 SUB 0.12fF $ **FLOATING
C4032 S.t133 SUB 0.02fF
C4033 S.n3655 SUB 0.14fF $ **FLOATING
C4034 S.n3657 SUB 2.58fF $ **FLOATING
C4035 S.n3658 SUB 2.13fF $ **FLOATING
C4036 S.t623 SUB 0.02fF
C4037 S.n3659 SUB 0.24fF $ **FLOATING
C4038 S.n3660 SUB 0.90fF $ **FLOATING
C4039 S.n3661 SUB 0.05fF $ **FLOATING
C4040 S.t1019 SUB 0.02fF
C4041 S.n3662 SUB 0.12fF $ **FLOATING
C4042 S.n3663 SUB 0.14fF $ **FLOATING
C4043 S.n3665 SUB 0.77fF $ **FLOATING
C4044 S.n3666 SUB 2.27fF $ **FLOATING
C4045 S.n3667 SUB 1.86fF $ **FLOATING
C4046 S.n3668 SUB 0.12fF $ **FLOATING
C4047 S.t862 SUB 0.02fF
C4048 S.n3669 SUB 0.14fF $ **FLOATING
C4049 S.t544 SUB 0.02fF
C4050 S.n3671 SUB 0.24fF $ **FLOATING
C4051 S.n3672 SUB 0.35fF $ **FLOATING
C4052 S.n3673 SUB 0.60fF $ **FLOATING
C4053 S.n3674 SUB 1.37fF $ **FLOATING
C4054 S.n3675 SUB 0.70fF $ **FLOATING
C4055 S.n3676 SUB 1.13fF $ **FLOATING
C4056 S.n3677 SUB 0.35fF $ **FLOATING
C4057 S.n3678 SUB 2.00fF $ **FLOATING
C4058 S.t235 SUB 0.02fF
C4059 S.n3679 SUB 0.24fF $ **FLOATING
C4060 S.n3680 SUB 0.90fF $ **FLOATING
C4061 S.n3681 SUB 0.05fF $ **FLOATING
C4062 S.t11 SUB 0.02fF
C4063 S.n3682 SUB 0.12fF $ **FLOATING
C4064 S.n3683 SUB 0.14fF $ **FLOATING
C4065 S.n3685 SUB 1.87fF $ **FLOATING
C4066 S.n3686 SUB 1.86fF $ **FLOATING
C4067 S.t154 SUB 0.02fF
C4068 S.n3687 SUB 0.24fF $ **FLOATING
C4069 S.n3688 SUB 0.35fF $ **FLOATING
C4070 S.n3689 SUB 0.60fF $ **FLOATING
C4071 S.n3690 SUB 0.12fF $ **FLOATING
C4072 S.t486 SUB 0.02fF
C4073 S.n3691 SUB 0.14fF $ **FLOATING
C4074 S.n3693 SUB 1.14fF $ **FLOATING
C4075 S.n3694 SUB 0.22fF $ **FLOATING
C4076 S.n3695 SUB 0.25fF $ **FLOATING
C4077 S.n3696 SUB 0.09fF $ **FLOATING
C4078 S.n3697 SUB 1.86fF $ **FLOATING
C4079 S.t959 SUB 0.02fF
C4080 S.n3698 SUB 0.24fF $ **FLOATING
C4081 S.n3699 SUB 0.90fF $ **FLOATING
C4082 S.n3700 SUB 0.05fF $ **FLOATING
C4083 S.t768 SUB 0.02fF
C4084 S.n3701 SUB 0.12fF $ **FLOATING
C4085 S.n3702 SUB 0.14fF $ **FLOATING
C4086 S.n3704 SUB 14.09fF $ **FLOATING
C4087 S.n3705 SUB 1.86fF $ **FLOATING
C4088 S.n3706 SUB 2.64fF $ **FLOATING
C4089 S.t115 SUB 0.02fF
C4090 S.n3707 SUB 0.24fF $ **FLOATING
C4091 S.n3708 SUB 0.35fF $ **FLOATING
C4092 S.n3709 SUB 0.60fF $ **FLOATING
C4093 S.n3710 SUB 0.12fF $ **FLOATING
C4094 S.t452 SUB 0.02fF
C4095 S.n3711 SUB 0.14fF $ **FLOATING
C4096 S.n3713 SUB 2.77fF $ **FLOATING
C4097 S.n3714 SUB 2.28fF $ **FLOATING
C4098 S.t797 SUB 0.02fF
C4099 S.n3715 SUB 0.12fF $ **FLOATING
C4100 S.n3716 SUB 0.14fF $ **FLOATING
C4101 S.t905 SUB 0.02fF
C4102 S.n3718 SUB 0.24fF $ **FLOATING
C4103 S.n3719 SUB 0.90fF $ **FLOATING
C4104 S.n3720 SUB 0.05fF $ **FLOATING
C4105 S.n3721 SUB 1.86fF $ **FLOATING
C4106 S.n3722 SUB 2.64fF $ **FLOATING
C4107 S.t848 SUB 0.02fF
C4108 S.n3723 SUB 0.24fF $ **FLOATING
C4109 S.n3724 SUB 0.35fF $ **FLOATING
C4110 S.n3725 SUB 0.60fF $ **FLOATING
C4111 S.n3726 SUB 0.12fF $ **FLOATING
C4112 S.t41 SUB 0.02fF
C4113 S.n3727 SUB 0.14fF $ **FLOATING
C4114 S.n3729 SUB 2.77fF $ **FLOATING
C4115 S.n3730 SUB 2.28fF $ **FLOATING
C4116 S.t416 SUB 0.02fF
C4117 S.n3731 SUB 0.12fF $ **FLOATING
C4118 S.n3732 SUB 0.14fF $ **FLOATING
C4119 S.t531 SUB 0.02fF
C4120 S.n3734 SUB 0.24fF $ **FLOATING
C4121 S.n3735 SUB 0.90fF $ **FLOATING
C4122 S.n3736 SUB 0.05fF $ **FLOATING
C4123 S.n3737 SUB 2.77fF $ **FLOATING
C4124 S.n3738 SUB 1.86fF $ **FLOATING
C4125 S.n3739 SUB 0.12fF $ **FLOATING
C4126 S.t786 SUB 0.02fF
C4127 S.n3740 SUB 0.14fF $ **FLOATING
C4128 S.t473 SUB 0.02fF
C4129 S.n3742 SUB 0.24fF $ **FLOATING
C4130 S.n3743 SUB 0.35fF $ **FLOATING
C4131 S.n3744 SUB 0.60fF $ **FLOATING
C4132 S.n3745 SUB 2.64fF $ **FLOATING
C4133 S.n3746 SUB 2.28fF $ **FLOATING
C4134 S.t1132 SUB 0.02fF
C4135 S.n3747 SUB 0.12fF $ **FLOATING
C4136 S.n3748 SUB 0.14fF $ **FLOATING
C4137 S.t144 SUB 0.02fF
C4138 S.n3750 SUB 0.24fF $ **FLOATING
C4139 S.n3751 SUB 0.90fF $ **FLOATING
C4140 S.n3752 SUB 0.05fF $ **FLOATING
C4141 S.n3753 SUB 1.86fF $ **FLOATING
C4142 S.n3754 SUB 2.65fF $ **FLOATING
C4143 S.t73 SUB 0.02fF
C4144 S.n3755 SUB 0.24fF $ **FLOATING
C4145 S.n3756 SUB 0.35fF $ **FLOATING
C4146 S.n3757 SUB 0.60fF $ **FLOATING
C4147 S.n3758 SUB 0.12fF $ **FLOATING
C4148 S.t404 SUB 0.02fF
C4149 S.n3759 SUB 0.14fF $ **FLOATING
C4150 S.n3761 SUB 5.11fF $ **FLOATING
C4151 S.t747 SUB 0.02fF
C4152 S.n3762 SUB 0.12fF $ **FLOATING
C4153 S.n3763 SUB 0.14fF $ **FLOATING
C4154 S.t871 SUB 0.02fF
C4155 S.n3765 SUB 0.24fF $ **FLOATING
C4156 S.n3766 SUB 0.90fF $ **FLOATING
C4157 S.n3767 SUB 0.05fF $ **FLOATING
C4158 S.n3768 SUB 2.70fF $ **FLOATING
C4159 S.n3769 SUB 1.58fF $ **FLOATING
C4160 S.n3770 SUB 0.12fF $ **FLOATING
C4161 S.t153 SUB 0.02fF
C4162 S.n3771 SUB 0.14fF $ **FLOATING
C4163 S.t694 SUB 0.02fF
C4164 S.n3773 SUB 0.24fF $ **FLOATING
C4165 S.n3774 SUB 0.35fF $ **FLOATING
C4166 S.n3775 SUB 0.60fF $ **FLOATING
C4167 S.n3776 SUB 0.07fF $ **FLOATING
C4168 S.n3777 SUB 0.01fF $ **FLOATING
C4169 S.n3778 SUB 0.23fF $ **FLOATING
C4170 S.n3779 SUB 1.15fF $ **FLOATING
C4171 S.n3780 SUB 1.33fF $ **FLOATING
C4172 S.n3781 SUB 2.28fF $ **FLOATING
C4173 S.t487 SUB 0.02fF
C4174 S.n3782 SUB 0.12fF $ **FLOATING
C4175 S.n3783 SUB 0.14fF $ **FLOATING
C4176 S.t1136 SUB 0.02fF
C4177 S.n3785 SUB 0.24fF $ **FLOATING
C4178 S.n3786 SUB 0.90fF $ **FLOATING
C4179 S.n3787 SUB 0.05fF $ **FLOATING
C4180 S.t10 SUB 32.35fF
C4181 S.t387 SUB 0.02fF
C4182 S.n3788 SUB 0.12fF $ **FLOATING
C4183 S.n3789 SUB 0.14fF $ **FLOATING
C4184 S.t577 SUB 0.02fF
C4185 S.n3791 SUB 0.24fF $ **FLOATING
C4186 S.n3792 SUB 0.90fF $ **FLOATING
C4187 S.n3793 SUB 0.05fF $ **FLOATING
C4188 S.t883 SUB 0.02fF
C4189 S.n3794 SUB 0.24fF $ **FLOATING
C4190 S.n3795 SUB 0.35fF $ **FLOATING
C4191 S.n3796 SUB 0.60fF $ **FLOATING
C4192 S.n3797 SUB 0.31fF $ **FLOATING
C4193 S.n3798 SUB 1.08fF $ **FLOATING
C4194 S.n3799 SUB 0.15fF $ **FLOATING
C4195 S.n3800 SUB 2.08fF $ **FLOATING
C4196 S.n3801 SUB 2.91fF $ **FLOATING
C4197 S.n3802 SUB 1.86fF $ **FLOATING
C4198 S.n3803 SUB 0.12fF $ **FLOATING
C4199 S.t682 SUB 0.02fF
C4200 S.n3804 SUB 0.14fF $ **FLOATING
C4201 S.t226 SUB 0.02fF
C4202 S.n3806 SUB 0.24fF $ **FLOATING
C4203 S.n3807 SUB 0.35fF $ **FLOATING
C4204 S.n3808 SUB 0.60fF $ **FLOATING
C4205 S.n3809 SUB 0.91fF $ **FLOATING
C4206 S.n3810 SUB 0.31fF $ **FLOATING
C4207 S.n3811 SUB 0.91fF $ **FLOATING
C4208 S.n3812 SUB 1.08fF $ **FLOATING
C4209 S.n3813 SUB 0.15fF $ **FLOATING
C4210 S.n3814 SUB 4.90fF $ **FLOATING
C4211 S.t787 SUB 0.02fF
C4212 S.n3815 SUB 0.12fF $ **FLOATING
C4213 S.n3816 SUB 0.14fF $ **FLOATING
C4214 S.t899 SUB 0.02fF
C4215 S.n3818 SUB 0.24fF $ **FLOATING
C4216 S.n3819 SUB 0.90fF $ **FLOATING
C4217 S.n3820 SUB 0.05fF $ **FLOATING
C4218 S.n3821 SUB 1.86fF $ **FLOATING
C4219 S.n3822 SUB 2.64fF $ **FLOATING
C4220 S.t1010 SUB 0.02fF
C4221 S.n3823 SUB 0.24fF $ **FLOATING
C4222 S.n3824 SUB 0.35fF $ **FLOATING
C4223 S.n3825 SUB 0.60fF $ **FLOATING
C4224 S.n3826 SUB 0.12fF $ **FLOATING
C4225 S.t361 SUB 0.02fF
C4226 S.n3827 SUB 0.14fF $ **FLOATING
C4227 S.n3829 SUB 1.86fF $ **FLOATING
C4228 S.n3830 SUB 2.64fF $ **FLOATING
C4229 S.t508 SUB 0.02fF
C4230 S.n3831 SUB 0.24fF $ **FLOATING
C4231 S.n3832 SUB 0.35fF $ **FLOATING
C4232 S.n3833 SUB 0.60fF $ **FLOATING
C4233 S.t183 SUB 0.02fF
C4234 S.n3834 SUB 0.24fF $ **FLOATING
C4235 S.n3835 SUB 0.90fF $ **FLOATING
C4236 S.n3836 SUB 0.05fF $ **FLOATING
C4237 S.t1104 SUB 0.02fF
C4238 S.n3837 SUB 0.12fF $ **FLOATING
C4239 S.n3838 SUB 0.14fF $ **FLOATING
C4240 S.n3840 SUB 0.12fF $ **FLOATING
C4241 S.t829 SUB 0.02fF
C4242 S.n3841 SUB 0.14fF $ **FLOATING
C4243 S.n3843 SUB 2.28fF $ **FLOATING
C4244 S.n3844 SUB 2.91fF $ **FLOATING
C4245 S.n3845 SUB 5.10fF $ **FLOATING
C4246 S.t405 SUB 0.02fF
C4247 S.n3846 SUB 0.12fF $ **FLOATING
C4248 S.n3847 SUB 0.14fF $ **FLOATING
C4249 S.t596 SUB 0.02fF
C4250 S.n3849 SUB 0.24fF $ **FLOATING
C4251 S.n3850 SUB 0.90fF $ **FLOATING
C4252 S.n3851 SUB 0.05fF $ **FLOATING
C4253 S.n3852 SUB 1.86fF $ **FLOATING
C4254 S.n3853 SUB 2.64fF $ **FLOATING
C4255 S.t633 SUB 0.02fF
C4256 S.n3854 SUB 0.24fF $ **FLOATING
C4257 S.n3855 SUB 0.35fF $ **FLOATING
C4258 S.n3856 SUB 0.60fF $ **FLOATING
C4259 S.n3857 SUB 0.12fF $ **FLOATING
C4260 S.t1087 SUB 0.02fF
C4261 S.n3858 SUB 0.14fF $ **FLOATING
C4262 S.n3860 SUB 5.11fF $ **FLOATING
C4263 S.t1122 SUB 0.02fF
C4264 S.n3861 SUB 0.12fF $ **FLOATING
C4265 S.n3862 SUB 0.14fF $ **FLOATING
C4266 S.t201 SUB 0.02fF
C4267 S.n3864 SUB 0.24fF $ **FLOATING
C4268 S.n3865 SUB 0.90fF $ **FLOATING
C4269 S.n3866 SUB 0.05fF $ **FLOATING
C4270 S.n3867 SUB 1.86fF $ **FLOATING
C4271 S.n3868 SUB 2.64fF $ **FLOATING
C4272 S.t249 SUB 0.02fF
C4273 S.n3869 SUB 0.24fF $ **FLOATING
C4274 S.n3870 SUB 0.35fF $ **FLOATING
C4275 S.n3871 SUB 0.60fF $ **FLOATING
C4276 S.n3872 SUB 0.12fF $ **FLOATING
C4277 S.t700 SUB 0.02fF
C4278 S.n3873 SUB 0.14fF $ **FLOATING
C4279 S.n3875 SUB 5.11fF $ **FLOATING
C4280 S.t733 SUB 0.02fF
C4281 S.n3876 SUB 0.12fF $ **FLOATING
C4282 S.n3877 SUB 0.14fF $ **FLOATING
C4283 S.t923 SUB 0.02fF
C4284 S.n3879 SUB 0.24fF $ **FLOATING
C4285 S.n3880 SUB 0.90fF $ **FLOATING
C4286 S.n3881 SUB 0.05fF $ **FLOATING
C4287 S.n3882 SUB 1.86fF $ **FLOATING
C4288 S.n3883 SUB 0.12fF $ **FLOATING
C4289 S.t320 SUB 0.02fF
C4290 S.n3884 SUB 0.14fF $ **FLOATING
C4291 S.t974 SUB 0.02fF
C4292 S.n3886 SUB 0.24fF $ **FLOATING
C4293 S.n3887 SUB 0.35fF $ **FLOATING
C4294 S.n3888 SUB 0.60fF $ **FLOATING
C4295 S.n3889 SUB 2.64fF $ **FLOATING
C4296 S.n3890 SUB 4.85fF $ **FLOATING
C4297 S.t351 SUB 0.02fF
C4298 S.n3891 SUB 0.12fF $ **FLOATING
C4299 S.n3892 SUB 0.14fF $ **FLOATING
C4300 S.t545 SUB 0.02fF
C4301 S.n3894 SUB 0.24fF $ **FLOATING
C4302 S.n3895 SUB 0.90fF $ **FLOATING
C4303 S.n3896 SUB 0.05fF $ **FLOATING
C4304 S.n3897 SUB 1.86fF $ **FLOATING
C4305 S.n3898 SUB 2.64fF $ **FLOATING
C4306 S.t513 SUB 0.02fF
C4307 S.n3899 SUB 0.24fF $ **FLOATING
C4308 S.n3900 SUB 0.35fF $ **FLOATING
C4309 S.n3901 SUB 0.60fF $ **FLOATING
C4310 S.n3902 SUB 0.12fF $ **FLOATING
C4311 S.t240 SUB 0.02fF
C4312 S.n3903 SUB 0.14fF $ **FLOATING
C4313 S.n3905 SUB 5.38fF $ **FLOATING
C4314 S.t1079 SUB 0.02fF
C4315 S.n3906 SUB 0.12fF $ **FLOATING
C4316 S.n3907 SUB 0.14fF $ **FLOATING
C4317 S.t274 SUB 0.02fF
C4318 S.n3909 SUB 0.24fF $ **FLOATING
C4319 S.n3910 SUB 0.90fF $ **FLOATING
C4320 S.n3911 SUB 0.05fF $ **FLOATING
C4321 S.t42 SUB 31.97fF
C4322 S.t584 SUB 0.02fF
C4323 S.n3912 SUB 1.18fF $ **FLOATING
C4324 S.n3913 SUB 0.05fF $ **FLOATING
C4325 S.t1016 SUB 0.02fF
C4326 S.n3914 SUB 0.01fF $ **FLOATING
C4327 S.n3915 SUB 0.25fF $ **FLOATING
C4328 S.n3917 SUB 1.48fF $ **FLOATING
C4329 S.n3918 SUB 1.29fF $ **FLOATING
C4330 S.n3919 SUB 0.27fF $ **FLOATING
C4331 S.n3920 SUB 0.24fF $ **FLOATING
C4332 S.n3921 SUB 4.34fF $ **FLOATING
C4333 S.n3922 SUB 0.01fF $ **FLOATING
C4334 S.n3923 SUB 0.02fF $ **FLOATING
C4335 S.n3924 SUB 0.03fF $ **FLOATING
C4336 S.n3925 SUB 0.04fF $ **FLOATING
C4337 S.n3926 SUB 0.17fF $ **FLOATING
C4338 S.n3927 SUB 0.01fF $ **FLOATING
C4339 S.n3928 SUB 0.02fF $ **FLOATING
C4340 S.n3929 SUB 0.01fF $ **FLOATING
C4341 S.n3930 SUB 0.01fF $ **FLOATING
C4342 S.n3931 SUB 0.01fF $ **FLOATING
C4343 S.n3932 SUB 0.01fF $ **FLOATING
C4344 S.n3933 SUB 0.01fF $ **FLOATING
C4345 S.n3934 SUB 0.01fF $ **FLOATING
C4346 S.n3935 SUB 0.02fF $ **FLOATING
C4347 S.n3936 SUB 0.05fF $ **FLOATING
C4348 S.n3937 SUB 0.04fF $ **FLOATING
C4349 S.n3938 SUB 0.11fF $ **FLOATING
C4350 S.n3939 SUB 0.37fF $ **FLOATING
C4351 S.n3940 SUB 0.20fF $ **FLOATING
C4352 S.n3941 SUB 8.87fF $ **FLOATING
C4353 S.n3942 SUB 8.87fF $ **FLOATING
C4354 S.n3943 SUB 0.59fF $ **FLOATING
C4355 S.n3944 SUB 0.21fF $ **FLOATING
C4356 S.n3945 SUB 0.59fF $ **FLOATING
C4357 S.n3946 SUB 2.57fF $ **FLOATING
C4358 S.n3947 SUB 0.29fF $ **FLOATING
C4359 S.t156 SUB 14.50fF
C4360 S.n3948 SUB 15.77fF $ **FLOATING
C4361 S.n3949 SUB 0.76fF $ **FLOATING
C4362 S.n3950 SUB 0.27fF $ **FLOATING
C4363 S.n3951 SUB 3.96fF $ **FLOATING
C4364 S.n3952 SUB 1.34fF $ **FLOATING
C4365 S.t635 SUB 0.02fF
C4366 S.n3953 SUB 0.63fF $ **FLOATING
C4367 S.n3954 SUB 0.60fF $ **FLOATING
C4368 S.n3955 SUB 1.86fF $ **FLOATING
C4369 S.n3956 SUB 0.45fF $ **FLOATING
C4370 S.n3957 SUB 0.22fF $ **FLOATING
C4371 S.n3958 SUB 0.38fF $ **FLOATING
C4372 S.n3959 SUB 0.16fF $ **FLOATING
C4373 S.n3960 SUB 0.28fF $ **FLOATING
C4374 S.n3961 SUB 0.21fF $ **FLOATING
C4375 S.n3962 SUB 0.30fF $ **FLOATING
C4376 S.n3963 SUB 0.41fF $ **FLOATING
C4377 S.n3964 SUB 0.20fF $ **FLOATING
C4378 S.t354 SUB 0.02fF
C4379 S.n3965 SUB 0.24fF $ **FLOATING
C4380 S.n3966 SUB 0.35fF $ **FLOATING
C4381 S.n3967 SUB 0.60fF $ **FLOATING
C4382 S.n3968 SUB 0.12fF $ **FLOATING
C4383 S.t138 SUB 0.02fF
C4384 S.n3969 SUB 0.14fF $ **FLOATING
C4385 S.n3971 SUB 0.04fF $ **FLOATING
C4386 S.n3972 SUB 0.03fF $ **FLOATING
C4387 S.n3973 SUB 0.03fF $ **FLOATING
C4388 S.n3974 SUB 0.10fF $ **FLOATING
C4389 S.n3975 SUB 0.36fF $ **FLOATING
C4390 S.n3976 SUB 0.37fF $ **FLOATING
C4391 S.n3977 SUB 0.10fF $ **FLOATING
C4392 S.n3978 SUB 0.12fF $ **FLOATING
C4393 S.n3979 SUB 0.07fF $ **FLOATING
C4394 S.n3980 SUB 0.12fF $ **FLOATING
C4395 S.n3981 SUB 0.18fF $ **FLOATING
C4396 S.n3982 SUB 3.95fF $ **FLOATING
C4397 S.t864 SUB 0.02fF
C4398 S.n3983 SUB 0.24fF $ **FLOATING
C4399 S.n3984 SUB 0.90fF $ **FLOATING
C4400 S.n3985 SUB 0.05fF $ **FLOATING
C4401 S.t246 SUB 0.02fF
C4402 S.n3986 SUB 0.12fF $ **FLOATING
C4403 S.n3987 SUB 0.14fF $ **FLOATING
C4404 S.n3989 SUB 0.25fF $ **FLOATING
C4405 S.n3990 SUB 0.09fF $ **FLOATING
C4406 S.n3991 SUB 0.21fF $ **FLOATING
C4407 S.n3992 SUB 1.27fF $ **FLOATING
C4408 S.n3993 SUB 0.52fF $ **FLOATING
C4409 S.n3994 SUB 1.86fF $ **FLOATING
C4410 S.n3995 SUB 0.12fF $ **FLOATING
C4411 S.t724 SUB 0.02fF
C4412 S.n3996 SUB 0.14fF $ **FLOATING
C4413 S.t1004 SUB 0.02fF
C4414 S.n3998 SUB 0.24fF $ **FLOATING
C4415 S.n3999 SUB 0.35fF $ **FLOATING
C4416 S.n4000 SUB 0.60fF $ **FLOATING
C4417 S.n4001 SUB 1.56fF $ **FLOATING
C4418 S.n4002 SUB 2.42fF $ **FLOATING
C4419 S.t585 SUB 0.02fF
C4420 S.n4003 SUB 0.24fF $ **FLOATING
C4421 S.n4004 SUB 0.90fF $ **FLOATING
C4422 S.n4005 SUB 0.05fF $ **FLOATING
C4423 S.t835 SUB 0.02fF
C4424 S.n4006 SUB 0.12fF $ **FLOATING
C4425 S.n4007 SUB 0.14fF $ **FLOATING
C4426 S.n4009 SUB 1.87fF $ **FLOATING
C4427 S.n4010 SUB 0.06fF $ **FLOATING
C4428 S.n4011 SUB 0.03fF $ **FLOATING
C4429 S.n4012 SUB 0.03fF $ **FLOATING
C4430 S.n4013 SUB 0.98fF $ **FLOATING
C4431 S.n4014 SUB 0.02fF $ **FLOATING
C4432 S.n4015 SUB 0.01fF $ **FLOATING
C4433 S.n4016 SUB 0.02fF $ **FLOATING
C4434 S.n4017 SUB 0.08fF $ **FLOATING
C4435 S.n4018 SUB 0.36fF $ **FLOATING
C4436 S.n4019 SUB 1.83fF $ **FLOATING
C4437 S.t625 SUB 0.02fF
C4438 S.n4020 SUB 0.24fF $ **FLOATING
C4439 S.n4021 SUB 0.35fF $ **FLOATING
C4440 S.n4022 SUB 0.60fF $ **FLOATING
C4441 S.n4023 SUB 0.12fF $ **FLOATING
C4442 S.t344 SUB 0.02fF
C4443 S.n4024 SUB 0.14fF $ **FLOATING
C4444 S.n4026 SUB 0.69fF $ **FLOATING
C4445 S.n4027 SUB 0.22fF $ **FLOATING
C4446 S.n4028 SUB 0.22fF $ **FLOATING
C4447 S.n4029 SUB 0.69fF $ **FLOATING
C4448 S.n4030 SUB 1.14fF $ **FLOATING
C4449 S.n4031 SUB 0.22fF $ **FLOATING
C4450 S.n4032 SUB 0.25fF $ **FLOATING
C4451 S.n4033 SUB 0.09fF $ **FLOATING
C4452 S.n4034 SUB 1.86fF $ **FLOATING
C4453 S.t190 SUB 0.02fF
C4454 S.n4035 SUB 0.24fF $ **FLOATING
C4455 S.n4036 SUB 0.90fF $ **FLOATING
C4456 S.n4037 SUB 0.05fF $ **FLOATING
C4457 S.t460 SUB 0.02fF
C4458 S.n4038 SUB 0.12fF $ **FLOATING
C4459 S.n4039 SUB 0.14fF $ **FLOATING
C4460 S.n4041 SUB 14.09fF $ **FLOATING
C4461 S.n4042 SUB 1.70fF $ **FLOATING
C4462 S.n4043 SUB 0.65fF $ **FLOATING
C4463 S.n4044 SUB 0.68fF $ **FLOATING
C4464 S.n4045 SUB 0.71fF $ **FLOATING
C4465 S.n4046 SUB 0.36fF $ **FLOATING
C4466 S.t737 SUB 0.02fF
C4467 S.n4047 SUB 0.24fF $ **FLOATING
C4468 S.n4048 SUB 0.35fF $ **FLOATING
C4469 S.n4049 SUB 0.60fF $ **FLOATING
C4470 S.n4050 SUB 0.12fF $ **FLOATING
C4471 S.t526 SUB 0.02fF
C4472 S.n4051 SUB 0.14fF $ **FLOATING
C4473 S.n4053 SUB 0.31fF $ **FLOATING
C4474 S.n4054 SUB 0.22fF $ **FLOATING
C4475 S.n4055 SUB 0.65fF $ **FLOATING
C4476 S.n4056 SUB 0.94fF $ **FLOATING
C4477 S.n4057 SUB 0.22fF $ **FLOATING
C4478 S.n4058 SUB 0.20fF $ **FLOATING
C4479 S.n4059 SUB 0.20fF $ **FLOATING
C4480 S.n4060 SUB 0.06fF $ **FLOATING
C4481 S.n4061 SUB 0.09fF $ **FLOATING
C4482 S.n4062 SUB 0.09fF $ **FLOATING
C4483 S.n4063 SUB 1.66fF $ **FLOATING
C4484 S.t563 SUB 0.02fF
C4485 S.n4064 SUB 0.12fF $ **FLOATING
C4486 S.n4065 SUB 0.14fF $ **FLOATING
C4487 S.t139 SUB 0.02fF
C4488 S.n4067 SUB 0.24fF $ **FLOATING
C4489 S.n4068 SUB 0.90fF $ **FLOATING
C4490 S.n4069 SUB 0.05fF $ **FLOATING
C4491 S.n4070 SUB 1.86fF $ **FLOATING
C4492 S.n4071 SUB 0.12fF $ **FLOATING
C4493 S.t108 SUB 0.02fF
C4494 S.n4072 SUB 0.14fF $ **FLOATING
C4495 S.t403 SUB 0.02fF
C4496 S.n4074 SUB 0.12fF $ **FLOATING
C4497 S.n4075 SUB 0.14fF $ **FLOATING
C4498 S.t594 SUB 0.02fF
C4499 S.n4077 SUB 0.24fF $ **FLOATING
C4500 S.n4078 SUB 0.90fF $ **FLOATING
C4501 S.n4079 SUB 0.05fF $ **FLOATING
C4502 S.t890 SUB 0.02fF
C4503 S.n4080 SUB 0.24fF $ **FLOATING
C4504 S.n4081 SUB 0.35fF $ **FLOATING
C4505 S.n4082 SUB 0.60fF $ **FLOATING
C4506 S.n4083 SUB 0.31fF $ **FLOATING
C4507 S.n4084 SUB 1.08fF $ **FLOATING
C4508 S.n4085 SUB 0.15fF $ **FLOATING
C4509 S.n4086 SUB 2.08fF $ **FLOATING
C4510 S.n4087 SUB 2.91fF $ **FLOATING
C4511 S.n4088 SUB 1.86fF $ **FLOATING
C4512 S.n4089 SUB 0.12fF $ **FLOATING
C4513 S.t1068 SUB 0.02fF
C4514 S.n4090 SUB 0.14fF $ **FLOATING
C4515 S.t237 SUB 0.02fF
C4516 S.n4092 SUB 0.24fF $ **FLOATING
C4517 S.n4093 SUB 0.35fF $ **FLOATING
C4518 S.n4094 SUB 0.60fF $ **FLOATING
C4519 S.n4095 SUB 0.91fF $ **FLOATING
C4520 S.n4096 SUB 0.31fF $ **FLOATING
C4521 S.n4097 SUB 0.91fF $ **FLOATING
C4522 S.n4098 SUB 1.08fF $ **FLOATING
C4523 S.n4099 SUB 0.15fF $ **FLOATING
C4524 S.n4100 SUB 4.90fF $ **FLOATING
C4525 S.t55 SUB 0.02fF
C4526 S.n4101 SUB 0.12fF $ **FLOATING
C4527 S.n4102 SUB 0.14fF $ **FLOATING
C4528 S.t914 SUB 0.02fF
C4529 S.n4104 SUB 0.24fF $ **FLOATING
C4530 S.n4105 SUB 0.90fF $ **FLOATING
C4531 S.n4106 SUB 0.05fF $ **FLOATING
C4532 S.n4107 SUB 1.86fF $ **FLOATING
C4533 S.n4108 SUB 2.64fF $ **FLOATING
C4534 S.t966 SUB 0.02fF
C4535 S.n4109 SUB 0.24fF $ **FLOATING
C4536 S.n4110 SUB 0.35fF $ **FLOATING
C4537 S.n4111 SUB 0.60fF $ **FLOATING
C4538 S.n4112 SUB 0.12fF $ **FLOATING
C4539 S.t686 SUB 0.02fF
C4540 S.n4113 SUB 0.14fF $ **FLOATING
C4541 S.n4115 SUB 1.86fF $ **FLOATING
C4542 S.n4116 SUB 2.64fF $ **FLOATING
C4543 S.t519 SUB 0.02fF
C4544 S.n4117 SUB 0.24fF $ **FLOATING
C4545 S.n4118 SUB 0.35fF $ **FLOATING
C4546 S.n4119 SUB 0.60fF $ **FLOATING
C4547 S.t197 SUB 0.02fF
C4548 S.n4120 SUB 0.24fF $ **FLOATING
C4549 S.n4121 SUB 0.90fF $ **FLOATING
C4550 S.n4122 SUB 0.05fF $ **FLOATING
C4551 S.t1123 SUB 0.02fF
C4552 S.n4123 SUB 0.12fF $ **FLOATING
C4553 S.n4124 SUB 0.14fF $ **FLOATING
C4554 S.n4126 SUB 0.12fF $ **FLOATING
C4555 S.t840 SUB 0.02fF
C4556 S.n4127 SUB 0.14fF $ **FLOATING
C4557 S.n4129 SUB 2.28fF $ **FLOATING
C4558 S.n4130 SUB 2.91fF $ **FLOATING
C4559 S.n4131 SUB 5.10fF $ **FLOATING
C4560 S.t795 SUB 0.02fF
C4561 S.n4132 SUB 0.12fF $ **FLOATING
C4562 S.n4133 SUB 0.14fF $ **FLOATING
C4563 S.t536 SUB 0.02fF
C4564 S.n4135 SUB 0.24fF $ **FLOATING
C4565 S.n4136 SUB 0.90fF $ **FLOATING
C4566 S.n4137 SUB 0.05fF $ **FLOATING
C4567 S.n4138 SUB 1.86fF $ **FLOATING
C4568 S.n4139 SUB 2.64fF $ **FLOATING
C4569 S.t642 SUB 0.02fF
C4570 S.n4140 SUB 0.24fF $ **FLOATING
C4571 S.n4141 SUB 0.35fF $ **FLOATING
C4572 S.n4142 SUB 0.60fF $ **FLOATING
C4573 S.n4143 SUB 0.12fF $ **FLOATING
C4574 S.t365 SUB 0.02fF
C4575 S.n4144 SUB 0.14fF $ **FLOATING
C4576 S.n4146 SUB 5.11fF $ **FLOATING
C4577 S.t415 SUB 0.02fF
C4578 S.n4147 SUB 0.12fF $ **FLOATING
C4579 S.n4148 SUB 0.14fF $ **FLOATING
C4580 S.t216 SUB 0.02fF
C4581 S.n4150 SUB 0.24fF $ **FLOATING
C4582 S.n4151 SUB 0.90fF $ **FLOATING
C4583 S.n4152 SUB 0.05fF $ **FLOATING
C4584 S.n4153 SUB 1.86fF $ **FLOATING
C4585 S.n4154 SUB 2.64fF $ **FLOATING
C4586 S.t262 SUB 0.02fF
C4587 S.n4155 SUB 0.24fF $ **FLOATING
C4588 S.n4156 SUB 0.35fF $ **FLOATING
C4589 S.n4157 SUB 0.60fF $ **FLOATING
C4590 S.n4158 SUB 0.12fF $ **FLOATING
C4591 S.t1089 SUB 0.02fF
C4592 S.n4159 SUB 0.14fF $ **FLOATING
C4593 S.n4161 SUB 5.11fF $ **FLOATING
C4594 S.t1134 SUB 0.02fF
C4595 S.n4162 SUB 0.12fF $ **FLOATING
C4596 S.n4163 SUB 0.14fF $ **FLOATING
C4597 S.t941 SUB 0.02fF
C4598 S.n4165 SUB 0.24fF $ **FLOATING
C4599 S.n4166 SUB 0.90fF $ **FLOATING
C4600 S.n4167 SUB 0.05fF $ **FLOATING
C4601 S.n4168 SUB 1.86fF $ **FLOATING
C4602 S.n4169 SUB 0.12fF $ **FLOATING
C4603 S.t703 SUB 0.02fF
C4604 S.n4170 SUB 0.14fF $ **FLOATING
C4605 S.t984 SUB 0.02fF
C4606 S.n4172 SUB 0.24fF $ **FLOATING
C4607 S.n4173 SUB 0.35fF $ **FLOATING
C4608 S.n4174 SUB 0.60fF $ **FLOATING
C4609 S.n4175 SUB 2.64fF $ **FLOATING
C4610 S.n4176 SUB 5.12fF $ **FLOATING
C4611 S.t746 SUB 0.02fF
C4612 S.n4177 SUB 0.12fF $ **FLOATING
C4613 S.n4178 SUB 0.14fF $ **FLOATING
C4614 S.t561 SUB 0.02fF
C4615 S.n4180 SUB 0.24fF $ **FLOATING
C4616 S.n4181 SUB 0.90fF $ **FLOATING
C4617 S.n4182 SUB 0.05fF $ **FLOATING
C4618 S.n4183 SUB 1.86fF $ **FLOATING
C4619 S.n4184 SUB 2.64fF $ **FLOATING
C4620 S.t607 SUB 0.02fF
C4621 S.n4185 SUB 0.24fF $ **FLOATING
C4622 S.n4186 SUB 0.35fF $ **FLOATING
C4623 S.n4187 SUB 0.60fF $ **FLOATING
C4624 S.n4188 SUB 0.12fF $ **FLOATING
C4625 S.t325 SUB 0.02fF
C4626 S.n4189 SUB 0.14fF $ **FLOATING
C4627 S.n4191 SUB 4.84fF $ **FLOATING
C4628 S.t360 SUB 0.02fF
C4629 S.n4192 SUB 0.12fF $ **FLOATING
C4630 S.n4193 SUB 0.14fF $ **FLOATING
C4631 S.t169 SUB 0.02fF
C4632 S.n4195 SUB 0.24fF $ **FLOATING
C4633 S.n4196 SUB 0.90fF $ **FLOATING
C4634 S.n4197 SUB 0.05fF $ **FLOATING
C4635 S.n4198 SUB 1.86fF $ **FLOATING
C4636 S.n4199 SUB 2.64fF $ **FLOATING
C4637 S.t1024 SUB 0.02fF
C4638 S.n4200 SUB 0.24fF $ **FLOATING
C4639 S.n4201 SUB 0.35fF $ **FLOATING
C4640 S.n4202 SUB 0.60fF $ **FLOATING
C4641 S.n4203 SUB 0.12fF $ **FLOATING
C4642 S.t462 SUB 0.02fF
C4643 S.n4204 SUB 0.14fF $ **FLOATING
C4644 S.n4206 SUB 1.86fF $ **FLOATING
C4645 S.n4207 SUB 2.65fF $ **FLOATING
C4646 S.t821 SUB 0.02fF
C4647 S.n4208 SUB 0.24fF $ **FLOATING
C4648 S.n4209 SUB 0.35fF $ **FLOATING
C4649 S.n4210 SUB 0.60fF $ **FLOATING
C4650 S.t305 SUB 0.02fF
C4651 S.n4211 SUB 1.20fF $ **FLOATING
C4652 S.n4212 SUB 0.60fF $ **FLOATING
C4653 S.n4213 SUB 0.35fF $ **FLOATING
C4654 S.n4214 SUB 0.62fF $ **FLOATING
C4655 S.n4215 SUB 1.14fF $ **FLOATING
C4656 S.n4216 SUB 2.18fF $ **FLOATING
C4657 S.n4217 SUB 0.59fF $ **FLOATING
C4658 S.n4218 SUB 0.02fF $ **FLOATING
C4659 S.n4219 SUB 0.96fF $ **FLOATING
C4660 S.t85 SUB 14.50fF
C4661 S.n4220 SUB 14.37fF $ **FLOATING
C4662 S.n4222 SUB 0.37fF $ **FLOATING
C4663 S.n4223 SUB 0.23fF $ **FLOATING
C4664 S.n4224 SUB 2.86fF $ **FLOATING
C4665 S.n4225 SUB 2.43fF $ **FLOATING
C4666 S.n4226 SUB 2.50fF $ **FLOATING
C4667 S.n4227 SUB 3.90fF $ **FLOATING
C4668 S.n4228 SUB 0.25fF $ **FLOATING
C4669 S.n4229 SUB 0.01fF $ **FLOATING
C4670 S.t191 SUB 0.02fF
C4671 S.n4230 SUB 0.25fF $ **FLOATING
C4672 S.t1042 SUB 0.02fF
C4673 S.n4231 SUB 0.94fF $ **FLOATING
C4674 S.n4232 SUB 0.70fF $ **FLOATING
C4675 S.n4233 SUB 1.86fF $ **FLOATING
C4676 S.n4234 SUB 0.47fF $ **FLOATING
C4677 S.n4235 SUB 0.09fF $ **FLOATING
C4678 S.n4236 SUB 0.32fF $ **FLOATING
C4679 S.n4237 SUB 0.30fF $ **FLOATING
C4680 S.n4238 SUB 0.76fF $ **FLOATING
C4681 S.n4239 SUB 0.58fF $ **FLOATING
C4682 S.t1034 SUB 0.02fF
C4683 S.n4240 SUB 0.24fF $ **FLOATING
C4684 S.n4241 SUB 0.35fF $ **FLOATING
C4685 S.n4242 SUB 0.60fF $ **FLOATING
C4686 S.n4243 SUB 0.12fF $ **FLOATING
C4687 S.t982 SUB 0.02fF
C4688 S.n4244 SUB 0.14fF $ **FLOATING
C4689 S.n4246 SUB 1.42fF $ **FLOATING
C4690 S.n4247 SUB 2.13fF $ **FLOATING
C4691 S.t666 SUB 0.02fF
C4692 S.n4248 SUB 0.24fF $ **FLOATING
C4693 S.n4249 SUB 0.90fF $ **FLOATING
C4694 S.n4250 SUB 0.05fF $ **FLOATING
C4695 S.t155 SUB 0.02fF
C4696 S.n4251 SUB 0.12fF $ **FLOATING
C4697 S.n4252 SUB 0.14fF $ **FLOATING
C4698 S.n4254 SUB 0.77fF $ **FLOATING
C4699 S.n4255 SUB 2.27fF $ **FLOATING
C4700 S.n4256 SUB 1.86fF $ **FLOATING
C4701 S.n4257 SUB 0.12fF $ **FLOATING
C4702 S.t875 SUB 0.02fF
C4703 S.n4258 SUB 0.14fF $ **FLOATING
C4704 S.t560 SUB 0.02fF
C4705 S.n4260 SUB 0.24fF $ **FLOATING
C4706 S.n4261 SUB 0.35fF $ **FLOATING
C4707 S.n4262 SUB 0.60fF $ **FLOATING
C4708 S.n4263 SUB 1.37fF $ **FLOATING
C4709 S.n4264 SUB 0.70fF $ **FLOATING
C4710 S.n4265 SUB 1.13fF $ **FLOATING
C4711 S.n4266 SUB 0.35fF $ **FLOATING
C4712 S.n4267 SUB 2.00fF $ **FLOATING
C4713 S.t248 SUB 0.02fF
C4714 S.n4268 SUB 0.24fF $ **FLOATING
C4715 S.n4269 SUB 0.90fF $ **FLOATING
C4716 S.n4270 SUB 0.05fF $ **FLOATING
C4717 S.t884 SUB 0.02fF
C4718 S.n4271 SUB 0.12fF $ **FLOATING
C4719 S.n4272 SUB 0.14fF $ **FLOATING
C4720 S.n4274 SUB 1.87fF $ **FLOATING
C4721 S.n4275 SUB 1.86fF $ **FLOATING
C4722 S.t168 SUB 0.02fF
C4723 S.n4276 SUB 0.24fF $ **FLOATING
C4724 S.n4277 SUB 0.35fF $ **FLOATING
C4725 S.n4278 SUB 0.60fF $ **FLOATING
C4726 S.n4279 SUB 0.12fF $ **FLOATING
C4727 S.t497 SUB 0.02fF
C4728 S.n4280 SUB 0.14fF $ **FLOATING
C4729 S.n4282 SUB 1.14fF $ **FLOATING
C4730 S.n4283 SUB 0.22fF $ **FLOATING
C4731 S.n4284 SUB 0.25fF $ **FLOATING
C4732 S.n4285 SUB 0.09fF $ **FLOATING
C4733 S.n4286 SUB 1.86fF $ **FLOATING
C4734 S.t972 SUB 0.02fF
C4735 S.n4287 SUB 0.24fF $ **FLOATING
C4736 S.n4288 SUB 0.90fF $ **FLOATING
C4737 S.n4289 SUB 0.05fF $ **FLOATING
C4738 S.t785 SUB 0.02fF
C4739 S.n4290 SUB 0.12fF $ **FLOATING
C4740 S.n4291 SUB 0.14fF $ **FLOATING
C4741 S.n4293 SUB 14.09fF $ **FLOATING
C4742 S.n4294 SUB 1.86fF $ **FLOATING
C4743 S.n4295 SUB 2.64fF $ **FLOATING
C4744 S.t128 SUB 0.02fF
C4745 S.n4296 SUB 0.24fF $ **FLOATING
C4746 S.n4297 SUB 0.35fF $ **FLOATING
C4747 S.n4298 SUB 0.60fF $ **FLOATING
C4748 S.n4299 SUB 0.12fF $ **FLOATING
C4749 S.t464 SUB 0.02fF
C4750 S.n4300 SUB 0.14fF $ **FLOATING
C4751 S.n4302 SUB 2.77fF $ **FLOATING
C4752 S.n4303 SUB 2.28fF $ **FLOATING
C4753 S.t731 SUB 0.02fF
C4754 S.n4304 SUB 0.12fF $ **FLOATING
C4755 S.n4305 SUB 0.14fF $ **FLOATING
C4756 S.t920 SUB 0.02fF
C4757 S.n4307 SUB 0.24fF $ **FLOATING
C4758 S.n4308 SUB 0.90fF $ **FLOATING
C4759 S.n4309 SUB 0.05fF $ **FLOATING
C4760 S.n4310 SUB 1.86fF $ **FLOATING
C4761 S.n4311 SUB 2.64fF $ **FLOATING
C4762 S.t858 SUB 0.02fF
C4763 S.n4312 SUB 0.24fF $ **FLOATING
C4764 S.n4313 SUB 0.35fF $ **FLOATING
C4765 S.n4314 SUB 0.60fF $ **FLOATING
C4766 S.n4315 SUB 0.12fF $ **FLOATING
C4767 S.t58 SUB 0.02fF
C4768 S.n4316 SUB 0.14fF $ **FLOATING
C4769 S.n4318 SUB 2.77fF $ **FLOATING
C4770 S.n4319 SUB 2.28fF $ **FLOATING
C4771 S.t434 SUB 0.02fF
C4772 S.n4320 SUB 0.12fF $ **FLOATING
C4773 S.n4321 SUB 0.14fF $ **FLOATING
C4774 S.t543 SUB 0.02fF
C4775 S.n4323 SUB 0.24fF $ **FLOATING
C4776 S.n4324 SUB 0.90fF $ **FLOATING
C4777 S.n4325 SUB 0.05fF $ **FLOATING
C4778 S.n4326 SUB 1.86fF $ **FLOATING
C4779 S.n4327 SUB 2.64fF $ **FLOATING
C4780 S.t86 SUB 0.02fF
C4781 S.n4328 SUB 0.24fF $ **FLOATING
C4782 S.n4329 SUB 0.35fF $ **FLOATING
C4783 S.n4330 SUB 0.60fF $ **FLOATING
C4784 S.n4331 SUB 0.12fF $ **FLOATING
C4785 S.t421 SUB 0.02fF
C4786 S.n4332 SUB 0.14fF $ **FLOATING
C4787 S.n4334 SUB 2.77fF $ **FLOATING
C4788 S.n4335 SUB 2.28fF $ **FLOATING
C4789 S.t759 SUB 0.02fF
C4790 S.n4336 SUB 0.12fF $ **FLOATING
C4791 S.n4337 SUB 0.14fF $ **FLOATING
C4792 S.t882 SUB 0.02fF
C4793 S.n4339 SUB 0.24fF $ **FLOATING
C4794 S.n4340 SUB 0.90fF $ **FLOATING
C4795 S.n4341 SUB 0.05fF $ **FLOATING
C4796 S.n4342 SUB 2.70fF $ **FLOATING
C4797 S.n4343 SUB 1.58fF $ **FLOATING
C4798 S.n4344 SUB 0.12fF $ **FLOATING
C4799 S.t660 SUB 0.02fF
C4800 S.n4345 SUB 0.14fF $ **FLOATING
C4801 S.t94 SUB 0.02fF
C4802 S.n4347 SUB 0.24fF $ **FLOATING
C4803 S.n4348 SUB 0.35fF $ **FLOATING
C4804 S.n4349 SUB 0.60fF $ **FLOATING
C4805 S.n4350 SUB 0.07fF $ **FLOATING
C4806 S.n4351 SUB 0.01fF $ **FLOATING
C4807 S.n4352 SUB 0.23fF $ **FLOATING
C4808 S.n4353 SUB 1.15fF $ **FLOATING
C4809 S.n4354 SUB 1.33fF $ **FLOATING
C4810 S.n4355 SUB 2.28fF $ **FLOATING
C4811 S.t1006 SUB 0.02fF
C4812 S.n4356 SUB 0.12fF $ **FLOATING
C4813 S.n4357 SUB 0.14fF $ **FLOATING
C4814 S.t535 SUB 0.02fF
C4815 S.n4359 SUB 0.24fF $ **FLOATING
C4816 S.n4360 SUB 0.90fF $ **FLOATING
C4817 S.n4361 SUB 0.05fF $ **FLOATING
C4818 S.n4362 SUB 0.12fF $ **FLOATING
C4819 S.t801 SUB 0.02fF
C4820 S.n4363 SUB 0.14fF $ **FLOATING
C4821 S.t1150 SUB 0.02fF
C4822 S.n4364 SUB 0.12fF $ **FLOATING
C4823 S.n4365 SUB 0.14fF $ **FLOATING
C4824 S.n4366 SUB 2.64fF $ **FLOATING
C4825 S.n4367 SUB 1.86fF $ **FLOATING
C4826 S.n4368 SUB 2.77fF $ **FLOATING
C4827 S.n4369 SUB 0.24fF $ **FLOATING
C4828 S.t482 SUB 0.02fF
C4829 S.n4370 SUB 0.35fF $ **FLOATING
C4830 S.n4371 SUB 0.60fF $ **FLOATING
C4831 S.n4372 SUB 2.28fF $ **FLOATING
C4832 S.n4373 SUB 0.24fF $ **FLOATING
C4833 S.t157 SUB 0.02fF
C4834 S.n4374 SUB 0.90fF $ **FLOATING
C4835 S.n4375 SUB 0.05fF $ **FLOATING
C4836 S.t57 SUB 32.35fF
C4837 S.t506 SUB 0.02fF
C4838 S.n4376 SUB 0.24fF $ **FLOATING
C4839 S.n4377 SUB 0.90fF $ **FLOATING
C4840 S.n4378 SUB 0.05fF $ **FLOATING
C4841 S.t376 SUB 0.02fF
C4842 S.n4379 SUB 0.12fF $ **FLOATING
C4843 S.n4380 SUB 0.14fF $ **FLOATING
C4844 S.n4382 SUB 0.12fF $ **FLOATING
C4845 S.t1139 SUB 0.02fF
C4846 S.n4383 SUB 0.14fF $ **FLOATING
C4847 S.n4385 SUB 5.11fF $ **FLOATING
C4848 S.n4386 SUB 5.38fF $ **FLOATING
C4849 S.t1086 SUB 0.02fF
C4850 S.n4387 SUB 0.12fF $ **FLOATING
C4851 S.n4388 SUB 0.14fF $ **FLOATING
C4852 S.t739 SUB 0.02fF
C4853 S.n4390 SUB 0.24fF $ **FLOATING
C4854 S.n4391 SUB 0.90fF $ **FLOATING
C4855 S.n4392 SUB 0.05fF $ **FLOATING
C4856 S.t54 SUB 31.97fF
C4857 S.t203 SUB 0.02fF
C4858 S.n4393 SUB 1.18fF $ **FLOATING
C4859 S.n4394 SUB 0.05fF $ **FLOATING
C4860 S.t120 SUB 0.02fF
C4861 S.n4395 SUB 0.01fF $ **FLOATING
C4862 S.n4396 SUB 0.25fF $ **FLOATING
C4863 S.n4398 SUB 1.48fF $ **FLOATING
C4864 S.n4399 SUB 1.29fF $ **FLOATING
C4865 S.n4400 SUB 0.27fF $ **FLOATING
C4866 S.n4401 SUB 0.24fF $ **FLOATING
C4867 S.n4402 SUB 4.34fF $ **FLOATING
C4868 S.n4403 SUB 0.02fF $ **FLOATING
C4869 S.n4404 SUB 0.03fF $ **FLOATING
C4870 S.n4405 SUB 0.24fF $ **FLOATING
C4871 S.n4406 SUB 0.13fF $ **FLOATING
C4872 S.n4407 SUB 0.56fF $ **FLOATING
C4873 S.n4408 SUB 0.03fF $ **FLOATING
C4874 S.n4409 SUB 0.85fF $ **FLOATING
C4875 S.n4410 SUB 0.22fF $ **FLOATING
C4876 S.n4411 SUB 0.14fF $ **FLOATING
C4877 S.n4412 SUB 8.87fF $ **FLOATING
C4878 S.n4413 SUB 8.87fF $ **FLOATING
C4879 S.n4414 SUB 0.59fF $ **FLOATING
C4880 S.n4415 SUB 0.21fF $ **FLOATING
C4881 S.n4416 SUB 0.59fF $ **FLOATING
C4882 S.n4417 SUB 2.57fF $ **FLOATING
C4883 S.n4418 SUB 0.29fF $ **FLOATING
C4884 S.t126 SUB 14.50fF
C4885 S.n4419 SUB 15.77fF $ **FLOATING
C4886 S.n4420 SUB 0.76fF $ **FLOATING
C4887 S.n4421 SUB 0.27fF $ **FLOATING
C4888 S.n4422 SUB 3.96fF $ **FLOATING
C4889 S.n4423 SUB 1.13fF $ **FLOATING
C4890 S.t266 SUB 0.02fF
C4891 S.n4424 SUB 0.63fF $ **FLOATING
C4892 S.n4425 SUB 0.60fF $ **FLOATING
C4893 S.n4426 SUB 0.25fF $ **FLOATING
C4894 S.n4427 SUB 0.09fF $ **FLOATING
C4895 S.n4428 SUB 0.21fF $ **FLOATING
C4896 S.n4429 SUB 1.27fF $ **FLOATING
C4897 S.n4430 SUB 0.52fF $ **FLOATING
C4898 S.n4431 SUB 1.86fF $ **FLOATING
C4899 S.n4432 SUB 0.12fF $ **FLOATING
C4900 S.t1105 SUB 0.02fF
C4901 S.n4433 SUB 0.14fF $ **FLOATING
C4902 S.t273 SUB 0.02fF
C4903 S.n4435 SUB 0.24fF $ **FLOATING
C4904 S.n4436 SUB 0.35fF $ **FLOATING
C4905 S.n4437 SUB 0.60fF $ **FLOATING
C4906 S.n4438 SUB 1.56fF $ **FLOATING
C4907 S.n4439 SUB 2.42fF $ **FLOATING
C4908 S.t714 SUB 0.02fF
C4909 S.n4440 SUB 0.24fF $ **FLOATING
C4910 S.n4441 SUB 0.90fF $ **FLOATING
C4911 S.n4442 SUB 0.05fF $ **FLOATING
C4912 S.t96 SUB 0.02fF
C4913 S.n4443 SUB 0.12fF $ **FLOATING
C4914 S.n4444 SUB 0.14fF $ **FLOATING
C4915 S.n4446 SUB 1.87fF $ **FLOATING
C4916 S.n4447 SUB 0.06fF $ **FLOATING
C4917 S.n4448 SUB 0.03fF $ **FLOATING
C4918 S.n4449 SUB 0.03fF $ **FLOATING
C4919 S.n4450 SUB 0.98fF $ **FLOATING
C4920 S.n4451 SUB 0.02fF $ **FLOATING
C4921 S.n4452 SUB 0.01fF $ **FLOATING
C4922 S.n4453 SUB 0.02fF $ **FLOATING
C4923 S.n4454 SUB 0.08fF $ **FLOATING
C4924 S.n4455 SUB 0.36fF $ **FLOATING
C4925 S.n4456 SUB 1.83fF $ **FLOATING
C4926 S.t639 SUB 0.02fF
C4927 S.n4457 SUB 0.24fF $ **FLOATING
C4928 S.n4458 SUB 0.35fF $ **FLOATING
C4929 S.n4459 SUB 0.60fF $ **FLOATING
C4930 S.n4460 SUB 0.12fF $ **FLOATING
C4931 S.t359 SUB 0.02fF
C4932 S.n4461 SUB 0.14fF $ **FLOATING
C4933 S.n4463 SUB 0.69fF $ **FLOATING
C4934 S.n4464 SUB 0.22fF $ **FLOATING
C4935 S.n4465 SUB 0.22fF $ **FLOATING
C4936 S.n4466 SUB 0.69fF $ **FLOATING
C4937 S.n4467 SUB 1.14fF $ **FLOATING
C4938 S.n4468 SUB 0.22fF $ **FLOATING
C4939 S.n4469 SUB 0.25fF $ **FLOATING
C4940 S.n4470 SUB 0.09fF $ **FLOATING
C4941 S.n4471 SUB 1.86fF $ **FLOATING
C4942 S.t205 SUB 0.02fF
C4943 S.n4472 SUB 0.24fF $ **FLOATING
C4944 S.n4473 SUB 0.90fF $ **FLOATING
C4945 S.n4474 SUB 0.05fF $ **FLOATING
C4946 S.t472 SUB 0.02fF
C4947 S.n4475 SUB 0.12fF $ **FLOATING
C4948 S.n4476 SUB 0.14fF $ **FLOATING
C4949 S.n4478 SUB 14.09fF $ **FLOATING
C4950 S.n4479 SUB 2.36fF $ **FLOATING
C4951 S.n4480 SUB 0.45fF $ **FLOATING
C4952 S.n4481 SUB 0.22fF $ **FLOATING
C4953 S.n4482 SUB 0.38fF $ **FLOATING
C4954 S.n4483 SUB 0.16fF $ **FLOATING
C4955 S.n4484 SUB 0.28fF $ **FLOATING
C4956 S.n4485 SUB 0.21fF $ **FLOATING
C4957 S.n4486 SUB 0.30fF $ **FLOATING
C4958 S.n4487 SUB 0.20fF $ **FLOATING
C4959 S.t647 SUB 0.02fF
C4960 S.n4488 SUB 0.24fF $ **FLOATING
C4961 S.n4489 SUB 0.35fF $ **FLOATING
C4962 S.n4490 SUB 0.60fF $ **FLOATING
C4963 S.n4491 SUB 0.12fF $ **FLOATING
C4964 S.t384 SUB 0.02fF
C4965 S.n4492 SUB 0.14fF $ **FLOATING
C4966 S.n4494 SUB 0.19fF $ **FLOATING
C4967 S.n4495 SUB 1.56fF $ **FLOATING
C4968 S.n4496 SUB 2.18fF $ **FLOATING
C4969 S.n4497 SUB 0.32fF $ **FLOATING
C4970 S.n4498 SUB 2.36fF $ **FLOATING
C4971 S.t432 SUB 0.02fF
C4972 S.n4499 SUB 0.12fF $ **FLOATING
C4973 S.n4500 SUB 0.14fF $ **FLOATING
C4974 S.t1107 SUB 0.02fF
C4975 S.n4502 SUB 0.24fF $ **FLOATING
C4976 S.n4503 SUB 0.90fF $ **FLOATING
C4977 S.n4504 SUB 0.05fF $ **FLOATING
C4978 S.n4505 SUB 1.86fF $ **FLOATING
C4979 S.n4506 SUB 0.12fF $ **FLOATING
C4980 S.t117 SUB 0.02fF
C4981 S.n4507 SUB 0.14fF $ **FLOATING
C4982 S.t418 SUB 0.02fF
C4983 S.n4509 SUB 0.12fF $ **FLOATING
C4984 S.n4510 SUB 0.14fF $ **FLOATING
C4985 S.t604 SUB 0.02fF
C4986 S.n4512 SUB 0.24fF $ **FLOATING
C4987 S.n4513 SUB 0.90fF $ **FLOATING
C4988 S.n4514 SUB 0.05fF $ **FLOATING
C4989 S.t903 SUB 0.02fF
C4990 S.n4515 SUB 0.24fF $ **FLOATING
C4991 S.n4516 SUB 0.35fF $ **FLOATING
C4992 S.n4517 SUB 0.60fF $ **FLOATING
C4993 S.n4518 SUB 0.31fF $ **FLOATING
C4994 S.n4519 SUB 1.08fF $ **FLOATING
C4995 S.n4520 SUB 0.15fF $ **FLOATING
C4996 S.n4521 SUB 2.08fF $ **FLOATING
C4997 S.n4522 SUB 2.91fF $ **FLOATING
C4998 S.n4523 SUB 1.86fF $ **FLOATING
C4999 S.n4524 SUB 0.12fF $ **FLOATING
C5000 S.t1085 SUB 0.02fF
C5001 S.n4525 SUB 0.14fF $ **FLOATING
C5002 S.t253 SUB 0.02fF
C5003 S.n4527 SUB 0.24fF $ **FLOATING
C5004 S.n4528 SUB 0.35fF $ **FLOATING
C5005 S.n4529 SUB 0.60fF $ **FLOATING
C5006 S.n4530 SUB 0.91fF $ **FLOATING
C5007 S.n4531 SUB 0.31fF $ **FLOATING
C5008 S.n4532 SUB 0.91fF $ **FLOATING
C5009 S.n4533 SUB 1.08fF $ **FLOATING
C5010 S.n4534 SUB 0.15fF $ **FLOATING
C5011 S.n4535 SUB 4.90fF $ **FLOATING
C5012 S.t72 SUB 0.02fF
C5013 S.n4536 SUB 0.12fF $ **FLOATING
C5014 S.n4537 SUB 0.14fF $ **FLOATING
C5015 S.t928 SUB 0.02fF
C5016 S.n4539 SUB 0.24fF $ **FLOATING
C5017 S.n4540 SUB 0.90fF $ **FLOATING
C5018 S.n4541 SUB 0.05fF $ **FLOATING
C5019 S.n4542 SUB 1.86fF $ **FLOATING
C5020 S.n4543 SUB 2.64fF $ **FLOATING
C5021 S.t976 SUB 0.02fF
C5022 S.n4544 SUB 0.24fF $ **FLOATING
C5023 S.n4545 SUB 0.35fF $ **FLOATING
C5024 S.n4546 SUB 0.60fF $ **FLOATING
C5025 S.n4547 SUB 0.12fF $ **FLOATING
C5026 S.t699 SUB 0.02fF
C5027 S.n4548 SUB 0.14fF $ **FLOATING
C5028 S.n4550 SUB 1.86fF $ **FLOATING
C5029 S.n4551 SUB 2.64fF $ **FLOATING
C5030 S.t528 SUB 0.02fF
C5031 S.n4552 SUB 0.24fF $ **FLOATING
C5032 S.n4553 SUB 0.35fF $ **FLOATING
C5033 S.n4554 SUB 0.60fF $ **FLOATING
C5034 S.t213 SUB 0.02fF
C5035 S.n4555 SUB 0.24fF $ **FLOATING
C5036 S.n4556 SUB 0.90fF $ **FLOATING
C5037 S.n4557 SUB 0.05fF $ **FLOATING
C5038 S.t1137 SUB 0.02fF
C5039 S.n4558 SUB 0.12fF $ **FLOATING
C5040 S.n4559 SUB 0.14fF $ **FLOATING
C5041 S.n4561 SUB 0.12fF $ **FLOATING
C5042 S.t852 SUB 0.02fF
C5043 S.n4562 SUB 0.14fF $ **FLOATING
C5044 S.n4564 SUB 2.28fF $ **FLOATING
C5045 S.n4565 SUB 2.91fF $ **FLOATING
C5046 S.n4566 SUB 5.10fF $ **FLOATING
C5047 S.t810 SUB 0.02fF
C5048 S.n4567 SUB 0.12fF $ **FLOATING
C5049 S.n4568 SUB 0.14fF $ **FLOATING
C5050 S.t549 SUB 0.02fF
C5051 S.n4570 SUB 0.24fF $ **FLOATING
C5052 S.n4571 SUB 0.90fF $ **FLOATING
C5053 S.n4572 SUB 0.05fF $ **FLOATING
C5054 S.n4573 SUB 1.86fF $ **FLOATING
C5055 S.n4574 SUB 2.64fF $ **FLOATING
C5056 S.t601 SUB 0.02fF
C5057 S.n4575 SUB 0.24fF $ **FLOATING
C5058 S.n4576 SUB 0.35fF $ **FLOATING
C5059 S.n4577 SUB 0.60fF $ **FLOATING
C5060 S.n4578 SUB 0.12fF $ **FLOATING
C5061 S.t319 SUB 0.02fF
C5062 S.n4579 SUB 0.14fF $ **FLOATING
C5063 S.n4581 SUB 5.11fF $ **FLOATING
C5064 S.t430 SUB 0.02fF
C5065 S.n4582 SUB 0.12fF $ **FLOATING
C5066 S.n4583 SUB 0.14fF $ **FLOATING
C5067 S.t159 SUB 0.02fF
C5068 S.n4585 SUB 0.24fF $ **FLOATING
C5069 S.n4586 SUB 0.90fF $ **FLOATING
C5070 S.n4587 SUB 0.05fF $ **FLOATING
C5071 S.n4588 SUB 1.86fF $ **FLOATING
C5072 S.n4589 SUB 2.64fF $ **FLOATING
C5073 S.t276 SUB 0.02fF
C5074 S.n4590 SUB 0.24fF $ **FLOATING
C5075 S.n4591 SUB 0.35fF $ **FLOATING
C5076 S.n4592 SUB 0.60fF $ **FLOATING
C5077 S.n4593 SUB 0.12fF $ **FLOATING
C5078 S.t1103 SUB 0.02fF
C5079 S.n4594 SUB 0.14fF $ **FLOATING
C5080 S.n4596 SUB 5.11fF $ **FLOATING
C5081 S.t1149 SUB 0.02fF
C5082 S.n4597 SUB 0.12fF $ **FLOATING
C5083 S.n4598 SUB 0.14fF $ **FLOATING
C5084 S.t958 SUB 0.02fF
C5085 S.n4600 SUB 0.24fF $ **FLOATING
C5086 S.n4601 SUB 0.90fF $ **FLOATING
C5087 S.n4602 SUB 0.05fF $ **FLOATING
C5088 S.n4603 SUB 1.86fF $ **FLOATING
C5089 S.n4604 SUB 2.65fF $ **FLOATING
C5090 S.t994 SUB 0.02fF
C5091 S.n4605 SUB 0.24fF $ **FLOATING
C5092 S.n4606 SUB 0.35fF $ **FLOATING
C5093 S.n4607 SUB 0.60fF $ **FLOATING
C5094 S.n4608 SUB 0.12fF $ **FLOATING
C5095 S.t715 SUB 0.02fF
C5096 S.n4609 SUB 0.14fF $ **FLOATING
C5097 S.n4611 SUB 5.12fF $ **FLOATING
C5098 S.t760 SUB 0.02fF
C5099 S.n4612 SUB 0.12fF $ **FLOATING
C5100 S.n4613 SUB 0.14fF $ **FLOATING
C5101 S.t576 SUB 0.02fF
C5102 S.n4615 SUB 0.24fF $ **FLOATING
C5103 S.n4616 SUB 0.90fF $ **FLOATING
C5104 S.n4617 SUB 0.05fF $ **FLOATING
C5105 S.n4618 SUB 1.86fF $ **FLOATING
C5106 S.n4619 SUB 2.64fF $ **FLOATING
C5107 S.t621 SUB 0.02fF
C5108 S.n4620 SUB 0.24fF $ **FLOATING
C5109 S.n4621 SUB 0.35fF $ **FLOATING
C5110 S.n4622 SUB 0.60fF $ **FLOATING
C5111 S.n4623 SUB 0.12fF $ **FLOATING
C5112 S.t333 SUB 0.02fF
C5113 S.n4624 SUB 0.14fF $ **FLOATING
C5114 S.n4626 SUB 5.11fF $ **FLOATING
C5115 S.t375 SUB 0.02fF
C5116 S.n4627 SUB 0.12fF $ **FLOATING
C5117 S.n4628 SUB 0.14fF $ **FLOATING
C5118 S.t182 SUB 0.02fF
C5119 S.n4630 SUB 0.24fF $ **FLOATING
C5120 S.n4631 SUB 0.90fF $ **FLOATING
C5121 S.n4632 SUB 0.05fF $ **FLOATING
C5122 S.n4633 SUB 1.86fF $ **FLOATING
C5123 S.n4634 SUB 2.64fF $ **FLOATING
C5124 S.t233 SUB 0.02fF
C5125 S.n4635 SUB 0.24fF $ **FLOATING
C5126 S.n4636 SUB 0.35fF $ **FLOATING
C5127 S.n4637 SUB 0.60fF $ **FLOATING
C5128 S.n4638 SUB 0.12fF $ **FLOATING
C5129 S.t1062 SUB 0.02fF
C5130 S.n4639 SUB 0.14fF $ **FLOATING
C5131 S.n4641 SUB 4.84fF $ **FLOATING
C5132 S.t1098 SUB 0.02fF
C5133 S.n4642 SUB 0.12fF $ **FLOATING
C5134 S.n4643 SUB 0.14fF $ **FLOATING
C5135 S.t904 SUB 0.02fF
C5136 S.n4645 SUB 0.24fF $ **FLOATING
C5137 S.n4646 SUB 0.90fF $ **FLOATING
C5138 S.n4647 SUB 0.05fF $ **FLOATING
C5139 S.n4648 SUB 1.86fF $ **FLOATING
C5140 S.n4649 SUB 2.64fF $ **FLOATING
C5141 S.t414 SUB 0.02fF
C5142 S.n4650 SUB 0.24fF $ **FLOATING
C5143 S.n4651 SUB 0.35fF $ **FLOATING
C5144 S.n4652 SUB 0.60fF $ **FLOATING
C5145 S.n4653 SUB 0.12fF $ **FLOATING
C5146 S.t977 SUB 0.02fF
C5147 S.n4654 SUB 0.14fF $ **FLOATING
C5148 S.n4656 SUB 1.86fF $ **FLOATING
C5149 S.n4657 SUB 2.65fF $ **FLOATING
C5150 S.t458 SUB 0.02fF
C5151 S.n4658 SUB 0.24fF $ **FLOATING
C5152 S.n4659 SUB 0.35fF $ **FLOATING
C5153 S.n4660 SUB 0.60fF $ **FLOATING
C5154 S.t188 SUB 0.02fF
C5155 S.n4661 SUB 1.20fF $ **FLOATING
C5156 S.n4662 SUB 0.41fF $ **FLOATING
C5157 S.n4663 SUB 0.44fF $ **FLOATING
C5158 S.n4664 SUB 0.36fF $ **FLOATING
C5159 S.n4665 SUB 0.20fF $ **FLOATING
C5160 S.n4666 SUB 0.25fF $ **FLOATING
C5161 S.n4667 SUB 1.27fF $ **FLOATING
C5162 S.n4668 SUB 0.35fF $ **FLOATING
C5163 S.n4669 SUB 0.62fF $ **FLOATING
C5164 S.n4670 SUB 1.14fF $ **FLOATING
C5165 S.n4671 SUB 2.18fF $ **FLOATING
C5166 S.n4672 SUB 0.59fF $ **FLOATING
C5167 S.n4673 SUB 0.02fF $ **FLOATING
C5168 S.n4674 SUB 0.96fF $ **FLOATING
C5169 S.t100 SUB 14.50fF
C5170 S.n4675 SUB 14.37fF $ **FLOATING
C5171 S.n4677 SUB 0.37fF $ **FLOATING
C5172 S.n4678 SUB 0.23fF $ **FLOATING
C5173 S.n4679 SUB 2.79fF $ **FLOATING
C5174 S.n4680 SUB 1.98fF $ **FLOATING
C5175 S.n4681 SUB 4.03fF $ **FLOATING
C5176 S.n4682 SUB 0.25fF $ **FLOATING
C5177 S.n4683 SUB 0.01fF $ **FLOATING
C5178 S.t37 SUB 0.02fF
C5179 S.n4684 SUB 0.25fF $ **FLOATING
C5180 S.t932 SUB 0.02fF
C5181 S.n4685 SUB 0.94fF $ **FLOATING
C5182 S.n4686 SUB 0.70fF $ **FLOATING
C5183 S.n4687 SUB 0.77fF $ **FLOATING
C5184 S.n4688 SUB 2.24fF $ **FLOATING
C5185 S.n4689 SUB 1.86fF $ **FLOATING
C5186 S.n4690 SUB 0.12fF $ **FLOATING
C5187 S.t844 SUB 0.02fF
C5188 S.n4691 SUB 0.14fF $ **FLOATING
C5189 S.t911 SUB 0.02fF
C5190 S.n4693 SUB 0.24fF $ **FLOATING
C5191 S.n4694 SUB 0.35fF $ **FLOATING
C5192 S.n4695 SUB 0.60fF $ **FLOATING
C5193 S.n4696 SUB 1.37fF $ **FLOATING
C5194 S.n4697 SUB 0.70fF $ **FLOATING
C5195 S.n4698 SUB 1.13fF $ **FLOATING
C5196 S.n4699 SUB 0.35fF $ **FLOATING
C5197 S.n4700 SUB 2.00fF $ **FLOATING
C5198 S.t554 SUB 0.02fF
C5199 S.n4701 SUB 0.24fF $ **FLOATING
C5200 S.n4702 SUB 0.90fF $ **FLOATING
C5201 S.n4703 SUB 0.05fF $ **FLOATING
C5202 S.t1127 SUB 0.02fF
C5203 S.n4704 SUB 0.12fF $ **FLOATING
C5204 S.n4705 SUB 0.14fF $ **FLOATING
C5205 S.n4707 SUB 1.87fF $ **FLOATING
C5206 S.n4708 SUB 1.86fF $ **FLOATING
C5207 S.t180 SUB 0.02fF
C5208 S.n4709 SUB 0.24fF $ **FLOATING
C5209 S.n4710 SUB 0.35fF $ **FLOATING
C5210 S.n4711 SUB 0.60fF $ **FLOATING
C5211 S.n4712 SUB 0.12fF $ **FLOATING
C5212 S.t510 SUB 0.02fF
C5213 S.n4713 SUB 0.14fF $ **FLOATING
C5214 S.n4715 SUB 1.14fF $ **FLOATING
C5215 S.n4716 SUB 0.22fF $ **FLOATING
C5216 S.n4717 SUB 0.25fF $ **FLOATING
C5217 S.n4718 SUB 0.09fF $ **FLOATING
C5218 S.n4719 SUB 1.86fF $ **FLOATING
C5219 S.t981 SUB 0.02fF
C5220 S.n4720 SUB 0.24fF $ **FLOATING
C5221 S.n4721 SUB 0.90fF $ **FLOATING
C5222 S.n4722 SUB 0.05fF $ **FLOATING
C5223 S.t743 SUB 0.02fF
C5224 S.n4723 SUB 0.12fF $ **FLOATING
C5225 S.n4724 SUB 0.14fF $ **FLOATING
C5226 S.n4726 SUB 14.09fF $ **FLOATING
C5227 S.n4727 SUB 1.86fF $ **FLOATING
C5228 S.n4728 SUB 2.64fF $ **FLOATING
C5229 S.t143 SUB 0.02fF
C5230 S.n4729 SUB 0.24fF $ **FLOATING
C5231 S.n4730 SUB 0.35fF $ **FLOATING
C5232 S.n4731 SUB 0.60fF $ **FLOATING
C5233 S.n4732 SUB 0.12fF $ **FLOATING
C5234 S.t476 SUB 0.02fF
C5235 S.n4733 SUB 0.14fF $ **FLOATING
C5236 S.n4735 SUB 2.77fF $ **FLOATING
C5237 S.n4736 SUB 2.28fF $ **FLOATING
C5238 S.t749 SUB 0.02fF
C5239 S.n4737 SUB 0.12fF $ **FLOATING
C5240 S.n4738 SUB 0.14fF $ **FLOATING
C5241 S.t939 SUB 0.02fF
C5242 S.n4740 SUB 0.24fF $ **FLOATING
C5243 S.n4741 SUB 0.90fF $ **FLOATING
C5244 S.n4742 SUB 0.05fF $ **FLOATING
C5245 S.n4743 SUB 1.86fF $ **FLOATING
C5246 S.n4744 SUB 2.64fF $ **FLOATING
C5247 S.t868 SUB 0.02fF
C5248 S.n4745 SUB 0.24fF $ **FLOATING
C5249 S.n4746 SUB 0.35fF $ **FLOATING
C5250 S.n4747 SUB 0.60fF $ **FLOATING
C5251 S.n4748 SUB 0.12fF $ **FLOATING
C5252 S.t78 SUB 0.02fF
C5253 S.n4749 SUB 0.14fF $ **FLOATING
C5254 S.n4751 SUB 2.77fF $ **FLOATING
C5255 S.n4752 SUB 2.28fF $ **FLOATING
C5256 S.t363 SUB 0.02fF
C5257 S.n4753 SUB 0.12fF $ **FLOATING
C5258 S.n4754 SUB 0.14fF $ **FLOATING
C5259 S.t558 SUB 0.02fF
C5260 S.n4756 SUB 0.24fF $ **FLOATING
C5261 S.n4757 SUB 0.90fF $ **FLOATING
C5262 S.n4758 SUB 0.05fF $ **FLOATING
C5263 S.n4759 SUB 1.86fF $ **FLOATING
C5264 S.n4760 SUB 2.65fF $ **FLOATING
C5265 S.t491 SUB 0.02fF
C5266 S.n4761 SUB 0.24fF $ **FLOATING
C5267 S.n4762 SUB 0.35fF $ **FLOATING
C5268 S.n4763 SUB 0.60fF $ **FLOATING
C5269 S.n4764 SUB 0.12fF $ **FLOATING
C5270 S.t813 SUB 0.02fF
C5271 S.n4765 SUB 0.14fF $ **FLOATING
C5272 S.n4767 SUB 2.77fF $ **FLOATING
C5273 S.n4768 SUB 2.28fF $ **FLOATING
C5274 S.t28 SUB 0.02fF
C5275 S.n4769 SUB 0.12fF $ **FLOATING
C5276 S.n4770 SUB 0.14fF $ **FLOATING
C5277 S.t167 SUB 0.02fF
C5278 S.n4772 SUB 0.24fF $ **FLOATING
C5279 S.n4773 SUB 0.90fF $ **FLOATING
C5280 S.n4774 SUB 0.05fF $ **FLOATING
C5281 S.n4775 SUB 1.86fF $ **FLOATING
C5282 S.n4776 SUB 2.64fF $ **FLOATING
C5283 S.t101 SUB 0.02fF
C5284 S.n4777 SUB 0.24fF $ **FLOATING
C5285 S.n4778 SUB 0.35fF $ **FLOATING
C5286 S.n4779 SUB 0.60fF $ **FLOATING
C5287 S.n4780 SUB 0.12fF $ **FLOATING
C5288 S.t438 SUB 0.02fF
C5289 S.n4781 SUB 0.14fF $ **FLOATING
C5290 S.n4783 SUB 2.77fF $ **FLOATING
C5291 S.n4784 SUB 2.28fF $ **FLOATING
C5292 S.t778 SUB 0.02fF
C5293 S.n4785 SUB 0.12fF $ **FLOATING
C5294 S.n4786 SUB 0.14fF $ **FLOATING
C5295 S.t892 SUB 0.02fF
C5296 S.n4788 SUB 0.24fF $ **FLOATING
C5297 S.n4789 SUB 0.90fF $ **FLOATING
C5298 S.n4790 SUB 0.05fF $ **FLOATING
C5299 S.n4791 SUB 1.86fF $ **FLOATING
C5300 S.n4792 SUB 2.64fF $ **FLOATING
C5301 S.t833 SUB 0.02fF
C5302 S.n4793 SUB 0.24fF $ **FLOATING
C5303 S.n4794 SUB 0.35fF $ **FLOATING
C5304 S.n4795 SUB 0.60fF $ **FLOATING
C5305 S.n4796 SUB 0.12fF $ **FLOATING
C5306 S.t9 SUB 0.02fF
C5307 S.n4797 SUB 0.14fF $ **FLOATING
C5308 S.n4799 SUB 2.77fF $ **FLOATING
C5309 S.n4800 SUB 2.28fF $ **FLOATING
C5310 S.t393 SUB 0.02fF
C5311 S.n4801 SUB 0.12fF $ **FLOATING
C5312 S.n4802 SUB 0.14fF $ **FLOATING
C5313 S.t517 SUB 0.02fF
C5314 S.n4804 SUB 0.24fF $ **FLOATING
C5315 S.n4805 SUB 0.90fF $ **FLOATING
C5316 S.n4806 SUB 0.05fF $ **FLOATING
C5317 S.n4807 SUB 0.12fF $ **FLOATING
C5318 S.t31 SUB 0.02fF
C5319 S.n4808 SUB 0.14fF $ **FLOATING
C5320 S.t617 SUB 0.02fF
C5321 S.n4810 SUB 0.24fF $ **FLOATING
C5322 S.n4811 SUB 0.35fF $ **FLOATING
C5323 S.n4812 SUB 0.60fF $ **FLOATING
C5324 S.n4813 SUB 1.58fF $ **FLOATING
C5325 S.n4814 SUB 0.03fF $ **FLOATING
C5326 S.n4815 SUB 0.14fF $ **FLOATING
C5327 S.n4816 SUB 0.58fF $ **FLOATING
C5328 S.n4817 SUB 0.12fF $ **FLOATING
C5329 S.n4818 SUB 0.53fF $ **FLOATING
C5330 S.n4819 SUB 0.41fF $ **FLOATING
C5331 S.n4820 SUB 0.24fF $ **FLOATING
C5332 S.n4821 SUB 0.24fF $ **FLOATING
C5333 S.n4822 SUB 0.67fF $ **FLOATING
C5334 S.n4823 SUB 1.95fF $ **FLOATING
C5335 S.t373 SUB 0.02fF
C5336 S.n4824 SUB 0.12fF $ **FLOATING
C5337 S.n4825 SUB 0.14fF $ **FLOATING
C5338 S.t1029 SUB 0.02fF
C5339 S.n4827 SUB 0.24fF $ **FLOATING
C5340 S.n4828 SUB 0.90fF $ **FLOATING
C5341 S.n4829 SUB 0.05fF $ **FLOATING
C5342 S.t8 SUB 32.35fF
C5343 S.t127 SUB 0.02fF
C5344 S.n4830 SUB 0.24fF $ **FLOATING
C5345 S.n4831 SUB 0.90fF $ **FLOATING
C5346 S.n4832 SUB 0.05fF $ **FLOATING
C5347 S.t1115 SUB 0.02fF
C5348 S.n4833 SUB 0.12fF $ **FLOATING
C5349 S.n4834 SUB 0.14fF $ **FLOATING
C5350 S.n4836 SUB 0.12fF $ **FLOATING
C5351 S.t767 SUB 0.02fF
C5352 S.n4837 SUB 0.14fF $ **FLOATING
C5353 S.n4839 SUB 5.11fF $ **FLOATING
C5354 S.n4840 SUB 5.38fF $ **FLOATING
C5355 S.t709 SUB 0.02fF
C5356 S.n4841 SUB 0.12fF $ **FLOATING
C5357 S.n4842 SUB 0.14fF $ **FLOATING
C5358 S.t152 SUB 0.02fF
C5359 S.n4844 SUB 0.24fF $ **FLOATING
C5360 S.n4845 SUB 0.90fF $ **FLOATING
C5361 S.n4846 SUB 0.05fF $ **FLOATING
C5362 S.t71 SUB 31.97fF
C5363 S.t942 SUB 0.02fF
C5364 S.n4847 SUB 1.18fF $ **FLOATING
C5365 S.n4848 SUB 0.05fF $ **FLOATING
C5366 S.t650 SUB 0.02fF
C5367 S.n4849 SUB 0.01fF $ **FLOATING
C5368 S.n4850 SUB 0.25fF $ **FLOATING
C5369 S.n4852 SUB 1.48fF $ **FLOATING
C5370 S.n4853 SUB 1.24fF $ **FLOATING
C5371 S.n4854 SUB 0.27fF $ **FLOATING
C5372 S.n4855 SUB 0.24fF $ **FLOATING
C5373 S.n4856 SUB 4.34fF $ **FLOATING
C5374 S.t218 SUB 0.02fF
C5375 S.n4857 SUB 1.20fF $ **FLOATING
C5376 S.n4858 SUB 0.35fF $ **FLOATING
C5377 S.n4859 SUB 0.46fF $ **FLOATING
C5378 S.n4860 SUB 1.12fF $ **FLOATING
C5379 S.n4861 SUB 1.86fF $ **FLOATING
C5380 S.n4862 SUB 0.12fF $ **FLOATING
C5381 S.t1041 SUB 0.02fF
C5382 S.n4863 SUB 0.14fF $ **FLOATING
C5383 S.t178 SUB 0.02fF
C5384 S.n4865 SUB 0.24fF $ **FLOATING
C5385 S.n4866 SUB 0.35fF $ **FLOATING
C5386 S.n4867 SUB 0.60fF $ **FLOATING
C5387 S.n4868 SUB 2.64fF $ **FLOATING
C5388 S.n4869 SUB 3.89fF $ **FLOATING
C5389 S.t166 SUB 0.02fF
C5390 S.n4870 SUB 0.24fF $ **FLOATING
C5391 S.n4871 SUB 0.90fF $ **FLOATING
C5392 S.n4872 SUB 0.05fF $ **FLOATING
C5393 S.t1054 SUB 0.02fF
C5394 S.n4873 SUB 0.12fF $ **FLOATING
C5395 S.n4874 SUB 0.14fF $ **FLOATING
C5396 S.n4876 SUB 1.86fF $ **FLOATING
C5397 S.n4877 SUB 2.64fF $ **FLOATING
C5398 S.t572 SUB 0.02fF
C5399 S.n4878 SUB 0.24fF $ **FLOATING
C5400 S.n4879 SUB 0.35fF $ **FLOATING
C5401 S.n4880 SUB 0.60fF $ **FLOATING
C5402 S.n4881 SUB 0.12fF $ **FLOATING
C5403 S.t311 SUB 0.02fF
C5404 S.n4882 SUB 0.14fF $ **FLOATING
C5405 S.n4884 SUB 5.11fF $ **FLOATING
C5406 S.t557 SUB 0.02fF
C5407 S.n4885 SUB 0.24fF $ **FLOATING
C5408 S.n4886 SUB 0.90fF $ **FLOATING
C5409 S.n4887 SUB 0.05fF $ **FLOATING
C5410 S.t328 SUB 0.02fF
C5411 S.n4888 SUB 0.12fF $ **FLOATING
C5412 S.n4889 SUB 0.14fF $ **FLOATING
C5413 S.n4891 SUB 1.86fF $ **FLOATING
C5414 S.n4892 SUB 2.64fF $ **FLOATING
C5415 S.t957 SUB 0.02fF
C5416 S.n4893 SUB 0.24fF $ **FLOATING
C5417 S.n4894 SUB 0.35fF $ **FLOATING
C5418 S.n4895 SUB 0.60fF $ **FLOATING
C5419 S.n4896 SUB 0.12fF $ **FLOATING
C5420 S.t681 SUB 0.02fF
C5421 S.n4897 SUB 0.14fF $ **FLOATING
C5422 S.n4899 SUB 5.11fF $ **FLOATING
C5423 S.t938 SUB 0.02fF
C5424 S.n4900 SUB 0.24fF $ **FLOATING
C5425 S.n4901 SUB 0.90fF $ **FLOATING
C5426 S.n4902 SUB 0.05fF $ **FLOATING
C5427 S.t710 SUB 0.02fF
C5428 S.n4903 SUB 0.12fF $ **FLOATING
C5429 S.n4904 SUB 0.14fF $ **FLOATING
C5430 S.n4906 SUB 1.86fF $ **FLOATING
C5431 S.n4907 SUB 2.64fF $ **FLOATING
C5432 S.t230 SUB 0.02fF
C5433 S.n4908 SUB 0.24fF $ **FLOATING
C5434 S.n4909 SUB 0.35fF $ **FLOATING
C5435 S.n4910 SUB 0.60fF $ **FLOATING
C5436 S.n4911 SUB 0.12fF $ **FLOATING
C5437 S.t1061 SUB 0.02fF
C5438 S.n4912 SUB 0.14fF $ **FLOATING
C5439 S.n4914 SUB 5.11fF $ **FLOATING
C5440 S.t212 SUB 0.02fF
C5441 S.n4915 SUB 0.24fF $ **FLOATING
C5442 S.n4916 SUB 0.90fF $ **FLOATING
C5443 S.n4917 SUB 0.05fF $ **FLOATING
C5444 S.t1095 SUB 0.02fF
C5445 S.n4918 SUB 0.12fF $ **FLOATING
C5446 S.n4919 SUB 0.14fF $ **FLOATING
C5447 S.n4921 SUB 1.86fF $ **FLOATING
C5448 S.n4922 SUB 2.64fF $ **FLOATING
C5449 S.t546 SUB 0.02fF
C5450 S.n4923 SUB 0.24fF $ **FLOATING
C5451 S.n4924 SUB 0.35fF $ **FLOATING
C5452 S.n4925 SUB 0.60fF $ **FLOATING
C5453 S.n4926 SUB 0.12fF $ **FLOATING
C5454 S.t301 SUB 0.02fF
C5455 S.n4927 SUB 0.14fF $ **FLOATING
C5456 S.n4929 SUB 5.11fF $ **FLOATING
C5457 S.t534 SUB 0.02fF
C5458 S.n4930 SUB 0.24fF $ **FLOATING
C5459 S.n4931 SUB 0.90fF $ **FLOATING
C5460 S.n4932 SUB 0.05fF $ **FLOATING
C5461 S.t374 SUB 0.02fF
C5462 S.n4933 SUB 0.12fF $ **FLOATING
C5463 S.n4934 SUB 0.14fF $ **FLOATING
C5464 S.n4936 SUB 1.86fF $ **FLOATING
C5465 S.n4937 SUB 2.64fF $ **FLOATING
C5466 S.t927 SUB 0.02fF
C5467 S.n4938 SUB 0.24fF $ **FLOATING
C5468 S.n4939 SUB 0.35fF $ **FLOATING
C5469 S.n4940 SUB 0.60fF $ **FLOATING
C5470 S.n4941 SUB 0.12fF $ **FLOATING
C5471 S.t671 SUB 0.02fF
C5472 S.n4942 SUB 0.14fF $ **FLOATING
C5473 S.n4944 SUB 5.11fF $ **FLOATING
C5474 S.t909 SUB 0.02fF
C5475 S.n4945 SUB 0.24fF $ **FLOATING
C5476 S.n4946 SUB 0.90fF $ **FLOATING
C5477 S.n4947 SUB 0.05fF $ **FLOATING
C5478 S.t758 SUB 0.02fF
C5479 S.n4948 SUB 0.12fF $ **FLOATING
C5480 S.n4949 SUB 0.14fF $ **FLOATING
C5481 S.n4951 SUB 1.86fF $ **FLOATING
C5482 S.n4952 SUB 2.64fF $ **FLOATING
C5483 S.t204 SUB 0.02fF
C5484 S.n4953 SUB 0.24fF $ **FLOATING
C5485 S.n4954 SUB 0.35fF $ **FLOATING
C5486 S.n4955 SUB 0.60fF $ **FLOATING
C5487 S.n4956 SUB 0.12fF $ **FLOATING
C5488 S.t1048 SUB 0.02fF
C5489 S.n4957 SUB 0.14fF $ **FLOATING
C5490 S.n4959 SUB 5.11fF $ **FLOATING
C5491 S.t186 SUB 0.02fF
C5492 S.n4960 SUB 0.24fF $ **FLOATING
C5493 S.n4961 SUB 0.90fF $ **FLOATING
C5494 S.n4962 SUB 0.05fF $ **FLOATING
C5495 S.t1147 SUB 0.02fF
C5496 S.n4963 SUB 0.12fF $ **FLOATING
C5497 S.n4964 SUB 0.14fF $ **FLOATING
C5498 S.n4966 SUB 1.86fF $ **FLOATING
C5499 S.n4967 SUB 2.64fF $ **FLOATING
C5500 S.t600 SUB 0.02fF
C5501 S.n4968 SUB 0.24fF $ **FLOATING
C5502 S.n4969 SUB 0.35fF $ **FLOATING
C5503 S.n4970 SUB 0.60fF $ **FLOATING
C5504 S.n4971 SUB 0.12fF $ **FLOATING
C5505 S.t317 SUB 0.02fF
C5506 S.n4972 SUB 0.14fF $ **FLOATING
C5507 S.n4974 SUB 1.92fF $ **FLOATING
C5508 S.n4975 SUB 2.51fF $ **FLOATING
C5509 S.t109 SUB 0.02fF
C5510 S.n4976 SUB 0.24fF $ **FLOATING
C5511 S.n4977 SUB 0.35fF $ **FLOATING
C5512 S.n4978 SUB 0.60fF $ **FLOATING
C5513 S.t935 SUB 0.02fF
C5514 S.n4979 SUB 0.24fF $ **FLOATING
C5515 S.n4980 SUB 0.90fF $ **FLOATING
C5516 S.n4981 SUB 0.05fF $ **FLOATING
C5517 S.t1106 SUB 0.02fF
C5518 S.n4982 SUB 0.12fF $ **FLOATING
C5519 S.n4983 SUB 0.14fF $ **FLOATING
C5520 S.n4985 SUB 0.12fF $ **FLOATING
C5521 S.t842 SUB 0.02fF
C5522 S.n4986 SUB 0.14fF $ **FLOATING
C5523 S.n4988 SUB 2.28fF $ **FLOATING
C5524 S.n4989 SUB 1.75fF $ **FLOATING
C5525 S.n4990 SUB 5.10fF $ **FLOATING
C5526 S.t586 SUB 0.02fF
C5527 S.n4991 SUB 0.24fF $ **FLOATING
C5528 S.n4992 SUB 0.90fF $ **FLOATING
C5529 S.n4993 SUB 0.05fF $ **FLOATING
C5530 S.t431 SUB 0.02fF
C5531 S.n4994 SUB 0.12fF $ **FLOATING
C5532 S.n4995 SUB 0.14fF $ **FLOATING
C5533 S.n4997 SUB 1.92fF $ **FLOATING
C5534 S.n4998 SUB 0.12fF $ **FLOATING
C5535 S.t97 SUB 0.02fF
C5536 S.n4999 SUB 0.14fF $ **FLOATING
C5537 S.n5001 SUB 14.09fF $ **FLOATING
C5538 S.n5002 SUB 0.04fF $ **FLOATING
C5539 S.n5003 SUB 0.09fF $ **FLOATING
C5540 S.n5004 SUB 0.29fF $ **FLOATING
C5541 S.n5005 SUB 0.25fF $ **FLOATING
C5542 S.n5006 SUB 0.12fF $ **FLOATING
C5543 S.n5007 SUB 0.05fF $ **FLOATING
C5544 S.n5008 SUB 0.17fF $ **FLOATING
C5545 S.n5009 SUB 1.24fF $ **FLOATING
C5546 S.n5010 SUB 2.74fF $ **FLOATING
C5547 S.n5011 SUB 0.12fF $ **FLOATING
C5548 S.t1092 SUB 0.02fF
C5549 S.n5012 SUB 0.14fF $ **FLOATING
C5550 S.t369 SUB 0.02fF
C5551 S.n5014 SUB 0.24fF $ **FLOATING
C5552 S.n5015 SUB 0.35fF $ **FLOATING
C5553 S.n5016 SUB 0.60fF $ **FLOATING
C5554 S.n5017 SUB 2.59fF $ **FLOATING
C5555 S.n5018 SUB 2.03fF $ **FLOATING
C5556 S.t332 SUB 0.02fF
C5557 S.n5019 SUB 0.12fF $ **FLOATING
C5558 S.n5020 SUB 0.14fF $ **FLOATING
C5559 S.t88 SUB 0.02fF
C5560 S.n5022 SUB 0.24fF $ **FLOATING
C5561 S.n5023 SUB 0.90fF $ **FLOATING
C5562 S.n5024 SUB 0.05fF $ **FLOATING
C5563 S.t612 SUB 0.02fF
C5564 S.n5025 SUB 0.94fF $ **FLOATING
C5565 S.n5026 SUB 0.70fF $ **FLOATING
C5566 S.n5027 SUB 0.01fF $ **FLOATING
C5567 S.t433 SUB 0.02fF
C5568 S.n5028 SUB 0.25fF $ **FLOATING
C5569 S.t929 SUB 0.02fF
C5570 S.n5029 SUB 1.20fF $ **FLOATING
C5571 S.n5030 SUB 1.94fF $ **FLOATING
C5572 S.n5031 SUB 0.06fF $ **FLOATING
C5573 S.n5032 SUB 0.10fF $ **FLOATING
C5574 S.n5033 SUB 0.60fF $ **FLOATING
C5575 S.n5034 SUB 2.18fF $ **FLOATING
C5576 S.n5035 SUB 0.92fF $ **FLOATING
C5577 S.n5036 SUB 0.83fF $ **FLOATING
C5578 S.n5037 SUB 0.02fF $ **FLOATING
C5579 S.n5038 SUB 0.96fF $ **FLOATING
C5580 S.t62 SUB 14.50fF
C5581 S.n5039 SUB 14.07fF $ **FLOATING
C5582 S.n5041 SUB 1.21fF $ **FLOATING
C5583 S.n5042 SUB 1.43fF $ **FLOATING
C5584 S.n5043 SUB 2.87fF $ **FLOATING
C5585 S.n5044 SUB 2.39fF $ **FLOATING
C5586 S.n5045 SUB 3.81fF $ **FLOATING
C5587 S.n5046 SUB 0.25fF $ **FLOATING
C5588 S.n5047 SUB 1.92fF $ **FLOATING
C5589 S.n5048 SUB 2.51fF $ **FLOATING
C5590 S.t841 SUB 0.02fF
C5591 S.n5049 SUB 0.24fF $ **FLOATING
C5592 S.n5050 SUB 0.35fF $ **FLOATING
C5593 S.n5051 SUB 0.60fF $ **FLOATING
C5594 S.n5052 SUB 0.12fF $ **FLOATING
C5595 S.t466 SUB 0.02fF
C5596 S.n5053 SUB 0.14fF $ **FLOATING
C5597 S.n5055 SUB 2.39fF $ **FLOATING
C5598 S.n5056 SUB 2.28fF $ **FLOATING
C5599 S.t736 SUB 0.02fF
C5600 S.n5057 SUB 0.12fF $ **FLOATING
C5601 S.n5058 SUB 0.14fF $ **FLOATING
C5602 S.t556 SUB 0.02fF
C5603 S.n5060 SUB 0.24fF $ **FLOATING
C5604 S.n5061 SUB 0.90fF $ **FLOATING
C5605 S.n5062 SUB 0.05fF $ **FLOATING
C5606 S.n5063 SUB 1.92fF $ **FLOATING
C5607 S.n5064 SUB 2.51fF $ **FLOATING
C5608 S.t465 SUB 0.02fF
C5609 S.n5065 SUB 0.24fF $ **FLOATING
C5610 S.n5066 SUB 0.35fF $ **FLOATING
C5611 S.n5067 SUB 0.60fF $ **FLOATING
C5612 S.n5068 SUB 0.12fF $ **FLOATING
C5613 S.t65 SUB 0.02fF
C5614 S.n5069 SUB 0.14fF $ **FLOATING
C5615 S.n5071 SUB 2.39fF $ **FLOATING
C5616 S.n5072 SUB 2.28fF $ **FLOATING
C5617 S.t352 SUB 0.02fF
C5618 S.n5073 SUB 0.12fF $ **FLOATING
C5619 S.n5074 SUB 0.14fF $ **FLOATING
C5620 S.t164 SUB 0.02fF
C5621 S.n5076 SUB 0.24fF $ **FLOATING
C5622 S.n5077 SUB 0.90fF $ **FLOATING
C5623 S.n5078 SUB 0.05fF $ **FLOATING
C5624 S.n5079 SUB 1.92fF $ **FLOATING
C5625 S.n5080 SUB 2.51fF $ **FLOATING
C5626 S.t63 SUB 0.02fF
C5627 S.n5081 SUB 0.24fF $ **FLOATING
C5628 S.n5082 SUB 0.35fF $ **FLOATING
C5629 S.n5083 SUB 0.60fF $ **FLOATING
C5630 S.n5084 SUB 0.12fF $ **FLOATING
C5631 S.t806 SUB 0.02fF
C5632 S.n5085 SUB 0.14fF $ **FLOATING
C5633 S.n5087 SUB 2.39fF $ **FLOATING
C5634 S.n5088 SUB 2.28fF $ **FLOATING
C5635 S.t1076 SUB 0.02fF
C5636 S.n5089 SUB 0.12fF $ **FLOATING
C5637 S.n5090 SUB 0.14fF $ **FLOATING
C5638 S.t889 SUB 0.02fF
C5639 S.n5092 SUB 0.24fF $ **FLOATING
C5640 S.n5093 SUB 0.90fF $ **FLOATING
C5641 S.n5094 SUB 0.05fF $ **FLOATING
C5642 S.n5095 SUB 1.92fF $ **FLOATING
C5643 S.n5096 SUB 2.51fF $ **FLOATING
C5644 S.t805 SUB 0.02fF
C5645 S.n5097 SUB 0.24fF $ **FLOATING
C5646 S.n5098 SUB 0.35fF $ **FLOATING
C5647 S.n5099 SUB 0.60fF $ **FLOATING
C5648 S.n5100 SUB 0.12fF $ **FLOATING
C5649 S.t423 SUB 0.02fF
C5650 S.n5101 SUB 0.14fF $ **FLOATING
C5651 S.n5103 SUB 2.39fF $ **FLOATING
C5652 S.n5104 SUB 2.28fF $ **FLOATING
C5653 S.t695 SUB 0.02fF
C5654 S.n5105 SUB 0.12fF $ **FLOATING
C5655 S.n5106 SUB 0.14fF $ **FLOATING
C5656 S.t518 SUB 0.02fF
C5657 S.n5108 SUB 0.24fF $ **FLOATING
C5658 S.n5109 SUB 0.90fF $ **FLOATING
C5659 S.n5110 SUB 0.05fF $ **FLOATING
C5660 S.n5111 SUB 1.92fF $ **FLOATING
C5661 S.n5112 SUB 2.51fF $ **FLOATING
C5662 S.t422 SUB 0.02fF
C5663 S.n5113 SUB 0.24fF $ **FLOATING
C5664 S.n5114 SUB 0.35fF $ **FLOATING
C5665 S.n5115 SUB 0.60fF $ **FLOATING
C5666 S.n5116 SUB 0.12fF $ **FLOATING
C5667 S.t1140 SUB 0.02fF
C5668 S.n5117 SUB 0.14fF $ **FLOATING
C5669 S.n5119 SUB 2.39fF $ **FLOATING
C5670 S.n5120 SUB 2.28fF $ **FLOATING
C5671 S.t380 SUB 0.02fF
C5672 S.n5121 SUB 0.12fF $ **FLOATING
C5673 S.n5122 SUB 0.14fF $ **FLOATING
C5674 S.t125 SUB 0.02fF
C5675 S.n5124 SUB 0.24fF $ **FLOATING
C5676 S.n5125 SUB 0.90fF $ **FLOATING
C5677 S.n5126 SUB 0.05fF $ **FLOATING
C5678 S.n5127 SUB 1.92fF $ **FLOATING
C5679 S.n5128 SUB 2.51fF $ **FLOATING
C5680 S.t1138 SUB 0.02fF
C5681 S.n5129 SUB 0.24fF $ **FLOATING
C5682 S.n5130 SUB 0.35fF $ **FLOATING
C5683 S.n5131 SUB 0.60fF $ **FLOATING
C5684 S.n5132 SUB 0.12fF $ **FLOATING
C5685 S.t750 SUB 0.02fF
C5686 S.n5133 SUB 0.14fF $ **FLOATING
C5687 S.n5135 SUB 2.39fF $ **FLOATING
C5688 S.n5136 SUB 2.28fF $ **FLOATING
C5689 S.t1097 SUB 0.02fF
C5690 S.n5137 SUB 0.12fF $ **FLOATING
C5691 S.n5138 SUB 0.14fF $ **FLOATING
C5692 S.t857 SUB 0.02fF
C5693 S.n5140 SUB 0.24fF $ **FLOATING
C5694 S.n5141 SUB 0.90fF $ **FLOATING
C5695 S.n5142 SUB 0.05fF $ **FLOATING
C5696 S.n5143 SUB 2.38fF $ **FLOATING
C5697 S.n5144 SUB 1.96fF $ **FLOATING
C5698 S.n5145 SUB 0.12fF $ **FLOATING
C5699 S.t368 SUB 0.02fF
C5700 S.n5146 SUB 0.14fF $ **FLOATING
C5701 S.t751 SUB 0.02fF
C5702 S.n5148 SUB 0.24fF $ **FLOATING
C5703 S.n5149 SUB 0.35fF $ **FLOATING
C5704 S.n5150 SUB 0.60fF $ **FLOATING
C5705 S.n5151 SUB 2.52fF $ **FLOATING
C5706 S.n5152 SUB 2.28fF $ **FLOATING
C5707 S.t711 SUB 0.02fF
C5708 S.n5153 SUB 0.12fF $ **FLOATING
C5709 S.n5154 SUB 0.14fF $ **FLOATING
C5710 S.t480 SUB 0.02fF
C5711 S.n5156 SUB 0.24fF $ **FLOATING
C5712 S.n5157 SUB 0.90fF $ **FLOATING
C5713 S.n5158 SUB 0.05fF $ **FLOATING
C5714 S.n5159 SUB 0.04fF $ **FLOATING
C5715 S.n5160 SUB 0.09fF $ **FLOATING
C5716 S.n5161 SUB 0.29fF $ **FLOATING
C5717 S.n5162 SUB 0.25fF $ **FLOATING
C5718 S.n5163 SUB 0.12fF $ **FLOATING
C5719 S.n5164 SUB 0.05fF $ **FLOATING
C5720 S.n5165 SUB 0.17fF $ **FLOATING
C5721 S.n5166 SUB 1.13fF $ **FLOATING
C5722 S.n5167 SUB 1.85fF $ **FLOATING
C5723 S.n5168 SUB 0.12fF $ **FLOATING
C5724 S.t1038 SUB 0.02fF
C5725 S.n5169 SUB 0.14fF $ **FLOATING
C5726 S.t364 SUB 0.02fF
C5727 S.n5171 SUB 0.24fF $ **FLOATING
C5728 S.n5172 SUB 0.35fF $ **FLOATING
C5729 S.n5173 SUB 0.60fF $ **FLOATING
C5730 S.n5174 SUB 2.52fF $ **FLOATING
C5731 S.n5175 SUB 1.92fF $ **FLOATING
C5732 S.t282 SUB 0.02fF
C5733 S.n5176 SUB 0.12fF $ **FLOATING
C5734 S.n5177 SUB 0.14fF $ **FLOATING
C5735 S.t507 SUB 0.02fF
C5736 S.n5179 SUB 0.24fF $ **FLOATING
C5737 S.n5180 SUB 0.90fF $ **FLOATING
C5738 S.n5181 SUB 0.05fF $ **FLOATING
C5739 S.t64 SUB 32.35fF
C5740 S.t385 SUB 0.02fF
C5741 S.n5182 SUB 0.12fF $ **FLOATING
C5742 S.n5183 SUB 0.14fF $ **FLOATING
C5743 S.t224 SUB 0.02fF
C5744 S.n5185 SUB 0.24fF $ **FLOATING
C5745 S.n5186 SUB 0.90fF $ **FLOATING
C5746 S.n5187 SUB 0.05fF $ **FLOATING
C5747 S.t550 SUB 0.02fF
C5748 S.n5188 SUB 0.24fF $ **FLOATING
C5749 S.n5189 SUB 0.35fF $ **FLOATING
C5750 S.n5190 SUB 0.60fF $ **FLOATING
C5751 S.n5191 SUB 0.30fF $ **FLOATING
C5752 S.n5192 SUB 1.08fF $ **FLOATING
C5753 S.n5193 SUB 0.15fF $ **FLOATING
C5754 S.n5194 SUB 2.08fF $ **FLOATING
C5755 S.n5195 SUB 1.77fF $ **FLOATING
C5756 S.n5196 SUB 1.86fF $ **FLOATING
C5757 S.n5197 SUB 0.12fF $ **FLOATING
C5758 S.t782 SUB 0.02fF
C5759 S.n5198 SUB 0.14fF $ **FLOATING
C5760 S.t1026 SUB 0.02fF
C5761 S.n5200 SUB 0.24fF $ **FLOATING
C5762 S.n5201 SUB 0.35fF $ **FLOATING
C5763 S.n5202 SUB 0.60fF $ **FLOATING
C5764 S.n5203 SUB 0.91fF $ **FLOATING
C5765 S.n5204 SUB 0.31fF $ **FLOATING
C5766 S.n5205 SUB 0.91fF $ **FLOATING
C5767 S.n5206 SUB 1.08fF $ **FLOATING
C5768 S.n5207 SUB 0.15fF $ **FLOATING
C5769 S.n5208 SUB 4.90fF $ **FLOATING
C5770 S.t493 SUB 0.02fF
C5771 S.n5209 SUB 0.24fF $ **FLOATING
C5772 S.n5210 SUB 0.90fF $ **FLOATING
C5773 S.n5211 SUB 0.05fF $ **FLOATING
C5774 S.t873 SUB 0.02fF
C5775 S.n5212 SUB 0.12fF $ **FLOATING
C5776 S.n5213 SUB 0.14fF $ **FLOATING
C5777 S.t200 SUB 0.02fF
C5778 S.n5215 SUB 0.94fF $ **FLOATING
C5779 S.n5216 SUB 0.70fF $ **FLOATING
C5780 S.n5217 SUB 1.74fF $ **FLOATING
C5781 S.n5218 SUB 3.01fF $ **FLOATING
C5782 S.t296 SUB 0.02fF
C5783 S.n5219 SUB 0.24fF $ **FLOATING
C5784 S.n5220 SUB 0.35fF $ **FLOATING
C5785 S.n5221 SUB 0.60fF $ **FLOATING
C5786 S.n5222 SUB 0.12fF $ **FLOATING
C5787 S.t36 SUB 0.02fF
C5788 S.n5223 SUB 0.14fF $ **FLOATING
C5789 S.n5225 SUB 0.18fF $ **FLOATING
C5790 S.n5226 SUB 0.20fF $ **FLOATING
C5791 S.n5227 SUB 0.22fF $ **FLOATING
C5792 S.n5228 SUB 0.65fF $ **FLOATING
C5793 S.n5229 SUB 0.90fF $ **FLOATING
C5794 S.n5230 SUB 0.22fF $ **FLOATING
C5795 S.n5231 SUB 0.09fF $ **FLOATING
C5796 S.n5232 SUB 0.20fF $ **FLOATING
C5797 S.n5233 SUB 0.07fF $ **FLOATING
C5798 S.n5234 SUB 0.06fF $ **FLOATING
C5799 S.n5235 SUB 0.07fF $ **FLOATING
C5800 S.n5236 SUB 1.97fF $ **FLOATING
C5801 S.t870 SUB 0.02fF
C5802 S.n5237 SUB 0.24fF $ **FLOATING
C5803 S.n5238 SUB 0.90fF $ **FLOATING
C5804 S.n5239 SUB 0.05fF $ **FLOATING
C5805 S.t82 SUB 0.02fF
C5806 S.n5240 SUB 0.12fF $ **FLOATING
C5807 S.n5241 SUB 0.14fF $ **FLOATING
C5808 S.n5243 SUB 14.09fF $ **FLOATING
C5809 S.n5244 SUB 0.25fF $ **FLOATING
C5810 S.n5245 SUB 0.09fF $ **FLOATING
C5811 S.n5246 SUB 0.20fF $ **FLOATING
C5812 S.n5247 SUB 0.77fF $ **FLOATING
C5813 S.n5248 SUB 1.91fF $ **FLOATING
C5814 S.n5249 SUB 1.86fF $ **FLOATING
C5815 S.n5250 SUB 0.12fF $ **FLOATING
C5816 S.t129 SUB 0.02fF
C5817 S.n5251 SUB 0.14fF $ **FLOATING
C5818 S.t676 SUB 0.02fF
C5819 S.n5253 SUB 0.24fF $ **FLOATING
C5820 S.n5254 SUB 0.35fF $ **FLOATING
C5821 S.n5255 SUB 0.60fF $ **FLOATING
C5822 S.n5256 SUB 2.64fF $ **FLOATING
C5823 S.n5257 SUB 2.96fF $ **FLOATING
C5824 S.t678 SUB 0.02fF
C5825 S.n5258 SUB 0.12fF $ **FLOATING
C5826 S.n5259 SUB 0.14fF $ **FLOATING
C5827 S.t39 SUB 0.02fF
C5828 S.n5261 SUB 0.24fF $ **FLOATING
C5829 S.n5262 SUB 0.90fF $ **FLOATING
C5830 S.n5263 SUB 0.05fF $ **FLOATING
C5831 S.t913 SUB 0.02fF
C5832 S.n5264 SUB 0.01fF $ **FLOATING
C5833 S.n5265 SUB 0.25fF $ **FLOATING
C5834 S.t35 SUB 32.35fF
C5835 S.n5266 SUB 0.25fF $ **FLOATING
C5836 S.n5267 SUB 2.89fF $ **FLOATING
C5837 S.n5268 SUB 13.46fF $ **FLOATING
C5838 S.n5269 SUB 0.59fF $ **FLOATING
C5839 S.n5270 SUB 0.44fF $ **FLOATING
C5840 S.n5271 SUB 0.59fF $ **FLOATING
C5841 S.n5272 SUB 2.57fF $ **FLOATING
C5842 S.n5273 SUB 0.29fF $ **FLOATING
C5843 S.t87 SUB 14.50fF
C5844 S.n5274 SUB 15.77fF $ **FLOATING
C5845 S.n5275 SUB 0.76fF $ **FLOATING
C5846 S.n5276 SUB 0.27fF $ **FLOATING
C5847 S.n5277 SUB 13.46fF $ **FLOATING
C5848 S.n5278 SUB 4.45fF $ **FLOATING
C5849 S.n5279 SUB 2.30fF $ **FLOATING
C5850 S.n5280 SUB 4.52fF $ **FLOATING
C5851 S.n5281 SUB 14.62fF $ **FLOATING
C5852 S.n5282 SUB 1.71fF $ **FLOATING
C5853 S.n5283 SUB 22.66fF $ **FLOATING
C5854 S.n5285 SUB 2.36fF $ **FLOATING
C5855 S.n5286 SUB 0.76fF $ **FLOATING
C5856 S.n5287 SUB 0.52fF $ **FLOATING
C5857 S.n5288 SUB 11.50fF $ **FLOATING
C5858 S.n5289 SUB 2.50fF $ **FLOATING
C5859 S.t503 SUB 0.02fF
C5860 S.n5290 SUB 1.26fF $ **FLOATING
C5861 S.t725 SUB 0.02fF
C5862 S.n5291 SUB 0.44fF $ **FLOATING
C5863 S.n5292 SUB 14.09fF $ **FLOATING
C5864 S.n5293 SUB 0.03fF $ **FLOATING
C5865 S.n5294 SUB 0.02fF $ **FLOATING
C5866 S.n5295 SUB 0.03fF $ **FLOATING
C5867 S.n5296 SUB 0.03fF $ **FLOATING
C5868 S.n5297 SUB 0.02fF $ **FLOATING
C5869 S.n5298 SUB 0.02fF $ **FLOATING
C5870 S.n5299 SUB 0.62fF $ **FLOATING
C5871 S.n5300 SUB 0.24fF $ **FLOATING
C5872 S.n5301 SUB 0.15fF $ **FLOATING
C5873 S.n5302 SUB 0.18fF $ **FLOATING
C5874 S.n5303 SUB 1.22fF $ **FLOATING
C5875 S.n5304 SUB 0.23fF $ **FLOATING
C5876 S.n5305 SUB 1.22fF $ **FLOATING
C5877 S.n5306 SUB 0.23fF $ **FLOATING
C5878 S.n5307 SUB 1.22fF $ **FLOATING
C5879 S.n5308 SUB 0.23fF $ **FLOATING
C5880 S.n5309 SUB 1.22fF $ **FLOATING
C5881 S.n5310 SUB 0.23fF $ **FLOATING
C5882 S.n5311 SUB 1.22fF $ **FLOATING
C5883 S.n5312 SUB 0.23fF $ **FLOATING
C5884 S.n5313 SUB 1.22fF $ **FLOATING
C5885 S.n5314 SUB 0.23fF $ **FLOATING
C5886 S.n5315 SUB 1.22fF $ **FLOATING
C5887 S.n5316 SUB 0.23fF $ **FLOATING
C5888 S.n5317 SUB 1.22fF $ **FLOATING
C5889 S.n5318 SUB 0.23fF $ **FLOATING
C5890 S.n5320 SUB 1.45fF $ **FLOATING
C5891 S.n5321 SUB 0.39fF $ **FLOATING
C5892 S.n5323 SUB 1.45fF $ **FLOATING
C5893 S.n5324 SUB 0.39fF $ **FLOATING
C5894 S.n5326 SUB 1.45fF $ **FLOATING
C5895 S.n5327 SUB 0.39fF $ **FLOATING
C5896 S.n5329 SUB 1.45fF $ **FLOATING
C5897 S.n5330 SUB 0.39fF $ **FLOATING
C5898 S.n5332 SUB 1.45fF $ **FLOATING
C5899 S.n5333 SUB 0.39fF $ **FLOATING
C5900 S.n5335 SUB 1.45fF $ **FLOATING
C5901 S.n5336 SUB 0.39fF $ **FLOATING
C5902 S.n5338 SUB 1.45fF $ **FLOATING
C5903 S.n5339 SUB 0.39fF $ **FLOATING
C5904 S.n5341 SUB 1.66fF $ **FLOATING
C5905 S.n5342 SUB 0.39fF $ **FLOATING
C5906 S.n5343 SUB 90.90fF $ **FLOATING
C5907 S.n5344 SUB 4.63fF $ **FLOATING
C5908 S.t1028 SUB 0.02fF
C5909 S.n5345 SUB 0.88fF $ **FLOATING
C5910 S.t250 SUB 0.02fF
C5911 S.n5346 SUB 0.02fF $ **FLOATING
C5912 S.n5347 SUB 0.37fF $ **FLOATING
C5913 S.t1055 SUB 0.02fF
C5914 S.n5348 SUB 0.88fF $ **FLOATING
C5915 S.n5349 SUB 0.92fF $ **FLOATING
C5916 S.n5350 SUB 4.04fF $ **FLOATING
C5917 S.n5351 SUB 1.83fF $ **FLOATING
C5918 S.t772 SUB 0.02fF
C5919 S.n5352 SUB 0.88fF $ **FLOATING
C5920 S.t812 SUB 0.02fF
C5921 S.n5353 SUB 0.88fF $ **FLOATING
C5922 S.n5354 SUB 2.10fF $ **FLOATING
C5923 S.n5355 SUB 1.18fF $ **FLOATING
C5924 S.n5356 SUB 0.32fF $ **FLOATING
C5925 S.n5357 SUB 0.31fF $ **FLOATING
C5926 S.t645 SUB 0.02fF
C5927 S.n5358 SUB 0.02fF $ **FLOATING
C5928 S.n5359 SUB 0.37fF $ **FLOATING
C5929 S.n5360 SUB 0.20fF $ **FLOATING
C5930 S.n5361 SUB 2.16fF $ **FLOATING
C5931 S.n5362 SUB 1.26fF $ **FLOATING
C5932 S.n5363 SUB 0.31fF $ **FLOATING
C5933 S.t489 SUB 0.02fF
C5934 S.n5364 SUB 0.88fF $ **FLOATING
C5935 S.t391 SUB 0.02fF
C5936 S.n5365 SUB 0.88fF $ **FLOATING
C5937 S.n5366 SUB 3.80fF $ **FLOATING
C5938 S.n5367 SUB 2.76fF $ **FLOATING
C5939 S.t270 SUB 0.02fF
C5940 S.n5368 SUB 0.02fF $ **FLOATING
C5941 S.n5369 SUB 0.37fF $ **FLOATING
C5942 S.n5370 SUB 2.40fF $ **FLOATING
C5943 S.t732 SUB 0.02fF
C5944 S.n5371 SUB 0.88fF $ **FLOATING
C5945 S.t663 SUB 0.02fF
C5946 S.n5372 SUB 0.88fF $ **FLOATING
C5947 S.n5373 SUB 0.95fF $ **FLOATING
C5948 S.n5374 SUB 3.56fF $ **FLOATING
C5949 S.n5375 SUB 2.76fF $ **FLOATING
C5950 S.t869 SUB 0.02fF
C5951 S.n5376 SUB 0.02fF $ **FLOATING
C5952 S.n5377 SUB 0.37fF $ **FLOATING
C5953 S.n5378 SUB 2.40fF $ **FLOATING
C5954 S.t350 SUB 0.02fF
C5955 S.n5379 SUB 0.88fF $ **FLOATING
C5956 S.t293 SUB 0.02fF
C5957 S.n5380 SUB 0.88fF $ **FLOATING
C5958 S.n5381 SUB 0.95fF $ **FLOATING
C5959 S.n5382 SUB 3.56fF $ **FLOATING
C5960 S.n5383 SUB 2.76fF $ **FLOATING
C5961 S.t492 SUB 0.02fF
C5962 S.n5384 SUB 0.02fF $ **FLOATING
C5963 S.n5385 SUB 0.37fF $ **FLOATING
C5964 S.n5386 SUB 2.40fF $ **FLOATING
C5965 S.t1077 SUB 0.02fF
C5966 S.n5387 SUB 0.88fF $ **FLOATING
C5967 S.t1021 SUB 0.02fF
C5968 S.n5388 SUB 0.88fF $ **FLOATING
C5969 S.n5389 SUB 0.95fF $ **FLOATING
C5970 S.n5390 SUB 3.56fF $ **FLOATING
C5971 S.n5391 SUB 2.76fF $ **FLOATING
C5972 S.t102 SUB 0.02fF
C5973 S.n5392 SUB 0.02fF $ **FLOATING
C5974 S.n5393 SUB 0.37fF $ **FLOATING
C5975 S.n5394 SUB 2.40fF $ **FLOATING
C5976 S.t690 SUB 0.02fF
C5977 S.n5395 SUB 0.88fF $ **FLOATING
C5978 S.t648 SUB 0.02fF
C5979 S.n5396 SUB 0.88fF $ **FLOATING
C5980 S.n5397 SUB 0.95fF $ **FLOATING
C5981 S.n5398 SUB 3.56fF $ **FLOATING
C5982 S.n5399 SUB 2.76fF $ **FLOATING
C5983 S.t834 SUB 0.02fF
C5984 S.n5400 SUB 0.02fF $ **FLOATING
C5985 S.n5401 SUB 0.37fF $ **FLOATING
C5986 S.n5402 SUB 2.40fF $ **FLOATING
C5987 S.t313 SUB 0.02fF
C5988 S.n5403 SUB 0.88fF $ **FLOATING
C5989 S.t300 SUB 0.02fF
C5990 S.n5404 SUB 0.88fF $ **FLOATING
C5991 S.n5405 SUB 0.95fF $ **FLOATING
C5992 S.n5406 SUB 3.56fF $ **FLOATING
C5993 S.n5407 SUB 2.76fF $ **FLOATING
C5994 S.t514 SUB 0.02fF
C5995 S.n5408 SUB 0.02fF $ **FLOATING
C5996 S.n5409 SUB 0.37fF $ **FLOATING
C5997 S.n5410 SUB 2.40fF $ **FLOATING
C5998 S.t1045 SUB 0.02fF
C5999 S.n5411 SUB 0.88fF $ **FLOATING
C6000 S.t1031 SUB 0.02fF
C6001 S.n5412 SUB 0.88fF $ **FLOATING
C6002 S.n5413 SUB 0.95fF $ **FLOATING
C6003 S.n5414 SUB 3.56fF $ **FLOATING
C6004 S.n5415 SUB 2.76fF $ **FLOATING
C6005 S.t122 SUB 0.02fF
C6006 S.n5416 SUB 0.02fF $ **FLOATING
C6007 S.n5417 SUB 0.37fF $ **FLOATING
C6008 S.n5418 SUB 0.95fF $ **FLOATING
C6009 S.n5419 SUB 3.56fF $ **FLOATING
C6010 S.n5420 SUB 2.77fF $ **FLOATING
C6011 S.t656 SUB 0.02fF
C6012 S.n5421 SUB 0.88fF $ **FLOATING
C6013 S.t668 SUB 0.02fF
C6014 S.n5422 SUB 0.88fF $ **FLOATING
C6015 S.n5423 SUB 2.40fF $ **FLOATING
C6016 S.t853 SUB 0.02fF
C6017 S.n5424 SUB 0.02fF $ **FLOATING
C6018 S.n5425 SUB 0.37fF $ **FLOATING
C6019 S.n5426 SUB 3.91fF $ **FLOATING
C6020 S.n5427 SUB 2.75fF $ **FLOATING
C6021 S.n5428 SUB 0.03fF $ **FLOATING
C6022 S.n5429 SUB 0.02fF $ **FLOATING
C6023 S.n5430 SUB 0.03fF $ **FLOATING
C6024 S.n5431 SUB 0.03fF $ **FLOATING
C6025 S.n5432 SUB 0.02fF $ **FLOATING
C6026 S.n5433 SUB 0.02fF $ **FLOATING
C6027 S.n5434 SUB 0.62fF $ **FLOATING
C6028 S.n5435 SUB 0.24fF $ **FLOATING
C6029 S.n5436 SUB 0.15fF $ **FLOATING
C6030 S.n5437 SUB 0.18fF $ **FLOATING
C6031 S.t284 SUB 0.02fF
C6032 S.n5438 SUB 0.88fF $ **FLOATING
C6033 S.t297 SUB 0.02fF
C6034 S.n5439 SUB 0.88fF $ **FLOATING
C6035 S.t477 SUB 0.02fF
C6036 S.n5440 SUB 0.02fF $ **FLOATING
C6037 S.n5441 SUB 0.37fF $ **FLOATING
C6038 S.t283 SUB 111.86fF
C6039 S.n5442 SUB 0.46fF $ **FLOATING
C6040 S.n5443 SUB 4.38fF $ **FLOATING
C6041 S.n5444 SUB 2.49fF $ **FLOATING
C6042 S.n5445 SUB 6.90fF $ **FLOATING
C6043 S.n5446 SUB 15.90fF $ **FLOATING
C6044 S.n5447 SUB 8.87fF $ **FLOATING
C6045 S.n5448 SUB 8.87fF $ **FLOATING
C6046 S.n5449 SUB 0.59fF $ **FLOATING
C6047 S.n5450 SUB 0.21fF $ **FLOATING
C6048 S.n5451 SUB 0.59fF $ **FLOATING
C6049 S.n5452 SUB 2.57fF $ **FLOATING
C6050 S.n5453 SUB 0.29fF $ **FLOATING
C6051 S.t118 SUB 14.50fF
C6052 S.n5454 SUB 15.77fF $ **FLOATING
C6053 S.n5455 SUB 0.76fF $ **FLOATING
C6054 S.n5456 SUB 0.27fF $ **FLOATING
C6055 S.n5457 SUB 4.22fF $ **FLOATING
C6056 S.n5458 SUB 2.77fF $ **FLOATING
C6057 S.n5459 SUB 1.87fF $ **FLOATING
C6058 S.n5460 SUB 0.06fF $ **FLOATING
C6059 S.n5461 SUB 0.03fF $ **FLOATING
C6060 S.n5462 SUB 0.03fF $ **FLOATING
C6061 S.n5463 SUB 0.98fF $ **FLOATING
C6062 S.n5464 SUB 0.02fF $ **FLOATING
C6063 S.n5465 SUB 0.01fF $ **FLOATING
C6064 S.n5466 SUB 0.02fF $ **FLOATING
C6065 S.n5467 SUB 0.08fF $ **FLOATING
C6066 S.n5468 SUB 0.36fF $ **FLOATING
C6067 S.n5469 SUB 1.83fF $ **FLOATING
C6068 S.t119 SUB 0.02fF
C6069 S.n5470 SUB 0.24fF $ **FLOATING
C6070 S.n5471 SUB 0.35fF $ **FLOATING
C6071 S.n5472 SUB 0.60fF $ **FLOATING
C6072 S.n5473 SUB 0.12fF $ **FLOATING
C6073 S.t1012 SUB 0.02fF
C6074 S.n5474 SUB 0.14fF $ **FLOATING
C6075 S.n5476 SUB 0.69fF $ **FLOATING
C6076 S.n5477 SUB 0.22fF $ **FLOATING
C6077 S.n5478 SUB 0.22fF $ **FLOATING
C6078 S.n5479 SUB 0.69fF $ **FLOATING
C6079 S.n5480 SUB 1.14fF $ **FLOATING
C6080 S.n5481 SUB 0.22fF $ **FLOATING
C6081 S.n5482 SUB 0.25fF $ **FLOATING
C6082 S.n5483 SUB 0.09fF $ **FLOATING
C6083 S.n5484 SUB 1.86fF $ **FLOATING
C6084 S.t636 SUB 0.02fF
C6085 S.n5485 SUB 0.24fF $ **FLOATING
C6086 S.n5486 SUB 0.90fF $ **FLOATING
C6087 S.n5487 SUB 0.05fF $ **FLOATING
C6088 S.t1060 SUB 0.02fF
C6089 S.n5488 SUB 0.12fF $ **FLOATING
C6090 S.n5489 SUB 0.14fF $ **FLOATING
C6091 S.n5491 SUB 14.09fF $ **FLOATING
C6092 S.n5492 SUB 0.09fF $ **FLOATING
C6093 S.n5493 SUB 0.20fF $ **FLOATING
C6094 S.n5494 SUB 0.07fF $ **FLOATING
C6095 S.n5495 SUB 0.06fF $ **FLOATING
C6096 S.n5496 SUB 0.07fF $ **FLOATING
C6097 S.n5497 SUB 0.18fF $ **FLOATING
C6098 S.n5498 SUB 0.19fF $ **FLOATING
C6099 S.n5499 SUB 1.02fF $ **FLOATING
C6100 S.n5500 SUB 0.53fF $ **FLOATING
C6101 S.n5501 SUB 2.31fF $ **FLOATING
C6102 S.n5502 SUB 0.12fF $ **FLOATING
C6103 S.t285 SUB 0.02fF
C6104 S.n5503 SUB 0.14fF $ **FLOATING
C6105 S.t511 SUB 0.02fF
C6106 S.n5505 SUB 0.24fF $ **FLOATING
C6107 S.n5506 SUB 0.35fF $ **FLOATING
C6108 S.n5507 SUB 0.60fF $ **FLOATING
C6109 S.n5508 SUB 1.71fF $ **FLOATING
C6110 S.n5509 SUB 2.41fF $ **FLOATING
C6111 S.t298 SUB 0.02fF
C6112 S.n5510 SUB 0.12fF $ **FLOATING
C6113 S.n5511 SUB 0.14fF $ **FLOATING
C6114 S.t1013 SUB 0.02fF
C6115 S.n5513 SUB 0.24fF $ **FLOATING
C6116 S.n5514 SUB 0.90fF $ **FLOATING
C6117 S.n5515 SUB 0.05fF $ **FLOATING
C6118 S.n5516 SUB 2.91fF $ **FLOATING
C6119 S.n5517 SUB 1.86fF $ **FLOATING
C6120 S.n5518 SUB 0.12fF $ **FLOATING
C6121 S.t1096 SUB 0.02fF
C6122 S.n5519 SUB 0.14fF $ **FLOATING
C6123 S.t269 SUB 0.02fF
C6124 S.n5521 SUB 0.24fF $ **FLOATING
C6125 S.n5522 SUB 0.35fF $ **FLOATING
C6126 S.n5523 SUB 0.60fF $ **FLOATING
C6127 S.n5524 SUB 0.91fF $ **FLOATING
C6128 S.n5525 SUB 0.31fF $ **FLOATING
C6129 S.n5526 SUB 0.91fF $ **FLOATING
C6130 S.n5527 SUB 1.08fF $ **FLOATING
C6131 S.n5528 SUB 0.15fF $ **FLOATING
C6132 S.n5529 SUB 4.90fF $ **FLOATING
C6133 S.t84 SUB 0.02fF
C6134 S.n5530 SUB 0.12fF $ **FLOATING
C6135 S.n5531 SUB 0.14fF $ **FLOATING
C6136 S.t946 SUB 0.02fF
C6137 S.n5533 SUB 0.24fF $ **FLOATING
C6138 S.n5534 SUB 0.90fF $ **FLOATING
C6139 S.n5535 SUB 0.05fF $ **FLOATING
C6140 S.n5536 SUB 1.86fF $ **FLOATING
C6141 S.n5537 SUB 2.64fF $ **FLOATING
C6142 S.t988 SUB 0.02fF
C6143 S.n5538 SUB 0.24fF $ **FLOATING
C6144 S.n5539 SUB 0.35fF $ **FLOATING
C6145 S.n5540 SUB 0.60fF $ **FLOATING
C6146 S.n5541 SUB 0.12fF $ **FLOATING
C6147 S.t708 SUB 0.02fF
C6148 S.n5542 SUB 0.14fF $ **FLOATING
C6149 S.n5544 SUB 2.91fF $ **FLOATING
C6150 S.n5545 SUB 5.10fF $ **FLOATING
C6151 S.t820 SUB 0.02fF
C6152 S.n5546 SUB 0.12fF $ **FLOATING
C6153 S.n5547 SUB 0.14fF $ **FLOATING
C6154 S.t565 SUB 0.02fF
C6155 S.n5549 SUB 0.24fF $ **FLOATING
C6156 S.n5550 SUB 0.90fF $ **FLOATING
C6157 S.n5551 SUB 0.05fF $ **FLOATING
C6158 S.n5552 SUB 1.86fF $ **FLOATING
C6159 S.n5553 SUB 2.64fF $ **FLOATING
C6160 S.t611 SUB 0.02fF
C6161 S.n5554 SUB 0.24fF $ **FLOATING
C6162 S.n5555 SUB 0.35fF $ **FLOATING
C6163 S.n5556 SUB 0.60fF $ **FLOATING
C6164 S.n5557 SUB 0.12fF $ **FLOATING
C6165 S.t330 SUB 0.02fF
C6166 S.n5558 SUB 0.14fF $ **FLOATING
C6167 S.n5560 SUB 5.11fF $ **FLOATING
C6168 S.t449 SUB 0.02fF
C6169 S.n5561 SUB 0.12fF $ **FLOATING
C6170 S.n5562 SUB 0.14fF $ **FLOATING
C6171 S.t172 SUB 0.02fF
C6172 S.n5564 SUB 0.24fF $ **FLOATING
C6173 S.n5565 SUB 0.90fF $ **FLOATING
C6174 S.n5566 SUB 0.05fF $ **FLOATING
C6175 S.n5567 SUB 1.86fF $ **FLOATING
C6176 S.n5568 SUB 2.64fF $ **FLOATING
C6177 S.t223 SUB 0.02fF
C6178 S.n5569 SUB 0.24fF $ **FLOATING
C6179 S.n5570 SUB 0.35fF $ **FLOATING
C6180 S.n5571 SUB 0.60fF $ **FLOATING
C6181 S.n5572 SUB 0.12fF $ **FLOATING
C6182 S.t1056 SUB 0.02fF
C6183 S.n5573 SUB 0.14fF $ **FLOATING
C6184 S.n5575 SUB 5.11fF $ **FLOATING
C6185 S.t26 SUB 0.02fF
C6186 S.n5576 SUB 0.12fF $ **FLOATING
C6187 S.n5577 SUB 0.14fF $ **FLOATING
C6188 S.t897 SUB 0.02fF
C6189 S.n5579 SUB 0.24fF $ **FLOATING
C6190 S.n5580 SUB 0.90fF $ **FLOATING
C6191 S.n5581 SUB 0.05fF $ **FLOATING
C6192 S.n5582 SUB 1.86fF $ **FLOATING
C6193 S.n5583 SUB 2.64fF $ **FLOATING
C6194 S.t1008 SUB 0.02fF
C6195 S.n5584 SUB 0.24fF $ **FLOATING
C6196 S.n5585 SUB 0.35fF $ **FLOATING
C6197 S.n5586 SUB 0.60fF $ **FLOATING
C6198 S.n5587 SUB 0.12fF $ **FLOATING
C6199 S.t730 SUB 0.02fF
C6200 S.n5588 SUB 0.14fF $ **FLOATING
C6201 S.n5590 SUB 5.11fF $ **FLOATING
C6202 S.t775 SUB 0.02fF
C6203 S.n5591 SUB 0.12fF $ **FLOATING
C6204 S.n5592 SUB 0.14fF $ **FLOATING
C6205 S.t593 SUB 0.02fF
C6206 S.n5594 SUB 0.24fF $ **FLOATING
C6207 S.n5595 SUB 0.90fF $ **FLOATING
C6208 S.n5596 SUB 0.05fF $ **FLOATING
C6209 S.n5597 SUB 1.86fF $ **FLOATING
C6210 S.n5598 SUB 2.64fF $ **FLOATING
C6211 S.t631 SUB 0.02fF
C6212 S.n5599 SUB 0.24fF $ **FLOATING
C6213 S.n5600 SUB 0.35fF $ **FLOATING
C6214 S.n5601 SUB 0.60fF $ **FLOATING
C6215 S.n5602 SUB 0.12fF $ **FLOATING
C6216 S.t347 SUB 0.02fF
C6217 S.n5603 SUB 0.14fF $ **FLOATING
C6218 S.n5605 SUB 5.11fF $ **FLOATING
C6219 S.t394 SUB 0.02fF
C6220 S.n5606 SUB 0.12fF $ **FLOATING
C6221 S.n5607 SUB 0.14fF $ **FLOATING
C6222 S.t196 SUB 0.02fF
C6223 S.n5609 SUB 0.24fF $ **FLOATING
C6224 S.n5610 SUB 0.90fF $ **FLOATING
C6225 S.n5611 SUB 0.05fF $ **FLOATING
C6226 S.n5612 SUB 1.86fF $ **FLOATING
C6227 S.n5613 SUB 2.64fF $ **FLOATING
C6228 S.t247 SUB 0.02fF
C6229 S.n5614 SUB 0.24fF $ **FLOATING
C6230 S.n5615 SUB 0.35fF $ **FLOATING
C6231 S.n5616 SUB 0.60fF $ **FLOATING
C6232 S.n5617 SUB 0.12fF $ **FLOATING
C6233 S.t1075 SUB 0.02fF
C6234 S.n5618 SUB 0.14fF $ **FLOATING
C6235 S.n5620 SUB 5.11fF $ **FLOATING
C6236 S.t1114 SUB 0.02fF
C6237 S.n5621 SUB 0.12fF $ **FLOATING
C6238 S.n5622 SUB 0.14fF $ **FLOATING
C6239 S.t918 SUB 0.02fF
C6240 S.n5624 SUB 0.24fF $ **FLOATING
C6241 S.n5625 SUB 0.90fF $ **FLOATING
C6242 S.n5626 SUB 0.05fF $ **FLOATING
C6243 S.n5627 SUB 1.86fF $ **FLOATING
C6244 S.n5628 SUB 2.64fF $ **FLOATING
C6245 S.t970 SUB 0.02fF
C6246 S.n5629 SUB 0.24fF $ **FLOATING
C6247 S.n5630 SUB 0.35fF $ **FLOATING
C6248 S.n5631 SUB 0.60fF $ **FLOATING
C6249 S.n5632 SUB 0.12fF $ **FLOATING
C6250 S.t693 SUB 0.02fF
C6251 S.n5633 SUB 0.14fF $ **FLOATING
C6252 S.n5635 SUB 4.84fF $ **FLOATING
C6253 S.t723 SUB 0.02fF
C6254 S.n5636 SUB 0.12fF $ **FLOATING
C6255 S.n5637 SUB 0.14fF $ **FLOATING
C6256 S.t542 SUB 0.02fF
C6257 S.n5639 SUB 0.24fF $ **FLOATING
C6258 S.n5640 SUB 0.90fF $ **FLOATING
C6259 S.n5641 SUB 0.05fF $ **FLOATING
C6260 S.n5642 SUB 0.10fF $ **FLOATING
C6261 S.n5643 SUB 0.12fF $ **FLOATING
C6262 S.n5644 SUB 0.09fF $ **FLOATING
C6263 S.n5645 SUB 0.12fF $ **FLOATING
C6264 S.n5646 SUB 0.18fF $ **FLOATING
C6265 S.n5647 SUB 1.86fF $ **FLOATING
C6266 S.n5648 SUB 0.12fF $ **FLOATING
C6267 S.t401 SUB 0.02fF
C6268 S.n5649 SUB 0.14fF $ **FLOATING
C6269 S.t30 SUB 0.02fF
C6270 S.n5651 SUB 1.20fF $ **FLOATING
C6271 S.n5652 SUB 0.06fF $ **FLOATING
C6272 S.n5653 SUB 0.10fF $ **FLOATING
C6273 S.n5654 SUB 0.60fF $ **FLOATING
C6274 S.n5655 SUB 0.35fF $ **FLOATING
C6275 S.n5656 SUB 0.62fF $ **FLOATING
C6276 S.n5657 SUB 1.14fF $ **FLOATING
C6277 S.n5658 SUB 2.18fF $ **FLOATING
C6278 S.n5659 SUB 0.59fF $ **FLOATING
C6279 S.n5660 SUB 0.02fF $ **FLOATING
C6280 S.n5661 SUB 0.96fF $ **FLOATING
C6281 S.t29 SUB 14.50fF
C6282 S.n5662 SUB 14.37fF $ **FLOATING
C6283 S.n5664 SUB 0.37fF $ **FLOATING
C6284 S.n5665 SUB 0.23fF $ **FLOATING
C6285 S.n5666 SUB 2.86fF $ **FLOATING
C6286 S.n5667 SUB 2.39fF $ **FLOATING
C6287 S.n5668 SUB 2.44fF $ **FLOATING
C6288 S.n5669 SUB 4.24fF $ **FLOATING
C6289 S.n5670 SUB 0.25fF $ **FLOATING
C6290 S.n5671 SUB 0.01fF $ **FLOATING
C6291 S.t1037 SUB 0.02fF
C6292 S.n5672 SUB 0.25fF $ **FLOATING
C6293 S.t800 SUB 0.02fF
C6294 S.n5673 SUB 0.94fF $ **FLOATING
C6295 S.n5674 SUB 0.70fF $ **FLOATING
C6296 S.n5675 SUB 1.87fF $ **FLOATING
C6297 S.n5676 SUB 1.86fF $ **FLOATING
C6298 S.t779 SUB 0.02fF
C6299 S.n5677 SUB 0.24fF $ **FLOATING
C6300 S.n5678 SUB 0.35fF $ **FLOATING
C6301 S.n5679 SUB 0.60fF $ **FLOATING
C6302 S.n5680 SUB 0.12fF $ **FLOATING
C6303 S.t691 SUB 0.02fF
C6304 S.n5681 SUB 0.14fF $ **FLOATING
C6305 S.n5683 SUB 1.14fF $ **FLOATING
C6306 S.n5684 SUB 0.22fF $ **FLOATING
C6307 S.n5685 SUB 0.25fF $ **FLOATING
C6308 S.n5686 SUB 0.09fF $ **FLOATING
C6309 S.n5687 SUB 1.86fF $ **FLOATING
C6310 S.t420 SUB 0.02fF
C6311 S.n5688 SUB 0.24fF $ **FLOATING
C6312 S.n5689 SUB 0.90fF $ **FLOATING
C6313 S.n5690 SUB 0.05fF $ **FLOATING
C6314 S.t1023 SUB 0.02fF
C6315 S.n5691 SUB 0.12fF $ **FLOATING
C6316 S.n5692 SUB 0.14fF $ **FLOATING
C6317 S.n5694 SUB 0.76fF $ **FLOATING
C6318 S.n5695 SUB 0.44fF $ **FLOATING
C6319 S.n5696 SUB 1.56fF $ **FLOATING
C6320 S.n5697 SUB 0.12fF $ **FLOATING
C6321 S.t589 SUB 0.02fF
C6322 S.n5698 SUB 0.14fF $ **FLOATING
C6323 S.t1063 SUB 0.02fF
C6324 S.n5700 SUB 0.24fF $ **FLOATING
C6325 S.n5701 SUB 0.35fF $ **FLOATING
C6326 S.n5702 SUB 0.60fF $ **FLOATING
C6327 S.n5703 SUB 0.01fF $ **FLOATING
C6328 S.n5704 SUB 0.07fF $ **FLOATING
C6329 S.n5705 SUB 0.01fF $ **FLOATING
C6330 S.n5706 SUB 0.01fF $ **FLOATING
C6331 S.n5707 SUB 0.01fF $ **FLOATING
C6332 S.n5708 SUB 0.24fF $ **FLOATING
C6333 S.n5709 SUB 1.15fF $ **FLOATING
C6334 S.n5710 SUB 1.33fF $ **FLOATING
C6335 S.n5711 SUB 1.97fF $ **FLOATING
C6336 S.t402 SUB 0.02fF
C6337 S.n5712 SUB 0.24fF $ **FLOATING
C6338 S.n5713 SUB 0.90fF $ **FLOATING
C6339 S.n5714 SUB 0.05fF $ **FLOATING
C6340 S.t894 SUB 0.02fF
C6341 S.n5715 SUB 0.12fF $ **FLOATING
C6342 S.n5716 SUB 0.14fF $ **FLOATING
C6343 S.n5718 SUB 14.09fF $ **FLOATING
C6344 S.n5719 SUB 1.86fF $ **FLOATING
C6345 S.n5720 SUB 0.12fF $ **FLOATING
C6346 S.t131 SUB 0.02fF
C6347 S.n5721 SUB 0.14fF $ **FLOATING
C6348 S.t917 SUB 0.02fF
C6349 S.n5723 SUB 0.24fF $ **FLOATING
C6350 S.n5724 SUB 0.35fF $ **FLOATING
C6351 S.n5725 SUB 0.60fF $ **FLOATING
C6352 S.n5726 SUB 0.31fF $ **FLOATING
C6353 S.n5727 SUB 1.08fF $ **FLOATING
C6354 S.n5728 SUB 0.15fF $ **FLOATING
C6355 S.n5729 SUB 2.08fF $ **FLOATING
C6356 S.t649 SUB 0.02fF
C6357 S.n5730 SUB 0.12fF $ **FLOATING
C6358 S.n5731 SUB 0.14fF $ **FLOATING
C6359 S.t619 SUB 0.02fF
C6360 S.n5733 SUB 0.24fF $ **FLOATING
C6361 S.n5734 SUB 0.90fF $ **FLOATING
C6362 S.n5735 SUB 0.05fF $ **FLOATING
C6363 S.n5736 SUB 1.86fF $ **FLOATING
C6364 S.n5737 SUB 2.64fF $ **FLOATING
C6365 S.t541 SUB 0.02fF
C6366 S.n5738 SUB 0.24fF $ **FLOATING
C6367 S.n5739 SUB 0.35fF $ **FLOATING
C6368 S.n5740 SUB 0.60fF $ **FLOATING
C6369 S.n5741 SUB 0.12fF $ **FLOATING
C6370 S.t860 SUB 0.02fF
C6371 S.n5742 SUB 0.14fF $ **FLOATING
C6372 S.n5744 SUB 2.28fF $ **FLOATING
C6373 S.t5 SUB 0.02fF
C6374 S.n5745 SUB 0.12fF $ **FLOATING
C6375 S.n5746 SUB 0.14fF $ **FLOATING
C6376 S.t231 SUB 0.02fF
C6377 S.n5748 SUB 0.24fF $ **FLOATING
C6378 S.n5749 SUB 0.90fF $ **FLOATING
C6379 S.n5750 SUB 0.05fF $ **FLOATING
C6380 S.n5751 SUB 1.86fF $ **FLOATING
C6381 S.n5752 SUB 2.64fF $ **FLOATING
C6382 S.t151 SUB 0.02fF
C6383 S.n5753 SUB 0.24fF $ **FLOATING
C6384 S.n5754 SUB 0.35fF $ **FLOATING
C6385 S.n5755 SUB 0.60fF $ **FLOATING
C6386 S.n5756 SUB 0.12fF $ **FLOATING
C6387 S.t484 SUB 0.02fF
C6388 S.n5757 SUB 0.14fF $ **FLOATING
C6389 S.n5759 SUB 2.77fF $ **FLOATING
C6390 S.n5760 SUB 2.28fF $ **FLOATING
C6391 S.t765 SUB 0.02fF
C6392 S.n5761 SUB 0.12fF $ **FLOATING
C6393 S.n5762 SUB 0.14fF $ **FLOATING
C6394 S.t960 SUB 0.02fF
C6395 S.n5764 SUB 0.24fF $ **FLOATING
C6396 S.n5765 SUB 0.90fF $ **FLOATING
C6397 S.n5766 SUB 0.05fF $ **FLOATING
C6398 S.n5767 SUB 1.86fF $ **FLOATING
C6399 S.n5768 SUB 2.64fF $ **FLOATING
C6400 S.t881 SUB 0.02fF
C6401 S.n5769 SUB 0.24fF $ **FLOATING
C6402 S.n5770 SUB 0.35fF $ **FLOATING
C6403 S.n5771 SUB 0.60fF $ **FLOATING
C6404 S.n5772 SUB 0.12fF $ **FLOATING
C6405 S.t93 SUB 0.02fF
C6406 S.n5773 SUB 0.14fF $ **FLOATING
C6407 S.n5775 SUB 2.77fF $ **FLOATING
C6408 S.n5776 SUB 2.28fF $ **FLOATING
C6409 S.t383 SUB 0.02fF
C6410 S.n5777 SUB 0.12fF $ **FLOATING
C6411 S.n5778 SUB 0.14fF $ **FLOATING
C6412 S.t574 SUB 0.02fF
C6413 S.n5780 SUB 0.24fF $ **FLOATING
C6414 S.n5781 SUB 0.90fF $ **FLOATING
C6415 S.n5782 SUB 0.05fF $ **FLOATING
C6416 S.n5783 SUB 1.86fF $ **FLOATING
C6417 S.n5784 SUB 2.64fF $ **FLOATING
C6418 S.t504 SUB 0.02fF
C6419 S.n5785 SUB 0.24fF $ **FLOATING
C6420 S.n5786 SUB 0.35fF $ **FLOATING
C6421 S.n5787 SUB 0.60fF $ **FLOATING
C6422 S.n5788 SUB 0.12fF $ **FLOATING
C6423 S.t827 SUB 0.02fF
C6424 S.n5789 SUB 0.14fF $ **FLOATING
C6425 S.n5791 SUB 2.77fF $ **FLOATING
C6426 S.n5792 SUB 2.28fF $ **FLOATING
C6427 S.t1101 SUB 0.02fF
C6428 S.n5793 SUB 0.12fF $ **FLOATING
C6429 S.n5794 SUB 0.14fF $ **FLOATING
C6430 S.t179 SUB 0.02fF
C6431 S.n5796 SUB 0.24fF $ **FLOATING
C6432 S.n5797 SUB 0.90fF $ **FLOATING
C6433 S.n5798 SUB 0.05fF $ **FLOATING
C6434 S.n5799 SUB 1.86fF $ **FLOATING
C6435 S.n5800 SUB 2.64fF $ **FLOATING
C6436 S.t114 SUB 0.02fF
C6437 S.n5801 SUB 0.24fF $ **FLOATING
C6438 S.n5802 SUB 0.35fF $ **FLOATING
C6439 S.n5803 SUB 0.60fF $ **FLOATING
C6440 S.n5804 SUB 0.12fF $ **FLOATING
C6441 S.t451 SUB 0.02fF
C6442 S.n5805 SUB 0.14fF $ **FLOATING
C6443 S.n5807 SUB 2.77fF $ **FLOATING
C6444 S.n5808 SUB 2.28fF $ **FLOATING
C6445 S.t794 SUB 0.02fF
C6446 S.n5809 SUB 0.12fF $ **FLOATING
C6447 S.n5810 SUB 0.14fF $ **FLOATING
C6448 S.t902 SUB 0.02fF
C6449 S.n5812 SUB 0.24fF $ **FLOATING
C6450 S.n5813 SUB 0.90fF $ **FLOATING
C6451 S.n5814 SUB 0.05fF $ **FLOATING
C6452 S.n5815 SUB 1.86fF $ **FLOATING
C6453 S.n5816 SUB 2.64fF $ **FLOATING
C6454 S.t847 SUB 0.02fF
C6455 S.n5817 SUB 0.24fF $ **FLOATING
C6456 S.n5818 SUB 0.35fF $ **FLOATING
C6457 S.n5819 SUB 0.60fF $ **FLOATING
C6458 S.n5820 SUB 0.12fF $ **FLOATING
C6459 S.t38 SUB 0.02fF
C6460 S.n5821 SUB 0.14fF $ **FLOATING
C6461 S.n5823 SUB 2.77fF $ **FLOATING
C6462 S.n5824 SUB 2.28fF $ **FLOATING
C6463 S.t413 SUB 0.02fF
C6464 S.n5825 SUB 0.12fF $ **FLOATING
C6465 S.n5826 SUB 0.14fF $ **FLOATING
C6466 S.t529 SUB 0.02fF
C6467 S.n5828 SUB 0.24fF $ **FLOATING
C6468 S.n5829 SUB 0.90fF $ **FLOATING
C6469 S.n5830 SUB 0.05fF $ **FLOATING
C6470 S.n5831 SUB 1.86fF $ **FLOATING
C6471 S.n5832 SUB 2.64fF $ **FLOATING
C6472 S.t470 SUB 0.02fF
C6473 S.n5833 SUB 0.24fF $ **FLOATING
C6474 S.n5834 SUB 0.35fF $ **FLOATING
C6475 S.n5835 SUB 0.60fF $ **FLOATING
C6476 S.n5836 SUB 0.12fF $ **FLOATING
C6477 S.t784 SUB 0.02fF
C6478 S.n5837 SUB 0.14fF $ **FLOATING
C6479 S.n5839 SUB 2.77fF $ **FLOATING
C6480 S.n5840 SUB 2.28fF $ **FLOATING
C6481 S.t1129 SUB 0.02fF
C6482 S.n5841 SUB 0.12fF $ **FLOATING
C6483 S.n5842 SUB 0.14fF $ **FLOATING
C6484 S.t140 SUB 0.02fF
C6485 S.n5844 SUB 0.24fF $ **FLOATING
C6486 S.n5845 SUB 0.90fF $ **FLOATING
C6487 S.n5846 SUB 0.05fF $ **FLOATING
C6488 S.t4 SUB 32.35fF
C6489 S.t745 SUB 0.02fF
C6490 S.n5847 SUB 0.12fF $ **FLOATING
C6491 S.n5848 SUB 0.14fF $ **FLOATING
C6492 S.t866 SUB 0.02fF
C6493 S.n5850 SUB 0.24fF $ **FLOATING
C6494 S.n5851 SUB 0.90fF $ **FLOATING
C6495 S.n5852 SUB 0.05fF $ **FLOATING
C6496 S.t70 SUB 0.02fF
C6497 S.n5853 SUB 0.24fF $ **FLOATING
C6498 S.n5854 SUB 0.35fF $ **FLOATING
C6499 S.n5855 SUB 0.60fF $ **FLOATING
C6500 S.n5856 SUB 2.63fF $ **FLOATING
C6501 S.n5857 SUB 3.24fF $ **FLOATING
C6502 S.n5858 SUB 0.10fF $ **FLOATING
C6503 S.n5859 SUB 0.35fF $ **FLOATING
C6504 S.n5860 SUB 0.46fF $ **FLOATING
C6505 S.n5861 SUB 1.12fF $ **FLOATING
C6506 S.n5862 SUB 1.85fF $ **FLOATING
C6507 S.n5863 SUB 0.12fF $ **FLOATING
C6508 S.t334 SUB 0.02fF
C6509 S.n5864 SUB 0.14fF $ **FLOATING
C6510 S.t924 SUB 0.02fF
C6511 S.n5866 SUB 0.24fF $ **FLOATING
C6512 S.n5867 SUB 0.35fF $ **FLOATING
C6513 S.n5868 SUB 0.60fF $ **FLOATING
C6514 S.n5869 SUB 1.25fF $ **FLOATING
C6515 S.n5870 SUB 2.36fF $ **FLOATING
C6516 S.n5871 SUB 4.16fF $ **FLOATING
C6517 S.t340 SUB 0.02fF
C6518 S.n5872 SUB 0.12fF $ **FLOATING
C6519 S.n5873 SUB 0.14fF $ **FLOATING
C6520 S.t661 SUB 0.02fF
C6521 S.n5875 SUB 0.24fF $ **FLOATING
C6522 S.n5876 SUB 0.90fF $ **FLOATING
C6523 S.n5877 SUB 0.05fF $ **FLOATING
C6524 S.t25 SUB 31.97fF
C6525 S.t1130 SUB 0.02fF
C6526 S.n5878 SUB 0.01fF $ **FLOATING
C6527 S.n5879 SUB 0.25fF $ **FLOATING
C6528 S.t580 SUB 0.02fF
C6529 S.n5881 SUB 1.18fF $ **FLOATING
C6530 S.n5882 SUB 0.05fF $ **FLOATING
C6531 S.t999 SUB 0.02fF
C6532 S.n5883 SUB 0.63fF $ **FLOATING
C6533 S.n5884 SUB 0.60fF $ **FLOATING
C6534 S.n5885 SUB 1.48fF $ **FLOATING
C6535 S.n5886 SUB 0.02fF $ **FLOATING
C6536 S.n5887 SUB 0.01fF $ **FLOATING
C6537 S.n5888 SUB 0.01fF $ **FLOATING
C6538 S.n5889 SUB 0.01fF $ **FLOATING
C6539 S.n5890 SUB 0.01fF $ **FLOATING
C6540 S.n5891 SUB 0.02fF $ **FLOATING
C6541 S.n5892 SUB 0.02fF $ **FLOATING
C6542 S.n5893 SUB 0.04fF $ **FLOATING
C6543 S.n5894 SUB 0.16fF $ **FLOATING
C6544 S.n5895 SUB 0.10fF $ **FLOATING
C6545 S.n5896 SUB 0.16fF $ **FLOATING
C6546 S.n5897 SUB 0.14fF $ **FLOATING
C6547 S.n5898 SUB 0.27fF $ **FLOATING
C6548 S.n5899 SUB 0.24fF $ **FLOATING
C6549 S.n5900 SUB 4.64fF $ **FLOATING
C6550 S.n5901 SUB 9.18fF $ **FLOATING
C6551 S.n5902 SUB 9.19fF $ **FLOATING
C6552 S.n5903 SUB 9.19fF $ **FLOATING
C6553 S.n5904 SUB 9.19fF $ **FLOATING
C6554 S.n5905 SUB 9.19fF $ **FLOATING
C6555 S.n5906 SUB 9.17fF $ **FLOATING
C6556 S.n5907 SUB 9.19fF $ **FLOATING
C6557 S.n5908 SUB 9.19fF $ **FLOATING
C6558 S.n5909 SUB 9.28fF $ **FLOATING
C6559 S.n5910 SUB 17.58fF $ **FLOATING
.ends

