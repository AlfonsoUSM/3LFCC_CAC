* NGSPICE file created from mag_files/POSTLAYOUT/nmos_flat_36x36.ext - technology: sky130A

.subckt mag_files/POSTLAYOUT/nmos_flat_36x36
X0 D G S.t2590 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=3.50005e+15p pd=2.37328e+10u as=0p ps=0u w=4.38e+06u l=500000u
X1 D G S.t2589 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 D G S.t2588 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D G S.t2587 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 D G S.t2586 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 S.t2585 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 D G S.t2584 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 D G S.t2583 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 D G S.t2582 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 S.t2581 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 D G S.t2580 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 D G S.t2579 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 D G S.t2578 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 S.t2577 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 D G S.t2576 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D G S.t2575 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 D G S.t2574 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 S.t2573 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 S.t2572 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 S.t2571 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 D G S.t2570 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 S.t2569 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 S.t2568 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D G S.t2567 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 S.t2566 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 D G S.t2565 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D G S.t2564 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 D G S.t2563 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D G S.t2562 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 D G S.t2561 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 D G S.t2560 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 D G S.t2559 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 D G S.t2558 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 D G S.t2557 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 D G S.t2556 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 D G S.t2555 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 S.t2554 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 D G S.t2553 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 D G S.t2552 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 D G S.t2551 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D G S.t2550 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 D G S.t2549 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 D G S.t2548 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 D G S.t2547 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 D G S.t2546 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 D G S.t2545 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 S.t2544 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 D G S.t2543 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 D G S.t2542 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 D G S.t2541 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 D G S.t2540 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D G S.t2539 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 D G S.t2538 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 D G S.t2537 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 D G S.t2536 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 S.t2535 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 D G S.t2534 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 D G S.t2533 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 S.t2532 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D G S.t2531 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 D G S.t2530 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 S.t2529 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 D G S.t2528 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 S.t2527 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 D G S.t2526 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 D G S.t2525 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 D G S.t2524 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 S.t2523 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 D G S.t2522 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 S.t2521 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 D G S.t2520 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D G S.t2519 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 D G S.t2518 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 D G S.t2517 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 S.t2516 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 D G S.t2515 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 S.t2514 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 D G S.t2513 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 D G S.t2512 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 D G S.t2511 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 D G S.t2510 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 S.t2509 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 S.t2508 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 S.t2507 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 D G S.t2506 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 D G S.t2505 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 S.t2504 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 D G S.t2503 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 S.t2502 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 D G S.t2501 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D G S.t2500 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 D G S.t2499 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 D G S.t2498 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 S.t2497 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 S.t2496 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 D G S.t2495 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D G S.t2494 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 S.t2493 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 D G S.t2492 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 D G S.t2491 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 D G S.t2490 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 D G S.t2489 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 D G S.t2488 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 D G S.t2487 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 S.t2486 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 D G S.t2485 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 D G S.t2484 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 D G S.t2483 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 D G S.t2482 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 D G S.t2481 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D G S.t2480 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 S.t2479 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 D G S.t2478 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 S.t2477 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 D G S.t2476 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 D G S.t2475 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 S.t2474 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 D G S.t2473 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 S.t2472 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 S.t2471 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 D G S.t2470 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 D G S.t2469 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 S.t2468 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 S.t2467 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 D G S.t2466 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 D G S.t2465 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 S.t2464 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 D G S.t2463 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 S.t2462 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 D G S.t2461 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 S.t2460 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 D G S.t2459 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 S.t2458 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t2457 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 D G S.t2456 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t2455 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 D G S.t2454 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 S.t2453 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 S.t2452 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 D G S.t2451 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 D G S.t2450 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 S.t2449 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 S.t2448 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 S.t2447 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 S.t2446 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 D G S.t2445 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 D G S.t2444 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 D G S.t2443 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 D G S.t2442 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 S.t2441 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 D G S.t2440 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 D G S.t2439 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 S.t2438 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 D G S.t2437 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 S.t2436 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 D G S.t2435 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 D G S.t2434 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 S.t2433 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 S.t2432 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 D G S.t2431 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 D G S.t2430 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 S.t2429 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 S.t2428 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 S.t2427 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 S.t2426 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 D G S.t2425 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 S.t2424 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 S.t2423 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 S.t2422 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 D G S.t2421 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 S.t2420 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 S.t2419 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 S.t2418 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 S.t2417 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 D G S.t2416 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 S.t2415 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 D G S.t2414 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 S.t2413 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 S.t2412 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 D G S.t2411 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 S.t2410 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 D G S.t2409 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 S.t2408 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 S.t2407 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 S.t2406 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 S.t2405 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 D G S.t2404 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 S.t2403 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 D G S.t2402 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 S.t2401 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 D G S.t2400 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 D G S.t2399 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 S.t2398 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 D G S.t2397 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 D G S.t2396 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 S.t2395 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 D G S.t2394 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 D G S.t2393 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 S.t2392 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 S.t2391 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 D G S.t2390 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 S.t2389 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 S.t2388 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 S.t2387 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 D G S.t2386 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 S.t2385 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 D G S.t2384 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 S.t2383 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 S.t2382 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 D G S.t2381 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 S.t2380 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 S.t2379 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 S.t2378 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 S.t2377 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 D G S.t2376 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 S.t2375 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 S.t2374 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 S.t2373 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 S.t2372 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 D G S.t2371 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 D G S.t2370 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 S.t2369 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 S.t2368 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 S.t2367 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 S.t2366 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 S.t2365 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 S.t2364 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 D G S.t2363 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 D G S.t2362 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 D G S.t2361 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 S.t2360 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 S.t2359 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 D G S.t2358 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 S.t2357 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 S.t2356 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 D G S.t2355 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 S.t2354 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 S.t2353 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 S.t2352 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 D G S.t2351 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 S.t2350 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 D G S.t2349 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 S.t2348 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 D G S.t2347 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 S.t2346 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 S.t2345 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 D G S.t2344 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 D G S.t2343 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 S.t2342 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 S.t2341 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 S.t2340 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 D G S.t2339 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 D G S.t2338 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 S.t2337 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 S.t2336 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 S.t2335 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 D G S.t2334 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 S.t2333 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 S.t2332 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 D G S.t2331 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 D G S.t2330 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 S.t2329 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 S.t2328 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 D G S.t2327 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 S.t2326 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 S.t2325 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 D G S.t2324 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 S.t2323 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 S.t2322 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 S.t2321 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 D G S.t2320 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 S.t2319 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 S.t2318 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 S.t2317 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 D G S.t2316 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 S.t2315 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 S.t2314 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 S.t2313 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 S.t2312 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 S.t2311 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 S.t2310 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 S.t2309 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 S.t2308 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D G S.t2307 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 S.t2306 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 S.t2305 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 D G S.t2304 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 D G S.t2303 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 D G S.t2302 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 D G S.t2301 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 D G S.t2300 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 S.t2299 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 D G S.t2298 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 D G S.t2297 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 D G S.t2296 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 D G S.t2295 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 D G S.t2294 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 S.t2293 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 S.t2292 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 S.t2291 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 D G S.t2290 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 S.t2289 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 D G S.t2288 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 S.t2287 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 D G S.t2286 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 S.t2285 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 D G S.t2284 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 D G S.t2283 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 D G S.t2282 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 S.t2281 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 S.t2280 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 D G S.t2279 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 S.t2278 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 S.t2277 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 D G S.t2276 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 D G S.t2275 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 S.t2274 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 D G S.t2273 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 S.t2272 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 S.t2271 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 S.t2270 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 S.t2269 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 D G S.t2268 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 S.t2267 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 D G S.t2266 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 D G S.t2265 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 D G S.t2264 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 D G S.t2263 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 D G S.t2262 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 D G S.t2261 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 D G S.t2260 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 D G S.t2259 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 S.t2258 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 D G S.t2257 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 S.t2256 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 D G S.t2255 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 S.t2254 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 S.t2253 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 D G S.t2252 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 S.t2251 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 S.t2250 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 D G S.t2249 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 D G S.t2248 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 S.t2247 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 S.t2246 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 D G S.t2245 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 S.t2244 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 D G S.t2243 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 D G S.t2242 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t2241 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 D G S.t2240 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 D G S.t2239 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 D G S.t2238 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 S.t2237 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 S.t2236 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 D G S.t2235 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 D G S.t2234 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 S.t2233 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 D G S.t2232 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 S.t2231 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 D G S.t2230 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 D G S.t2229 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 S.t2228 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 S.t2227 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 D G S.t2226 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 D G S.t2225 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 S.t2224 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 D G S.t2223 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 D G S.t2222 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 D G S.t2221 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 S.t2220 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 D G S.t2219 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 S.t2218 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 D G S.t2217 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 D G S.t2216 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 S.t2215 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 D G S.t2214 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 D G S.t2213 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 S.t2212 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 S.t2211 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 S.t2210 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 D G S.t2209 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 D G S.t2208 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 S.t2207 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 D G S.t2206 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 S.t2205 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 S.t2204 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 D G S.t2203 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 D G S.t2202 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 S.t2201 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 D G S.t2200 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 S.t2199 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 D G S.t2198 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 S.t2197 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 D G S.t2196 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 S.t2195 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 D G S.t2194 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 S.t2193 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 D G S.t2192 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 S.t2191 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 S.t2190 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 D G S.t2189 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 D G S.t2188 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 S.t2187 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 S.t2186 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 S.t2185 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 D G S.t2184 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 S.t2183 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 S.t2182 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 D G S.t2181 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 D G S.t2180 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 S.t2179 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 S.t2178 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 D G S.t2177 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 S.t2176 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 D G S.t2175 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 D G S.t2174 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 D G S.t2173 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 S.t2172 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 S.t2171 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 D G S.t2170 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 S.t2169 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 S.t2168 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 S.t2167 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 D G S.t2166 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 S.t2165 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 D G S.t2164 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 D G S.t2163 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 D G S.t2162 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 S.t2161 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 D G S.t2160 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 S.t2159 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 D G S.t2158 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 D G S.t2157 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 D G S.t2156 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 S.t2155 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 D G S.t2154 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 S.t2153 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 S.t2152 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 S.t2151 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 D G S.t2150 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 S.t2149 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 D G S.t2148 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 S.t2147 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 D G S.t2146 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 D G S.t2145 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 S.t2144 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 S.t2143 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 S.t2142 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 S.t2141 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 D G S.t2140 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 S.t2139 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 D G S.t2138 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 S.t2137 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 S.t2136 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 D G S.t2135 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 S.t2134 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 D G S.t2133 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 D G S.t2132 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 S.t2131 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 S.t2130 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 D G S.t2129 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 S.t2128 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t2127 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 D G S.t2126 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 S.t2125 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 S.t2124 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 S.t2123 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 S.t2122 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 D G S.t2121 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 S.t2120 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 D G S.t2119 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 S.t2118 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 D G S.t2117 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 S.t2116 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 D G S.t2115 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 S.t2114 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 S.t2113 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 D G S.t2112 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 D G S.t2111 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 D G S.t2110 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 D G S.t2109 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 S.t2108 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 D G S.t2107 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 D G S.t2106 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 D G S.t2105 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 S.t2104 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 S.t2103 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 S.t2102 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 S.t2101 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 D G S.t2100 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 S.t2099 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 S.t2098 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 D G S.t2097 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t2096 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 S.t2095 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 D G S.t2094 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 D G S.t2093 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 S.t2092 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 D G S.t2091 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 S.t2090 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 D G S.t2089 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 D G S.t2088 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 S.t2087 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 S.t2086 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 D G S.t2085 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 D G S.t2084 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 D G S.t2083 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 S.t2082 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 D G S.t2081 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t2080 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 D G S.t2079 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 D G S.t2078 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 D G S.t2077 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 D G S.t2076 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 S.t2075 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 S.t2074 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 D G S.t2073 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 D G S.t2072 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 D G S.t2071 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 S.t2070 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 S.t2069 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 D G S.t2068 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 S.t2067 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 S.t2066 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 D G S.t2065 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 D G S.t2064 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 D G S.t2063 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 D G S.t2062 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 S.t2061 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 S.t2060 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D G S.t2059 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 D G S.t2058 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 D G S.t2057 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 D G S.t2056 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 D G S.t2055 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 D G S.t2054 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 D G S.t2053 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 S.t2052 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 S.t2051 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 D G S.t2050 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 S.t2049 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 D G S.t2048 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 S.t2047 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 S.t2046 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t2045 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 D G S.t2044 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 S.t2043 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 S.t2042 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 D G S.t2041 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 S.t2040 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 D G S.t2039 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 D G S.t2038 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 S.t2037 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 D G S.t2036 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 S.t2035 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 S.t2034 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 D G S.t2033 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 S.t2032 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 D G S.t2031 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 S.t2030 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 S.t2029 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 D G S.t2028 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 S.t2027 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 D G S.t2026 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 S.t2025 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 D G S.t2024 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 D G S.t2023 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 D G S.t2022 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 S.t2021 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 S.t2020 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 S.t2019 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 D G S.t2018 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 S.t2017 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 D G S.t2016 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 S.t2015 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 D G S.t2014 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 D G S.t2013 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 S.t2012 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 D G S.t2011 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 D G S.t2010 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 S.t2009 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 D G S.t2008 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 S.t2007 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 D G S.t2006 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 D G S.t2005 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 S.t2004 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 D G S.t2003 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 D G S.t2002 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 D G S.t2001 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 D G S.t2000 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 D G S.t1999 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 D G S.t1998 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 D G S.t1997 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 S.t1996 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 S.t1995 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 S.t1994 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 S.t1993 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 D G S.t1992 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 D G S.t1991 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 S.t1990 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D G S.t1989 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 D G S.t1988 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 S.t1987 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 S.t1986 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 S.t1985 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 D G S.t1984 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 D G S.t1983 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 D G S.t1982 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 D G S.t1981 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 D G S.t1980 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 D G S.t1979 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 D G S.t1978 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 S.t1977 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 S.t1976 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 S.t1975 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 S.t1974 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 D G S.t1973 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 D G S.t1972 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 D G S.t1971 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 D G S.t1970 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 S.t1969 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 D G S.t1968 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 S.t1967 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 S.t1966 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 D G S.t1965 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 D G S.t1964 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 S.t1963 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 S.t1962 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 S.t1961 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 S.t1960 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 S.t1959 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 S.t1958 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 D G S.t1957 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 S.t1956 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 S.t1955 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 S.t1954 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 S.t1953 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 D G S.t1952 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 D G S.t1951 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 D G S.t1950 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 S.t1949 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 D G S.t1948 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 D G S.t1947 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 D G S.t1946 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 S.t1945 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 S.t1944 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 D G S.t1943 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 S.t1942 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 D G S.t1941 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 D G S.t1940 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 D G S.t1939 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 D G S.t1938 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 D G S.t1937 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 S.t1936 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 S.t1935 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 D G S.t1934 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 D G S.t1933 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 D G S.t1932 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 S.t1931 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 S.t1930 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 S.t1929 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 S.t1928 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 D G S.t1927 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 S.t1926 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 S.t1925 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 S.t1924 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 D G S.t1923 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 D G S.t1922 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 S.t1921 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 S.t1920 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 D G S.t1919 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 D G S.t1918 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 D G S.t1917 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 S.t1916 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 S.t1915 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 S.t1914 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 D G S.t1913 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 D G S.t1912 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 S.t1911 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 S.t1910 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 S.t1909 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 D G S.t1908 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 S.t1907 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 S.t1906 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 S.t1905 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 D G S.t1904 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 S.t1903 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 S.t1902 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 D G S.t1901 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 S.t1900 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 D G S.t1899 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 S.t1898 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 D G S.t1897 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 S.t1896 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 S.t1895 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 S.t1894 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 S.t1893 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 S.t1892 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 S.t1891 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 S.t1890 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 S.t1889 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 S.t1888 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 D G S.t1887 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 S.t1886 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 D G S.t1885 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 S.t1884 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 D G S.t1883 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 D G S.t1882 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 S.t1881 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 S.t1880 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 D G S.t1879 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 S.t1878 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 S.t1877 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 S.t1876 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 D G S.t1875 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 D G S.t1874 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 D G S.t1873 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 D G S.t1872 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 S.t1871 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 S.t1870 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 D G S.t1869 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 D G S.t1868 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 S.t1867 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 S.t1866 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 D G S.t1865 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 S.t1864 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 D G S.t1863 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 D G S.t1862 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 S.t1861 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 S.t1860 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 S.t1859 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 S.t1858 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 D G S.t1857 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 S.t1856 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 S.t1855 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 S.t1854 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 S.t1853 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 S.t1852 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 S.t1851 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 S.t1850 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 S.t1849 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 S.t1848 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 S.t1847 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 S.t1846 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 S.t1845 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 S.t1844 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 D G S.t1843 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 D G S.t1842 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 S.t1841 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 S.t1840 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 S.t1839 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 D G S.t1838 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 S.t1837 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 D G S.t1836 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 S.t1835 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 S.t1834 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 S.t1833 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 S.t1832 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 S.t1831 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 S.t1830 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 D G S.t1829 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 S.t1828 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 S.t1827 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 S.t1826 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 D G S.t1825 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 S.t1824 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 S.t1823 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 D G S.t1822 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 D G S.t1821 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 S.t1820 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 S.t1819 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 S.t1818 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 D G S.t1817 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 S.t1816 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 S.t1815 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 D G S.t1814 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 D G S.t1813 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 D G S.t1812 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 S.t1811 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 D G S.t1810 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 D G S.t1809 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 S.t1808 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 S.t1807 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 S.t1806 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 D G S.t1805 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 S.t1804 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 S.t1803 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 S.t1802 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 D G S.t1801 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 S.t1800 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 S.t1799 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 S.t1798 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 D G S.t1797 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 D G S.t1796 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 D G S.t1795 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 D G S.t1794 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 S.t1793 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 S.t1792 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 S.t1791 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 D G S.t1790 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 D G S.t1789 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 D G S.t1788 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 S.t1787 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 D G S.t1786 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 D G S.t1785 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 D G S.t1784 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 S.t1783 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 D G S.t1782 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 S.t1781 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 S.t1780 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 D G S.t1779 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 D G S.t1778 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 D G S.t1777 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 S.t1776 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 D G S.t1775 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 D G S.t1774 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 D G S.t1773 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 S.t1772 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 D G S.t1771 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 D G S.t1770 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 D G S.t1769 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 D G S.t1768 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 S.t1767 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 S.t1766 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 D G S.t1765 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 D G S.t1764 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 D G S.t1763 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 S.t1762 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 D G S.t1761 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 S.t1760 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 S.t1759 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 S.t1758 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 D G S.t1757 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 D G S.t1756 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 S.t1755 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 S.t1754 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 S.t1753 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 S.t1752 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 D G S.t1751 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 D G S.t1750 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 S.t1749 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 S.t1748 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 S.t1747 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 S.t1746 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 D G S.t1745 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 D G S.t1744 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 D G S.t1743 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 D G S.t1742 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 D G S.t1741 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 D G S.t1740 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 S.t1739 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 D G S.t1738 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 S.t1737 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 S.t1736 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 D G S.t1735 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 D G S.t1734 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 S.t1733 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 S.t1732 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 D G S.t1731 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 S.t1730 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 D G S.t1729 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 D G S.t1728 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 S.t1727 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 S.t1726 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 D G S.t1725 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 D G S.t1724 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 S.t1723 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 D G S.t1722 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 D G S.t1721 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 D G S.t1720 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 D G S.t1719 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 D G S.t1718 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 D G S.t1717 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 D G S.t1716 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 D G S.t1715 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 D G S.t1714 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 D G S.t1713 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 D G S.t1712 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 S.t1711 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 D G S.t1710 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 D G S.t1709 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 S.t1708 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 D G S.t1707 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 S.t1706 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 D G S.t1705 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 D G S.t1704 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 D G S.t1703 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 D G S.t1702 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 D G S.t1701 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 D G S.t1700 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 D G S.t1699 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 D G S.t1698 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 S.t1697 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 S.t1696 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 S.t1695 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 D G S.t1694 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 S.t1693 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 D G S.t1692 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 D G S.t1691 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 D G S.t1690 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 D G S.t1689 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 D G S.t1688 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 D G S.t1687 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 D G S.t1686 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 D G S.t1685 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 D G S.t1684 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 D G S.t1683 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 D G S.t1682 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 D G S.t1681 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 D G S.t1680 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 D G S.t1679 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 S.t1678 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 S.t1677 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 D G S.t1676 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 D G S.t1675 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 D G S.t1674 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 D G S.t1673 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 S.t1672 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 S.t1671 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 D G S.t1670 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 D G S.t1669 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 D G S.t1668 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 D G S.t1667 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 D G S.t1666 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 D G S.t1665 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 S.t1664 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 D G S.t1663 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 D G S.t1662 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 S.t1661 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 D G S.t1660 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 S.t1659 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 D G S.t1658 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 D G S.t1657 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 D G S.t1656 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 D G S.t1655 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 S.t1654 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 S.t1653 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 D G S.t1652 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 S.t1651 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 D G S.t1650 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 D G S.t1649 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 S.t1648 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 D G S.t1647 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 S.t1646 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 D G S.t1645 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 D G S.t1644 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 S.t1643 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 D G S.t1642 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 S.t1641 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 D G S.t1640 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 S.t1639 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 S.t1638 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 D G S.t1637 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 S.t1636 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 D G S.t1635 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 D G S.t1634 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 S.t1633 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 S.t1632 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 D G S.t1631 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 D G S.t1630 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 S.t1629 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 D G S.t1628 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 S.t1627 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 S.t1626 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 D G S.t1625 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 D G S.t1624 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 S.t1623 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 S.t1622 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 D G S.t1621 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 S.t1620 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 S.t1619 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 D G S.t1618 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 S.t1617 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 D G S.t1616 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 D G S.t1615 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 S.t1614 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 D G S.t1613 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 D G S.t1612 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 D G S.t1611 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 D G S.t1610 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 D G S.t1609 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 S.t1608 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 D G S.t1607 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 S.t1606 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 D G S.t1605 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 D G S.t1604 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 S.t1603 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 S.t1602 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 S.t1601 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 D G S.t1600 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 D G S.t1599 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 S.t1598 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 D G S.t1597 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 D G S.t1596 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 D G S.t1595 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 S.t1594 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 S.t1593 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 S.t1592 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 D G S.t1591 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 S.t1590 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 S.t1589 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 S.t1588 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 D G S.t1587 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 S.t1586 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 S.t1585 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 S.t1584 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 D G S.t1583 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 D G S.t1582 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 S.t1581 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 S.t1580 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 S.t1579 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 S.t1578 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 D G S.t1577 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 S.t1576 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 D G S.t1575 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 S.t1574 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 D G S.t1573 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 S.t1572 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 D G S.t1571 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 D G S.t1570 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 S.t1569 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 S.t1568 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 D G S.t1567 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 S.t1566 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 S.t1565 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 S.t1564 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 S.t1563 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 S.t1562 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 S.t1561 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 D G S.t1560 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 S.t1559 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 D G S.t1558 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 S.t1557 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 D G S.t1556 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 S.t1555 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 S.t1554 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 S.t1553 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 D G S.t1552 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 S.t1551 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 D G S.t1550 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 S.t1549 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 S.t1548 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 D G S.t1547 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 D G S.t1546 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 S.t1545 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 S.t1544 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 S.t1543 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 D G S.t1542 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 S.t1541 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 S.t1540 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 D G S.t1539 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 D G S.t1538 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 S.t1537 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 S.t1536 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 S.t1535 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 S.t1534 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 D G S.t1533 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 D G S.t1532 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 S.t1531 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 D G S.t1530 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 S.t1529 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 S.t1528 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 D G S.t1527 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 S.t1526 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 S.t1525 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 S.t1524 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 S.t1523 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 S.t1522 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 S.t1521 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 S.t1520 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 S.t1519 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 S.t1518 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 S.t1517 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 S.t1516 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 S.t1515 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 D G S.t1514 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 D G S.t1513 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 S.t1512 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 S.t1511 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 S.t1510 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 S.t1509 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 S.t1508 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 S.t1507 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 D G S.t1506 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 D G S.t1505 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 S.t1504 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 D G S.t1503 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 S.t1502 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 D G S.t1501 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 S.t1500 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 S.t1499 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 D G S.t1498 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 D G S.t1497 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 S.t1496 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 S.t1495 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 S.t1494 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 D G S.t1493 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 D G S.t1492 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 S.t1491 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 D G S.t1490 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 D G S.t1489 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 D G S.t1488 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 D G S.t1487 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1104 D G S.t1486 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1105 D G S.t1485 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1106 D G S.t1484 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1107 S.t1483 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1108 D G S.t1482 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1109 S.t1481 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1110 S.t1480 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1111 D G S.t1479 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1112 S.t1478 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1113 S.t1477 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1114 S.t1476 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1115 S.t1475 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1116 D G S.t1474 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1117 D G S.t1473 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1118 D G S.t1472 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1119 D G S.t1471 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1120 S.t1470 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1121 S.t1469 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1122 D G S.t1468 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1123 S.t1467 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1124 D G S.t1466 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1125 S.t1465 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1126 D G S.t1464 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1127 D G S.t1463 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1128 D G S.t1462 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1129 D G S.t1461 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1130 S.t1460 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1131 S.t1459 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1132 S.t1458 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1133 S.t1457 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1134 D G S.t1456 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1135 S.t1455 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1136 S.t1454 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1137 S.t1453 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1138 S.t1452 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1139 D G S.t1451 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1140 S.t1450 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1141 D G S.t1449 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1142 D G S.t1448 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1143 D G S.t1447 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1144 S.t1446 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1145 S.t1445 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1146 D G S.t1444 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1147 S.t1443 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1148 D G S.t1442 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1149 D G S.t1441 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1150 D G S.t1440 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1151 D G S.t1439 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1152 S.t1438 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1153 S.t1437 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1154 D G S.t1436 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1155 D G S.t1435 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1156 D G S.t1434 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1157 D G S.t1433 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1158 D G S.t1432 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1159 D G S.t1431 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1160 D G S.t1430 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1161 D G S.t1429 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1162 D G S.t1428 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1163 S.t1427 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1164 D G S.t1426 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1165 S.t1425 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1166 D G S.t1424 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1167 S.t1423 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1168 D G S.t1422 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1169 S.t1421 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1170 D G S.t1420 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1171 D G S.t1419 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1172 S.t1418 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1173 D G S.t1417 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1174 S.t1416 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1175 S.t1415 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1176 S.t1414 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1177 S.t1413 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1178 D G S.t1412 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1179 D G S.t1411 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1180 S.t1410 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1181 D G S.t1409 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1182 S.t1408 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1183 D G S.t1407 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1184 D G S.t1406 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1185 D G S.t1405 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1186 D G S.t1404 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1187 D G S.t1403 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1188 D G S.t1402 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1189 D G S.t1401 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1190 S.t1400 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1191 D G S.t1399 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1192 S.t1398 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1193 S.t1397 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1194 S.t1396 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1195 S.t1395 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1196 S.t1394 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1197 D G S.t1393 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1198 S.t1392 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1199 D G S.t1391 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1200 D G S.t1390 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1201 S.t1389 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1202 S.t1388 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1203 S.t1387 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1204 D G S.t1386 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1205 S.t1385 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1206 D G S.t1384 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1207 D G S.t1383 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1208 S.t1382 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1209 D G S.t1381 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1210 D G S.t1380 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1211 D G S.t1379 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1212 S.t1378 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1213 S.t1377 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1214 S.t1376 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1215 S.t1375 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1216 D G S.t1374 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1217 D G S.t1373 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1218 D G S.t1372 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1219 S.t1371 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1220 D G S.t1370 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1221 S.t1369 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1222 S.t1368 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1223 S.t1367 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1224 S.t1366 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1225 D G S.t1365 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1226 D G S.t1364 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1227 D G S.t1363 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1228 S.t1362 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1229 D G S.t1361 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1230 D G S.t1360 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1231 D G S.t1359 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1232 S.t1358 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1233 D G S.t1357 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1234 D G S.t1356 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1235 D G S.t1355 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1236 S.t1354 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1237 D G S.t1353 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1238 S.t1352 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1239 D G S.t1351 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1240 D G S.t1350 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1241 S.t1349 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1242 D G S.t1348 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1243 D G S.t1347 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1244 S.t1346 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1245 D G S.t1345 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1246 S.t1344 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1247 D G S.t1343 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1248 D G S.t1342 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1249 S.t1341 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1250 D G S.t1340 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1251 S.t1339 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1252 D G S.t1338 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1253 S.t1337 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1254 D G S.t1336 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1255 S.t1335 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1256 S.t1334 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1257 S.t1333 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1258 D G S.t1332 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1259 D G S.t1331 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1260 S.t1330 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1261 D G S.t1329 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1262 S.t1328 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1263 D G S.t1327 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1264 D G S.t1326 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1265 S.t1325 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1266 D G S.t1324 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1267 S.t1323 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1268 S.t1322 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1269 S.t1321 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1270 D G S.t1320 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1271 D G S.t1319 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1272 S.t1318 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1273 S.t1317 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1274 S.t1316 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1275 D G S.t1315 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1276 S.t1314 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1277 D G S.t1313 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1278 S.t1312 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1279 D G S.t1311 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1280 D G S.t1310 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1281 S.t1309 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1282 D G S.t1308 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1283 S.t1307 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1284 S.t1306 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1285 S.t1305 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1286 D G S.t1304 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1287 S.t1303 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1288 S.t1302 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1289 D G S.t1301 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1290 S.t1300 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1291 S.t1299 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1292 D G S.t1298 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1293 S.t1297 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1294 S.t1296 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1295 D G S.t1295 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1296 D G S.t1294 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1297 D G S.t1293 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1298 S.t1292 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1299 S.t1291 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1300 D G S.t1290 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1301 S.t1289 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1302 D G S.t1288 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1303 S.t1287 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1304 D G S.t1286 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1305 S.t1285 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1306 S.t1284 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1307 D G S.t1283 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1308 D G S.t1282 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1309 D G S.t1281 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1310 S.t1280 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1311 S.t1279 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1312 D G S.t1278 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1313 S.t1277 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1314 D G S.t1276 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1315 D G S.t1275 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1316 D G S.t1274 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1317 S.t1273 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1318 S.t1272 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1319 S.t1271 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1320 D G S.t1270 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1321 D G S.t1269 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1322 D G S.t1268 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1323 D G S.t1267 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1324 S.t1266 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1325 D G S.t1265 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1326 S.t1264 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1327 D G S.t1263 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1328 D G S.t1262 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1329 S.t1261 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1330 D G S.t1260 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1331 S.t1259 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1332 S.t1258 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1333 D G S.t1257 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1334 S.t1256 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1335 S.t1255 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1336 D G S.t1254 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1337 D G S.t1253 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1338 S.t1252 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1339 D G S.t1251 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1340 D G S.t1250 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1341 S.t1249 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1342 D G S.t1248 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1343 D G S.t1247 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1344 D G S.t1246 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1345 S.t1245 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1346 D G S.t1244 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1347 S.t1243 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1348 S.t1242 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1349 D G S.t1241 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1350 D G S.t1240 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1351 D G S.t1239 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1352 S.t1238 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1353 S.t1237 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1354 S.t1236 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1355 D G S.t1235 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1356 S.t1234 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1357 S.t1233 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1358 D G S.t1232 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1359 S.t1231 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1360 S.t1230 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1361 D G S.t1229 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1362 S.t1228 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1363 D G S.t1227 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1364 D G S.t1226 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1365 D G S.t1225 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1366 S.t1224 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1367 S.t1223 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1368 D G S.t1222 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1369 D G S.t1221 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1370 S.t1220 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1371 D G S.t1219 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1372 S.t1218 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1373 S.t1217 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1374 D G S.t1216 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1375 D G S.t1215 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1376 S.t1214 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1377 D G S.t1213 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1378 S.t1212 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1379 D G S.t1211 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1380 D G S.t1210 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1381 S.t1209 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1382 D G S.t1208 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1383 D G S.t1207 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1384 S.t1206 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1385 S.t1205 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1386 S.t1204 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1387 D G S.t1203 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1388 S.t1202 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1389 D G S.t1201 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1390 D G S.t1200 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1391 D G S.t1199 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1392 D G S.t1198 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1393 D G S.t1197 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1394 D G S.t1196 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1395 D G S.t1195 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1396 D G S.t1194 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1397 D G S.t1193 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1398 D G S.t1192 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1399 S.t1191 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1400 S.t1190 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1401 S.t1189 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1402 D G S.t1188 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1403 S.t1187 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1404 S.t1186 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1405 D G S.t1185 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1406 D G S.t1184 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1407 D G S.t1183 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1408 S.t1182 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1409 D G S.t1181 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1410 S.t1180 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1411 S.t1179 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1412 S.t1178 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1413 D G S.t1177 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1414 D G S.t1176 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1415 S.t1175 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1416 S.t1174 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1417 D G S.t1173 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1418 D G S.t1172 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1419 S.t1171 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1420 D G S.t1170 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1421 D G S.t1169 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1422 S.t1168 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1423 D G S.t1167 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1424 D G S.t1166 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1425 S.t1165 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1426 S.t1164 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1427 D G S.t1163 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1428 S.t1162 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1429 D G S.t1161 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1430 S.t1160 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1431 D G S.t1159 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1432 D G S.t1158 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1433 S.t1157 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1434 D G S.t1156 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1435 D G S.t1155 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1436 S.t1154 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1437 S.t1153 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1438 S.t1152 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1439 D G S.t1151 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1440 D G S.t1150 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1441 D G S.t1149 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1442 D G S.t1148 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1443 D G S.t1147 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1444 S.t1146 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1445 S.t1145 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1446 S.t1144 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1447 D G S.t1143 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1448 S.t1142 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1449 D G S.t1141 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1450 S.t1140 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1451 D G S.t1139 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1452 D G S.t1138 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1453 S.t1137 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1454 D G S.t1136 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1455 D G S.t1135 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1456 D G S.t1134 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1457 S.t1133 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1458 S.t1132 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1459 D G S.t1131 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1460 S.t1130 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1461 D G S.t1129 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1462 S.t1128 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1463 D G S.t1127 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1464 S.t1126 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1465 D G S.t1125 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1466 S.t1124 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1467 S.t1123 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1468 S.t1122 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1469 D G S.t1121 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1470 S.t1120 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1471 S.t1119 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1472 D G S.t1118 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1473 D G S.t1117 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1474 D G S.t1116 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1475 D G S.t1115 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1476 S.t1114 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1477 S.t1113 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1478 S.t1112 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1479 D G S.t1111 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1480 D G S.t1110 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1481 D G S.t1109 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1482 S.t1108 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1483 D G S.t1107 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1484 S.t1106 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1485 S.t1105 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1486 S.t1104 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1487 D G S.t1103 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1488 S.t1102 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1489 S.t1101 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1490 S.t1100 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1491 S.t1099 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1492 S.t1098 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1493 D G S.t1097 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1494 S.t1096 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1495 S.t1095 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1496 S.t1094 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1497 S.t1093 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1498 D G S.t1092 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1499 S.t1091 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1500 D G S.t1090 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1501 D G S.t1089 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1502 S.t1088 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1503 S.t1087 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1504 D G S.t1086 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1505 D G S.t1085 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1506 S.t1084 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1507 D G S.t1083 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1508 D G S.t1082 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1509 S.t1081 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1510 D G S.t1080 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1511 D G S.t1079 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1512 S.t1078 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1513 S.t1077 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1514 D G S.t1076 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1515 D G S.t1075 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1516 D G S.t1074 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1517 S.t1073 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1518 D G S.t1072 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1519 S.t1071 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1520 S.t1070 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1521 D G S.t1069 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1522 S.t1068 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1523 S.t1067 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1524 S.t1066 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1525 S.t1065 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1526 D G S.t1064 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1527 S.t1063 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1528 D G S.t1062 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1529 D G S.t1061 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1530 S.t1060 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1531 S.t1059 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1532 D G S.t1058 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1533 D G S.t1057 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1534 S.t1056 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1535 S.t1055 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1536 S.t1054 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1537 S.t1053 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1538 S.t1052 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1539 S.t1051 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1540 S.t1050 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1541 S.t1049 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1542 D G S.t1048 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1543 S.t1047 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1544 S.t1046 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1545 D G S.t1045 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1546 S.t1044 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1547 S.t1043 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1548 D G S.t1042 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1549 S.t1041 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1550 S.t1040 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1551 D G S.t1039 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1552 S.t1038 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1553 D G S.t1037 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1554 D G S.t1036 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1555 S.t1035 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1556 S.t1034 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1557 S.t1033 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1558 S.t1032 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1559 S.t1031 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1560 D G S.t1030 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1561 S.t1029 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1562 S.t1028 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1563 S.t1027 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1564 S.t1026 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1565 S.t1025 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1566 D G S.t1024 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1567 S.t1023 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1568 S.t1022 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1569 D G S.t1021 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1570 D G S.t1020 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1571 S.t1019 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1572 S.t1018 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1573 S.t1017 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1574 S.t1016 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1575 D G S.t1015 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1576 S.t1014 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1577 S.t1013 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1578 S.t1012 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1579 S.t1011 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1580 S.t1010 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1581 S.t1009 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1582 D G S.t1008 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1583 S.t1007 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1584 D G S.t1006 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1585 D G S.t1005 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1586 S.t1004 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1587 S.t1003 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1588 D G S.t1002 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1589 S.t1001 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1590 D G S.t1000 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1591 S.t999 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1592 S.t998 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1593 D G S.t997 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1594 D G S.t996 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1595 S.t995 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1596 D G S.t994 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1597 D G S.t993 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1598 S.t992 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1599 S.t991 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1600 D G S.t990 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1601 S.t989 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1602 S.t988 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1603 S.t987 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1604 S.t986 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1605 S.t985 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1606 S.t984 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1607 S.t983 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1608 S.t982 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1609 D G S.t981 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1610 S.t980 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1611 D G S.t979 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1612 S.t978 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1613 D G S.t977 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1614 S.t976 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1615 S.t975 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1616 S.t974 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1617 D G S.t973 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1618 D G S.t972 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1619 D G S.t971 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1620 D G S.t970 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1621 S.t969 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1622 S.t968 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1623 S.t967 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1624 S.t966 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1625 S.t965 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1626 S.t964 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1627 D G S.t963 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1628 S.t962 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1629 D G S.t961 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1630 S.t960 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1631 S.t959 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1632 S.t958 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1633 D G S.t957 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1634 D G S.t956 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1635 S.t955 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1636 S.t954 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1637 S.t953 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1638 D G S.t952 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1639 D G S.t951 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1640 D G S.t950 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1641 S.t949 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1642 S.t948 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1643 D G S.t947 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1644 D G S.t946 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1645 D G S.t945 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1646 S.t944 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1647 D G S.t943 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1648 S.t942 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1649 S.t941 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1650 D G S.t940 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1651 D G S.t939 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1652 D G S.t938 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1653 S.t937 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1654 D G S.t936 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1655 S.t935 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1656 D G S.t934 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1657 D G S.t933 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1658 S.t932 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1659 S.t931 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1660 D G S.t930 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1661 S.t929 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1662 S.t928 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1663 D G S.t927 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1664 S.t926 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1665 D G S.t925 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1666 D G S.t924 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1667 S.t923 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1668 D G S.t922 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1669 D G S.t921 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1670 D G S.t920 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1671 D G S.t919 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1672 S.t918 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1673 D G S.t917 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1674 D G S.t916 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1675 D G S.t915 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1676 S.t914 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1677 S.t913 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1678 D G S.t912 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1679 S.t911 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1680 D G S.t910 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1681 D G S.t909 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1682 S.t908 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1683 D G S.t907 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1684 S.t906 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1685 D G S.t905 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1686 D G S.t904 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1687 D G S.t903 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1688 D G S.t902 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1689 S.t901 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1690 S.t900 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1691 D G S.t899 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1692 S.t898 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1693 D G S.t897 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1694 D G S.t896 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1695 D G S.t895 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1696 D G S.t894 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1697 S.t893 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1698 S.t892 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1699 D G S.t891 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1700 D G S.t890 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1701 D G S.t889 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1702 D G S.t888 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1703 D G S.t887 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1704 D G S.t886 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1705 S.t885 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1706 D G S.t884 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1707 S.t883 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1708 S.t882 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1709 D G S.t881 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1710 D G S.t880 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1711 D G S.t879 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1712 D G S.t878 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1713 D G S.t877 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1714 S.t876 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1715 S.t875 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1716 D G S.t874 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1717 D G S.t873 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1718 D G S.t872 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1719 D G S.t871 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1720 S.t870 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1721 D G S.t869 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1722 D G S.t868 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1723 D G S.t867 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1724 D G S.t866 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1725 D G S.t865 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1726 S.t864 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1727 D G S.t863 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1728 S.t862 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1729 D G S.t861 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1730 D G S.t860 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1731 S.t859 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1732 S.t858 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1733 D G S.t857 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1734 D G S.t856 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1735 D G S.t855 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1736 S.t854 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1737 D G S.t853 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1738 D G S.t852 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1739 S.t851 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1740 D G S.t850 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1741 D G S.t849 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1742 D G S.t848 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1743 D G S.t847 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1744 D G S.t846 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1745 D G S.t845 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1746 D G S.t844 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1747 D G S.t843 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1748 D G S.t842 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1749 D G S.t841 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1750 D G S.t840 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1751 D G S.t839 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1752 S.t838 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1753 S.t837 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1754 D G S.t836 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1755 D G S.t835 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1756 S.t834 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1757 D G S.t833 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1758 D G S.t832 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1759 S.t831 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1760 D G S.t830 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1761 D G S.t829 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1762 D G S.t828 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1763 S.t827 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1764 D G S.t826 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1765 D G S.t825 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1766 D G S.t824 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1767 S.t823 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1768 S.t822 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1769 D G S.t821 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1770 D G S.t820 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1771 D G S.t819 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1772 S.t818 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1773 S.t817 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1774 D G S.t816 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1775 D G S.t815 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1776 D G S.t814 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1777 D G S.t813 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1778 S.t812 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1779 D G S.t811 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1780 S.t810 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1781 D G S.t809 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1782 S.t808 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1783 D G S.t807 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1784 S.t806 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1785 D G S.t805 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1786 D G S.t804 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1787 S.t803 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1788 S.t802 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1789 D G S.t801 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1790 D G S.t800 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1791 S.t799 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1792 D G S.t798 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1793 S.t797 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1794 S.t796 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1795 D G S.t795 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1796 D G S.t794 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1797 D G S.t793 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1798 S.t792 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1799 D G S.t791 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1800 S.t790 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1801 D G S.t789 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1802 D G S.t788 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1803 S.t787 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1804 D G S.t786 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1805 D G S.t785 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1806 D G S.t784 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1807 S.t783 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1808 S.t782 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1809 S.t781 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1810 S.t780 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1811 D G S.t779 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1812 D G S.t778 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1813 S.t777 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1814 S.t776 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1815 D G S.t775 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1816 D G S.t774 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1817 S.t773 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1818 S.t772 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1819 S.t771 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1820 D G S.t770 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1821 S.t769 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1822 S.t768 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1823 D G S.t767 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1824 D G S.t766 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1825 S.t765 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1826 D G S.t764 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1827 D G S.t763 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1828 S.t762 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1829 D G S.t761 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1830 S.t760 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1831 D G S.t759 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1832 S.t758 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1833 D G S.t757 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1834 S.t756 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1835 S.t755 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1836 D G S.t754 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1837 S.t753 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1838 S.t752 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1839 S.t751 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1840 D G S.t750 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1841 S.t749 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1842 D G S.t748 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1843 D G S.t747 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1844 D G S.t746 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1845 D G S.t745 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1846 S.t744 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1847 D G S.t743 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1848 S.t742 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1849 D G S.t741 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1850 D G S.t740 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1851 S.t739 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1852 S.t738 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1853 S.t737 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1854 D G S.t736 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1855 S.t735 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1856 D G S.t734 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1857 D G S.t733 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1858 D G S.t732 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1859 S.t731 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1860 S.t730 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1861 S.t729 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1862 S.t728 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1863 S.t727 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1864 S.t726 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1865 S.t725 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1866 S.t724 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1867 S.t723 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1868 S.t722 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1869 S.t721 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1870 S.t720 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1871 S.t719 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1872 D G S.t718 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1873 S.t717 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1874 D G S.t716 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1875 D G S.t715 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1876 S.t714 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1877 S.t713 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1878 S.t712 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1879 S.t711 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1880 S.t710 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1881 D G S.t709 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1882 S.t708 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1883 S.t707 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1884 D G S.t706 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1885 D G S.t705 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1886 S.t704 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1887 D G S.t703 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1888 D G S.t702 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1889 S.t701 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1890 S.t700 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1891 D G S.t699 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1892 S.t698 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1893 S.t697 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1894 D G S.t696 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1895 S.t695 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1896 D G S.t694 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1897 S.t693 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1898 S.t692 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1899 S.t691 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1900 S.t690 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1901 S.t689 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1902 D G S.t688 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1903 S.t687 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1904 S.t686 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1905 D G S.t685 S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1906 D G S.t684 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1907 S.t683 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1908 S.t682 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1909 S.t681 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1910 S.t680 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1911 D G S.t679 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1912 D G S.t678 S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1913 D G S.t677 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1914 S.t676 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1915 S.t675 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1916 S.t674 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1917 D G S.t673 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1918 S.t672 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1919 S.t671 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1920 D G S.t670 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1921 S.t669 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1922 S.t668 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1923 S.t667 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1924 D G S.t666 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1925 S.t665 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1926 S.t664 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1927 S.t663 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1928 S.t662 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1929 S.t661 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1930 S.t660 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1931 S.t659 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1932 S.t658 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1933 S.t657 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1934 S.t656 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1935 S.t655 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1936 S.t654 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1937 D G S.t653 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1938 S.t652 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1939 S.t651 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1940 S.t650 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1941 S.t649 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1942 S.t648 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1943 D G S.t647 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1944 D G S.t646 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1945 D G S.t645 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1946 D G S.t644 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1947 D G S.t643 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1948 D G S.t642 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1949 S.t641 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1950 D G S.t640 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1951 D G S.t639 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1952 D G S.t638 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1953 S.t637 G D S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1954 S.t636 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1955 D G S.t635 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1956 D G S.t634 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1957 S.t633 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1958 S.t632 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1959 S.t631 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1960 D G S.t630 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1961 D G S.t629 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1962 S.t628 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1963 S.t627 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1964 S.t626 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1965 D G S.t625 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1966 D G S.t624 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1967 D G S.t623 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1968 S.t622 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1969 D G S.t621 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1970 S.t620 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1971 S.t619 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1972 S.t618 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1973 D G S.t617 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1974 S.t616 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1975 S.t615 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1976 S.t614 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1977 D G S.t613 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1978 D G S.t612 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1979 D G S.t611 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1980 D G S.t610 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1981 D G S.t609 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1982 D G S.t608 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1983 S.t607 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1984 S.t606 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1985 D G S.t605 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1986 D G S.t604 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1987 S.t603 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1988 D G S.t602 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1989 S.t601 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1990 S.t600 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1991 S.t599 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1992 D G S.t598 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1993 S.t597 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1994 S.t596 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1995 S.t595 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1996 S.t594 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1997 S.t593 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1998 D G S.t592 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1999 D G S.t591 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2000 D G S.t590 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2001 D G S.t589 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2002 D G S.t588 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2003 D G S.t587 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2004 D G S.t586 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2005 D G S.t585 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2006 S.t584 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2007 D G S.t583 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2008 S.t582 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2009 S.t581 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2010 D G S.t580 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2011 D G S.t579 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2012 D G S.t578 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2013 D G S.t577 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2014 D G S.t576 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2015 S.t575 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2016 D G S.t574 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2017 D G S.t573 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2018 D G S.t572 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2019 D G S.t571 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2020 D G S.t570 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2021 D G S.t569 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2022 S.t568 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2023 S.t567 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2024 D G S.t566 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2025 D G S.t565 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2026 D G S.t564 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2027 D G S.t563 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2028 S.t562 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2029 D G S.t561 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2030 S.t560 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2031 S.t559 G D S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2032 D G S.t558 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2033 D G S.t557 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2034 S.t556 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2035 S.t555 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2036 D G S.t554 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2037 D G S.t553 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2038 S.t552 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2039 S.t551 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2040 S.t550 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2041 S.t549 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2042 S.t548 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2043 D G S.t547 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2044 D G S.t546 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2045 S.t545 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2046 S.t544 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2047 D G S.t543 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2048 S.t542 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2049 S.t541 G D S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2050 D G S.t540 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2051 D G S.t539 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2052 S.t538 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2053 D G S.t537 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2054 D G S.t536 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2055 S.t535 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2056 D G S.t534 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2057 S.t533 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2058 D G S.t532 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2059 D G S.t531 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2060 D G S.t530 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2061 S.t529 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2062 D G S.t528 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2063 S.t527 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2064 S.t526 G D S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2065 S.t525 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2066 S.t524 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2067 S.t523 G D S.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2068 D G S.t521 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2069 S.t520 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2070 D G S.t519 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2071 D G S.t518 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2072 D G S.t517 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2073 S.t516 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2074 D G S.t515 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2075 D G S.t514 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2076 S.t513 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2077 D G S.t512 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2078 S.t511 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2079 S.t510 G D S.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2080 D G S.t508 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2081 S.t507 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2082 D G S.t506 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2083 D G S.t505 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2084 S.t504 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2085 S.t503 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2086 D G S.t502 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2087 D G S.t501 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2088 D G S.t500 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2089 D G S.t499 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2090 S.t498 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2091 D G S.t497 S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2092 S.t496 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2093 S.t495 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2094 D G S.t494 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2095 D G S.t493 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2096 S.t492 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2097 D G S.t491 S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2098 D G S.t490 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2099 S.t489 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2100 D G S.t488 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2101 D G S.t487 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2102 D G S.t486 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2103 S.t485 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2104 S.t484 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2105 S.t483 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2106 D G S.t482 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2107 D G S.t481 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2108 S.t480 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2109 D G S.t479 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2110 D G S.t478 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2111 D G S.t477 S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2112 S.t476 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2113 S.t475 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2114 S.t474 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2115 S.t473 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2116 S.t472 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2117 S.t471 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2118 D G S.t470 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2119 S.t469 G D S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2120 D G S.t468 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2121 S.t467 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2122 D G S.t466 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2123 S.t465 G D S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2124 D G S.t464 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2125 S.t463 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2126 S.t462 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2127 D G S.t461 S.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2128 D G S.t459 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2129 S.t458 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2130 S.t457 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2131 S.t456 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2132 D G S.t455 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2133 S.t454 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2134 S.t453 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2135 D G S.t452 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2136 S.t451 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2137 S.t450 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2138 S.t449 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2139 D G S.t448 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2140 S.t447 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2141 D G S.t446 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2142 D G S.t445 S.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2143 S.t443 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2144 S.t442 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2145 S.t441 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2146 S.t440 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2147 D G S.t439 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2148 S.t438 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2149 D G S.t437 S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2150 S.t436 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2151 S.t435 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2152 D G S.t434 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2153 S.t433 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2154 D G S.t432 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2155 D G S.t431 S.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2156 D G S.t429 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2157 D G S.t428 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2158 S.t427 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2159 S.t426 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2160 D G S.t425 S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2161 S.t424 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2162 S.t423 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2163 D G S.t422 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2164 D G S.t421 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2165 D G S.t420 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2166 S.t419 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2167 S.t418 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2168 D G S.t417 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2169 S.t416 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2170 D G S.t415 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2171 S.t414 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2172 D G S.t413 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2173 S.t412 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2174 D G S.t411 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2175 D G S.t410 S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2176 D G S.t409 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2177 D G S.t408 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2178 D G S.t407 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2179 D G S.t406 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2180 D G S.t405 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2181 S.t404 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2182 D G S.t403 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2183 S.t402 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2184 D G S.t401 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2185 S.t400 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2186 S.t399 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2187 D G S.t398 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2188 S.t397 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2189 D G S.t396 S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2190 D G S.t395 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2191 D G S.t394 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2192 S.t393 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2193 D G S.t392 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2194 S.t391 G D S.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2195 D G S.t389 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2196 D G S.t388 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2197 D G S.t387 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2198 D G S.t386 S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2199 S.t385 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2200 D G S.t384 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2201 S.t383 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2202 D G S.t382 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2203 S.t381 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2204 S.t380 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2205 D G S.t379 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2206 S.t378 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2207 D G S.t377 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2208 S.t376 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2209 D G S.t375 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2210 S.t374 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2211 S.t373 G D S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2212 S.t372 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2213 D G S.t371 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2214 S.t370 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2215 D G S.t369 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2216 S.t368 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2217 S.t367 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2218 D G S.t366 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2219 S.t365 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2220 D G S.t364 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2221 S.t363 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2222 D G S.t362 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2223 S.t361 G D S.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2224 D G S.t359 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2225 S.t358 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2226 D G S.t357 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2227 S.t356 G D S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2228 D G S.t355 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2229 S.t354 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2230 S.t353 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2231 S.t352 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2232 D G S.t351 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2233 S.t350 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2234 D G S.t349 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2235 S.t348 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2236 D G S.t347 S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2237 S.t346 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2238 S.t345 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2239 D G S.t344 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2240 D G S.t343 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2241 D G S.t342 S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2242 D G S.t341 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2243 D G S.t340 S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2244 D G S.t339 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2245 S.t338 G D S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2246 D G S.t337 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2247 S.t336 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2248 D G S.t335 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2249 D G S.t334 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2250 S.t333 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2251 D G S.t332 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2252 D G S.t331 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2253 D G S.t330 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2254 D G S.t329 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2255 S.t328 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2256 S.t327 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2257 S.t326 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2258 S.t325 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2259 D G S.t324 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2260 D G S.t323 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2261 D G S.t322 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2262 D G S.t321 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2263 D G S.t319 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2264 D G S.t318 S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2265 D G S.t317 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2266 D G S.t316 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2267 D G S.t315 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2268 D G S.t314 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2269 S.t313 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2270 S.t312 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2271 S.t311 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2272 D G S.t310 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2273 D G S.t309 S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2274 D G S.t308 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2275 D G S.t307 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2276 S.t306 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2277 D G S.t305 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2278 D G S.t304 S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2279 S.t303 G D S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2280 S.t302 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2281 S.t301 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2282 D G S.t300 S.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2283 S.t298 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2284 D G S.t297 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2285 D G S.t296 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2286 D G S.t295 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2287 S.t294 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2288 S.t293 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2289 S.t292 G D S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2290 S.t291 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2291 S.t290 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2292 D G S.t289 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2293 S.t288 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2294 D G S.t287 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2295 D G S.t286 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2296 D G S.t285 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2297 D G S.t284 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2298 S.t283 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2299 D G S.t282 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2300 D G S.t281 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2301 D G S.t280 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2302 S.t279 G D S.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2303 S.t277 G D S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2304 S.t276 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2305 D G S.t275 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2306 D G S.t274 S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2307 S.t273 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2308 S.t272 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2309 D G S.t271 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2310 S.t270 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2311 D G S.t269 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2312 S.t268 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2313 D G S.t267 S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2314 S.t266 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2315 S.t265 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2316 S.t264 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2317 D G S.t263 S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2318 D G S.t262 S.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2319 S.t260 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2320 S.t259 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2321 S.t258 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2322 D G S.t257 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2323 D G S.t256 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2324 D G S.t255 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2325 S.t254 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2326 S.t253 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2327 D G S.t252 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2328 D G S.t251 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2329 S.t250 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2330 D G S.t249 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2331 D G S.t248 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2332 S.t247 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2333 S.t246 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2334 S.t245 G D S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2335 S.t244 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2336 S.t243 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2337 D G S.t242 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2338 S.t241 G D S.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2339 S.t239 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2340 S.t238 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2341 D G S.t237 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2342 S.t236 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2343 D G S.t235 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2344 S.t234 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2345 D G S.t233 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2346 S.t232 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2347 D G S.t231 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2348 S.t230 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2349 S.t229 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2350 S.t228 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2351 S.t227 G D S.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2352 S.t225 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2353 S.t224 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2354 S.t223 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2355 D G S.t222 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2356 S.t221 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2357 S.t220 G D S.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2358 S.t218 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2359 D G S.t217 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2360 S.t216 G D S.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2361 D G S.t214 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2362 S.t213 G D S.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2363 D G S.t211 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2364 S.t210 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2365 S.t209 G D S.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2366 D G S.t207 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2367 D G S.t206 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2368 D G S.t205 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2369 D G S.t204 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2370 S.t203 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2371 D G S.t202 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2372 S.t201 G D S.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2373 S.t199 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2374 D G S.t198 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2375 D G S.t197 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2376 S.t196 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2377 D G S.t195 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2378 D G S.t194 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2379 S.t193 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2380 S.t192 G D S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2381 S.t191 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2382 D G S.t190 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2383 S.t189 G D S.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2384 S.t187 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2385 S.t186 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2386 S.t185 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2387 S.t184 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2388 S.t183 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2389 S.t182 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2390 D G S.t181 S.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2391 S.t179 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2392 D G S.t178 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2393 D G S.t177 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2394 S.t176 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2395 S.t175 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2396 S.t174 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2397 D G S.t173 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2398 S.t172 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2399 D G S.t171 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2400 S.t170 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2401 S.t169 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2402 S.t168 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2403 S.t167 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2404 D G S.t166 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2405 S.t165 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2406 S.t164 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2407 S.t163 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2408 S.t162 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2409 D G S.t161 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2410 D G S.t160 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2411 S.t159 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2412 S.t158 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2413 S.t157 G D S.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2414 S.t155 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2415 S.t154 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2416 D G S.t153 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2417 S.t152 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2418 S.t151 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2419 D G S.t150 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2420 S.t149 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2421 D G S.t148 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2422 S.t147 G D S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2423 S.t146 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2424 S.t145 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2425 D G S.t144 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2426 D G S.t143 S.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2427 S.t141 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2428 D G S.t140 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2429 S.t139 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2430 S.t138 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2431 S.t137 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2432 S.t136 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2433 S.t135 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2434 S.t134 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2435 S.t133 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2436 D G S.t132 S.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2437 S.t130 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2438 S.t129 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2439 S.t127 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2440 D G S.t126 S.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2441 D G S.t124 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2442 S.t123 G D S.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2443 S.t121 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2444 S.t120 G D S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2445 D G S.t118 S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2446 D G S.t117 S.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2447 D G S.t115 S.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2448 S.t113 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2449 D G S.t112 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2450 D G S.t111 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2451 S.t110 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2452 S.t108 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2453 S.t107 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2454 S.t106 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2455 D G S.t105 S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2456 D G S.t104 S.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2457 D G S.t102 S.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2458 D G S.t100 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2459 S.t99 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2460 D G S.t98 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2461 D G S.t97 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2462 S.t96 G D S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2463 D G S.t95 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2464 D G S.t94 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2465 D G S.t93 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2466 S.t92 G D S.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2467 D G S.t90 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2468 D G S.t89 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2469 S.t88 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2470 D G S.t87 S.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2471 D G S.t85 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2472 S.t83 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2473 S.t82 G D S.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2474 D G S.t80 S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2475 S.t79 G D S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2476 D G S.t77 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2477 D G S.t76 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2478 S.t75 G D S.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2479 S.t73 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2480 S.t71 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2481 S.t70 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2482 S.t68 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2483 S.t66 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2484 D G S.t65 S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2485 S.t64 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2486 S.t62 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2487 S.t60 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2488 S.t58 G D S.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2489 S.t56 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2490 S.t54 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2491 D G S.t52 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2492 D G S.t50 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2493 D G S.t49 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2494 D G S.t48 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2495 S.t47 G D S.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2496 D G S.t45 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2497 S.t43 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2498 S.t41 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2499 D G S.t39 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2500 D G S.t38 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2501 S.t36 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2502 S.t34 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2503 S.t32 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2504 S.t31 G D S.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2505 S.t29 G D S.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2506 S.t27 G D S.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2507 D G S.t25 S.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2508 D G S.t23 S.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2509 S.t21 G D S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2510 S.t19 G D S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2511 D G S.t17 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2512 D G S.t15 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2513 S.t13 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2514 S.t11 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2515 D G S.t9 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2516 D G S.t7 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2517 S.t5 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2518 D G S.t3 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2519 D G S.t1 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 S.n867 S.n865 169.353
R1 S.n990 S.n989 169.353
R2 S.n1834 S.n1833 169.353
R3 S.n2717 S.n2716 169.353
R4 S.n3558 S.n3557 169.353
R5 S.n4390 S.n4389 169.353
R6 S.n5196 S.n5195 169.353
R7 S.n5993 S.n5992 169.353
R8 S.n6764 S.n6763 169.353
R9 S.n7526 S.n7525 169.353
R10 S.n8262 S.n8261 169.353
R11 S.n8989 S.n8988 169.353
R12 S.n9690 S.n9689 169.353
R13 S.n10382 S.n10381 169.353
R14 S.n11041 S.n11040 169.353
R15 S.n12284 S.n12283 169.353
R16 S.n13154 S.n13153 169.353
R17 S.n867 S.n866 169.353
R18 S.n13152 S.n13151 137.98
R19 S.n12282 S.n12281 137.98
R20 S.n11039 S.n11038 137.98
R21 S.n10380 S.n10379 137.98
R22 S.n9688 S.n9687 137.98
R23 S.n8987 S.n8986 137.98
R24 S.n8260 S.n8259 137.98
R25 S.n7524 S.n7523 137.98
R26 S.n6762 S.n6761 137.98
R27 S.n5991 S.n5990 137.98
R28 S.n5194 S.n5193 137.98
R29 S.n4388 S.n4387 137.98
R30 S.n3556 S.n3555 137.98
R31 S.n2715 S.n2714 137.98
R32 S.n1832 S.n1831 137.98
R33 S.n988 S.n987 137.98
R34 S.n864 S.n863 137.98
R35 S.n465 S.n464 135.611
R36 S.n1035 S.n1034 135.611
R37 S.n2326 S.n2325 135.611
R38 S.n3200 S.n3199 135.611
R39 S.n4065 S.n4064 135.611
R40 S.n4873 S.n4872 135.611
R41 S.n5672 S.n5671 135.611
R42 S.n6445 S.n6444 135.611
R43 S.n7209 S.n7208 135.611
R44 S.n7780 S.n7779 135.611
R45 S.n8494 S.n8493 135.611
R46 S.n9379 S.n9378 135.611
R47 S.n10073 S.n10072 135.611
R48 S.n10744 S.n10743 135.611
R49 S.n11387 S.n11386 135.611
R50 S.n11958 S.n11957 135.611
R51 S.n12610 S.n12609 135.611
R52 S.n476 S.n475 91.65
R53 S.n12621 S.n12620 91.65
R54 S.n9391 S.n9390 91.65
R55 S.n10084 S.n10083 91.65
R56 S.n10756 S.n10755 91.65
R57 S.n11398 S.n11397 91.65
R58 S.n11970 S.n11969 91.65
R59 S.n7792 S.n7791 91.65
R60 S.n8505 S.n8504 91.65
R61 S.n6457 S.n6456 91.65
R62 S.n7220 S.n7219 91.65
R63 S.n4885 S.n4884 91.65
R64 S.n5683 S.n5682 91.65
R65 S.n3212 S.n3211 91.65
R66 S.n4076 S.n4075 91.65
R67 S.n1047 S.n1046 91.65
R68 S.n2337 S.n2336 91.65
R69 S.n12273 S.n12272 91.389
R70 S.n882 S.n881 91.389
R71 S.n1798 S.n1797 91.389
R72 S.n2686 S.n2685 91.389
R73 S.n3527 S.n3526 91.389
R74 S.n4359 S.n4358 91.389
R75 S.n5165 S.n5164 91.389
R76 S.n5962 S.n5961 91.389
R77 S.n6733 S.n6732 91.389
R78 S.n7495 S.n7494 91.389
R79 S.n8231 S.n8230 91.389
R80 S.n8958 S.n8957 91.389
R81 S.n9659 S.n9658 91.389
R82 S.n10351 S.n10350 91.389
R83 S.n11020 S.n11019 91.389
R84 S.n11660 S.n11659 91.389
R85 S.n13143 S.n13142 91.389
R86 S.n951 S.n950 87.222
R87 S.n948 S.n947 87.222
R88 S.n201 S.n200 87.222
R89 S.n975 S.n974 87.222
R90 S.n216 S.n215 87.222
R91 S.n922 S.n921 87.222
R92 S.n939 S.n938 87.222
R93 S.n189 S.n188 87.222
R94 S.n971 S.n970 87.222
R95 S.n177 S.n176 87.222
R96 S.n967 S.n966 87.222
R97 S.n164 S.n163 87.222
R98 S.n963 S.n962 87.222
R99 S.n151 S.n150 87.222
R100 S.n959 S.n958 87.222
R101 S.n138 S.n137 87.222
R102 S.n955 S.n954 87.222
R103 S.n12542 S.n12541 86.961
R104 S.n12482 S.n12481 86.961
R105 S.n12486 S.n12485 86.961
R106 S.n12490 S.n12489 86.961
R107 S.n12494 S.n12493 86.961
R108 S.n12498 S.n12497 86.961
R109 S.n12502 S.n12501 86.961
R110 S.n12506 S.n12505 86.961
R111 S.n12510 S.n12509 86.961
R112 S.n12514 S.n12513 86.961
R113 S.n12518 S.n12517 86.961
R114 S.n12522 S.n12521 86.961
R115 S.n12526 S.n12525 86.961
R116 S.n12530 S.n12529 86.961
R117 S.n12534 S.n12533 86.961
R118 S.n12538 S.n12537 86.961
R119 S.n12478 S.n12477 86.961
R120 S.t28 S.t278 57.619
R121 S.n869 S.t61 50.285
R122 S.n467 S.t20 50.285
R123 S.n992 S.t33 50.285
R124 S.n1037 S.t509 50.285
R125 S.n1836 S.t63 50.285
R126 S.n2328 S.t215 50.285
R127 S.n2719 S.t10 50.285
R128 S.n3202 S.t46 50.285
R129 S.n3560 S.t78 50.285
R130 S.n4067 S.t522 50.285
R131 S.n4392 S.t53 50.285
R132 S.n4875 S.t226 50.285
R133 S.n5198 S.t4 50.285
R134 S.n5674 S.t74 50.285
R135 S.n5995 S.t69 50.285
R136 S.n6447 S.t125 50.285
R137 S.n6766 S.t42 50.285
R138 S.n7211 S.t219 50.285
R139 S.n7528 S.t299 50.285
R140 S.n7782 S.t156 50.285
R141 S.n8264 S.t84 50.285
R142 S.n8496 S.t188 50.285
R143 S.n8991 S.t67 50.285
R144 S.n9381 S.t212 50.285
R145 S.n9692 S.t101 50.285
R146 S.n10075 S.t30 50.285
R147 S.n10384 S.t91 50.285
R148 S.n10746 S.t6 50.285
R149 S.n11043 S.t261 50.285
R150 S.n11389 S.t208 50.285
R151 S.n12286 S.t114 50.285
R152 S.n11960 S.t57 50.285
R153 S.n13156 S.t180 50.285
R154 S.n12612 S.t128 50.285
R155 S.t116 S.n830 48.609
R156 S.t430 S.n736 48.609
R157 S.t320 S.n1792 48.609
R158 S.t142 S.n1317 48.609
R159 S.t200 S.n2282 48.609
R160 S.t55 S.n2599 48.609
R161 S.t240 S.n3117 48.609
R162 S.t444 S.n3455 48.609
R163 S.t109 S.n3929 48.609
R164 S.t51 S.n4302 48.609
R165 S.t360 S.n4729 48.609
R166 S.t81 S.n5092 48.609
R167 S.t390 S.n5506 48.609
R168 S.t460 S.n5873 48.609
R169 S.t119 S.n6271 48.609
R170 S.t8 S.n6628 48.609
R171 S.t37 S.n7013 48.609
R172 S.t40 S.n7374 48.609
R173 S.t59 S.n7743 48.609
R174 S.t22 S.n7927 48.609
R175 S.t131 S.n8450 48.609
R176 S.t0 S.n8623 48.609
R177 S.t24 S.n9145 48.609
R178 S.t26 S.n9490 48.609
R179 S.t86 S.n9817 48.609
R180 S.t16 S.n10166 48.609
R181 S.t103 S.n10477 48.609
R182 S.t122 S.n10819 48.609
R183 S.t12 S.n11102 48.609
R184 S.t18 S.n11440 48.609
R185 S.t44 S.n11699 48.609
R186 S.t2 S.n12016 48.609
R187 S.t72 S.n12571 48.609
R188 S.t14 S.n12670 48.609
R189 S.t35 S.n12479 48.609
R190 S.n1794 S.t2223 3.904
R191 S.n1796 S.n1795 3.904
R192 S.n12542 S.t1057 3.904
R193 S.n12540 S.t642 3.904
R194 S.n12634 S.n12633 3.904
R195 S.n12645 S.t747 3.904
R196 S.n12642 S.t181 3.904
R197 S.n12637 S.n12636 3.904
R198 S.n12558 S.n12557 3.904
R199 S.n12569 S.t1532 3.904
R200 S.n12566 S.t80 3.904
R201 S.n12561 S.n12560 3.904
R202 S.n11996 S.n11995 3.904
R203 S.n12014 S.t1991 3.904
R204 S.n12011 S.t887 3.904
R205 S.n11999 S.n11998 3.904
R206 S.n12273 S.t2543 3.904
R207 S.n12275 S.t1248 3.904
R208 S.n12544 S.t1645 3.904
R209 S.n12545 S.t1110 3.904
R210 S.n477 S.t1276 3.904
R211 S.n840 S.n839 3.904
R212 S.n853 S.t117 3.904
R213 S.n856 S.t1313 3.904
R214 S.n843 S.n842 3.904
R215 S.n949 S.t1595 3.904
R216 S.n945 S.t1901 3.904
R217 S.n817 S.n816 3.904
R218 S.n828 S.t2105 3.904
R219 S.n825 S.t2483 3.904
R220 S.n820 S.n819 3.904
R221 S.n1776 S.n1775 3.904
R222 S.n1790 S.t2135 3.904
R223 S.n1787 S.t2487 3.904
R224 S.n1773 S.n1772 3.904
R225 S.n12622 S.t1472 3.904
R226 S.n12578 S.n12577 3.904
R227 S.n12593 S.t316 3.904
R228 S.n12596 S.t1978 3.904
R229 S.n12575 S.n12574 3.904
R230 S.n11979 S.n11978 3.904
R231 S.n11990 S.t2302 3.904
R232 S.n11987 S.t1092 3.904
R233 S.n11976 S.n11975 3.904
R234 S.n11682 S.n11681 3.904
R235 S.n11697 S.t2434 3.904
R236 S.n11694 S.t1419 3.904
R237 S.n11679 S.n11678 3.904
R238 S.n11427 S.n11426 3.904
R239 S.n11438 S.t1712 3.904
R240 S.n11435 S.t512 3.904
R241 S.n11424 S.n11423 3.904
R242 S.n11085 S.n11084 3.904
R243 S.n11100 S.t1897 3.904
R244 S.n11097 S.t956 3.904
R245 S.n11082 S.n11081 3.904
R246 S.n10806 S.n10805 3.904
R247 S.n10817 S.t1270 3.904
R248 S.n10814 S.t2409 3.904
R249 S.n10803 S.n10802 3.904
R250 S.n10460 S.n10459 3.904
R251 S.n10475 S.t1310 3.904
R252 S.n10472 S.t343 3.904
R253 S.n10457 S.n10456 3.904
R254 S.n10153 S.n10152 3.904
R255 S.n10164 S.t673 3.904
R256 S.n10161 S.t1872 3.904
R257 S.n10150 S.n10149 3.904
R258 S.n9800 S.n9799 3.904
R259 S.n9815 S.t1024 3.904
R260 S.n9812 S.t2301 3.904
R261 S.n9797 S.n9796 3.904
R262 S.n9477 S.n9476 3.904
R263 S.n9488 S.t77 3.904
R264 S.n9485 S.t1538 3.904
R265 S.n9474 S.n9473 3.904
R266 S.n9128 S.n9127 3.904
R267 S.n9143 S.t415 3.904
R268 S.n9140 S.t1705 3.904
R269 S.n9125 S.n9124 3.904
R270 S.n8610 S.n8609 3.904
R271 S.n8621 S.t2028 3.904
R272 S.n8618 S.t994 3.904
R273 S.n8607 S.n8606 3.904
R274 S.n8433 S.n8432 3.904
R275 S.n8448 S.t2347 3.904
R276 S.n8445 S.t1143 3.904
R277 S.n8430 S.n8429 3.904
R278 S.n7914 S.n7913 3.904
R279 S.n7925 S.t1462 3.904
R280 S.n7922 S.t384 3.904
R281 S.n7911 S.n7910 3.904
R282 S.n7726 S.n7725 3.904
R283 S.n7741 S.t1918 3.904
R284 S.n7738 S.t573 3.904
R285 S.n7723 S.n7722 3.904
R286 S.n7361 S.n7360 3.904
R287 S.n7372 S.t865 3.904
R288 S.n7369 S.t1331 3.904
R289 S.n7358 S.n7357 3.904
R290 S.n6996 S.n6995 3.904
R291 S.n7011 S.t173 3.904
R292 S.n7008 S.t413 3.904
R293 S.n6993 S.n6992 3.904
R294 S.n6615 S.n6614 3.904
R295 S.n6626 S.t1769 3.904
R296 S.n6623 S.t1770 3.904
R297 S.n6612 S.n6611 3.904
R298 S.n6254 S.n6253 3.904
R299 S.n6269 S.t623 3.904
R300 S.n6266 S.t2520 3.904
R301 S.n6251 S.n6250 3.904
R302 S.n5860 S.n5859 3.904
R303 S.n5871 S.t1383 3.904
R304 S.n5868 S.t1734 3.904
R305 S.n5857 S.n5856 3.904
R306 S.n5489 S.n5488 3.904
R307 S.n5504 S.t605 3.904
R308 S.n5501 S.t2489 3.904
R309 S.n5486 S.n5485 3.904
R310 S.n5079 S.n5078 3.904
R311 S.n5090 S.t1355 3.904
R312 S.n5087 S.t1703 3.904
R313 S.n5076 S.n5075 3.904
R314 S.n4712 S.n4711 3.904
R315 S.n4727 S.t585 3.904
R316 S.n4724 S.t2459 3.904
R317 S.n4709 S.n4708 3.904
R318 S.n4289 S.n4288 3.904
R319 S.n4300 S.t1327 3.904
R320 S.n4297 S.t1674 3.904
R321 S.n4286 S.n4285 3.904
R322 S.n3912 S.n3911 3.904
R323 S.n3927 S.t564 3.904
R324 S.n3924 S.t2584 3.904
R325 S.n3909 S.n3908 3.904
R326 S.n3442 S.n3441 3.904
R327 S.n3453 S.t1431 3.904
R328 S.n3450 S.t1637 3.904
R329 S.n3439 S.n3438 3.904
R330 S.n3100 S.n3099 3.904
R331 S.n3115 S.t534 3.904
R332 S.n3112 S.t2550 3.904
R333 S.n3097 S.n3096 3.904
R334 S.n2586 S.n2585 3.904
R335 S.n2597 S.t1405 3.904
R336 S.n2594 S.t1609 3.904
R337 S.n2583 S.n2582 3.904
R338 S.n2263 S.n2262 3.904
R339 S.n2280 S.t2164 3.904
R340 S.n2277 S.t2517 3.904
R341 S.n2260 S.n2259 3.904
R342 S.n1306 S.n1305 3.904
R343 S.n1315 S.t1381 3.904
R344 S.n1312 S.t734 3.904
R345 S.n1303 S.n1302 3.904
R346 S.n723 S.n722 3.904
R347 S.n734 S.t1353 3.904
R348 S.n731 S.t706 3.904
R349 S.n726 S.n725 3.904
R350 S.n195 S.t491 3.904
R351 S.n420 S.n419 3.904
R352 S.n431 S.t1424 3.904
R353 S.n428 S.t1624 3.904
R354 S.n423 S.n422 3.904
R355 S.n1665 S.n1664 3.904
R356 S.n1678 S.t1442 3.904
R357 S.n1675 S.t1657 3.904
R358 S.n1662 S.n1661 3.904
R359 S.n9392 S.t841 3.904
R360 S.n9152 S.n9151 3.904
R361 S.n9166 S.t2248 3.904
R362 S.n9169 S.t880 3.904
R363 S.n9149 S.n9148 3.904
R364 S.n8514 S.n8513 3.904
R365 S.n8525 S.t1208 3.904
R366 S.n8522 S.t269 3.904
R367 S.n8511 S.n8510 3.904
R368 S.n8286 S.n8285 3.904
R369 S.n8301 S.t1628 3.904
R370 S.n8298 S.t297 3.904
R371 S.n8283 S.n8282 3.904
R372 S.n7818 S.n7817 3.904
R373 S.n7829 S.t629 3.904
R374 S.n7826 S.t2221 3.904
R375 S.n7815 S.n7814 3.904
R376 S.n7579 S.n7578 3.904
R377 S.n7594 S.t1090 3.904
R378 S.n7591 S.t2355 3.904
R379 S.n7576 S.n7575 3.904
R380 S.n7265 S.n7264 3.904
R381 S.n7276 S.t178 3.904
R382 S.n7273 S.t1600 3.904
R383 S.n7262 S.n7261 3.904
R384 S.n6849 S.n6848 3.904
R385 S.n6864 S.t505 3.904
R386 S.n6861 S.t1796 3.904
R387 S.n6846 S.n6845 3.904
R388 S.n6519 S.n6518 3.904
R389 S.n6530 S.t2117 3.904
R390 S.n6527 S.t572 3.904
R391 S.n6516 S.n6515 3.904
R392 S.n6107 S.n6106 3.904
R393 S.n6122 S.t1939 3.904
R394 S.n6119 S.t1021 3.904
R395 S.n6104 S.n6103 3.904
R396 S.n5764 S.n5763 3.904
R397 S.n5775 S.t1340 3.904
R398 S.n5772 S.t2466 3.904
R399 S.n5761 S.n5760 3.904
R400 S.n5342 S.n5341 3.904
R401 S.n5357 S.t1373 3.904
R402 S.n5354 S.t410 3.904
R403 S.n5339 S.n5338 3.904
R404 S.n4983 S.n4982 3.904
R405 S.n4994 S.t715 3.904
R406 S.n4991 S.t1923 3.904
R407 S.n4980 S.n4979 3.904
R408 S.n4565 S.n4564 3.904
R409 S.n4580 S.t748 3.904
R410 S.n4577 S.t2343 3.904
R411 S.n4562 S.n4561 3.904
R412 S.n4193 S.n4192 3.904
R413 S.n4204 S.t160 3.904
R414 S.n4201 S.t1347 3.904
R415 S.n4190 S.n4189 3.904
R416 S.n3765 S.n3764 3.904
R417 S.n3780 S.t308 3.904
R418 S.n3777 S.t1778 3.904
R419 S.n3762 S.n3761 3.904
R420 S.n3346 S.n3345 3.904
R421 S.n3357 S.t2088 3.904
R422 S.n3354 S.t979 3.904
R423 S.n3343 S.n3342 3.904
R424 S.n2953 S.n2952 3.904
R425 S.n2968 S.t2327 3.904
R426 S.n2965 S.t1722 3.904
R427 S.n2950 S.n2949 3.904
R428 S.n2490 S.n2489 3.904
R429 S.n2501 S.t574 3.904
R430 S.n2498 S.t947 3.904
R431 S.n2487 S.n2486 3.904
R432 S.n2110 S.n2109 3.904
R433 S.n2127 S.t1456 3.904
R434 S.n2124 S.t1689 3.904
R435 S.n2107 S.n2106 3.904
R436 S.n1209 S.n1208 3.904
R437 S.n1218 S.t554 3.904
R438 S.n1215 S.t2565 3.904
R439 S.n1206 S.n1205 3.904
R440 S.n973 S.t2268 3.904
R441 S.n440 S.n439 3.904
R442 S.n451 S.t557 3.904
R443 S.n448 S.t915 3.904
R444 S.n443 S.n442 3.904
R445 S.n10085 S.t281 3.904
R446 S.n9828 S.n9827 3.904
R447 S.n9843 S.t1957 3.904
R448 S.n9846 S.t611 3.904
R449 S.n9831 S.n9830 3.904
R450 S.n9398 S.n9397 3.904
R451 S.n9409 S.t936 3.904
R452 S.n9406 S.t2484 3.904
R453 S.n9401 S.n9400 3.904
R454 S.n9005 S.n9004 3.904
R455 S.n9025 S.t1390 3.904
R456 S.n9022 S.t2525 3.904
R457 S.n9008 S.n9007 3.904
R458 S.n8531 S.n8530 3.904
R459 S.n8542 S.t330 3.904
R460 S.n8539 S.t1932 3.904
R461 S.n8534 S.n8533 3.904
R462 S.n8310 S.n8309 3.904
R463 S.n8330 S.t761 3.904
R464 S.n8327 S.t2078 3.904
R465 S.n8313 S.n8312 3.904
R466 S.n7835 S.n7834 3.904
R467 S.n7846 S.t2381 3.904
R468 S.n7843 S.t1360 3.904
R469 S.n7838 S.n7837 3.904
R470 S.n7603 S.n7602 3.904
R471 S.n7623 S.t211 3.904
R472 S.n7620 S.t1497 3.904
R473 S.n7606 S.n7605 3.904
R474 S.n7282 S.n7281 3.904
R475 S.n7293 S.t1843 3.904
R476 S.n7290 S.t736 3.904
R477 S.n7285 S.n7284 3.904
R478 S.n6873 S.n6872 3.904
R479 S.n6893 S.t2148 3.904
R480 S.n6890 S.t930 3.904
R481 S.n6876 S.n6875 3.904
R482 S.n6536 S.n6535 3.904
R483 S.n6547 S.t1246 3.904
R484 S.n6544 S.t2217 3.904
R485 S.n6539 S.n6538 3.904
R486 S.n6131 S.n6130 3.904
R487 S.n6151 S.t1082 3.904
R488 S.n6148 S.t118 3.904
R489 S.n6134 S.n6133 3.904
R490 S.n5781 S.n5780 3.904
R491 S.n5792 S.t461 3.904
R492 S.n5789 S.t1597 3.904
R493 S.n5784 S.n5783 3.904
R494 S.n5366 S.n5365 3.904
R495 S.n5386 S.t500 3.904
R496 S.n5383 S.t2058 3.904
R497 S.n5369 S.n5368 3.904
R498 S.n5000 S.n4999 3.904
R499 S.n5011 S.t2370 3.904
R500 S.n5008 S.t1061 3.904
R501 S.n5003 S.n5002 3.904
R502 S.n4589 S.n4588 3.904
R503 S.n4609 S.t2540 3.904
R504 S.n4606 S.t1487 3.904
R505 S.n4592 S.n4591 3.904
R506 S.n4210 S.n4209 3.904
R507 S.n4221 S.t1821 3.904
R508 S.n4218 S.t98 3.904
R509 S.n4213 S.n4212 3.904
R510 S.n3789 S.n3788 3.904
R511 S.n3809 S.t1489 3.904
R512 S.n3806 S.t881 3.904
R513 S.n3792 S.n3791 3.904
R514 S.n3363 S.n3362 3.904
R515 S.n3374 S.t2245 3.904
R516 S.n3371 S.t49 3.904
R517 S.n3366 S.n3365 3.904
R518 S.n2977 S.n2976 3.904
R519 S.n2997 S.t1468 3.904
R520 S.n2994 S.t850 3.904
R521 S.n2980 S.n2979 3.904
R522 S.n2507 S.n2506 3.904
R523 S.n2518 S.t2219 3.904
R524 S.n2515 S.t2586 3.904
R525 S.n2510 S.n2509 3.904
R526 S.n2136 S.n2135 3.904
R527 S.n2156 S.t598 3.904
R528 S.n2153 S.t815 3.904
R529 S.n2139 S.n2138 3.904
R530 S.n1224 S.n1223 3.904
R531 S.n1237 S.t2192 3.904
R532 S.n1234 S.t1692 3.904
R533 S.n1227 S.n1226 3.904
R534 S.n1243 S.n1242 3.904
R535 S.n1257 S.t1332 3.904
R536 S.n1254 S.t820 3.904
R537 S.n1246 S.n1245 3.904
R538 S.n455 S.n454 3.904
R539 S.n756 S.t1434 3.904
R540 S.n759 S.t791 3.904
R541 S.n762 S.n761 3.904
R542 S.n770 S.n769 3.904
R543 S.n785 S.t2194 3.904
R544 S.n782 S.t2555 3.904
R545 S.n773 S.n772 3.904
R546 S.n209 S.t1409 3.904
R547 S.n2174 S.n2173 3.904
R548 S.n2191 S.t2249 3.904
R549 S.n2188 S.t2463 3.904
R550 S.n2171 S.n2170 3.904
R551 S.n3014 S.n3013 3.904
R552 S.n3029 S.t608 3.904
R553 S.n3026 S.t2494 3.904
R554 S.n3011 S.n3010 3.904
R555 S.n3826 S.n3825 3.904
R556 S.n3841 S.t624 3.904
R557 S.n3838 S.t2526 3.904
R558 S.n3823 S.n3822 3.904
R559 S.n4626 S.n4625 3.904
R560 S.n4641 S.t646 3.904
R561 S.n4638 S.t2558 3.904
R562 S.n4623 S.n4622 3.904
R563 S.n5403 S.n5402 3.904
R564 S.n5418 S.t2276 3.904
R565 S.n5415 S.t1197 3.904
R566 S.n5400 S.n5399 3.904
R567 S.n6168 S.n6167 3.904
R568 S.n6183 S.t205 3.904
R569 S.n6180 S.t1790 3.904
R570 S.n6165 S.n6164 3.904
R571 S.n6910 S.n6909 3.904
R572 S.n6925 S.t1288 3.904
R573 S.n6922 S.t2570 3.904
R574 S.n6907 S.n6906 3.904
R575 S.n7640 S.n7639 3.904
R576 S.n7655 S.t1879 3.904
R577 S.n7652 S.t634 3.904
R578 S.n7637 S.n7636 3.904
R579 S.n8347 S.n8346 3.904
R580 S.n8362 S.t2414 3.904
R581 S.n8359 S.t1216 3.904
R582 S.n8344 S.n8343 3.904
R583 S.n9042 S.n9041 3.904
R584 S.n9057 S.t517 3.904
R585 S.n9054 S.t1813 3.904
R586 S.n9039 S.n9038 3.904
R587 S.n9714 S.n9713 3.904
R588 S.n9729 S.t1097 3.904
R589 S.n9726 S.t2265 3.904
R590 S.n9711 S.n9710 3.904
R591 S.n10487 S.n10486 3.904
R592 S.n10501 S.t1402 3.904
R593 S.n10504 S.t305 3.904
R594 S.n10484 S.n10483 3.904
R595 S.n10757 S.t2498 3.904
R596 S.n10093 S.n10092 3.904
R597 S.n10104 S.t638 3.904
R598 S.n10101 S.t1940 3.904
R599 S.n10090 S.n10089 3.904
R600 S.n9417 S.n9416 3.904
R601 S.n9428 S.t2575 3.904
R602 S.n9425 S.t1610 3.904
R603 S.n9414 S.n9413 3.904
R604 S.n8550 S.n8549 3.904
R605 S.n8561 S.t2126 3.904
R606 S.n8558 S.t1072 3.904
R607 S.n8547 S.n8546 3.904
R608 S.n7854 S.n7853 3.904
R609 S.n7865 S.t1527 3.904
R610 S.n7862 S.t487 3.904
R611 S.n7851 S.n7850 3.904
R612 S.n7301 S.n7300 3.904
R613 S.n7312 S.t981 3.904
R614 S.n7309 S.t2386 3.904
R615 S.n7298 S.n7297 3.904
R616 S.n6555 S.n6554 3.904
R617 S.n6566 S.t364 3.904
R618 S.n6563 S.t1357 3.904
R619 S.n6552 S.n6551 3.904
R620 S.n5800 S.n5799 3.904
R621 S.n5811 S.t2106 3.904
R622 S.n5808 S.t733 3.904
R623 S.n5797 S.n5796 3.904
R624 S.n5019 S.n5018 3.904
R625 S.n5030 S.t1513 3.904
R626 S.n5027 S.t1805 3.904
R627 S.n5016 S.n5015 3.904
R628 S.n4229 S.n4228 3.904
R629 S.n4240 S.t1412 3.904
R630 S.n4237 S.t1774 3.904
R631 S.n4226 S.n4225 3.904
R632 S.n3382 S.n3381 3.904
R633 S.n3393 S.t1386 3.904
R634 S.n3390 S.t1743 3.904
R635 S.n3379 S.n3378 3.904
R636 S.n2526 S.n2525 3.904
R637 S.n2537 S.t1359 3.904
R638 S.n2534 S.t1709 3.904
R639 S.n2523 S.n2522 3.904
R640 S.n1721 S.n1720 3.904
R641 S.n1740 S.t1361 3.904
R642 S.n1737 S.t1714 3.904
R643 S.n1724 S.n1723 3.904
R644 S.n680 S.n679 3.904
R645 S.n695 S.t570 3.904
R646 S.n692 S.t2440 3.904
R647 S.n683 S.n682 3.904
R648 S.n225 S.n224 3.904
R649 S.n887 S.t1338 3.904
R650 S.n890 S.t1683 3.904
R651 S.n893 S.n892 3.904
R652 S.n220 S.t543 3.904
R653 S.n11399 S.t2243 3.904
R654 S.n11116 S.n11115 3.904
R655 S.n11124 S.t1107 3.904
R656 S.n11127 S.t2537 3.904
R657 S.n11113 S.n11112 3.904
R658 S.n10770 S.n10769 3.904
R659 S.n10778 S.t339 3.904
R660 S.n10775 S.t1621 3.904
R661 S.n10767 S.n10766 3.904
R662 S.n10405 S.n10404 3.904
R663 S.n10423 S.t530 3.904
R664 S.n10420 S.t1970 3.904
R665 S.n10402 S.n10401 3.904
R666 S.n10117 S.n10116 3.904
R667 S.n10125 S.t2295 3.904
R668 S.n10122 S.t1080 3.904
R669 S.n10114 S.n10113 3.904
R670 S.n9745 S.n9744 3.904
R671 S.n9763 S.t222 3.904
R672 S.n9760 S.t1506 3.904
R673 S.n9742 S.n9741 3.904
R674 S.n9441 S.n9440 3.904
R675 S.n9449 S.t1857 3.904
R676 S.n9446 S.t746 3.904
R677 S.n9438 S.n9437 3.904
R678 S.n9073 S.n9072 3.904
R679 S.n9091 S.t2162 3.904
R680 S.n9088 S.t946 3.904
R681 S.n9070 S.n9069 3.904
R682 S.n8574 S.n8573 3.904
R683 S.n8582 S.t1260 3.904
R684 S.n8579 S.t195 3.904
R685 S.n8571 S.n8570 3.904
R686 S.n8378 S.n8377 3.904
R687 S.n8396 S.t1550 3.904
R688 S.n8393 S.t335 3.904
R689 S.n8375 S.n8374 3.904
R690 S.n7878 S.n7877 3.904
R691 S.n7886 S.t666 3.904
R692 S.n7883 S.t2132 3.904
R693 S.n7875 S.n7874 3.904
R694 S.n7671 S.n7670 3.904
R695 S.n7689 S.t1015 3.904
R696 S.n7686 S.t2290 3.904
R697 S.n7668 S.n7667 3.904
R698 S.n7325 S.n7324 3.904
R699 S.n7333 S.t48 3.904
R700 S.n7330 S.t1530 3.904
R701 S.n7322 S.n7321 3.904
R702 S.n6941 S.n6940 3.904
R703 S.n6959 S.t405 3.904
R704 S.n6956 S.t1694 3.904
R705 S.n6938 S.n6937 3.904
R706 S.n6579 S.n6578 3.904
R707 S.n6587 S.t2016 3.904
R708 S.n6584 S.t479 3.904
R709 S.n6576 S.n6575 3.904
R710 S.n6199 S.n6198 3.904
R711 S.n6217 S.t1979 3.904
R712 S.n6214 S.t921 3.904
R713 S.n6196 S.n6195 3.904
R714 S.n5824 S.n5823 3.904
R715 S.n5832 S.t1239 3.904
R716 S.n5829 S.t973 3.904
R717 S.n5821 S.n5820 3.904
R718 S.n5434 S.n5433 3.904
R719 S.n5452 S.t2324 3.904
R720 S.n5449 S.t1717 3.904
R721 S.n5431 S.n5430 3.904
R722 S.n5043 S.n5042 3.904
R723 S.n5051 S.t571 3.904
R724 S.n5048 S.t940 3.904
R725 S.n5040 S.n5039 3.904
R726 S.n4657 S.n4656 3.904
R727 S.n4675 S.t2303 3.904
R728 S.n4672 S.t1685 3.904
R729 S.n4654 S.n4653 3.904
R730 S.n4253 S.n4252 3.904
R731 S.n4261 S.t547 3.904
R732 S.n4258 S.t904 3.904
R733 S.n4250 S.n4249 3.904
R734 S.n3857 S.n3856 3.904
R735 S.n3875 S.t2283 3.904
R736 S.n3872 S.t1650 3.904
R737 S.n3854 S.n3853 3.904
R738 S.n3406 S.n3405 3.904
R739 S.n3414 S.t515 3.904
R740 S.n3411 S.t867 3.904
R741 S.n3403 S.n3402 3.904
R742 S.n3045 S.n3044 3.904
R743 S.n3063 S.t2261 3.904
R744 S.n3060 S.t1618 3.904
R745 S.n3042 S.n3041 3.904
R746 S.n2550 S.n2549 3.904
R747 S.n2558 S.t482 3.904
R748 S.n2555 S.t839 3.904
R749 S.n2547 S.n2546 3.904
R750 S.n2207 S.n2206 3.904
R751 S.n2225 S.t1391 3.904
R752 S.n2222 S.t1750 3.904
R753 S.n2204 S.n2203 3.904
R754 S.n1270 S.n1269 3.904
R755 S.n1278 S.t592 3.904
R756 S.n1275 S.t2465 3.904
R757 S.n1267 S.n1266 3.904
R758 S.n1749 S.n1748 3.904
R759 S.n1768 S.t488 3.904
R760 S.n1765 S.t843 3.904
R761 S.n1752 S.n1751 3.904
R762 S.n700 S.n699 3.904
R763 S.n714 S.t2214 3.904
R764 S.n711 S.t1575 3.904
R765 S.n703 S.n702 3.904
R766 S.n1289 S.n1288 3.904
R767 S.n1298 S.t2239 3.904
R768 S.n1295 S.t1596 3.904
R769 S.n1286 S.n1285 3.904
R770 S.n2234 S.n2233 3.904
R771 S.n2246 S.t519 3.904
R772 S.n2243 S.t871 3.904
R773 S.n2237 S.n2236 3.904
R774 S.n2564 S.n2563 3.904
R775 S.n2578 S.t2263 3.904
R776 S.n2575 S.t2482 3.904
R777 S.n2567 S.n2566 3.904
R778 S.n3072 S.n3071 3.904
R779 S.n3083 S.t1404 3.904
R780 S.n3080 S.t909 3.904
R781 S.n3075 S.n3074 3.904
R782 S.n3420 S.n3419 3.904
R783 S.n3434 S.t2160 3.904
R784 S.n3431 S.t2512 3.904
R785 S.n3423 S.n3422 3.904
R786 S.n3884 S.n3883 3.904
R787 S.n3895 S.t1429 3.904
R788 S.n3892 S.t779 3.904
R789 S.n3887 S.n3886 3.904
R790 S.n4267 S.n4266 3.904
R791 S.n4281 S.t2189 3.904
R792 S.n4278 S.t2547 3.904
R793 S.n4270 S.n4269 3.904
R794 S.n4684 S.n4683 3.904
R795 S.n4695 S.t1448 3.904
R796 S.n4692 S.t811 3.904
R797 S.n4687 S.n4686 3.904
R798 S.n5057 S.n5056 3.904
R799 S.n5071 S.t2216 3.904
R800 S.n5068 S.t2580 3.904
R801 S.n5060 S.n5059 3.904
R802 S.n5461 S.n5460 3.904
R803 S.n5472 S.t1466 3.904
R804 S.n5469 S.t846 3.904
R805 S.n5464 S.n5463 3.904
R806 S.n5838 S.n5837 3.904
R807 S.n5852 S.t2242 3.904
R808 S.n5849 S.t39 3.904
R809 S.n5841 S.n5840 3.904
R810 S.n6226 S.n6225 3.904
R811 S.n6237 S.t1485 3.904
R812 S.n6234 S.t874 3.904
R813 S.n6229 S.n6228 3.904
R814 S.n6593 S.n6592 3.904
R815 S.n6607 S.t1163 3.904
R816 S.n6604 S.t95 3.904
R817 S.n6596 S.n6595 3.904
R818 S.n6968 S.n6967 3.904
R819 S.n6979 S.t2196 3.904
R820 S.n6976 S.t819 3.904
R821 S.n6971 S.n6970 3.904
R822 S.n7339 S.n7338 3.904
R823 S.n7353 S.t1741 3.904
R824 S.n7350 S.t670 3.904
R825 S.n7342 S.n7341 3.904
R826 S.n7698 S.n7697 3.904
R827 S.n7709 S.t111 3.904
R828 S.n7706 S.t1436 3.904
R829 S.n7701 S.n7700 3.904
R830 S.n7892 S.n7891 3.904
R831 S.n7906 S.t2320 3.904
R832 S.n7903 S.t1267 3.904
R833 S.n7895 S.n7894 3.904
R834 S.n8405 S.n8404 3.904
R835 S.n8416 S.t688 3.904
R836 S.n8413 S.t1992 3.904
R837 S.n8408 S.n8407 3.904
R838 S.n8588 S.n8587 3.904
R839 S.n8602 S.t377 3.904
R840 S.n8599 S.t1863 3.904
R841 S.n8591 S.n8590 3.904
R842 S.n9100 S.n9099 3.904
R843 S.n9111 S.t1298 3.904
R844 S.n9108 S.t2583 3.904
R845 S.n9103 S.n9102 3.904
R846 S.n9455 S.n9454 3.904
R847 S.n9469 S.t990 3.904
R848 S.n9466 S.t2399 3.904
R849 S.n9458 S.n9457 3.904
R850 S.n9772 S.n9771 3.904
R851 S.n9783 S.t1887 3.904
R852 S.n9780 S.t645 3.904
R853 S.n9775 S.n9774 3.904
R854 S.n10131 S.n10130 3.904
R855 S.n10145 S.t1533 3.904
R856 S.n10142 S.t204 3.904
R857 S.n10134 S.n10133 3.904
R858 S.n10432 S.n10431 3.904
R859 S.n10443 S.t2173 3.904
R860 S.n10440 S.t1226 3.904
R861 S.n10435 S.n10434 3.904
R862 S.n10784 S.n10783 3.904
R863 S.n10798 S.t1997 3.904
R864 S.n10795 S.t754 3.904
R865 S.n10787 S.n10786 3.904
R866 S.n11057 S.n11056 3.904
R867 S.n11068 S.t231 3.904
R868 S.n11065 S.t1666 3.904
R869 S.n11060 S.n11059 3.904
R870 S.n11405 S.n11404 3.904
R871 S.n11419 S.t2588 3.904
R872 S.n11416 S.t1384 3.904
R873 S.n11408 S.n11407 3.904
R874 S.n11711 S.n11710 3.904
R875 S.n11719 S.t784 3.904
R876 S.n11722 S.t2275 3.904
R877 S.n11714 S.n11713 3.904
R878 S.n11971 S.t1952 3.904
R879 S.n927 S.t2184 3.904
R880 S.n790 S.n789 3.904
R881 S.n807 S.t459 3.904
R882 S.n804 S.t809 3.904
R883 S.n793 S.n792 3.904
R884 S.n1687 S.n1686 3.904
R885 S.n1706 S.t579 3.904
R886 S.n1703 S.t788 3.904
R887 S.n1690 S.n1689 3.904
R888 S.n664 S.n663 3.904
R889 S.n675 S.t2163 3.904
R890 S.n672 S.t1662 3.904
R891 S.n667 S.n666 3.904
R892 S.n647 S.n646 3.904
R893 S.n658 S.t521 3.904
R894 S.n655 S.t2534 3.904
R895 S.n650 S.n649 3.904
R896 S.n183 S.t2226 3.904
R897 S.n379 S.n378 3.904
R898 S.n390 S.t621 3.904
R899 S.n387 S.t855 3.904
R900 S.n382 S.n381 3.904
R901 S.n1606 S.n1605 3.904
R902 S.n1619 S.t639 3.904
R903 S.n1616 S.t888 3.904
R904 S.n1603 S.n1602 3.904
R905 S.n7793 S.t1439 3.904
R906 S.n7750 S.n7749 3.904
R907 S.n7764 S.t285 3.904
R908 S.n7767 S.t1463 3.904
R909 S.n7747 S.n7746 3.904
R910 S.n7229 S.n7228 3.904
R911 S.n7240 S.t1786 3.904
R912 S.n7237 S.t826 3.904
R913 S.n7226 S.n7225 3.904
R914 S.n6788 S.n6787 3.904
R915 S.n6803 S.t2238 3.904
R916 S.n6800 S.t869 3.904
R917 S.n6785 S.n6784 3.904
R918 S.n6483 S.n6482 3.904
R919 S.n6494 S.t1195 3.904
R920 S.n6491 S.t2288 3.904
R921 S.n6480 S.n6479 3.904
R922 S.n6046 S.n6045 3.904
R923 S.n6061 S.t1155 3.904
R924 S.n6058 S.t217 3.904
R925 S.n6043 S.n6042 3.904
R926 S.n5728 S.n5727 3.904
R927 S.n5739 S.t558 3.904
R928 S.n5736 S.t1691 3.904
R929 S.n5725 S.n5724 3.904
R930 S.n5281 S.n5280 3.904
R931 S.n5296 S.t587 3.904
R932 S.n5293 S.t2157 3.904
R933 S.n5278 S.n5277 3.904
R934 S.n4947 S.n4946 3.904
R935 S.n4958 S.t2451 3.904
R936 S.n4955 S.t1136 3.904
R937 S.n4944 S.n4943 3.904
R938 S.n4504 S.n4503 3.904
R939 S.n4519 S.t2488 3.904
R940 S.n4516 S.t1547 3.904
R941 S.n4501 S.n4500 3.904
R942 S.n4157 S.n4156 3.904
R943 S.n4168 S.t1908 3.904
R944 S.n4165 S.t565 3.904
R945 S.n4154 S.n4153 3.904
R946 S.n3704 S.n3703 3.904
R947 S.n3719 S.t1933 3.904
R948 S.n3716 S.t1005 3.904
R949 S.n3701 S.n3700 3.904
R950 S.n3310 S.n3309 3.904
R951 S.n3321 S.t1326 3.904
R952 S.n3318 S.t2456 3.904
R953 S.n3307 S.n3306 3.904
R954 S.n2892 S.n2891 3.904
R955 S.n2907 S.t1363 3.904
R956 S.n2904 S.t396 3.904
R957 S.n2889 S.n2888 3.904
R958 S.n2454 S.n2453 3.904
R959 S.n2465 S.t703 3.904
R960 S.n2462 S.t1913 3.904
R961 S.n2451 S.n2450 3.904
R962 S.n2047 S.n2046 3.904
R963 S.n2064 S.t1172 3.904
R964 S.n2061 S.t2338 3.904
R965 S.n2044 S.n2043 3.904
R966 S.n1175 S.n1174 3.904
R967 S.n1184 S.t143 3.904
R968 S.n1181 S.t1795 3.904
R969 S.n1172 S.n1171 3.904
R970 S.n969 S.t1365 3.904
R971 S.n399 S.n398 3.904
R972 S.n410 S.t2279 3.904
R973 S.n407 S.t2499 3.904
R974 S.n402 S.n401 3.904
R975 S.n8506 S.t1147 3.904
R976 S.n8461 S.n8460 3.904
R977 S.n8476 S.t2503 3.904
R978 S.n8479 S.t1173 3.904
R979 S.n8464 S.n8463 3.904
R980 S.n7799 S.n7798 3.904
R981 S.n7810 S.t1492 3.904
R982 S.n7807 S.t576 3.904
R983 S.n7802 S.n7801 3.904
R984 S.n7542 S.n7541 3.904
R985 S.n7562 S.t1948 3.904
R986 S.n7559 S.t604 3.904
R987 S.n7545 S.n7544 3.904
R988 S.n7246 S.n7245 3.904
R989 S.n7257 S.t920 3.904
R990 S.n7254 S.t2470 3.904
R991 S.n7249 S.n7248 3.904
R992 S.n6812 S.n6811 3.904
R993 S.n6832 S.t1379 3.904
R994 S.n6829 S.t126 3.904
R995 S.n6815 S.n6814 3.904
R996 S.n6500 S.n6499 3.904
R997 S.n6511 S.t468 3.904
R998 S.n6508 S.t1435 3.904
R999 S.n6503 S.n6502 3.904
R1000 S.n6070 S.n6069 3.904
R1001 S.n6090 S.t280 3.904
R1002 S.n6087 S.t1882 3.904
R1003 S.n6073 S.n6072 3.904
R1004 S.n5745 S.n5744 3.904
R1005 S.n5756 S.t2198 3.904
R1006 S.n5753 S.t821 3.904
R1007 S.n5748 S.n5747 3.904
R1008 S.n5305 S.n5304 3.904
R1009 S.n5325 S.t2235 3.904
R1010 S.n5322 S.t1294 3.904
R1011 S.n5308 S.n5307 3.904
R1012 S.n4964 S.n4963 3.904
R1013 S.n4975 S.t1582 3.904
R1014 S.n4972 S.t257 3.904
R1015 S.n4967 S.n4966 3.904
R1016 S.n4528 S.n4527 3.904
R1017 S.n4548 S.t1612 3.904
R1018 S.n4545 S.t685 3.904
R1019 S.n4531 S.n4530 3.904
R1020 S.n4174 S.n4173 3.904
R1021 S.n4185 S.t1048 3.904
R1022 S.n4182 S.t2208 3.904
R1023 S.n4177 S.n4176 3.904
R1024 S.n3728 S.n3727 3.904
R1025 S.n3748 S.t1074 3.904
R1026 S.n3745 S.t105 3.904
R1027 S.n3731 S.n3730 3.904
R1028 S.n3327 S.n3326 3.904
R1029 S.n3338 S.t445 3.904
R1030 S.n3335 S.t1587 3.904
R1031 S.n3330 S.n3329 3.904
R1032 S.n2916 S.n2915 3.904
R1033 S.n2936 S.t612 3.904
R1034 S.n2933 S.t2048 3.904
R1035 S.n2919 S.n2918 3.904
R1036 S.n2471 S.n2470 3.904
R1037 S.n2482 S.t2362 3.904
R1038 S.n2479 S.t1814 3.904
R1039 S.n2474 S.n2473 3.904
R1040 S.n2073 S.n2072 3.904
R1041 S.n2093 S.t2316 3.904
R1042 S.n2090 S.t2563 3.904
R1043 S.n2076 S.n2075 3.904
R1044 S.n1190 S.n1189 3.904
R1045 S.n1201 S.t1420 3.904
R1046 S.n1198 S.t925 3.904
R1047 S.n1193 S.n1192 3.904
R1048 S.n1628 S.n1627 3.904
R1049 S.n1648 S.t2298 3.904
R1050 S.n1645 S.t2530 3.904
R1051 S.n1631 S.n1630 3.904
R1052 S.n631 S.n630 3.904
R1053 S.n642 S.t1393 3.904
R1054 S.n639 S.t891 3.904
R1055 S.n634 S.n633 3.904
R1056 S.n614 S.n613 3.904
R1057 S.n625 S.t2252 3.904
R1058 S.n622 S.t1765 3.904
R1059 S.n617 S.n616 3.904
R1060 S.n170 S.t696 3.904
R1061 S.n338 S.n337 3.904
R1062 S.n349 S.t1742 3.904
R1063 S.n346 S.t386 3.904
R1064 S.n341 S.n340 3.904
R1065 S.n1547 S.n1546 3.904
R1066 S.n1560 S.t2213 3.904
R1067 S.n1557 S.t996 3.904
R1068 S.n1544 S.n1543 3.904
R1069 S.n6458 S.t1498 3.904
R1070 S.n6278 S.n6277 3.904
R1071 S.n6292 S.t351 3.904
R1072 S.n6295 S.t1838 3.904
R1073 S.n6275 S.n6274 3.904
R1074 S.n5692 S.n5691 3.904
R1075 S.n5703 S.t2150 3.904
R1076 S.n5700 S.t927 3.904
R1077 S.n5689 S.n5688 3.904
R1078 S.n5220 S.n5219 3.904
R1079 S.n5235 S.t2304 3.904
R1080 S.n5232 S.t1240 3.904
R1081 S.n5217 S.n5216 3.904
R1082 S.n4911 S.n4910 3.904
R1083 S.n4922 S.t1542 3.904
R1084 S.n4919 S.t323 3.904
R1085 S.n4908 S.n4907 3.904
R1086 S.n4443 S.n4442 3.904
R1087 S.n4458 S.t1713 3.904
R1088 S.n4455 S.t757 3.904
R1089 S.n4440 S.n4439 3.904
R1090 S.n4121 S.n4120 3.904
R1091 S.n4132 S.t1121 3.904
R1092 S.n4129 S.t2284 3.904
R1093 S.n4118 S.n4117 3.904
R1094 S.n3643 S.n3642 3.904
R1095 S.n3658 S.t1149 3.904
R1096 S.n3655 S.t206 3.904
R1097 S.n3640 S.n3639 3.904
R1098 S.n3274 S.n3273 3.904
R1099 S.n3285 S.t546 3.904
R1100 S.n3282 S.t1682 3.904
R1101 S.n3271 S.n3270 3.904
R1102 S.n2831 S.n2830 3.904
R1103 S.n2846 S.t577 3.904
R1104 S.n2843 S.t2146 3.904
R1105 S.n2828 S.n2827 3.904
R1106 S.n2418 S.n2417 3.904
R1107 S.n2429 S.t2437 3.904
R1108 S.n2426 S.t1127 3.904
R1109 S.n2415 S.n2414 3.904
R1110 S.n1984 S.n1983 3.904
R1111 S.n2001 S.t263 3.904
R1112 S.n1998 S.t1539 3.904
R1113 S.n1981 S.n1980 3.904
R1114 S.n1141 S.n1140 3.904
R1115 S.n1150 S.t1899 3.904
R1116 S.n1147 S.t795 3.904
R1117 S.n1138 S.n1137 3.904
R1118 S.n965 S.t580 3.904
R1119 S.n358 S.n357 3.904
R1120 S.n369 S.t1482 3.904
R1121 S.n366 S.t1728 3.904
R1122 S.n361 S.n360 3.904
R1123 S.n7221 S.t1700 3.904
R1124 S.n7024 S.n7023 3.904
R1125 S.n7039 S.t591 3.904
R1126 S.n7042 S.t1745 3.904
R1127 S.n7027 S.n7026 3.904
R1128 S.n6464 S.n6463 3.904
R1129 S.n6475 S.t2057 3.904
R1130 S.n6472 S.t635 3.904
R1131 S.n6467 S.n6466 3.904
R1132 S.n6009 S.n6008 3.904
R1133 S.n6029 S.t2008 3.904
R1134 S.n6026 S.t972 3.904
R1135 S.n6012 S.n6011 3.904
R1136 S.n5709 S.n5708 3.904
R1137 S.n5720 S.t1290 3.904
R1138 S.n5717 S.t2567 3.904
R1139 S.n5712 S.n5711 3.904
R1140 S.n5244 S.n5243 3.904
R1141 S.n5264 S.t1449 3.904
R1142 S.n5261 S.t514 3.904
R1143 S.n5247 S.n5246 3.904
R1144 S.n4928 S.n4927 3.904
R1145 S.n4939 S.t801 3.904
R1146 S.n4936 S.t1984 3.904
R1147 S.n4931 S.n4930 3.904
R1148 S.n4467 S.n4466 3.904
R1149 S.n4487 S.t844 3.904
R1150 S.n4484 S.t2411 3.904
R1151 S.n4470 S.n4469 3.904
R1152 S.n4138 S.n4137 3.904
R1153 S.n4149 S.t242 3.904
R1154 S.n4146 S.t1430 3.904
R1155 S.n4141 S.n4140 3.904
R1156 S.n3667 S.n3666 3.904
R1157 S.n3687 S.t271 3.904
R1158 S.n3684 S.t1874 3.904
R1159 S.n3670 S.n3669 3.904
R1160 S.n3291 S.n3290 3.904
R1161 S.n3302 S.t2188 3.904
R1162 S.n3299 S.t807 3.904
R1163 S.n3294 S.n3293 3.904
R1164 S.n2855 S.n2854 3.904
R1165 S.n2875 S.t2222 3.904
R1166 S.n2872 S.t1283 3.904
R1167 S.n2858 S.n2857 3.904
R1168 S.n2435 S.n2434 3.904
R1169 S.n2446 S.t1573 3.904
R1170 S.n2443 S.t249 3.904
R1171 S.n2438 S.n2437 3.904
R1172 S.n2010 S.n2009 3.904
R1173 S.n2030 S.t1927 3.904
R1174 S.n2027 S.t678 3.904
R1175 S.n2013 S.n2012 3.904
R1176 S.n1156 S.n1155 3.904
R1177 S.n1167 S.t1039 3.904
R1178 S.n1164 S.t2443 3.904
R1179 S.n1159 S.n1158 3.904
R1180 S.n1569 S.n1568 3.904
R1181 S.n1589 S.t1464 3.904
R1182 S.n1586 S.t89 3.904
R1183 S.n1572 S.n1571 3.904
R1184 S.n598 S.n597 3.904
R1185 S.n609 S.t431 3.904
R1186 S.n606 S.t90 3.904
R1187 S.n601 S.n600 3.904
R1188 S.n581 S.n580 3.904
R1189 S.n592 S.t1311 3.904
R1190 S.n589 S.t235 3.904
R1191 S.n584 S.n583 3.904
R1192 S.n157 S.t2425 3.904
R1193 S.n317 S.n316 3.904
R1194 S.n328 S.t814 3.904
R1195 S.n325 S.t2133 3.904
R1196 S.n320 S.n319 3.904
R1197 S.n1488 S.n1487 3.904
R1198 S.n1501 S.t1433 3.904
R1199 S.n1498 S.t198 3.904
R1200 S.n1485 S.n1484 3.904
R1201 S.n4886 S.t2065 3.904
R1202 S.n4736 S.n4735 3.904
R1203 S.n4750 S.t951 3.904
R1204 S.n4753 S.t2371 3.904
R1205 S.n4733 S.n4732 3.904
R1206 S.n4085 S.n4084 3.904
R1207 S.n4096 S.t202 3.904
R1208 S.n4093 S.t1490 3.904
R1209 S.n4082 S.n4081 3.904
R1210 S.n3582 S.n3581 3.904
R1211 S.n3597 S.t341 3.904
R1212 S.n3594 S.t1822 3.904
R1213 S.n3579 S.n3578 3.904
R1214 S.n3238 S.n3237 3.904
R1215 S.n3249 S.t2138 3.904
R1216 S.n3246 S.t912 3.904
R1217 S.n3235 S.n3234 3.904
R1218 S.n2770 S.n2769 3.904
R1219 S.n2785 S.t2297 3.904
R1220 S.n2782 S.t1374 3.904
R1221 S.n2767 S.n2766 3.904
R1222 S.n2382 S.n2381 3.904
R1223 S.n2393 S.t1656 3.904
R1224 S.n2390 S.t315 3.904
R1225 S.n2379 S.n2378 3.904
R1226 S.n1921 S.n1920 3.904
R1227 S.n1938 S.t1989 3.904
R1228 S.n1935 S.t750 3.904
R1229 S.n1918 S.n1917 3.904
R1230 S.n1107 S.n1106 3.904
R1231 S.n1116 S.t1111 3.904
R1232 S.n1113 S.t2542 3.904
R1233 S.n1104 S.n1103 3.904
R1234 S.n961 S.t1560 3.904
R1235 S.n47 S.n46 3.904
R1236 S.n50 S.t2461 3.904
R1237 S.n53 S.t1268 3.904
R1238 S.n56 S.n55 3.904
R1239 S.n5684 S.t1797 3.904
R1240 S.n5517 S.n5516 3.904
R1241 S.n5532 S.t647 3.904
R1242 S.n5535 S.t2107 3.904
R1243 S.n5520 S.n5519 3.904
R1244 S.n4892 S.n4891 3.904
R1245 S.n4903 S.t2404 3.904
R1246 S.n4900 S.t1203 3.904
R1247 S.n4895 S.n4894 3.904
R1248 S.n4406 S.n4405 3.904
R1249 S.n4426 S.t2589 3.904
R1250 S.n4423 S.t1514 3.904
R1251 S.n4409 S.n4408 3.904
R1252 S.n4102 S.n4101 3.904
R1253 S.n4113 S.t1869 3.904
R1254 S.n4110 S.t625 3.904
R1255 S.n4105 S.n4104 3.904
R1256 S.n3606 S.n3605 3.904
R1257 S.n3626 S.t1999 3.904
R1258 S.n3623 S.t1083 3.904
R1259 S.n3609 S.n3608 3.904
R1260 S.n3255 S.n3254 3.904
R1261 S.n3266 S.t1411 3.904
R1262 S.n3263 S.t2553 3.904
R1263 S.n3258 S.n3257 3.904
R1264 S.n2794 S.n2793 3.904
R1265 S.n2814 S.t1441 3.904
R1266 S.n2811 S.t501 3.904
R1267 S.n2797 S.n2796 3.904
R1268 S.n2399 S.n2398 3.904
R1269 S.n2410 S.t786 3.904
R1270 S.n2407 S.t1980 3.904
R1271 S.n2402 S.n2401 3.904
R1272 S.n1947 S.n1946 3.904
R1273 S.n1967 S.t1139 3.904
R1274 S.n1964 S.t2402 3.904
R1275 S.n1950 S.n1949 3.904
R1276 S.n1122 S.n1121 3.904
R1277 S.n1133 S.t233 3.904
R1278 S.n1130 S.t1670 3.904
R1279 S.n1125 S.n1124 3.904
R1280 S.n1510 S.n1509 3.904
R1281 S.n1530 S.t569 3.904
R1282 S.n1527 S.t1865 3.904
R1283 S.n1513 S.n1512 3.904
R1284 S.n565 S.n564 3.904
R1285 S.n576 S.t2175 3.904
R1286 S.n573 S.t1117 3.904
R1287 S.n568 S.n567 3.904
R1288 S.n548 S.n547 3.904
R1289 S.n559 S.t532 3.904
R1290 S.n556 S.t1972 3.904
R1291 S.n551 S.n550 3.904
R1292 S.n144 S.t1642 3.904
R1293 S.n276 S.n275 3.904
R1294 S.n287 S.t2561 3.904
R1295 S.n284 S.t1364 3.904
R1296 S.n279 S.n278 3.904
R1297 S.n1429 S.n1428 3.904
R1298 S.n1442 S.t630 3.904
R1299 S.n1439 S.t1934 3.904
R1300 S.n1426 S.n1425 3.904
R1301 S.n3213 S.t112 3.904
R1302 S.n3124 S.n3123 3.904
R1303 S.n3138 S.t1501 3.904
R1304 S.n3141 S.t448 3.904
R1305 S.n3121 S.n3120 3.904
R1306 S.n2346 S.n2345 3.904
R1307 S.n2357 S.t743 3.904
R1308 S.n2354 S.t2054 3.904
R1309 S.n2343 S.n2342 3.904
R1310 S.n1858 S.n1857 3.904
R1311 S.n1875 S.t1211 3.904
R1312 S.n1872 S.t2363 3.904
R1313 S.n1855 S.n1854 3.904
R1314 S.n1073 S.n1072 3.904
R1315 S.n1082 S.t190 3.904
R1316 S.n1079 S.t1773 3.904
R1317 S.n1070 S.n1069 3.904
R1318 S.n957 S.t774 3.904
R1319 S.n296 S.n295 3.904
R1320 S.n307 S.t1687 3.904
R1321 S.n304 S.t490 3.904
R1322 S.n299 S.n298 3.904
R1323 S.n4077 S.t2349 3.904
R1324 S.n3940 S.n3939 3.904
R1325 S.n3955 S.t1222 3.904
R1326 S.n3958 S.t161 3.904
R1327 S.n3943 S.n3942 3.904
R1328 S.n3219 S.n3218 3.904
R1329 S.n3230 S.t493 3.904
R1330 S.n3227 S.t1784 3.904
R1331 S.n3222 S.n3221 3.904
R1332 S.n2733 S.n2732 3.904
R1333 S.n2753 S.t640 3.904
R1334 S.n2750 S.t2093 3.904
R1335 S.n2736 S.n2735 3.904
R1336 S.n2363 S.n2362 3.904
R1337 S.n2374 S.t2394 3.904
R1338 S.n2371 S.t1194 3.904
R1339 S.n2366 S.n2365 3.904
R1340 S.n1884 S.n1883 3.904
R1341 S.n1904 S.t332 3.904
R1342 S.n1901 S.t1613 3.904
R1343 S.n1887 S.n1886 3.904
R1344 S.n1088 S.n1087 3.904
R1345 S.n1099 S.t1965 3.904
R1346 S.n1096 S.t899 3.904
R1347 S.n1091 S.n1090 3.904
R1348 S.n1451 S.n1450 3.904
R1349 S.n1471 S.t2286 3.904
R1350 S.n1454 S.t1075 3.904
R1351 S.n1457 S.n1456 3.904
R1352 S.n532 S.n531 3.904
R1353 S.n543 S.t1403 3.904
R1354 S.n540 S.t310 3.904
R1355 S.n535 S.n534 3.904
R1356 S.n515 S.n514 3.904
R1357 S.n526 S.t2260 3.904
R1358 S.n523 S.t1185 3.904
R1359 S.n518 S.n517 3.904
R1360 S.n131 S.t732 3.904
R1361 S.n235 S.n234 3.904
R1362 S.n246 S.t1789 3.904
R1363 S.n243 S.t434 3.904
R1364 S.n238 S.n237 3.904
R1365 S.n1368 S.n1367 3.904
R1366 S.n1383 S.t2351 3.904
R1367 S.n1380 S.t1042 3.904
R1368 S.n1365 S.n1364 3.904
R1369 S.n1048 S.t1002 3.904
R1370 S.n953 S.t2519 3.904
R1371 S.n255 S.n254 3.904
R1372 S.n266 S.t919 3.904
R1373 S.n263 S.t2225 3.904
R1374 S.n258 S.n257 3.904
R1375 S.n2338 S.t406 3.904
R1376 S.n2293 S.n2292 3.904
R1377 S.n2308 S.t2072 3.904
R1378 S.n2311 S.t705 3.904
R1379 S.n2296 S.n2295 3.904
R1380 S.n1054 S.n1053 3.904
R1381 S.n1065 S.t1069 3.904
R1382 S.n1062 S.t97 3.904
R1383 S.n1057 S.n1056 3.904
R1384 S.n1392 S.n1391 3.904
R1385 S.n1412 S.t1493 3.904
R1386 S.n1409 S.t148 3.904
R1387 S.n1395 S.n1394 3.904
R1388 S.n499 S.n498 3.904
R1389 S.n510 S.t478 3.904
R1390 S.n507 S.t2039 3.904
R1391 S.n502 S.n501 3.904
R1392 S.n482 S.n481 3.904
R1393 S.n493 S.t1356 3.904
R1394 S.n490 S.t389 3.904
R1395 S.n485 S.n484 3.904
R1396 S.n882 S.t1688 3.904
R1397 S.n884 S.t886 3.904
R1398 S.n740 S.n739 3.904
R1399 S.n750 S.t537 3.904
R1400 S.n753 S.t197 3.904
R1401 S.n743 S.n742 3.904
R1402 S.n1349 S.n1348 3.904
R1403 S.n1360 S.t1269 3.904
R1404 S.n1357 S.t1148 3.904
R1405 S.n1352 S.n1351 3.904
R1406 S.n1026 S.n1025 3.904
R1407 S.n1335 S.t506 3.904
R1408 S.n1338 S.t2384 3.904
R1409 S.n1341 S.n1340 3.904
R1410 S.n2636 S.n2635 3.904
R1411 S.n2648 S.t1301 3.904
R1412 S.n2651 S.t1640 3.904
R1413 S.n2639 S.n2638 3.904
R1414 S.n2315 S.n2314 3.904
R1415 S.n2621 S.t536 3.904
R1416 S.n2624 S.t745 3.904
R1417 S.n2627 S.n2626 3.904
R1418 S.n3163 S.n3162 3.904
R1419 S.n3175 S.t2177 3.904
R1420 S.n3178 S.t1680 3.904
R1421 S.n3166 S.n3165 3.904
R1422 S.n3145 S.n3144 3.904
R1423 S.n3148 S.t566 3.904
R1424 S.n3151 S.t770 3.904
R1425 S.n3154 S.n3153 3.904
R1426 S.n3980 S.n3979 3.904
R1427 S.n3992 S.t2206 3.904
R1428 S.n3995 S.t1707 3.904
R1429 S.n3983 S.n3982 3.904
R1430 S.n3962 S.n3961 3.904
R1431 S.n3965 S.t588 3.904
R1432 S.n3968 S.t800 3.904
R1433 S.n3971 S.n3970 3.904
R1434 S.n4775 S.n4774 3.904
R1435 S.n4787 S.t2232 3.904
R1436 S.n4790 S.t1740 3.904
R1437 S.n4778 S.n4777 3.904
R1438 S.n4757 S.n4756 3.904
R1439 S.n4760 S.t477 3.904
R1440 S.n4763 S.t830 3.904
R1441 S.n4766 S.n4765 3.904
R1442 S.n5557 S.n5556 3.904
R1443 S.n5569 S.t2257 3.904
R1444 S.n5572 S.t1615 3.904
R1445 S.n5560 S.n5559 3.904
R1446 S.n5539 S.n5538 3.904
R1447 S.n5542 S.t508 3.904
R1448 S.n5545 S.t860 3.904
R1449 S.n5548 S.n5547 3.904
R1450 S.n6317 S.n6316 3.904
R1451 S.n6329 S.t2282 3.904
R1452 S.n6332 S.t1644 3.904
R1453 S.n6320 S.n6319 3.904
R1454 S.n6299 S.n6298 3.904
R1455 S.n6302 S.t895 3.904
R1456 S.n6305 S.t896 3.904
R1457 S.n6308 S.n6307 3.904
R1458 S.n7064 S.n7063 3.904
R1459 S.n7076 S.t1836 3.904
R1460 S.n7079 S.t2062 3.904
R1461 S.n7067 S.n7066 3.904
R1462 S.n7046 S.n7045 3.904
R1463 S.n7049 S.t933 3.904
R1464 S.n7052 S.t452 3.904
R1465 S.n7055 S.n7054 3.904
R1466 S.n8075 S.n8074 3.904
R1467 S.n8087 S.t1868 3.904
R1468 S.n8090 S.t2094 3.904
R1469 S.n8078 S.n8077 3.904
R1470 S.n7771 S.n7770 3.904
R1471 S.n8060 S.t602 3.904
R1472 S.n8063 S.t481 3.904
R1473 S.n8066 S.n8065 3.904
R1474 S.n8787 S.n8786 3.904
R1475 S.n8799 S.t1591 3.904
R1476 S.n8802 S.t267 3.904
R1477 S.n8790 S.n8789 3.904
R1478 S.n8483 S.n8482 3.904
R1479 S.n8772 S.t1170 3.904
R1480 S.n8775 S.t85 3.904
R1481 S.n8778 S.n8777 3.904
R1482 S.n9191 S.n9190 3.904
R1483 S.n9203 S.t2063 3.904
R1484 S.n9206 S.t833 3.904
R1485 S.n9194 S.n9193 3.904
R1486 S.n9173 S.n9172 3.904
R1487 S.n9176 S.t1756 3.904
R1488 S.n9179 S.t677 3.904
R1489 S.n9182 S.n9181 3.904
R1490 S.n9868 S.n9867 3.904
R1491 S.n9880 S.t124 3.904
R1492 S.n9883 S.t1444 3.904
R1493 S.n9871 S.n9870 3.904
R1494 S.n9850 S.n9849 3.904
R1495 S.n9853 S.t2330 3.904
R1496 S.n9856 S.t1006 3.904
R1497 S.n9859 S.n9858 3.904
R1498 S.n10526 S.n10525 3.904
R1499 S.n10538 S.t428 3.904
R1500 S.n10541 S.t2002 3.904
R1501 S.n10529 S.n10528 3.904
R1502 S.n10508 S.n10507 3.904
R1503 S.n10511 S.t387 3.904
R1504 S.n10514 S.t1546 3.904
R1505 S.n10517 S.n10516 3.904
R1506 S.n11149 S.n11148 3.904
R1507 S.n11161 S.t1037 3.904
R1508 S.n11164 S.t7 3.904
R1509 S.n11152 S.n11151 3.904
R1510 S.n11131 S.n11130 3.904
R1511 S.n11134 S.t997 3.904
R1512 S.n11137 S.t2156 3.904
R1513 S.n11140 S.n11139 3.904
R1514 S.n11727 S.n11726 3.904
R1515 S.n11739 S.t1570 3.904
R1516 S.n11742 S.t653 3.904
R1517 S.n11730 S.n11729 3.904
R1518 S.n12019 S.n12018 3.904
R1519 S.n12029 S.t1447 3.904
R1520 S.n12032 S.t214 3.904
R1521 S.n12022 S.n12021 3.904
R1522 S.n12896 S.n12895 3.904
R1523 S.n12908 S.t1981 3.904
R1524 S.n12911 S.t1125 3.904
R1525 S.n12899 S.n12898 3.904
R1526 S.n12600 S.n12599 3.904
R1527 S.n12880 S.t902 3.904
R1528 S.n12883 S.t610 3.904
R1529 S.n12886 S.n12885 3.904
R1530 S.n12482 S.t1440 3.904
R1531 S.n12480 S.t1973 3.904
R1532 S.n1798 S.t321 3.904
R1533 S.n1800 S.t2562 3.904
R1534 S.n1321 S.n1320 3.904
R1535 S.n1329 S.t1647 3.904
R1536 S.n1332 S.t1329 3.904
R1537 S.n1324 S.n1323 3.904
R1538 S.n2659 S.n2658 3.904
R1539 S.n2678 S.t417 3.904
R1540 S.n2681 S.t2296 3.904
R1541 S.n2656 S.n2655 3.904
R1542 S.n12486 S.t578 3.904
R1543 S.n12484 S.t1118 3.904
R1544 S.n12933 S.n12932 3.904
R1545 S.n12930 S.t2545 3.904
R1546 S.n12927 S.t2264 3.904
R1547 S.n12924 S.n12923 3.904
R1548 S.n12919 S.n12918 3.904
R1549 S.n12939 S.t1131 3.904
R1550 S.n12942 S.t357 3.904
R1551 S.n12916 S.n12915 3.904
R1552 S.n12040 S.n12039 3.904
R1553 S.n12044 S.t679 3.904
R1554 S.n12047 S.t1883 3.904
R1555 S.n12037 S.n12036 3.904
R1556 S.n11750 S.n11749 3.904
R1557 S.n11755 S.t702 3.904
R1558 S.n11758 S.t2307 3.904
R1559 S.n11747 S.n11746 3.904
R1560 S.n11186 S.n11185 3.904
R1561 S.n11183 S.t93 3.904
R1562 S.n11180 S.t1293 3.904
R1563 S.n11177 S.n11176 3.904
R1564 S.n11172 S.n11171 3.904
R1565 S.n11192 S.t140 3.904
R1566 S.n11195 S.t1719 3.904
R1567 S.n11169 S.n11168 3.904
R1568 S.n10563 S.n10562 3.904
R1569 S.n10560 S.t2036 3.904
R1570 S.n10557 S.t684 3.904
R1571 S.n10554 S.n10553 3.904
R1572 S.n10549 S.n10548 3.904
R1573 S.n10569 S.t2077 3.904
R1574 S.n10572 S.t1150 3.904
R1575 S.n10546 S.n10545 3.904
R1576 S.n9905 S.n9904 3.904
R1577 S.n9902 S.t1471 3.904
R1578 S.n9899 S.t102 3.904
R1579 S.n9896 S.n9895 3.904
R1580 S.n9891 S.n9890 3.904
R1581 S.n9911 S.t1794 3.904
R1582 S.n9914 S.t583 3.904
R1583 S.n9888 S.n9887 3.904
R1584 S.n9228 S.n9227 3.904
R1585 S.n9225 S.t878 3.904
R1586 S.n9222 S.t2334 3.904
R1587 S.n9219 S.n9218 3.904
R1588 S.n9214 S.n9213 3.904
R1589 S.n9234 S.t1351 3.904
R1590 S.n9237 S.t2478 3.904
R1591 S.n9211 S.n9210 3.904
R1592 S.n8824 S.n8823 3.904
R1593 S.n8821 S.t295 3.904
R1594 S.n8818 S.t2158 3.904
R1595 S.n8815 S.n8814 3.904
R1596 S.n8810 S.n8809 3.904
R1597 S.n8830 S.t1030 3.904
R1598 S.n8833 S.t1263 3.904
R1599 S.n8807 S.n8806 3.904
R1600 S.n8112 S.n8111 3.904
R1601 S.n8109 S.t23 3.904
R1602 S.n8106 S.t2129 3.904
R1603 S.n8103 S.n8102 3.904
R1604 S.n8098 S.n8097 3.904
R1605 S.n8118 S.t1000 3.904
R1606 S.n8121 S.t1229 3.904
R1607 S.n8095 S.n8094 3.904
R1608 S.n7101 S.n7100 3.904
R1609 S.n7098 S.t2576 3.904
R1610 S.n7095 S.t2097 3.904
R1611 S.n7092 S.n7091 3.904
R1612 S.n7087 S.n7086 3.904
R1613 S.n7107 S.t970 3.904
R1614 S.n7110 S.t1200 3.904
R1615 S.n7084 S.n7083 3.904
R1616 S.n6354 S.n6353 3.904
R1617 S.n6351 S.t2541 3.904
R1618 S.n6348 S.t2538 3.904
R1619 S.n6345 S.n6344 3.904
R1620 S.n6340 S.n6339 3.904
R1621 S.n6360 S.t1426 3.904
R1622 S.n6363 S.t775 3.904
R1623 S.n6337 S.n6336 3.904
R1624 S.n5594 S.n5593 3.904
R1625 S.n5591 S.t2154 3.904
R1626 S.n5588 S.t2505 3.904
R1627 S.n5585 S.n5584 3.904
R1628 S.n5580 S.n5579 3.904
R1629 S.n5600 S.t1399 3.904
R1630 S.n5603 S.t903 3.904
R1631 S.n5577 S.n5576 3.904
R1632 S.n4812 S.n4811 3.904
R1633 S.n4809 S.t2259 3.904
R1634 S.n4806 S.t2475 3.904
R1635 S.n4803 S.n4802 3.904
R1636 S.n4798 S.n4797 3.904
R1637 S.n4818 S.t1370 3.904
R1638 S.n4821 S.t866 3.904
R1639 S.n4795 S.n4794 3.904
R1640 S.n4020 S.n4019 3.904
R1641 S.n4017 S.t2234 3.904
R1642 S.n4014 S.t2450 3.904
R1643 S.n4011 S.n4010 3.904
R1644 S.n4006 S.n4005 3.904
R1645 S.n3998 S.t1348 3.904
R1646 S.n4026 S.t836 3.904
R1647 S.n4003 S.n4002 3.904
R1648 S.n3498 S.n3497 3.904
R1649 S.n3495 S.t2209 3.904
R1650 S.n3492 S.t2421 3.904
R1651 S.n3191 S.n3190 3.904
R1652 S.n3186 S.n3185 3.904
R1653 S.n3504 S.t1315 3.904
R1654 S.n3507 S.t804 3.904
R1655 S.n3183 S.n3182 3.904
R1656 S.n2673 S.n2672 3.904
R1657 S.n2670 S.t2180 3.904
R1658 S.n2667 S.t2396 3.904
R1659 S.n2664 S.n2663 3.904
R1660 S.n2686 S.t1488 3.904
R1661 S.n2683 S.t1720 3.904
R1662 S.n2603 S.n2602 3.904
R1663 S.n2615 S.t296 3.904
R1664 S.n2618 S.t586 3.904
R1665 S.n2606 S.n2605 3.904
R1666 S.n3515 S.n3514 3.904
R1667 S.n3519 S.t437 3.904
R1668 S.n3522 S.t938 3.904
R1669 S.n3512 S.n3511 3.904
R1670 S.n12490 S.t2331 3.904
R1671 S.n12488 S.t237 3.904
R1672 S.n12677 S.n12676 3.904
R1673 S.n12682 S.t1825 3.904
R1674 S.n12685 S.t1406 3.904
R1675 S.n12674 S.n12673 3.904
R1676 S.n12950 S.n12949 3.904
R1677 S.n12954 S.t252 3.904
R1678 S.n12957 S.t2011 3.904
R1679 S.n12947 S.n12946 3.904
R1680 S.n12055 S.n12054 3.904
R1681 S.n12060 S.t2339 3.904
R1682 S.n12063 S.t1020 3.904
R1683 S.n12052 S.n12051 3.904
R1684 S.n11766 S.n11765 3.904
R1685 S.n11770 S.t2361 3.904
R1686 S.n11773 S.t1451 3.904
R1687 S.n11763 S.n11762 3.904
R1688 S.n11447 S.n11446 3.904
R1689 S.n11452 S.t1768 3.904
R1690 S.n11455 S.t409 3.904
R1691 S.n11444 S.n11443 3.904
R1692 S.n11203 S.n11202 3.904
R1693 S.n11207 S.t1810 3.904
R1694 S.n11210 S.t848 3.904
R1695 S.n11200 S.n11199 3.904
R1696 S.n10826 S.n10825 3.904
R1697 S.n10831 S.t1181 3.904
R1698 S.n10834 S.t2344 3.904
R1699 S.n10823 S.n10822 3.904
R1700 S.n10580 S.n10579 3.904
R1701 S.n10584 S.t1215 3.904
R1702 S.n10587 S.t274 3.904
R1703 S.n10577 S.n10576 3.904
R1704 S.n10173 S.n10172 3.904
R1705 S.n10178 S.t609 3.904
R1706 S.n10181 S.t1777 3.904
R1707 S.n10170 S.n10169 3.904
R1708 S.n9922 S.n9921 3.904
R1709 S.n9926 S.t1064 3.904
R1710 S.n9929 S.t2230 3.904
R1711 S.n9919 S.n9918 3.904
R1712 S.n9497 S.n9496 3.904
R1713 S.n9502 S.t2522 3.904
R1714 S.n9505 S.t1324 3.904
R1715 S.n9494 S.n9493 3.904
R1716 S.n9245 S.n9244 3.904
R1717 S.n9249 S.t166 3.904
R1718 S.n9252 S.t408 3.904
R1719 S.n9242 S.n9241 3.904
R1720 S.n8630 S.n8629 3.904
R1721 S.n8635 S.t1763 3.904
R1722 S.n8638 S.t1295 3.904
R1723 S.n8627 S.n8626 3.904
R1724 S.n8841 S.n8840 3.904
R1725 S.n8845 S.t132 3.904
R1726 S.n8848 S.t379 3.904
R1727 S.n8838 S.n8837 3.904
R1728 S.n7934 S.n7933 3.904
R1729 S.n7939 S.t1731 3.904
R1730 S.n7942 S.t1265 3.904
R1731 S.n7931 S.n7930 3.904
R1732 S.n8129 S.n8128 3.904
R1733 S.n8133 S.t94 3.904
R1734 S.n8136 S.t347 3.904
R1735 S.n8126 S.n8125 3.904
R1736 S.n7381 S.n7380 3.904
R1737 S.n7386 S.t1699 3.904
R1738 S.n7389 S.t1232 3.904
R1739 S.n7378 S.n7377 3.904
R1740 S.n7118 S.n7117 3.904
R1741 S.n7122 S.t38 3.904
R1742 S.n7125 S.t322 3.904
R1743 S.n7115 S.n7114 3.904
R1744 S.n6635 S.n6634 3.904
R1745 S.n6640 S.t1669 3.904
R1746 S.n6643 S.t1667 3.904
R1747 S.n6632 S.n6631 3.904
R1748 S.n6371 S.n6370 3.904
R1749 S.n6375 S.t561 3.904
R1750 S.n6378 S.t2579 3.904
R1751 S.n6368 S.n6367 3.904
R1752 S.n5880 S.n5879 3.904
R1753 S.n5885 S.t1428 3.904
R1754 S.n5888 S.t1630 3.904
R1755 S.n5877 S.n5876 3.904
R1756 S.n5611 S.n5610 3.904
R1757 S.n5615 S.t528 3.904
R1758 S.n5618 S.t2546 3.904
R1759 S.n5608 S.n5607 3.904
R1760 S.n5099 S.n5098 3.904
R1761 S.n5104 S.t1401 3.904
R1762 S.n5107 S.t1605 3.904
R1763 S.n5096 S.n5095 3.904
R1764 S.n4829 S.n4828 3.904
R1765 S.n4833 S.t497 3.904
R1766 S.n4836 S.t2511 3.904
R1767 S.n4826 S.n4825 3.904
R1768 S.n4309 S.n4308 3.904
R1769 S.n4314 S.t1372 3.904
R1770 S.n4317 S.t1583 3.904
R1771 S.n4306 S.n4305 3.904
R1772 S.n4034 S.n4033 3.904
R1773 S.n4038 S.t470 3.904
R1774 S.n4041 S.t2480 3.904
R1775 S.n4031 S.n4030 3.904
R1776 S.n3462 S.n3461 3.904
R1777 S.n3466 S.t1350 3.904
R1778 S.n3469 S.t1556 3.904
R1779 S.n3459 S.n3458 3.904
R1780 S.n3527 S.t2000 3.904
R1781 S.n3524 S.t877 3.904
R1782 S.n3474 S.n3473 3.904
R1783 S.n3486 S.t1461 3.904
R1784 S.n3489 S.t1675 3.904
R1785 S.n3477 S.n3476 3.904
R1786 S.n4049 S.n4048 3.904
R1787 S.n4351 S.t2119 3.904
R1788 S.n4354 S.t2073 3.904
R1789 S.n4046 S.n4045 3.904
R1790 S.n12494 S.t1473 3.904
R1791 S.n12492 S.t1904 3.904
R1792 S.n12693 S.n12692 3.904
R1793 S.n12698 S.t961 3.904
R1794 S.n12701 S.t539 3.904
R1795 S.n12690 S.n12689 3.904
R1796 S.n12965 S.n12964 3.904
R1797 S.n12969 S.t1919 3.904
R1798 S.n12972 S.t1159 3.904
R1799 S.n12962 S.n12961 3.904
R1800 S.n12071 S.n12070 3.904
R1801 S.n12076 S.t1479 3.904
R1802 S.n12079 S.t115 3.904
R1803 S.n12068 S.n12067 3.904
R1804 S.n11781 S.n11780 3.904
R1805 S.n11785 S.t1505 3.904
R1806 S.n11788 S.t590 3.904
R1807 S.n11778 S.n11777 3.904
R1808 S.n11463 S.n11462 3.904
R1809 S.n11468 S.t894 3.904
R1810 S.n11471 S.t2056 3.904
R1811 S.n11460 S.n11459 3.904
R1812 S.n11218 S.n11217 3.904
R1813 S.n11222 S.t943 3.904
R1814 S.n11225 S.t2491 3.904
R1815 S.n11215 S.n11214 3.904
R1816 S.n10842 S.n10841 3.904
R1817 S.n10847 S.t304 3.904
R1818 S.n10850 S.t1484 3.904
R1819 S.n10839 S.n10838 3.904
R1820 S.n10595 S.n10594 3.904
R1821 S.n10599 S.t486 3.904
R1822 S.n10602 S.t1937 3.904
R1823 S.n10592 S.n10591 3.904
R1824 S.n10189 S.n10188 3.904
R1825 S.n10194 S.t2262 3.904
R1826 S.n10197 S.t1342 3.904
R1827 S.n10186 S.n10185 3.904
R1828 S.n9937 S.n9936 3.904
R1829 S.n9941 S.t1862 3.904
R1830 S.n9944 S.t2085 3.904
R1831 S.n9934 S.n9933 3.904
R1832 S.n9513 S.n9512 3.904
R1833 S.n9518 S.t924 3.904
R1834 S.n9521 S.t446 3.904
R1835 S.n9510 S.n9509 3.904
R1836 S.n9260 S.n9259 3.904
R1837 S.n9264 S.t1829 3.904
R1838 S.n9267 S.t2055 3.904
R1839 S.n9257 S.n9256 3.904
R1840 S.n8646 S.n8645 3.904
R1841 S.n8651 S.t890 3.904
R1842 S.n8654 S.t411 3.904
R1843 S.n8643 S.n8642 3.904
R1844 S.n8856 S.n8855 3.904
R1845 S.n8860 S.t1801 3.904
R1846 S.n8863 S.t2031 3.904
R1847 S.n8853 S.n8852 3.904
R1848 S.n7950 S.n7949 3.904
R1849 S.n7955 S.t857 3.904
R1850 S.n7958 S.t382 3.904
R1851 S.n7947 S.n7946 3.904
R1852 S.n8144 S.n8143 3.904
R1853 S.n8148 S.t1771 3.904
R1854 S.n8151 S.t2005 3.904
R1855 S.n8141 S.n8140 3.904
R1856 S.n7397 S.n7396 3.904
R1857 S.n7402 S.t825 3.904
R1858 S.n7405 S.t349 3.904
R1859 S.n7394 S.n7393 3.904
R1860 S.n7133 S.n7132 3.904
R1861 S.n7137 S.t1735 3.904
R1862 S.n7140 S.t2121 3.904
R1863 S.n7130 S.n7129 3.904
R1864 S.n6651 S.n6650 3.904
R1865 S.n6656 S.t957 3.904
R1866 S.n6659 S.t793 3.904
R1867 S.n6648 S.n6647 3.904
R1868 S.n6386 S.n6385 3.904
R1869 S.n6390 S.t2200 3.904
R1870 S.n6393 S.t1702 3.904
R1871 S.n6383 S.n6382 3.904
R1872 S.n5896 S.n5895 3.904
R1873 S.n5901 S.t563 3.904
R1874 S.n5904 S.t764 3.904
R1875 S.n5893 S.n5892 3.904
R1876 S.n5626 S.n5625 3.904
R1877 S.n5630 S.t2170 3.904
R1878 S.n5633 S.t1673 3.904
R1879 S.n5623 S.n5622 3.904
R1880 S.n5115 S.n5114 3.904
R1881 S.n5120 S.t531 3.904
R1882 S.n5123 S.t741 3.904
R1883 S.n5112 S.n5111 3.904
R1884 S.n4844 S.n4843 3.904
R1885 S.n4848 S.t2145 3.904
R1886 S.n4851 S.t1634 3.904
R1887 S.n4841 S.n4840 3.904
R1888 S.n4346 S.n4345 3.904
R1889 S.n4343 S.t502 3.904
R1890 S.n4340 S.t716 3.904
R1891 S.n4054 S.n4053 3.904
R1892 S.n4359 S.t643 3.904
R1893 S.n4356 S.t2556 3.904
R1894 S.n4322 S.n4321 3.904
R1895 S.n4334 S.t52 3.904
R1896 S.n4337 S.t287 3.904
R1897 S.n4325 S.n4324 3.904
R1898 S.n4859 S.n4858 3.904
R1899 S.n5157 S.t1281 3.904
R1900 S.n5160 S.t694 3.904
R1901 S.n4856 S.n4855 3.904
R1902 S.n12498 S.t613 3.904
R1903 S.n12496 S.t1045 3.904
R1904 S.n12709 S.n12708 3.904
R1905 S.n12714 S.t15 3.904
R1906 S.n12717 S.t2181 3.904
R1907 S.n12706 S.n12705 3.904
R1908 S.n12980 S.n12979 3.904
R1909 S.n12984 S.t1058 3.904
R1910 S.n12987 S.t286 3.904
R1911 S.n12977 S.n12976 3.904
R1912 S.n12087 S.n12086 3.904
R1913 S.n12092 S.t617 3.904
R1914 S.n12095 S.t1788 3.904
R1915 S.n12084 S.n12083 3.904
R1916 S.n11796 S.n11795 3.904
R1917 S.n11800 S.t644 3.904
R1918 S.n11803 S.t2240 3.904
R1919 S.n11793 S.n11792 3.904
R1920 S.n11479 S.n11478 3.904
R1921 S.n11484 S.t2536 3.904
R1922 S.n11487 S.t1196 3.904
R1923 S.n11476 S.n11475 3.904
R1924 S.n11233 S.n11232 3.904
R1925 S.n11237 S.t194 3.904
R1926 S.n11240 S.t1616 3.904
R1927 S.n11230 S.n11229 3.904
R1928 S.n10858 S.n10857 3.904
R1929 S.n10863 S.t1968 3.904
R1930 S.n10866 S.t494 3.904
R1931 S.n10855 S.n10854 3.904
R1932 S.n10610 S.n10609 3.904
R1933 S.n10614 S.t1873 3.904
R1934 S.n10617 S.t1257 3.904
R1935 S.n10607 S.n10606 3.904
R1936 S.n10205 S.n10204 3.904
R1937 S.n10210 S.t17 3.904
R1938 S.n10213 S.t464 3.904
R1939 S.n10202 S.n10201 3.904
R1940 S.n9952 S.n9951 3.904
R1941 S.n9956 S.t993 3.904
R1942 S.n9959 S.t1225 3.904
R1943 S.n9949 S.n9948 3.904
R1944 S.n9529 S.n9528 3.904
R1945 S.n9534 S.t2564 3.904
R1946 S.n9537 S.t2089 3.904
R1947 S.n9526 S.n9525 3.904
R1948 S.n9275 S.n9274 3.904
R1949 S.n9279 S.t963 3.904
R1950 S.n9282 S.t1198 3.904
R1951 S.n9272 S.n9271 3.904
R1952 S.n8662 S.n8661 3.904
R1953 S.n8667 S.t2533 3.904
R1954 S.n8670 S.t2059 3.904
R1955 S.n8659 S.n8658 3.904
R1956 S.n8871 S.n8870 3.904
R1957 S.n8875 S.t934 3.904
R1958 S.n8878 S.t1176 3.904
R1959 S.n8868 S.n8867 3.904
R1960 S.n7966 S.n7965 3.904
R1961 S.n7971 S.t2501 3.904
R1962 S.n7974 S.t2033 3.904
R1963 S.n7963 S.n7962 3.904
R1964 S.n8159 S.n8158 3.904
R1965 S.n8163 S.t897 3.904
R1966 S.n8166 S.t1286 3.904
R1967 S.n8156 S.n8155 3.904
R1968 S.n7413 S.n7412 3.904
R1969 S.n7418 S.t76 3.904
R1970 S.n7421 S.t2006 3.904
R1971 S.n7410 S.n7409 3.904
R1972 S.n7148 S.n7147 3.904
R1973 S.n7152 S.t861 3.904
R1974 S.n7155 S.t1253 3.904
R1975 S.n7145 S.n7144 3.904
R1976 S.n6667 S.n6666 3.904
R1977 S.n6672 S.t9 3.904
R1978 S.n6675 S.t2444 3.904
R1979 S.n6664 S.n6663 3.904
R1980 S.n6401 S.n6400 3.904
R1981 S.n6405 S.t1343 3.904
R1982 S.n6408 S.t829 3.904
R1983 S.n6398 S.n6397 3.904
R1984 S.n5912 S.n5911 3.904
R1985 S.n5917 S.t2202 3.904
R1986 S.n5920 S.t2416 3.904
R1987 S.n5909 S.n5908 3.904
R1988 S.n5641 S.n5640 3.904
R1989 S.n5645 S.t1308 3.904
R1990 S.n5648 S.t798 3.904
R1991 S.n5638 S.n5637 3.904
R1992 S.n5152 S.n5151 3.904
R1993 S.n5149 S.t2174 3.904
R1994 S.n5146 S.t2393 3.904
R1995 S.n4864 S.n4863 3.904
R1996 S.n5165 S.t1809 3.904
R1997 S.n5162 S.t1715 3.904
R1998 S.n5128 S.n5127 3.904
R1999 S.n5140 S.t1250 3.904
R2000 S.n5143 S.t1432 3.904
R2001 S.n5131 S.n5130 3.904
R2002 S.n5656 S.n5655 3.904
R2003 S.n5954 S.t425 3.904
R2004 S.n5957 S.t1885 3.904
R2005 S.n5653 S.n5652 3.904
R2006 S.n12502 S.t2266 3.904
R2007 S.n12500 S.t153 3.904
R2008 S.n12725 S.n12724 3.904
R2009 S.n12730 S.t1724 3.904
R2010 S.n12733 S.t1320 3.904
R2011 S.n12722 S.n12721 3.904
R2012 S.n12995 S.n12994 3.904
R2013 S.n12999 S.t171 3.904
R2014 S.n13002 S.t1947 3.904
R2015 S.n12992 S.n12991 3.904
R2016 S.n12103 S.n12102 3.904
R2017 S.n12108 S.t2273 3.904
R2018 S.n12111 S.t917 3.904
R2019 S.n12100 S.n12099 3.904
R2020 S.n11811 S.n11810 3.904
R2021 S.n11815 S.t2397 3.904
R2022 S.n11818 S.t1380 3.904
R2023 S.n11808 S.n11807 3.904
R2024 S.n11495 S.n11494 3.904
R2025 S.n11500 S.t1663 3.904
R2026 S.n11503 S.t2166 3.904
R2027 S.n11492 S.n11491 3.904
R2028 S.n11248 S.n11247 3.904
R2029 S.n11252 S.t1036 3.904
R2030 S.n11255 S.t403 3.904
R2031 S.n11245 S.n11244 3.904
R2032 S.n10874 S.n10873 3.904
R2033 S.n10879 S.t1761 3.904
R2034 S.n10882 S.t2140 3.904
R2035 S.n10871 S.n10870 3.904
R2036 S.n10625 S.n10624 3.904
R2037 S.n10629 S.t1008 3.904
R2038 S.n10632 S.t375 3.904
R2039 S.n10622 S.n10621 3.904
R2040 S.n10221 S.n10220 3.904
R2041 S.n10226 S.t1725 3.904
R2042 S.n10229 S.t2109 3.904
R2043 S.n10218 S.n10217 3.904
R2044 S.n9967 S.n9966 3.904
R2045 S.n9971 S.t87 3.904
R2046 S.n9974 S.t342 3.904
R2047 S.n9964 S.n9963 3.904
R2048 S.n9545 S.n9544 3.904
R2049 S.n9550 S.t1690 3.904
R2050 S.n9553 S.t1227 3.904
R2051 S.n9542 S.n9541 3.904
R2052 S.n9290 S.n9289 3.904
R2053 S.n9294 S.t25 3.904
R2054 S.n9297 S.t318 3.904
R2055 S.n9287 S.n9286 3.904
R2056 S.n8678 S.n8677 3.904
R2057 S.n8683 S.t1660 3.904
R2058 S.n8686 S.t1199 3.904
R2059 S.n8675 S.n8674 3.904
R2060 S.n8886 S.n8885 3.904
R2061 S.n8890 S.t2574 3.904
R2062 S.n8893 S.t432 3.904
R2063 S.n8883 S.n8882 3.904
R2064 S.n7982 S.n7981 3.904
R2065 S.n7987 S.t1785 3.904
R2066 S.n7990 S.t1177 3.904
R2067 S.n7979 S.n7978 3.904
R2068 S.n8174 S.n8173 3.904
R2069 S.n8178 S.t2539 3.904
R2070 S.n8181 S.t398 3.904
R2071 S.n8171 S.n8170 3.904
R2072 S.n7429 S.n7428 3.904
R2073 S.n7434 S.t1757 3.904
R2074 S.n7437 S.t1156 3.904
R2075 S.n7426 S.n7425 3.904
R2076 S.n7163 S.n7162 3.904
R2077 S.n7167 S.t2506 3.904
R2078 S.n7170 S.t371 3.904
R2079 S.n7160 S.n7159 3.904
R2080 S.n6683 S.n6682 3.904
R2081 S.n6688 S.t1721 3.904
R2082 S.n6691 S.t1577 3.904
R2083 S.n6680 S.n6679 3.904
R2084 S.n6416 S.n6415 3.904
R2085 S.n6420 S.t466 3.904
R2086 S.n6423 S.t2476 3.904
R2087 S.n6413 S.n6412 3.904
R2088 S.n5949 S.n5948 3.904
R2089 S.n5946 S.t1345 3.904
R2090 S.n5943 S.t1552 3.904
R2091 S.n5661 S.n5660 3.904
R2092 S.n5962 S.t429 3.904
R2093 S.n5959 S.t872 3.904
R2094 S.n5925 S.n5924 3.904
R2095 S.n5937 S.t2376 3.904
R2096 S.n5940 S.t2515 3.904
R2097 S.n5928 S.n5927 3.904
R2098 S.n6431 S.n6430 3.904
R2099 S.n6725 S.t2112 3.904
R2100 S.n6728 S.t518 3.904
R2101 S.n6428 S.n6427 3.904
R2102 S.n12506 S.t1407 3.904
R2103 S.n12504 S.t1817 3.904
R2104 S.n12741 S.n12740 3.904
R2105 S.n12746 S.t852 3.904
R2106 S.n12749 S.t439 3.904
R2107 S.n12738 S.n12737 3.904
R2108 S.n13010 S.n13009 3.904
R2109 S.n13014 S.t1951 3.904
R2110 S.n13017 S.t1089 3.904
R2111 S.n13007 S.n13006 3.904
R2112 S.n12119 S.n12118 3.904
R2113 S.n12124 S.t1417 3.904
R2114 S.n12127 S.t1336 3.904
R2115 S.n12116 S.n12115 3.904
R2116 S.n11826 S.n11825 3.904
R2117 S.n11830 S.t177 3.904
R2118 S.n11833 S.t2083 3.904
R2119 S.n11823 S.n11822 3.904
R2120 S.n11511 S.n11510 3.904
R2121 S.n11516 S.t922 3.904
R2122 S.n11519 S.t1304 3.904
R2123 S.n11508 S.n11507 3.904
R2124 S.n11263 S.n11262 3.904
R2125 S.n11267 S.t144 3.904
R2126 S.n11270 S.t2053 3.904
R2127 S.n11260 S.n11259 3.904
R2128 S.n10890 S.n10889 3.904
R2129 S.n10895 S.t884 3.904
R2130 S.n10898 S.t1274 3.904
R2131 S.n10887 S.n10886 3.904
R2132 S.n10640 S.n10639 3.904
R2133 S.n10644 S.t104 3.904
R2134 S.n10647 S.t2026 3.904
R2135 S.n10637 S.n10636 3.904
R2136 S.n10237 S.n10236 3.904
R2137 S.n10242 S.t853 3.904
R2138 S.n10245 S.t1244 3.904
R2139 S.n10234 S.n10233 3.904
R2140 S.n9982 S.n9981 3.904
R2141 S.n9986 S.t1764 3.904
R2142 S.n9989 S.t2001 3.904
R2143 S.n9979 S.n9978 3.904
R2144 S.n9561 S.n9560 3.904
R2145 S.n9566 S.t816 3.904
R2146 S.n9569 S.t344 3.904
R2147 S.n9558 S.n9557 3.904
R2148 S.n9305 S.n9304 3.904
R2149 S.n9309 S.t1729 3.904
R2150 S.n9312 S.t2115 3.904
R2151 S.n9302 S.n9301 3.904
R2152 S.n8694 S.n8693 3.904
R2153 S.n8699 S.t952 3.904
R2154 S.n8702 S.t319 3.904
R2155 S.n8691 S.n8690 3.904
R2156 S.n8901 S.n8900 3.904
R2157 S.n8905 S.t1698 3.904
R2158 S.n8908 S.t2079 3.904
R2159 S.n8898 S.n8897 3.904
R2160 S.n7998 S.n7997 3.904
R2161 S.n8003 S.t916 3.904
R2162 S.n8006 S.t300 3.904
R2163 S.n7995 S.n7994 3.904
R2164 S.n8189 S.n8188 3.904
R2165 S.n8193 S.t1668 3.904
R2166 S.n8196 S.t2050 3.904
R2167 S.n8186 S.n8185 3.904
R2168 S.n7445 S.n7444 3.904
R2169 S.n7450 S.t879 3.904
R2170 S.n7453 S.t282 3.904
R2171 S.n7442 S.n7441 3.904
R2172 S.n7178 S.n7177 3.904
R2173 S.n7182 S.t1631 3.904
R2174 S.n7185 S.t2024 3.904
R2175 S.n7175 S.n7174 3.904
R2176 S.n6720 S.n6719 3.904
R2177 S.n6717 S.t849 3.904
R2178 S.n6714 S.t709 3.904
R2179 S.n6436 S.n6435 3.904
R2180 S.n6733 S.t1558 3.904
R2181 S.n6730 S.t2552 3.904
R2182 S.n6696 S.n6695 3.904
R2183 S.n6708 S.t317 3.904
R2184 S.n6711 S.t1141 3.904
R2185 S.n6699 S.n6698 3.904
R2186 S.n7193 S.n7192 3.904
R2187 S.n7487 S.t763 3.904
R2188 S.n7490 S.t971 3.904
R2189 S.n7190 S.n7189 3.904
R2190 S.n12510 S.t540 3.904
R2191 S.n12508 S.t1079 3.904
R2192 S.n12757 S.n12756 3.904
R2193 S.n12762 S.t2492 3.904
R2194 S.n12765 S.t2064 3.904
R2195 S.n12754 S.n12753 3.904
R2196 S.n13025 S.n13024 3.904
R2197 S.n13029 S.t939 3.904
R2198 S.n13032 S.t1251 3.904
R2199 S.n13022 S.n13021 3.904
R2200 S.n12135 S.n12134 3.904
R2201 S.n12140 S.t3 3.904
R2202 S.n12143 S.t455 3.904
R2203 S.n12132 S.n12131 3.904
R2204 S.n11841 S.n11840 3.904
R2205 S.n11845 S.t1842 3.904
R2206 S.n11848 S.t1221 3.904
R2207 S.n11838 S.n11837 3.904
R2208 S.n11527 S.n11526 3.904
R2209 S.n11532 S.t2559 3.904
R2210 S.n11535 S.t420 3.904
R2211 S.n11524 S.n11523 3.904
R2212 S.n11278 S.n11277 3.904
R2213 S.n11282 S.t1812 3.904
R2214 S.n11285 S.t1193 3.904
R2215 S.n11275 S.n11274 3.904
R2216 S.n10906 S.n10905 3.904
R2217 S.n10911 S.t2528 3.904
R2218 S.n10914 S.t392 3.904
R2219 S.n10903 S.n10902 3.904
R2220 S.n10655 S.n10654 3.904
R2221 S.n10659 S.t1779 3.904
R2222 S.n10662 S.t1169 3.904
R2223 S.n10652 S.n10651 3.904
R2224 S.n10253 S.n10252 3.904
R2225 S.n10258 S.t2495 3.904
R2226 S.n10261 S.t362 3.904
R2227 S.n10250 S.n10249 3.904
R2228 S.n9997 S.n9996 3.904
R2229 S.n10001 S.t889 3.904
R2230 S.n10004 S.t1278 3.904
R2231 S.n9994 S.n9993 3.904
R2232 S.n9577 S.n9576 3.904
R2233 S.n9582 S.t65 3.904
R2234 S.n9585 S.t2003 3.904
R2235 S.n9574 S.n9573 3.904
R2236 S.n9320 S.n9319 3.904
R2237 S.n9324 S.t856 3.904
R2238 S.n9327 S.t1247 3.904
R2239 S.n9317 S.n9316 3.904
R2240 S.n8710 S.n8709 3.904
R2241 S.n8715 S.t1 3.904
R2242 S.n8718 S.t1982 3.904
R2243 S.n8707 S.n8706 3.904
R2244 S.n8916 S.n8915 3.904
R2245 S.n8920 S.t824 3.904
R2246 S.n8923 S.t1219 3.904
R2247 S.n8913 S.n8912 3.904
R2248 S.n8014 S.n8013 3.904
R2249 S.n8019 S.t2557 3.904
R2250 S.n8022 S.t1964 3.904
R2251 S.n8011 S.n8010 3.904
R2252 S.n8204 S.n8203 3.904
R2253 S.n8208 S.t794 3.904
R2254 S.n8211 S.t1192 3.904
R2255 S.n8201 S.n8200 3.904
R2256 S.n7482 S.n7481 3.904
R2257 S.n7479 S.t2524 3.904
R2258 S.n7476 S.t1941 3.904
R2259 S.n7198 S.n7197 3.904
R2260 S.n7495 S.t150 3.904
R2261 S.n7492 S.t2091 3.904
R2262 S.n7458 S.n7457 3.904
R2263 S.n7470 S.t1486 3.904
R2264 S.n7473 S.t2445 3.904
R2265 S.n7461 S.n7460 3.904
R2266 S.n8219 S.n8218 3.904
R2267 S.n8223 S.t2442 3.904
R2268 S.n8226 S.t2111 3.904
R2269 S.n8216 S.n8215 3.904
R2270 S.n12514 S.t1943 3.904
R2271 S.n12512 S.t1649 3.904
R2272 S.n12773 S.n12772 3.904
R2273 S.n12778 S.t1655 3.904
R2274 S.n12781 S.t1201 3.904
R2275 S.n12770 S.n12769 3.904
R2276 S.n13040 S.n13039 3.904
R2277 S.n13044 S.t2578 3.904
R2278 S.n13047 S.t369 3.904
R2279 S.n13037 S.n13036 3.904
R2280 S.n12151 S.n12150 3.904
R2281 S.n12156 S.t1718 3.904
R2282 S.n12159 S.t2100 3.904
R2283 S.n12148 S.n12147 3.904
R2284 S.n11856 S.n11855 3.904
R2285 S.n11860 S.t977 3.904
R2286 S.n11863 S.t340 3.904
R2287 S.n11853 S.n11852 3.904
R2288 S.n11543 S.n11542 3.904
R2289 S.n11548 S.t1686 3.904
R2290 S.n11551 S.t2071 3.904
R2291 S.n11540 S.n11539 3.904
R2292 S.n11293 S.n11292 3.904
R2293 S.n11297 S.t945 3.904
R2294 S.n11300 S.t314 3.904
R2295 S.n11290 S.n11289 3.904
R2296 S.n10922 S.n10921 3.904
R2297 S.n10927 S.t1652 3.904
R2298 S.n10930 S.t2041 3.904
R2299 S.n10919 S.n10918 3.904
R2300 S.n10670 S.n10669 3.904
R2301 S.n10674 S.t907 3.904
R2302 S.n10677 S.t422 3.904
R2303 S.n10667 S.n10666 3.904
R2304 S.n10269 S.n10268 3.904
R2305 S.n10274 S.t1782 3.904
R2306 S.n10277 S.t2014 3.904
R2307 S.n10266 S.n10265 3.904
R2308 S.n10012 S.n10011 3.904
R2309 S.n10016 S.t2531 3.904
R2310 S.n10019 S.t394 3.904
R2311 S.n10009 S.n10008 3.904
R2312 S.n9593 S.n9592 3.904
R2313 S.n9598 S.t1751 3.904
R2314 S.n9601 S.t1151 3.904
R2315 S.n9590 S.n9589 3.904
R2316 S.n9335 S.n9334 3.904
R2317 S.n9339 S.t2500 3.904
R2318 S.n9342 S.t366 3.904
R2319 S.n9332 S.n9331 3.904
R2320 S.n8726 S.n8725 3.904
R2321 S.n8731 S.t1716 3.904
R2322 S.n8734 S.t1134 3.904
R2323 S.n8723 S.n8722 3.904
R2324 S.n8931 S.n8930 3.904
R2325 S.n8935 S.t2469 3.904
R2326 S.n8938 S.t337 3.904
R2327 S.n8928 S.n8927 3.904
R2328 S.n8030 S.n8029 3.904
R2329 S.n8034 S.t1684 3.904
R2330 S.n8037 S.t1109 3.904
R2331 S.n8027 S.n8026 3.904
R2332 S.n8231 S.t1319 3.904
R2333 S.n8228 S.t1262 3.904
R2334 S.n8042 S.n8041 3.904
R2335 S.n8054 S.t100 3.904
R2336 S.n8057 S.t1085 3.904
R2337 S.n8045 S.n8044 3.904
R2338 S.n8946 S.n8945 3.904
R2339 S.n8950 S.t1599 3.904
R2340 S.n8953 S.t718 3.904
R2341 S.n8943 S.n8942 3.904
R2342 S.n12518 S.t1086 3.904
R2343 S.n12516 S.t778 3.904
R2344 S.n12789 S.n12788 3.904
R2345 S.n12794 S.t785 3.904
R2346 S.n12797 S.t324 3.904
R2347 S.n12786 S.n12785 3.904
R2348 S.n13055 S.n13054 3.904
R2349 S.n13059 S.t1701 3.904
R2350 S.n13062 S.t2022 3.904
R2351 S.n13052 S.n13051 3.904
R2352 S.n12167 S.n12166 3.904
R2353 S.n12172 S.t847 3.904
R2354 S.n12175 S.t1235 3.904
R2355 S.n12164 S.n12163 3.904
R2356 S.n11871 S.n11870 3.904
R2357 S.n11875 S.t45 3.904
R2358 S.n11878 S.t1998 3.904
R2359 S.n11868 S.n11867 3.904
R2360 S.n11559 S.n11558 3.904
R2361 S.n11564 S.t813 3.904
R2362 S.n11567 S.t1210 3.904
R2363 S.n11556 S.n11555 3.904
R2364 S.n11308 S.n11307 3.904
R2365 S.n11312 S.t2582 3.904
R2366 S.n11315 S.t2110 3.904
R2367 S.n11305 S.n11304 3.904
R2368 S.n10938 S.n10937 3.904
R2369 S.n10943 S.t950 3.904
R2370 S.n10946 S.t1184 3.904
R2371 S.n10935 S.n10934 3.904
R2372 S.n10685 S.n10684 3.904
R2373 S.n10689 S.t2549 3.904
R2374 S.n10692 S.t2076 3.904
R2375 S.n10682 S.n10681 3.904
R2376 S.n10285 S.n10284 3.904
R2377 S.n10290 S.t910 3.904
R2378 S.n10293 S.t1161 3.904
R2379 S.n10282 S.n10281 3.904
R2380 S.n10027 S.n10026 3.904
R2381 S.n10031 S.t1658 3.904
R2382 S.n10034 S.t2044 3.904
R2383 S.n10024 S.n10023 3.904
R2384 S.n9609 S.n9608 3.904
R2385 S.n9614 S.t873 3.904
R2386 S.n9617 S.t275 3.904
R2387 S.n9606 S.n9605 3.904
R2388 S.n9350 S.n9349 3.904
R2389 S.n9354 S.t1625 3.904
R2390 S.n9357 S.t2018 3.904
R2391 S.n9347 S.n9346 3.904
R2392 S.n8742 S.n8741 3.904
R2393 S.n8746 S.t845 3.904
R2394 S.n8749 S.t255 3.904
R2395 S.n8739 S.n8738 3.904
R2396 S.n8958 S.t2430 3.904
R2397 S.n8955 S.t407 3.904
R2398 S.n8754 S.n8753 3.904
R2399 S.n8766 S.t1282 3.904
R2400 S.n8769 S.t2203 3.904
R2401 S.n8757 S.n8756 3.904
R2402 S.n9365 S.n9364 3.904
R2403 S.n9651 S.t759 3.904
R2404 S.n9654 S.t1912 3.904
R2405 S.n9362 S.n9361 3.904
R2406 S.n12522 S.t207 3.904
R2407 S.n12520 S.t2431 3.904
R2408 S.n12805 S.n12804 3.904
R2409 S.n12810 S.t2435 3.904
R2410 S.n12813 S.t1983 3.904
R2411 S.n12802 S.n12801 3.904
R2412 S.n13070 S.n13069 3.904
R2413 S.n13074 S.t828 3.904
R2414 S.n13077 S.t1166 3.904
R2415 S.n13067 S.n13066 3.904
R2416 S.n12183 S.n12182 3.904
R2417 S.n12188 S.t2490 3.904
R2418 S.n12191 S.t355 3.904
R2419 S.n12180 S.n12179 3.904
R2420 S.n11886 S.n11885 3.904
R2421 S.n11890 S.t1738 3.904
R2422 S.n11893 S.t1275 3.904
R2423 S.n11883 S.n11882 3.904
R2424 S.n11575 S.n11574 3.904
R2425 S.n11580 S.t50 3.904
R2426 S.n11583 S.t331 3.904
R2427 S.n11572 S.n11571 3.904
R2428 S.n11323 S.n11322 3.904
R2429 S.n11327 S.t1704 3.904
R2430 S.n11330 S.t1241 3.904
R2431 S.n11320 S.n11319 3.904
R2432 S.n10954 S.n10953 3.904
R2433 S.n10959 S.t2587 3.904
R2434 S.n10962 S.t309 3.904
R2435 S.n10951 S.n10950 3.904
R2436 S.n10700 S.n10699 3.904
R2437 S.n10704 S.t1679 3.904
R2438 S.n10707 S.t1213 3.904
R2439 S.n10697 S.n10696 3.904
R2440 S.n10301 S.n10300 3.904
R2441 S.n10306 S.t2551 3.904
R2442 S.n10309 S.t289 3.904
R2443 S.n10298 S.n10297 3.904
R2444 S.n10042 S.n10041 3.904
R2445 S.n10046 S.t789 3.904
R2446 S.n10049 S.t1188 3.904
R2447 S.n10039 S.n10038 3.904
R2448 S.n9646 S.n9645 3.904
R2449 S.n9643 S.t2518 3.904
R2450 S.n9640 S.t1938 3.904
R2451 S.n9370 S.n9369 3.904
R2452 S.n9659 S.t1103 3.904
R2453 S.n9656 S.t2084 3.904
R2454 S.n9622 S.n9621 3.904
R2455 S.n9634 S.t2400 3.904
R2456 S.n9637 S.t766 3.904
R2457 S.n9625 S.n9624 3.904
R2458 S.n10057 S.n10056 3.904
R2459 S.n10343 S.t2439 3.904
R2460 S.n10346 S.t553 3.904
R2461 S.n10054 S.n10053 3.904
R2462 S.n12526 S.t1875 3.904
R2463 S.n12524 S.t1567 3.904
R2464 S.n12821 S.n12820 3.904
R2465 S.n12826 S.t1571 3.904
R2466 S.n12829 S.t1135 3.904
R2467 S.n12818 S.n12817 3.904
R2468 S.n13085 S.n13084 3.904
R2469 S.n13089 S.t2473 3.904
R2470 S.n13092 S.t421 3.904
R2471 S.n13082 S.n13081 3.904
R2472 S.n12199 S.n12198 3.904
R2473 S.n12204 S.t1775 3.904
R2474 S.n12207 S.t2010 3.904
R2475 S.n12196 S.n12195 3.904
R2476 S.n11901 S.n11900 3.904
R2477 S.n11905 S.t863 3.904
R2478 S.n11908 S.t388 3.904
R2479 S.n11898 S.n11897 3.904
R2480 S.n11591 S.n11590 3.904
R2481 S.n11596 S.t1744 3.904
R2482 S.n11599 S.t1988 3.904
R2483 S.n11588 S.n11587 3.904
R2484 S.n11338 S.n11337 3.904
R2485 S.n11342 S.t835 3.904
R2486 S.n11345 S.t359 3.904
R2487 S.n11335 S.n11334 3.904
R2488 S.n10970 S.n10969 3.904
R2489 S.n10975 S.t1710 3.904
R2490 S.n10978 S.t1971 3.904
R2491 S.n10967 S.n10966 3.904
R2492 S.n10715 S.n10714 3.904
R2493 S.n10719 S.t805 3.904
R2494 S.n10722 S.t334 3.904
R2495 S.n10712 S.n10711 3.904
R2496 S.n10338 S.n10337 3.904
R2497 S.n10335 S.t1681 3.904
R2498 S.n10332 S.t1950 3.904
R2499 S.n10062 S.n10061 3.904
R2500 S.n10351 S.t2255 3.904
R2501 S.n10348 S.t1254 3.904
R2502 S.n10314 S.n10313 3.904
R2503 S.n10326 S.t1076 3.904
R2504 S.n10329 S.t2560 3.904
R2505 S.n10317 S.n10316 3.904
R2506 S.n10730 S.n10729 3.904
R2507 S.n11012 S.t2454 3.904
R2508 S.n11015 S.t1665 3.904
R2509 S.n10727 S.n10726 3.904
R2510 S.n12530 S.t1129 3.904
R2511 S.n12528 S.t699 3.904
R2512 S.n12837 S.n12836 3.904
R2513 S.n12842 S.t842 3.904
R2514 S.n12845 S.t256 3.904
R2515 S.n12834 S.n12833 3.904
R2516 S.n13100 S.n13099 3.904
R2517 S.n13104 S.t1604 3.904
R2518 S.n13107 S.t2068 3.904
R2519 S.n13097 S.n13096 3.904
R2520 S.n12215 S.n12214 3.904
R2521 S.n12220 S.t905 3.904
R2522 S.n12223 S.t1158 3.904
R2523 S.n12212 S.n12211 3.904
R2524 S.n11916 S.n11915 3.904
R2525 S.n11920 S.t2510 3.904
R2526 S.n11923 S.t2038 3.904
R2527 S.n11913 S.n11912 3.904
R2528 S.n11607 S.n11606 3.904
R2529 S.n11612 S.t868 3.904
R2530 S.n11615 S.t1138 3.904
R2531 S.n11604 S.n11603 3.904
R2532 S.n11353 S.n11352 3.904
R2533 S.n11357 S.t2481 3.904
R2534 S.n11360 S.t2013 3.904
R2535 S.n11350 S.n11349 3.904
R2536 S.n11007 S.n11006 3.904
R2537 S.n11004 S.t840 3.904
R2538 S.n11001 S.t1116 3.904
R2539 S.n10735 S.n10734 3.904
R2540 S.n11020 S.t248 3.904
R2541 S.n11017 S.t401 3.904
R2542 S.n10983 S.n10982 3.904
R2543 S.n10995 S.t2229 3.904
R2544 S.n10998 S.t1167 3.904
R2545 S.n10986 S.n10985 3.904
R2546 S.n11368 S.n11367 3.904
R2547 S.n11652 S.t1607 3.904
R2548 S.n11655 S.t307 3.904
R2549 S.n11365 S.n11364 3.904
R2550 S.n12534 S.t251 3.904
R2551 S.n12532 S.t2358 3.904
R2552 S.n12853 S.n12852 3.904
R2553 S.n12858 S.t2485 3.904
R2554 S.n12861 S.t1922 3.904
R2555 S.n12850 S.n12849 3.904
R2556 S.n13115 S.n13114 3.904
R2557 S.n13119 S.t740 3.904
R2558 S.n13122 S.t1207 3.904
R2559 S.n13112 S.n13111 3.904
R2560 S.n12231 S.n12230 3.904
R2561 S.n12236 S.t2548 3.904
R2562 S.n12239 S.t284 3.904
R2563 S.n12228 S.n12227 3.904
R2564 S.n11931 S.n11930 3.904
R2565 S.n11935 S.t1635 3.904
R2566 S.n11938 S.t1183 3.904
R2567 S.n11928 S.n11927 3.904
R2568 S.n11647 S.n11646 3.904
R2569 S.n11644 S.t2513 3.904
R2570 S.n11641 S.t262 3.904
R2571 S.n11373 S.n11372 3.904
R2572 S.n11660 S.t1422 3.904
R2573 S.n11657 S.t2081 3.904
R2574 S.n11618 S.n11617 3.904
R2575 S.n11635 S.t832 3.904
R2576 S.n11638 S.t2294 3.904
R2577 S.n11621 S.n11620 3.904
R2578 S.n12258 S.n12257 3.904
R2579 S.n12267 S.t767 3.904
R2580 S.n12270 S.t1474 3.904
R2581 S.n12261 S.n12260 3.904
R2582 S.n12538 S.t1917 3.904
R2583 S.n12536 S.t1503 3.904
R2584 S.n12866 S.n12865 3.904
R2585 S.n12874 S.t1611 3.904
R2586 S.n12877 S.t1062 3.904
R2587 S.n12869 S.n12868 3.904
R2588 S.n13129 S.n13128 3.904
R2589 S.n13137 S.t2390 3.904
R2590 S.n13140 S.t329 3.904
R2591 S.n13132 S.n13131 3.904
R2592 S.n11947 S.n11946 3.904
R2593 S.n12242 S.t1676 3.904
R2594 S.n12245 S.t1946 3.904
R2595 S.n12248 S.n12247 3.904
R2596 S.n12478 S.t499 3.904
R2597 S.n12476 S.t2300 3.904
R2598 S.n12657 S.n12656 3.904
R2599 S.n12668 S.t589 3.904
R2600 S.n12665 S.t1115 3.904
R2601 S.n12660 S.n12659 3.904
R2602 S.n13143 S.t2023 3.904
R2603 S.n13145 S.t395 3.904
R2604 S.n1021 S.n1020 3.904
R2605 S.n1023 S.t2590 3.904
R2606 S.n1794 S.n1793 3.643
R2607 S.n1796 S.t2151 3.643
R2608 S.n12543 S.t593 3.643
R2609 S.n12634 S.t2467 3.643
R2610 S.n12645 S.n12644 3.643
R2611 S.n12642 S.n12641 3.643
R2612 S.n12637 S.t822 3.643
R2613 S.n12558 S.t264 3.643
R2614 S.n12569 S.n12568 3.643
R2615 S.n12566 S.n12565 3.643
R2616 S.n12561 S.t1526 3.643
R2617 S.n11996 S.t1259 3.643
R2618 S.n12014 S.n12013 3.643
R2619 S.n12011 S.n12010 3.643
R2620 S.n11999 S.t2410 3.643
R2621 S.n12277 S.t2207 3.643
R2622 S.n476 S.t1521 3.643
R2623 S.n457 S.t1828 3.643
R2624 S.n840 S.t2427 3.643
R2625 S.n853 S.n852 3.643
R2626 S.n856 S.n855 3.643
R2627 S.n843 S.t475 3.643
R2628 S.n951 S.t1233 3.643
R2629 S.n952 S.t965 3.643
R2630 S.n948 S.t1277 3.643
R2631 S.n944 S.t1142 3.643
R2632 S.n817 S.t2422 3.643
R2633 S.n828 S.n827 3.643
R2634 S.n825 S.n824 3.643
R2635 S.n820 S.t1202 3.643
R2636 S.n1776 S.t2052 3.643
R2637 S.n1790 S.n1789 3.643
R2638 S.n1787 S.n1786 3.643
R2639 S.n1773 S.t34 3.643
R2640 S.n12621 S.t1108 3.643
R2641 S.n12602 S.t2236 3.643
R2642 S.n12578 S.t130 3.643
R2643 S.n12593 S.n12592 3.643
R2644 S.n12596 S.n12595 3.643
R2645 S.n12575 S.t664 3.643
R2646 S.n11979 S.t1601 3.643
R2647 S.n11990 S.n11989 3.643
R2648 S.n11987 S.n11986 3.643
R2649 S.n11976 S.t1924 3.643
R2650 S.n11682 S.t2278 3.643
R2651 S.n11697 S.n11696 3.643
R2652 S.n11694 S.n11693 3.643
R2653 S.n11679 S.t276 3.643
R2654 S.n11427 S.t1066 3.643
R2655 S.n11438 S.n11437 3.643
R2656 S.n11435 S.n11434 3.643
R2657 S.n11424 S.t1349 3.643
R2658 S.n11085 S.t1824 3.643
R2659 S.n11100 S.n11099 3.643
R2660 S.n11097 S.n11096 3.643
R2661 S.n11082 S.t2337 3.643
R2662 S.n10806 S.t472 3.643
R2663 S.n10817 S.n10816 3.643
R2664 S.n10814 S.n10813 3.643
R2665 S.n10803 S.t724 3.643
R2666 S.n10460 S.t1230 3.643
R2667 S.n10475 S.n10474 3.643
R2668 S.n10472 S.n10471 3.643
R2669 S.n10457 S.t1767 3.643
R2670 S.n10153 S.t2380 3.643
R2671 S.n10164 S.n10163 3.643
R2672 S.n10161 S.n10160 3.643
R2673 S.n10150 S.t170 3.643
R2674 S.n9800 S.t949 3.643
R2675 S.n9815 S.n9814 3.643
R2676 S.n9812 S.n9811 3.643
R2677 S.n9797 S.t1180 3.643
R2678 S.n9477 S.t1837 3.643
R2679 S.n9488 S.n9487 3.643
R2680 S.n9485 S.n9484 3.643
R2681 S.n9474 S.t2104 3.643
R2682 S.n9128 S.t338 3.643
R2683 S.n9143 S.n9142 3.643
R2684 S.n9140 S.n9139 3.643
R2685 S.n9125 S.t875 3.643
R2686 S.n8610 S.t1242 3.643
R2687 S.n8621 S.n8620 3.643
R2688 S.n8618 S.n8617 3.643
R2689 S.n8607 S.t1512 3.643
R2690 S.n8433 S.t2292 3.643
R2691 S.n8448 S.n8447 3.643
R2692 S.n8445 S.n8444 3.643
R2693 S.n8430 S.t293 3.643
R2694 S.n7914 S.t756 3.643
R2695 S.n7925 S.n7924 3.643
R2696 S.n7922 S.n7921 3.643
R2697 S.n7911 S.t954 3.643
R2698 S.n7726 S.t1696 3.643
R2699 S.n7741 S.n7740 3.643
R2700 S.n7738 S.n7737 3.643
R2701 S.n7723 S.t2251 3.643
R2702 S.n7361 S.t1133 3.643
R2703 S.n7372 S.n7371 3.643
R2704 S.n7369 S.n7368 3.643
R2705 S.n7358 S.t365 3.643
R2706 S.n6996 S.t2468 3.643
R2707 S.n7011 S.n7010 3.643
R2708 S.n7008 S.n7007 3.643
R2709 S.n6993 S.t533 3.643
R2710 S.n6615 S.t1104 3.643
R2711 S.n6626 S.n6625 3.643
R2712 S.n6623 S.n6622 3.643
R2713 S.n6612 S.t336 3.643
R2714 S.n6254 S.t419 3.643
R2715 S.n6269 S.n6268 3.643
R2716 S.n6266 S.n6265 3.643
R2717 S.n6251 S.t988 3.643
R2718 S.n5860 S.t676 3.643
R2719 S.n5871 S.n5870 3.643
R2720 S.n5868 S.n5867 3.643
R2721 S.n5857 S.t2441 3.643
R2722 S.n5489 S.t391 3.643
R2723 S.n5504 S.n5503 3.643
R2724 S.n5501 S.n5500 3.643
R2725 S.n5486 S.t953 3.643
R2726 S.n5079 S.t658 3.643
R2727 S.n5090 S.n5089 3.643
R2728 S.n5087 S.n5086 3.643
R2729 S.n5076 S.t2415 3.643
R2730 S.n4712 S.t361 3.643
R2731 S.n4727 S.n4726 3.643
R2732 S.n4724 S.n4723 3.643
R2733 S.n4709 S.t918 3.643
R2734 S.n4289 S.t636 3.643
R2735 S.n4300 S.n4299 3.643
R2736 S.n4297 S.n4296 3.643
R2737 S.n4286 S.t2389 3.643
R2738 S.n3912 S.t483 3.643
R2739 S.n3927 S.n3926 3.643
R2740 S.n3924 S.n3923 3.643
R2741 S.n3909 S.t1040 3.643
R2742 S.n3442 S.t619 3.643
R2743 S.n3453 S.n3452 3.643
R2744 S.n3450 S.n3449 3.643
R2745 S.n3439 S.t2369 3.643
R2746 S.n3100 S.t453 3.643
R2747 S.n3115 S.n3114 3.643
R2748 S.n3112 S.n3111 3.643
R2749 S.n3097 S.t1010 3.643
R2750 S.n2586 S.t599 3.643
R2751 S.n2597 S.n2596 3.643
R2752 S.n2594 S.n2593 3.643
R2753 S.n2583 S.t2352 3.643
R2754 S.n2263 S.t2082 3.643
R2755 S.n2280 S.n2279 3.643
R2756 S.n2277 S.n2276 3.643
R2757 S.n2260 S.t985 3.643
R2758 S.n1306 S.t581 3.643
R2759 S.n1315 S.n1314 3.643
R2760 S.n1312 S.n1311 3.643
R2761 S.n1303 S.t2333 3.643
R2762 S.n723 S.t559 3.643
R2763 S.n734 S.n733 3.643
R2764 S.n731 S.n730 3.643
R2765 S.n726 S.t2310 3.643
R2766 S.n201 S.t1557 3.643
R2767 S.n194 S.t2322 3.643
R2768 S.n420 S.t1204 3.643
R2769 S.n431 S.n430 3.643
R2770 S.n428 S.n427 3.643
R2771 S.n423 S.t1749 3.643
R2772 S.n1665 S.t1231 3.643
R2773 S.n1678 S.n1677 3.643
R2774 S.n1675 S.n1674 3.643
R2775 S.n1662 S.t1780 3.643
R2776 S.n9391 S.t1132 3.643
R2777 S.n9372 S.t1423 3.643
R2778 S.n9152 S.t2030 3.643
R2779 S.n9166 S.n9165 3.643
R2780 S.n9169 S.n9168 3.643
R2781 S.n9149 S.t2568 3.643
R2782 S.n8514 S.t560 3.643
R2783 S.n8525 S.n8524 3.643
R2784 S.n8522 S.n8521 3.643
R2785 S.n8511 S.t799 3.643
R2786 S.n8286 S.t1467 3.643
R2787 S.n8301 S.n8300 3.643
R2788 S.n8298 S.n8297 3.643
R2789 S.n8283 S.t1985 3.643
R2790 S.n7818 S.t2452 3.643
R2791 S.n7829 S.n7828 3.643
R2792 S.n7826 S.n7825 3.643
R2793 S.n7815 S.t239 3.643
R2794 S.n7579 S.t1029 3.643
R2795 S.n7594 S.n7593 3.643
R2796 S.n7591 S.n7590 3.643
R2797 S.n7576 S.t1525 3.643
R2798 S.n7265 S.t1910 3.643
R2799 S.n7276 S.n7275 3.643
R2800 S.n7273 S.n7272 3.643
R2801 S.n7262 S.t2186 3.643
R2802 S.n6849 S.t418 3.643
R2803 S.n6864 S.n6863 3.643
R2804 S.n6861 S.n6860 3.643
R2805 S.n6846 S.t976 3.643
R2806 S.n6519 S.t1328 3.643
R2807 S.n6530 S.n6529 3.643
R2808 S.n6527 S.n6526 3.643
R2809 S.n6516 S.t1572 3.643
R2810 S.n6107 S.t1886 3.643
R2811 S.n6122 S.n6121 3.643
R2812 S.n6119 S.n6118 3.643
R2813 S.n6104 S.t2377 3.643
R2814 S.n5764 S.t541 3.643
R2815 S.n5775 S.n5774 3.643
R2816 S.n5772 S.n5771 3.643
R2817 S.n5761 S.t776 3.643
R2818 S.n5342 S.t1297 3.643
R2819 S.n5357 S.n5356 3.643
R2820 S.n5354 S.n5353 3.643
R2821 S.n5339 S.t1833 3.643
R2822 S.n4983 S.t2433 3.643
R2823 S.n4994 S.n4993 3.643
R2824 S.n4991 S.n4990 3.643
R2825 S.n4980 S.t227 3.643
R2826 S.n4565 S.t687 3.643
R2827 S.n4580 S.n4579 3.643
R2828 S.n4577 S.n4576 3.643
R2829 S.n4562 S.t1237 3.643
R2830 S.n4193 S.t1993 3.643
R2831 S.n4204 S.n4203 3.643
R2832 S.n4201 S.n4200 3.643
R2833 S.n4190 S.t2167 3.643
R2834 S.n3765 S.t110 3.643
R2835 S.n3780 S.n3779 3.643
R2836 S.n3777 S.n3776 3.643
R2837 S.n3762 S.t650 3.643
R2838 S.n3346 S.t2403 3.643
R2839 S.n3357 S.n3356 3.643
R2840 S.n3354 S.n3353 3.643
R2841 S.n3343 S.t1672 3.643
R2842 S.n2953 S.t2143 3.643
R2843 S.n2968 S.n2967 3.643
R2844 S.n2965 S.n2964 3.643
R2845 S.n2950 S.t163 3.643
R2846 S.n2490 S.t2379 3.643
R2847 S.n2501 S.n2500 3.643
R2848 S.n2498 S.n2497 3.643
R2849 S.n2487 S.t1633 3.643
R2850 S.n2110 S.t1264 3.643
R2851 S.n2127 S.n2126 3.643
R2852 S.n2124 S.n2123 3.643
R2853 S.n2107 S.t121 3.643
R2854 S.n1209 S.t2359 3.643
R2855 S.n1218 S.n1217 3.643
R2856 S.n1215 S.n1214 3.643
R2857 S.n1206 S.t1608 3.643
R2858 S.n975 S.t695 3.643
R2859 S.n976 S.t1460 3.643
R2860 S.n440 S.t473 3.643
R2861 S.n451 S.n450 3.643
R2862 S.n448 S.n447 3.643
R2863 S.n443 S.t1032 3.643
R2864 S.n10084 S.t812 3.643
R2865 S.n10064 S.t1128 3.643
R2866 S.n9828 S.t1760 3.643
R2867 S.n9843 S.n9842 3.643
R2868 S.n9846 S.n9845 3.643
R2869 S.n9831 S.t1994 3.643
R2870 S.n9398 S.t254 3.643
R2871 S.n9409 S.n9408 3.643
R2872 S.n9406 S.n9405 3.643
R2873 S.n9401 S.t556 3.643
R2874 S.n9005 S.t1175 3.643
R2875 S.n9025 S.n9024 3.643
R2876 S.n9022 S.n9021 3.643
R2877 S.n9008 S.t1695 3.643
R2878 S.n8531 S.t2199 3.643
R2879 S.n8542 S.n8541 3.643
R2880 S.n8539 S.n8538 3.643
R2881 S.n8534 S.t2448 3.643
R2882 S.n8310 S.t697 3.643
R2883 S.n8330 S.n8329 3.643
R2884 S.n8327 S.n8326 3.643
R2885 S.n8313 S.t1256 3.643
R2886 S.n7835 S.t1584 3.643
R2887 S.n7846 S.n7845 3.643
R2888 S.n7843 S.n7842 3.643
R2889 S.n7838 S.t1906 3.643
R2890 S.n7603 S.t133 3.643
R2891 S.n7623 S.n7622 3.643
R2892 S.n7620 S.n7619 3.643
R2893 S.n7606 S.t665 3.643
R2894 S.n7282 S.t1051 3.643
R2895 S.n7293 S.n7292 3.643
R2896 S.n7290 S.n7289 3.643
R2897 S.n7285 S.t1323 3.643
R2898 S.n6873 S.t2067 3.643
R2899 S.n6893 S.n6892 3.643
R2900 S.n6890 S.n6889 3.643
R2901 S.n6876 S.t43 3.643
R2902 S.n6536 S.t449 3.643
R2903 S.n6547 S.n6546 3.643
R2904 S.n6544 S.n6543 3.643
R2905 S.n6539 S.t701 3.643
R2906 S.n6131 S.t1023 3.643
R2907 S.n6151 S.n6150 3.643
R2908 S.n6148 S.n6147 3.643
R2909 S.n6134 S.t1520 3.643
R2910 S.n5781 S.t2182 3.643
R2911 S.n5792 S.n5791 3.643
R2912 S.n5789 S.n5788 3.643
R2913 S.n5784 S.t2428 3.643
R2914 S.n5366 S.t414 3.643
R2915 S.n5386 S.n5385 3.643
R2916 S.n5383 S.n5382 3.643
R2917 S.n5369 S.t967 3.643
R2918 S.n5000 S.t1706 3.643
R2919 S.n5011 S.n5010 3.643
R2920 S.n5008 S.n5007 3.643
R2921 S.n5003 S.t1893 3.643
R2922 S.n4589 S.t2346 3.643
R2923 S.n4609 S.n4608 3.643
R2924 S.n4606 S.n4605 3.643
R2925 S.n4592 S.t354 3.643
R2926 S.n4210 S.t1561 3.643
R2927 S.n4221 S.n4220 3.643
R2928 S.n4218 S.n4217 3.643
R2929 S.n4213 S.t827 3.643
R2930 S.n3789 S.t1305 3.643
R2931 S.n3809 S.n3808 3.643
R2932 S.n3806 S.n3805 3.643
R2933 S.n3792 S.t1858 3.643
R2934 S.n3363 S.t1541 3.643
R2935 S.n3374 S.n3373 3.643
R2936 S.n3371 S.n3370 3.643
R2937 S.n3366 S.t797 3.643
R2938 S.n2977 S.t1279 3.643
R2939 S.n2997 S.n2996 3.643
R2940 S.n2994 S.n2993 3.643
R2941 S.n2980 S.t1826 3.643
R2942 S.n2507 S.t1523 3.643
R2943 S.n2518 S.n2517 3.643
R2944 S.n2515 S.n2514 3.643
R2945 S.n2510 S.t769 3.643
R2946 S.n2136 S.t381 3.643
R2947 S.n2156 S.n2155 3.643
R2948 S.n2153 S.n2152 3.643
R2949 S.n2139 S.t1792 3.643
R2950 S.n1224 S.t1502 3.643
R2951 S.n1237 S.n1236 3.643
R2952 S.n1234 S.n1233 3.643
R2953 S.n1227 S.t744 3.643
R2954 S.n1243 S.t641 3.643
R2955 S.n1257 S.n1256 3.643
R2956 S.n1254 S.n1253 3.643
R2957 S.n1246 S.t2395 3.643
R2958 S.n455 S.t622 3.643
R2959 S.n756 S.n755 3.643
R2960 S.n759 S.n758 3.643
R2961 S.n762 S.t2373 3.643
R2962 S.n770 S.t2123 3.643
R2963 S.n785 S.n784 3.643
R2964 S.n782 S.n781 3.643
R2965 S.n773 S.t135 3.643
R2966 S.n216 S.t2354 3.643
R2967 S.n208 S.t603 3.643
R2968 S.n2174 S.t2032 3.643
R2969 S.n2191 S.n2190 3.643
R2970 S.n2188 S.n2187 3.643
R2971 S.n2171 S.t923 3.643
R2972 S.n3014 S.t393 3.643
R2973 S.n3029 S.n3028 3.643
R2974 S.n3026 S.n3025 3.643
R2975 S.n3011 S.t958 3.643
R2976 S.n3826 S.t423 3.643
R2977 S.n3841 S.n3840 3.643
R2978 S.n3838 S.n3837 3.643
R2979 S.n3823 S.t991 3.643
R2980 S.n4626 S.t463 3.643
R2981 S.n4641 S.n4640 3.643
R2982 S.n4638 S.n4637 3.643
R2983 S.n4623 S.t1019 3.643
R2984 S.n5403 S.t2061 3.643
R2985 S.n5418 S.n5417 3.643
R2986 S.n5415 S.n5414 3.643
R2987 S.n5400 S.t32 3.643
R2988 S.n6168 S.t120 3.643
R2989 S.n6183 S.n6182 3.643
R2990 S.n6180 S.n6179 3.643
R2991 S.n6165 S.t660 3.643
R2992 S.n6910 S.t1205 3.643
R2993 S.n6925 S.n6924 3.643
R2994 S.n6922 S.n6921 3.643
R2995 S.n6907 S.t1737 3.643
R2996 S.n7640 S.t1802 3.643
R2997 S.n7655 S.n7654 3.643
R2998 S.n7652 S.n7651 3.643
R2999 S.n7637 S.t2319 3.643
R3000 S.n8347 S.t2356 3.643
R3001 S.n8362 S.n8361 3.643
R3002 S.n8359 S.n8358 3.643
R3003 S.n8344 S.t374 3.643
R3004 S.n9042 S.t433 3.643
R3005 S.n9057 S.n9056 3.643
R3006 S.n9054 S.n9053 3.643
R3007 S.n9039 S.t987 3.643
R3008 S.n9714 S.t883 3.643
R3009 S.n9729 S.n9728 3.643
R3010 S.n9726 S.n9725 3.643
R3011 S.n9711 S.t1144 3.643
R3012 S.n10487 S.t1186 3.643
R3013 S.n10501 S.n10500 3.643
R3014 S.n10504 S.n10503 3.643
R3015 S.n10484 S.t1708 3.643
R3016 S.n10756 S.t568 3.643
R3017 S.n10737 S.t810 3.643
R3018 S.n10093 S.t2460 3.643
R3019 S.n10104 S.n10103 3.643
R3020 S.n10101 S.n10100 3.643
R3021 S.n10090 S.t250 3.643
R3022 S.n9417 S.t1921 3.643
R3023 S.n9428 S.n9427 3.643
R3024 S.n9425 S.n9424 3.643
R3025 S.n9414 S.t2195 3.643
R3026 S.n8550 S.t1341 3.643
R3027 S.n8561 S.n8560 3.643
R3028 S.n8558 S.n8557 3.643
R3029 S.n8547 S.t1580 3.643
R3030 S.n7854 S.t717 3.643
R3031 S.n7865 S.n7864 3.643
R3032 S.n7862 S.n7861 3.643
R3033 S.n7851 S.t1047 3.643
R3034 S.n7301 S.t162 3.643
R3035 S.n7312 S.n7311 3.643
R3036 S.n7309 S.n7308 3.643
R3037 S.n7298 S.t443 3.643
R3038 S.n6555 S.t2092 3.643
R3039 S.n6566 S.n6565 3.643
R3040 S.n6563 S.n6562 3.643
R3041 S.n6552 S.t2360 3.643
R3042 S.n5800 S.t1445 3.643
R3043 S.n5811 S.n5810 3.643
R3044 S.n5808 S.n5807 3.643
R3045 S.n5797 S.t1562 3.643
R3046 S.n5019 S.t722 3.643
R3047 S.n5030 S.n5029 3.643
R3048 S.n5027 S.n5026 3.643
R3049 S.n5016 S.t2504 3.643
R3050 S.n4229 S.t698 3.643
R3051 S.n4240 S.n4239 3.643
R3052 S.n4237 S.n4236 3.643
R3053 S.n4226 S.t2474 3.643
R3054 S.n3382 S.t681 3.643
R3055 S.n3393 S.n3392 3.643
R3056 S.n3390 S.n3389 3.643
R3057 S.n3379 S.t2449 3.643
R3058 S.n2526 S.t662 3.643
R3059 S.n2537 S.n2536 3.643
R3060 S.n2534 S.n2533 3.643
R3061 S.n2523 S.t2420 3.643
R3062 S.n1721 S.t1291 3.643
R3063 S.n1740 S.n1739 3.643
R3064 S.n1737 S.n1736 3.643
R3065 S.n1724 S.t1832 3.643
R3066 S.n680 S.t2280 3.643
R3067 S.n695 S.n694 3.643
R3068 S.n692 S.n691 3.643
R3069 S.n683 S.t1517 3.643
R3070 S.n225 S.t1258 3.643
R3071 S.n887 S.n886 3.643
R3072 S.n890 S.n889 3.643
R3073 S.n893 S.t1804 3.643
R3074 S.n922 S.t1496 3.643
R3075 S.n219 S.t2256 3.643
R3076 S.n11398 S.t260 3.643
R3077 S.n11375 S.t567 3.643
R3078 S.n11116 S.t901 3.643
R3079 S.n11124 S.n11123 3.643
R3080 S.n11127 S.n11126 3.643
R3081 S.n11113 S.t1446 3.643
R3082 S.n10770 S.t2211 3.643
R3083 S.n10778 S.n10777 3.643
R3084 S.n10775 S.n10774 3.643
R3085 S.n10767 S.t2457 3.643
R3086 S.n10405 S.t311 3.643
R3087 S.n10423 S.n10422 3.643
R3088 S.n10420 S.n10419 3.643
R3089 S.n10402 S.t837 3.643
R3090 S.n10117 S.t1592 3.643
R3091 S.n10125 S.n10124 3.643
R3092 S.n10122 S.n10121 3.643
R3093 S.n10114 S.t1916 3.643
R3094 S.n9745 S.t147 3.643
R3095 S.n9763 S.n9762 3.643
R3096 S.n9760 S.n9759 3.643
R3097 S.n9742 S.t385 3.643
R3098 S.n9441 S.t1059 3.643
R3099 S.n9449 S.n9448 3.643
R3100 S.n9446 S.n9445 3.643
R3101 S.n9438 S.t1339 3.643
R3102 S.n9073 S.t2080 3.643
R3103 S.n9091 S.n9090 3.643
R3104 S.n9088 S.n9087 3.643
R3105 S.n9070 S.t68 3.643
R3106 S.n8574 S.t462 3.643
R3107 S.n8582 S.n8581 3.643
R3108 S.n8579 S.n8578 3.643
R3109 S.n8571 S.t713 3.643
R3110 S.n8378 S.t1500 3.643
R3111 S.n8396 S.n8395 3.643
R3112 S.n8393 S.n8392 3.643
R3113 S.n8375 S.t2025 3.643
R3114 S.n7878 S.t2372 3.643
R3115 S.n7886 S.n7885 3.643
R3116 S.n7883 S.n7882 3.643
R3117 S.n7875 S.t157 3.643
R3118 S.n7671 S.t932 3.643
R3119 S.n7689 S.n7688 3.643
R3120 S.n7686 S.n7685 3.643
R3121 S.n7668 S.t1458 3.643
R3122 S.n7325 S.t1823 3.643
R3123 S.n7333 S.n7332 3.643
R3124 S.n7330 S.n7329 3.643
R3125 S.n7322 S.t2087 3.643
R3126 S.n6941 S.t327 3.643
R3127 S.n6959 S.n6958 3.643
R3128 S.n6956 S.n6955 3.643
R3129 S.n6938 S.t862 3.643
R3130 S.n6579 S.t1375 3.643
R3131 S.n6587 S.n6586 3.643
R3132 S.n6584 S.n6583 3.643
R3133 S.n6576 S.t1504 3.643
R3134 S.n6199 S.t1791 3.643
R3135 S.n6217 S.n6216 3.643
R3136 S.n6214 S.n6213 3.643
R3137 S.n6196 S.t2315 3.643
R3138 S.n5824 S.t2398 3.643
R3139 S.n5832 S.n5831 3.643
R3140 S.n5829 S.n5828 3.643
R3141 S.n5821 S.t1664 3.643
R3142 S.n5434 S.t2139 3.643
R3143 S.n5452 S.n5451 3.643
R3144 S.n5449 S.n5448 3.643
R3145 S.n5431 S.t154 3.643
R3146 S.n5043 S.t2375 3.643
R3147 S.n5051 S.n5050 3.643
R3148 S.n5048 S.n5047 3.643
R3149 S.n5040 S.t1629 3.643
R3150 S.n4657 S.t2108 3.643
R3151 S.n4675 S.n4674 3.643
R3152 S.n4672 S.n4671 3.643
R3153 S.n4654 S.t113 3.643
R3154 S.n4253 S.t2357 3.643
R3155 S.n4261 S.n4260 3.643
R3156 S.n4258 S.n4257 3.643
R3157 S.n4250 S.t1603 3.643
R3158 S.n3857 S.t2075 3.643
R3159 S.n3875 S.n3874 3.643
R3160 S.n3872 S.n3871 3.643
R3161 S.n3854 S.t79 3.643
R3162 S.n3406 S.t2340 3.643
R3163 S.n3414 S.n3413 3.643
R3164 S.n3411 S.n3410 3.643
R3165 S.n3403 S.t1581 3.643
R3166 S.n3045 S.t2045 3.643
R3167 S.n3063 S.n3062 3.643
R3168 S.n3060 S.n3059 3.643
R3169 S.n3042 S.t11 3.643
R3170 S.n2550 S.t2317 3.643
R3171 S.n2558 S.n2557 3.643
R3172 S.n2555 S.n2554 3.643
R3173 S.n2547 S.t1554 3.643
R3174 S.n2207 S.t1317 3.643
R3175 S.n2225 S.n2224 3.643
R3176 S.n2222 S.n2221 3.643
R3177 S.n2204 S.t183 3.643
R3178 S.n1270 S.t2299 3.643
R3179 S.n1278 S.n1277 3.643
R3180 S.n1275 S.n1274 3.643
R3181 S.n1267 S.t1535 3.643
R3182 S.n1749 S.t404 3.643
R3183 S.n1768 S.n1767 3.643
R3184 S.n1765 S.n1764 3.643
R3185 S.n1752 S.t966 3.643
R3186 S.n700 S.t1425 3.643
R3187 S.n714 S.n713 3.643
R3188 S.n711 S.n710 3.643
R3189 S.n703 S.t656 3.643
R3190 S.n1289 S.t1443 3.643
R3191 S.n1298 S.n1297 3.643
R3192 S.n1295 S.n1294 3.643
R3193 S.n1286 S.t675 3.643
R3194 S.n2234 S.t438 3.643
R3195 S.n2246 S.n2245 3.643
R3196 S.n2243 S.n2242 3.643
R3197 S.n2237 S.t1847 3.643
R3198 S.n2564 S.t1457 3.643
R3199 S.n2578 S.n2577 3.643
R3200 S.n2575 S.n2574 3.643
R3201 S.n2567 S.t691 3.643
R3202 S.n3072 S.t1333 3.643
R3203 S.n3083 S.n3082 3.643
R3204 S.n3080 S.n3079 3.643
R3205 S.n3075 S.t1876 3.643
R3206 S.n3420 S.t1481 3.643
R3207 S.n3434 S.n3433 3.643
R3208 S.n3431 S.n3430 3.643
R3209 S.n3423 S.t714 3.643
R3210 S.n3884 S.t1214 3.643
R3211 S.n3895 S.n3894 3.643
R3212 S.n3892 S.n3891 3.643
R3213 S.n3887 S.t1758 3.643
R3214 S.n4267 S.t1499 3.643
R3215 S.n4281 S.n4280 3.643
R3216 S.n4278 S.n4277 3.643
R3217 S.n4270 S.t739 3.643
R3218 S.n4684 S.t1243 3.643
R3219 S.n4695 S.n4694 3.643
R3220 S.n4692 S.n4691 3.643
R3221 S.n4687 S.t1787 3.643
R3222 S.n5057 S.t1519 3.643
R3223 S.n5071 S.n5070 3.643
R3224 S.n5068 S.n5067 3.643
R3225 S.n5060 S.t762 3.643
R3226 S.n5461 S.t1273 3.643
R3227 S.n5472 S.n5471 3.643
R3228 S.n5469 S.n5468 3.643
R3229 S.n5464 S.t1818 3.643
R3230 S.n5838 S.t1536 3.643
R3231 S.n5852 S.n5851 3.643
R3232 S.n5849 S.n5848 3.643
R3233 S.n5841 S.t792 3.643
R3234 S.n6226 S.t1303 3.643
R3235 S.n6237 S.n6236 3.643
R3236 S.n6234 S.n6233 3.643
R3237 S.n6229 S.t1851 3.643
R3238 S.n6593 S.t1962 3.643
R3239 S.n6607 S.n6606 3.643
R3240 S.n6604 S.n6603 3.643
R3241 S.n6596 S.t1218 3.643
R3242 S.n6968 S.t1986 3.643
R3243 S.n6979 S.n6978 3.643
R3244 S.n6976 S.n6975 3.643
R3245 S.n6971 S.t2507 3.643
R3246 S.n7339 S.t1084 3.643
R3247 S.n7353 S.n7352 3.643
R3248 S.n7350 S.n7349 3.643
R3249 S.n7342 S.t1223 3.643
R3250 S.n7698 S.t2573 3.643
R3251 S.n7709 S.n7708 3.643
R3252 S.n7706 S.n7705 3.643
R3253 S.n7701 S.t600 3.643
R3254 S.n7892 S.t1515 3.643
R3255 S.n7906 S.n7905 3.643
R3256 S.n7903 S.n7902 3.643
R3257 S.n7895 S.t1820 3.643
R3258 S.n8405 S.t637 3.643
R3259 S.n8416 S.n8415 3.643
R3260 S.n8413 S.n8412 3.643
R3261 S.n8408 S.t1168 3.643
R3262 S.n8588 S.t2113 3.643
R3263 S.n8602 S.n8601 3.643
R3264 S.n8599 S.n8598 3.643
R3265 S.n8591 S.t2368 3.643
R3266 S.n9100 S.t1217 3.643
R3267 S.n9111 S.n9110 3.643
R3268 S.n9108 S.n9107 3.643
R3269 S.n9103 S.t1752 3.643
R3270 S.n9455 S.t174 3.643
R3271 S.n9469 S.n9468 3.643
R3272 S.n9466 S.n9465 3.643
R3273 S.n9458 S.t458 3.643
R3274 S.n9772 S.t1816 3.643
R3275 S.n9783 S.n9782 3.643
R3276 S.n9780 S.n9779 3.643
R3277 S.n9775 S.t2035 3.643
R3278 S.n10131 S.t728 3.643
R3279 S.n10145 S.n10144 3.643
R3280 S.n10142 S.n10141 3.643
R3281 S.n10134 S.t1056 3.643
R3282 S.n10432 S.t2095 3.643
R3283 S.n10443 S.n10442 3.643
R3284 S.n10440 S.n10439 3.643
R3285 S.n10435 S.t92 3.643
R3286 S.n10784 S.t1352 3.643
R3287 S.n10798 S.n10797 3.643
R3288 S.n10795 S.n10794 3.643
R3289 S.n10787 S.t1589 3.643
R3290 S.n11057 S.t2544 3.643
R3291 S.n11068 S.n11067 3.643
R3292 S.n11065 S.n11064 3.643
R3293 S.n11060 S.t584 3.643
R3294 S.n11405 S.t1926 3.643
R3295 S.n11419 S.n11418 3.643
R3296 S.n11416 S.n11415 3.643
R3297 S.n11408 S.t2210 3.643
R3298 S.n11711 S.t620 3.643
R3299 S.n11719 S.n11718 3.643
R3300 S.n11722 S.n11721 3.643
R3301 S.n11714 S.t1152 3.643
R3302 S.n11970 S.t2471 3.643
R3303 S.n11949 S.t258 3.643
R3304 S.n939 S.t633 3.643
R3305 S.n926 S.t1396 3.643
R3306 S.n790 S.t373 3.643
R3307 S.n807 S.n806 3.643
R3308 S.n804 S.n803 3.643
R3309 S.n793 S.t937 3.643
R3310 S.n1687 S.t348 3.643
R3311 S.n1706 S.n1705 3.643
R3312 S.n1703 S.n1702 3.643
R3313 S.n1690 S.t908 3.643
R3314 S.n664 S.t1483 3.643
R3315 S.n675 S.n674 3.643
R3316 S.n672 S.n671 3.643
R3317 S.n667 S.t720 3.643
R3318 S.n647 S.t2342 3.643
R3319 S.n658 S.n657 3.643
R3320 S.n655 S.n654 3.643
R3321 S.n650 S.t1585 3.643
R3322 S.n189 S.t772 3.643
R3323 S.n182 S.t1528 3.643
R3324 S.n379 S.t416 3.643
R3325 S.n390 S.n389 3.643
R3326 S.n387 S.n386 3.643
R3327 S.n382 S.t984 3.643
R3328 S.n1606 S.t451 3.643
R3329 S.n1619 S.n1618 3.643
R3330 S.n1616 S.n1615 3.643
R3331 S.n1603 S.t1007 3.643
R3332 S.n7792 S.t1677 3.643
R3333 S.n7773 S.t1974 3.643
R3334 S.n7750 S.t60 3.643
R3335 S.n7764 S.n7763 3.643
R3336 S.n7767 S.n7766 3.643
R3337 S.n7747 S.t626 3.643
R3338 S.n7229 S.t1122 3.643
R3339 S.n7240 S.n7239 3.643
R3340 S.n7237 S.n7236 3.643
R3341 S.n7226 S.t1410 3.643
R3342 S.n6788 S.t2020 3.643
R3343 S.n6803 S.n6802 3.643
R3344 S.n6800 S.n6799 3.643
R3345 S.n6785 S.t2554 3.643
R3346 S.n6483 S.t551 3.643
R3347 S.n6494 S.n6493 3.643
R3348 S.n6491 S.n6490 3.643
R3349 S.n6480 S.t783 3.643
R3350 S.n6046 S.t1096 3.643
R3351 S.n6061 S.n6060 3.643
R3352 S.n6058 S.n6057 3.643
R3353 S.n6043 S.t1588 3.643
R3354 S.n5728 S.t2267 3.643
R3355 S.n5739 S.n5738 3.643
R3356 S.n5736 S.n5735 3.643
R3357 S.n5725 S.t2523 3.643
R3358 S.n5281 S.t516 3.643
R3359 S.n5296 S.n5295 3.643
R3360 S.n5293 S.n5292 3.643
R3361 S.n5278 S.t1055 3.643
R3362 S.n4947 S.t1651 3.643
R3363 S.n4958 S.n4957 3.643
R3364 S.n4955 S.n4954 3.643
R3365 S.n4944 S.t1960 3.643
R3366 S.n4504 S.t2413 3.643
R3367 S.n4519 S.n4518 3.643
R3368 S.n4516 S.n4515 3.643
R3369 S.n4501 S.t457 3.643
R3370 S.n4157 S.t1105 3.643
R3371 S.n4168 S.n4167 3.643
R3372 S.n4165 S.n4164 3.643
R3373 S.n4154 S.t1395 3.643
R3374 S.n3704 S.t1878 3.643
R3375 S.n3719 S.n3718 3.643
R3376 S.n3716 S.n3715 3.643
R3377 S.n3701 S.t2367 3.643
R3378 S.n3310 S.t526 3.643
R3379 S.n3321 S.n3320 3.643
R3380 S.n3318 S.n3317 3.643
R3381 S.n3307 S.t768 3.643
R3382 S.n2892 S.t1287 3.643
R3383 S.n2907 S.n2906 3.643
R3384 S.n2904 S.n2903 3.643
R3385 S.n2889 S.t1819 3.643
R3386 S.n2454 S.t2571 3.643
R3387 S.n2465 S.n2464 3.643
R3388 S.n2462 S.n2461 3.643
R3389 S.n2451 S.t216 3.643
R3390 S.n2047 S.t999 3.643
R3391 S.n2064 S.n2063 3.643
R3392 S.n2061 S.n2060 3.643
R3393 S.n2044 S.t1224 3.643
R3394 S.n1175 S.t1566 3.643
R3395 S.n1184 S.n1183 3.643
R3396 S.n1181 S.n1180 3.643
R3397 S.n1172 S.t834 3.643
R3398 S.n971 S.t2423 3.643
R3399 S.n972 S.t668 3.643
R3400 S.n399 S.t2066 3.643
R3401 S.n410 S.n409 3.643
R3402 S.n407 S.n406 3.643
R3403 S.n402 S.t62 3.643
R3404 S.n8505 S.t1427 3.643
R3405 S.n8485 S.t1671 3.643
R3406 S.n8461 S.t2325 3.643
R3407 S.n8476 S.n8475 3.643
R3408 S.n8479 S.n8478 3.643
R3409 S.n8464 S.t325 3.643
R3410 S.n7799 S.t802 3.643
R3411 S.n7810 S.n7809 3.643
R3412 S.n7807 S.n7806 3.643
R3413 S.n7802 S.t1119 3.643
R3414 S.n7542 S.t1747 3.643
R3415 S.n7562 S.n7561 3.643
R3416 S.n7559 S.n7558 3.643
R3417 S.n7545 S.t2285 3.643
R3418 S.n7246 S.t244 3.643
R3419 S.n7257 S.n7256 3.643
R3420 S.n7254 S.n7253 3.643
R3421 S.n7249 S.t545 3.643
R3422 S.n6812 S.t1302 3.643
R3423 S.n6832 S.n6831 3.643
R3424 S.n6829 S.n6828 3.643
R3425 S.n6815 S.t1840 3.643
R3426 S.n6500 S.t2190 3.643
R3427 S.n6511 S.n6510 3.643
R3428 S.n6508 S.n6507 3.643
R3429 S.n6503 S.t2436 3.643
R3430 S.n6070 S.t221 3.643
R3431 S.n6090 S.n6089 3.643
R3432 S.n6087 S.n6086 3.643
R3433 S.n6073 S.t723 3.643
R3434 S.n5745 S.t1408 3.643
R3435 S.n5756 S.n5755 3.643
R3436 S.n5753 S.n5752 3.643
R3437 S.n5748 S.t1648 3.643
R3438 S.n5305 S.t2161 3.643
R3439 S.n5325 S.n5324 3.643
R3440 S.n5322 S.n5321 3.643
R3441 S.n5308 S.t168 3.643
R3442 S.n4964 S.t780 3.643
R3443 S.n4975 S.n4974 3.643
R3444 S.n4972 S.n4971 3.643
R3445 S.n4967 S.t1102 3.643
R3446 S.n4528 S.t1549 3.643
R3447 S.n4548 S.n4547 3.643
R3448 S.n4545 S.n4544 3.643
R3449 S.n4531 S.t2103 3.643
R3450 S.n4174 S.t229 3.643
R3451 S.n4185 S.n4184 3.643
R3452 S.n4182 S.n4181 3.643
R3453 S.n4177 S.t523 3.643
R3454 S.n3728 S.t1013 3.643
R3455 S.n3748 S.n3747 3.643
R3456 S.n3745 S.n3744 3.643
R3457 S.n3731 S.t1510 3.643
R3458 S.n3327 S.t2291 3.643
R3459 S.n3338 S.n3337 3.643
R3460 S.n3335 S.n3334 3.643
R3461 S.n3330 S.t2417 3.643
R3462 S.n2916 S.t400 3.643
R3463 S.n2936 S.n2935 3.643
R3464 S.n2933 S.n2932 3.643
R3465 S.n2919 S.t955 3.643
R3466 S.n2471 S.t727 3.643
R3467 S.n2482 S.n2481 3.643
R3468 S.n2479 S.n2478 3.643
R3469 S.n2474 S.t2509 3.643
R3470 S.n2073 S.t2128 3.643
R3471 S.n2093 S.n2092 3.643
R3472 S.n2090 S.n2089 3.643
R3473 S.n2076 S.t1025 3.643
R3474 S.n1190 S.t700 3.643
R3475 S.n1201 S.n1200 3.643
R3476 S.n1198 S.n1197 3.643
R3477 S.n1193 S.t2479 3.643
R3478 S.n1628 S.t2096 3.643
R3479 S.n1648 S.n1647 3.643
R3480 S.n1645 S.n1644 3.643
R3481 S.n1631 S.t107 3.643
R3482 S.n631 S.t683 3.643
R3483 S.n642 S.n641 3.643
R3484 S.n639 S.n638 3.643
R3485 S.n634 S.t2453 3.643
R3486 S.n614 S.t1544 3.643
R3487 S.n625 S.n624 3.643
R3488 S.n622 S.n621 3.643
R3489 S.n617 S.t803 3.643
R3490 S.n177 S.t2516 3.643
R3491 S.n169 S.t729 3.643
R3492 S.n338 S.t1534 3.643
R3493 S.n349 S.n348 3.643
R3494 S.n346 S.n345 3.643
R3495 S.n341 S.t2074 3.643
R3496 S.n1547 S.t2137 3.643
R3497 S.n1560 S.n1559 3.643
R3498 S.n1557 S.n1556 3.643
R3499 S.n1544 S.t138 3.643
R3500 S.n6457 S.t2271 3.643
R3501 S.n6438 S.t2529 3.643
R3502 S.n6278 S.t176 3.643
R3503 S.n6292 S.n6291 3.643
R3504 S.n6295 S.n6294 3.643
R3505 S.n6275 S.t686 3.643
R3506 S.n5692 S.t1475 3.643
R3507 S.n5703 S.n5702 3.643
R3508 S.n5700 S.n5699 3.643
R3509 S.n5689 S.t1755 3.643
R3510 S.n5220 S.t2114 3.643
R3511 S.n5235 S.n5234 3.643
R3512 S.n5232 S.n5231 3.643
R3513 S.n5217 S.t106 3.643
R3514 S.n4911 S.t882 3.643
R3515 S.n4922 S.n4921 3.643
R3516 S.n4919 S.n4918 3.643
R3517 S.n4908 S.t1171 3.643
R3518 S.n4443 S.t1627 3.643
R3519 S.n4458 S.n4457 3.643
R3520 S.n4455 S.n4454 3.643
R3521 S.n4440 S.t2193 3.643
R3522 S.n4121 S.t298 3.643
R3523 S.n4132 S.n4131 3.643
R3524 S.n4129 S.n4128 3.643
R3525 S.n4118 S.t601 3.643
R3526 S.n3643 S.t1088 3.643
R3527 S.n3658 S.n3657 3.643
R3528 S.n3655 S.n3654 3.643
R3529 S.n3640 S.t1579 3.643
R3530 S.n3274 S.t2258 3.643
R3531 S.n3285 S.n3284 3.643
R3532 S.n3282 S.n3281 3.643
R3533 S.n3271 S.t2508 3.643
R3534 S.n2831 S.t504 3.643
R3535 S.n2846 S.n2845 3.643
R3536 S.n2843 S.n2842 3.643
R3537 S.n2828 S.t1046 3.643
R3538 S.n2418 S.t1638 3.643
R3539 S.n2429 S.n2428 3.643
R3540 S.n2426 S.n2425 3.643
R3541 S.n2415 S.t1953 3.643
R3542 S.n1984 S.t201 3.643
R3543 S.n2001 S.n2000 3.643
R3544 S.n1998 S.n1997 3.643
R3545 S.n1981 S.t441 3.643
R3546 S.n1141 S.t1095 3.643
R3547 S.n1150 S.n1149 3.643
R3548 S.n1147 S.n1146 3.643
R3549 S.n1138 S.t1385 3.643
R3550 S.n967 S.t1639 3.643
R3551 S.n968 S.t2382 3.643
R3552 S.n358 S.t1299 3.643
R3553 S.n369 S.n368 3.643
R3554 S.n366 S.n365 3.643
R3555 S.n361 S.t1846 3.643
R3556 S.n7220 S.t1976 3.643
R3557 S.n7200 S.t2269 3.643
R3558 S.n7024 S.t368 3.643
R3559 S.n7039 S.n7038 3.643
R3560 S.n7042 S.n7041 3.643
R3561 S.n7027 S.t913 3.643
R3562 S.n6464 S.t1415 3.643
R3563 S.n6475 S.n6474 3.643
R3564 S.n6472 S.n6471 3.643
R3565 S.n6467 S.t1654 3.643
R3566 S.n6009 S.t1841 3.643
R3567 S.n6029 S.n6028 3.643
R3568 S.n6026 S.n6025 3.643
R3569 S.n6012 S.t2345 3.643
R3570 S.n5709 S.t614 3.643
R3571 S.n5720 S.n5719 3.643
R3572 S.n5717 S.n5716 3.643
R3573 S.n5712 S.t876 3.643
R3574 S.n5244 S.t1389 3.643
R3575 S.n5264 S.n5263 3.643
R3576 S.n5261 S.n5260 3.643
R3577 S.n5247 S.t1915 3.643
R3578 S.n4928 S.t2527 3.643
R3579 S.n4939 S.n4938 3.643
R3580 S.n4936 S.n4935 3.643
R3581 S.n4931 S.t294 3.643
R3582 S.n4467 S.t760 3.643
R3583 S.n4487 S.n4486 3.643
R3584 S.n4484 S.n4483 3.643
R3585 S.n4470 S.t1337 3.643
R3586 S.n4138 S.t1961 3.643
R3587 S.n4149 S.n4148 3.643
R3588 S.n4146 S.n4145 3.643
R3589 S.n4141 S.t2254 3.643
R3590 S.n3667 S.t210 3.643
R3591 S.n3687 S.n3686 3.643
R3592 S.n3684 S.n3683 3.643
R3593 S.n3670 S.t712 3.643
R3594 S.n3291 S.t1397 3.643
R3595 S.n3302 S.n3301 3.643
R3596 S.n3299 S.n3298 3.643
R3597 S.n3294 S.t1636 3.643
R3598 S.n2855 S.t2147 3.643
R3599 S.n2875 S.n2874 3.643
R3600 S.n2872 S.n2871 3.643
R3601 S.n2858 S.t155 3.643
R3602 S.n2435 S.t771 3.643
R3603 S.n2446 S.n2445 3.643
R3604 S.n2443 S.n2442 3.643
R3605 S.n2438 S.t1093 3.643
R3606 S.n2010 S.t1866 3.643
R3607 S.n2030 S.n2029 3.643
R3608 S.n2027 S.n2026 3.643
R3609 S.n2013 S.t2086 3.643
R3610 S.n1156 S.t326 3.643
R3611 S.n1167 S.n1166 3.643
R3612 S.n1164 S.n1163 3.643
R3613 S.n1159 S.t510 3.643
R3614 S.n1569 S.t1272 3.643
R3615 S.n1589 S.n1588 3.643
R3616 S.n1586 S.n1585 3.643
R3617 S.n1572 S.t1807 3.643
R3618 S.n598 S.t2406 3.643
R3619 S.n609 S.n608 3.643
R3620 S.n606 S.n605 3.643
R3621 S.n601 S.t1678 3.643
R3622 S.n581 S.t627 3.643
R3623 S.n592 S.n591 3.643
R3624 S.n589 S.n588 3.643
R3625 S.n584 S.t755 3.643
R3626 S.n164 S.t1942 3.643
R3627 S.n156 S.t1626 3.643
R3628 S.n317 S.t742 3.643
R3629 S.n328 S.n327 3.643
R3630 S.n325 S.n324 3.643
R3631 S.n320 S.t1309 3.643
R3632 S.n1488 S.t1366 3.643
R3633 S.n1501 S.n1500 3.643
R3634 S.n1498 S.n1497 3.643
R3635 S.n1485 S.t1895 3.643
R3636 S.n4885 S.t82 3.643
R3637 S.n4866 S.t376 3.643
R3638 S.n4736 S.t719 3.643
R3639 S.n4750 S.n4749 3.643
R3640 S.n4753 S.n4752 3.643
R3641 S.n4733 S.t1284 3.643
R3642 S.n4085 S.t2029 3.643
R3643 S.n4096 S.n4095 3.643
R3644 S.n4093 S.n4092 3.643
R3645 S.n4082 S.t2321 3.643
R3646 S.n3582 S.t165 3.643
R3647 S.n3597 S.n3596 3.643
R3648 S.n3594 S.n3593 3.643
R3649 S.n3579 S.t680 3.643
R3650 S.n3238 S.t1465 3.643
R3651 S.n3249 S.n3248 3.643
R3652 S.n3246 S.n3245 3.643
R3653 S.n3235 S.t1739 3.643
R3654 S.n2770 S.t2237 3.643
R3655 S.n2785 S.n2784 3.643
R3656 S.n2782 S.n2781 3.643
R3657 S.n2767 S.t238 3.643
R3658 S.n2382 S.t870 3.643
R3659 S.n2393 S.n2392 3.643
R3660 S.n2390 S.n2389 3.643
R3661 S.n2379 S.t1162 3.643
R3662 S.n1921 S.t1935 3.643
R3663 S.n1938 S.n1937 3.643
R3664 S.n1935 S.n1934 3.643
R3665 S.n1918 S.t2185 3.643
R3666 S.n1107 S.t292 3.643
R3667 S.n1116 S.n1115 3.643
R3668 S.n1113 S.n1112 3.643
R3669 S.n1104 S.t595 3.643
R3670 S.n963 S.t1081 3.643
R3671 S.n964 S.t914 3.643
R3672 S.n47 S.t2391 3.643
R3673 S.n50 S.n49 3.643
R3674 S.n53 S.n52 3.643
R3675 S.n56 S.t426 3.643
R3676 S.n5683 S.t2332 3.643
R3677 S.n5663 S.t75 3.643
R3678 S.n5517 S.t467 3.643
R3679 S.n5532 S.n5531 3.643
R3680 S.n5535 S.n5534 3.643
R3681 S.n5520 S.t1009 3.643
R3682 S.n4892 S.t1759 3.643
R3683 S.n4903 S.n4902 3.643
R3684 S.n4900 S.n4899 3.643
R3685 S.n4895 S.t2027 3.643
R3686 S.n4406 S.t2374 3.643
R3687 S.n4426 S.n4425 3.643
R3688 S.n4423 S.n4422 3.643
R3689 S.n4409 S.t399 3.643
R3690 S.n4102 S.t1174 3.643
R3691 S.n4113 S.n4112 3.643
R3692 S.n4110 S.n4109 3.643
R3693 S.n4105 S.t1459 3.643
R3694 S.n3606 S.t1945 3.643
R3695 S.n3626 S.n3625 3.643
R3696 S.n3623 S.n3622 3.643
R3697 S.n3609 S.t2446 3.643
R3698 S.n3255 S.t606 3.643
R3699 S.n3266 S.n3265 3.643
R3700 S.n3263 S.n3262 3.643
R3701 S.n3258 S.t864 3.643
R3702 S.n2794 S.t1378 3.643
R3703 S.n2814 S.n2813 3.643
R3704 S.n2811 S.n2810 3.643
R3705 S.n2797 S.t1905 3.643
R3706 S.n2399 S.t2514 3.643
R3707 S.n2410 S.n2409 3.643
R3708 S.n2407 S.n2406 3.643
R3709 S.n2402 S.t290 3.643
R3710 S.n1947 S.t1077 3.643
R3711 S.n1967 S.n1966 3.643
R3712 S.n1964 S.n1963 3.643
R3713 S.n1950 S.t1321 3.643
R3714 S.n1122 S.t1955 3.643
R3715 S.n1133 S.n1132 3.643
R3716 S.n1130 S.n1129 3.643
R3717 S.n1125 S.t2244 3.643
R3718 S.n1510 S.t492 3.643
R3719 S.n1530 S.n1529 3.643
R3720 S.n1527 S.n1526 3.643
R3721 S.n1513 S.t1035 3.643
R3722 S.n565 S.t1388 3.643
R3723 S.n576 S.n575 3.643
R3724 S.n573 S.n572 3.643
R3725 S.n568 S.t1620 3.643
R3726 S.n548 S.t2247 3.643
R3727 S.n559 S.n558 3.643
R3728 S.n556 S.n555 3.643
R3729 S.n551 S.t2497 3.643
R3730 S.n151 S.t1154 3.643
R3731 S.n143 S.t858 3.643
R3732 S.n276 S.t2477 3.643
R3733 S.n287 S.n286 3.643
R3734 S.n284 S.n283 3.643
R3735 S.n279 S.t527 3.643
R3736 S.n1429 S.t582 3.643
R3737 S.n1442 S.n1441 3.643
R3738 S.n1439 S.n1438 3.643
R3739 S.n1426 S.t1106 3.643
R3740 S.n3212 S.t669 3.643
R3741 S.n3193 S.t978 3.643
R3742 S.n3124 S.t1330 3.643
R3743 S.n3138 S.n3137 3.643
R3744 S.n3141 S.n3140 3.643
R3745 S.n3121 S.t1867 3.643
R3746 S.n2346 S.t56 3.643
R3747 S.n2357 S.n2356 3.643
R3748 S.n2354 S.n2353 3.643
R3749 S.n2343 S.t363 3.643
R3750 S.n1858 S.t1043 3.643
R3751 S.n1875 S.n1874 3.643
R3752 S.n1872 S.n1871 3.643
R3753 S.n1855 S.t1271 3.643
R3754 S.n1073 S.t2019 3.643
R3755 S.n1082 S.n1081 3.643
R3756 S.n1079 S.n1078 3.643
R3757 S.n1070 S.t2311 3.643
R3758 S.n959 S.t279 3.643
R3759 S.n960 S.t2502 3.643
R3760 S.n296 S.t1606 3.643
R3761 S.n307 S.n306 3.643
R3762 S.n304 S.n303 3.643
R3763 S.n299 S.t2172 3.643
R3764 S.n4076 S.t380 3.643
R3765 S.n4056 S.t667 3.643
R3766 S.n3940 S.t1053 3.643
R3767 S.n3955 S.n3954 3.643
R3768 S.n3958 S.n3957 3.643
R3769 S.n3943 S.t1540 3.643
R3770 S.n3219 S.t2323 3.643
R3771 S.n3230 S.n3229 3.643
R3772 S.n3227 S.n3226 3.643
R3773 S.n3222 S.t47 3.643
R3774 S.n2733 S.t450 3.643
R3775 S.n2753 S.n2752 3.643
R3776 S.n2750 S.n2749 3.643
R3777 S.n2736 S.t998 3.643
R3778 S.n2363 S.t1746 3.643
R3779 S.n2374 S.n2373 3.643
R3780 S.n2371 S.n2370 3.643
R3781 S.n2366 S.t2015 3.643
R3782 S.n1884 S.t272 3.643
R3783 S.n1904 S.n1903 3.643
R3784 S.n1901 S.n1900 3.643
R3785 S.n1887 S.t544 3.643
R3786 S.n1088 S.t1165 3.643
R3787 S.n1099 S.n1098 3.643
R3788 S.n1096 S.n1095 3.643
R3789 S.n1091 S.t1453 3.643
R3790 S.n1451 S.t2228 3.643
R3791 S.n1471 S.n1470 3.643
R3792 S.n1454 S.n1453 3.643
R3793 S.n1457 S.t230 3.643
R3794 S.n532 S.t597 3.643
R3795 S.n543 S.n542 3.643
R3796 S.n540 S.n539 3.643
R3797 S.n535 S.t854 3.643
R3798 S.n515 S.t1455 3.643
R3799 S.n526 S.n525 3.643
R3800 S.n523 S.n522 3.643
R3801 S.n518 S.t1727 3.643
R3802 S.n138 S.t350 3.643
R3803 S.n130 S.t29 3.643
R3804 S.n235 S.t1563 3.643
R3805 S.n246 S.n245 3.643
R3806 S.n243 S.n242 3.643
R3807 S.n238 S.t2125 3.643
R3808 S.n1368 S.t2178 3.643
R3809 S.n1383 S.n1382 3.643
R3810 S.n1380 S.n1379 3.643
R3811 S.n1365 S.t187 3.643
R3812 S.n1047 S.t1249 3.643
R3813 S.n1028 S.t1518 3.643
R3814 S.n955 S.t2007 3.643
R3815 S.n956 S.t1730 3.643
R3816 S.n255 S.t831 3.643
R3817 S.n266 S.n265 3.643
R3818 S.n263 S.n262 3.643
R3819 S.n258 S.t1398 3.643
R3820 S.n2337 S.t982 3.643
R3821 S.n2317 S.t1245 3.643
R3822 S.n2293 S.t1902 3.643
R3823 S.n2308 S.n2307 3.643
R3824 S.n2311 S.n2310 3.643
R3825 S.n2296 S.t2136 3.643
R3826 S.n1054 S.t367 3.643
R3827 S.n1065 S.n1064 3.643
R3828 S.n1062 S.n1061 3.643
R3829 S.n1057 S.t657 3.643
R3830 S.n1392 S.t1316 3.643
R3831 S.n1412 S.n1411 3.643
R3832 S.n1409 S.n1408 3.643
R3833 S.n1395 S.t1854 3.643
R3834 S.n499 S.t2313 3.643
R3835 S.n510 S.n509 3.643
R3836 S.n507 S.n506 3.643
R3837 S.n502 S.t21 3.643
R3838 S.n482 S.t659 3.643
R3839 S.n493 S.n492 3.643
R3840 S.n490 S.n489 3.643
R3841 S.n485 S.t962 3.643
R3842 S.n125 S.t1831 3.643
R3843 S.n102 S.t2099 3.643
R3844 S.n874 S.t1004 3.643
R3845 S.n740 S.t2289 3.643
R3846 S.n750 S.n749 3.643
R3847 S.n753 S.n752 3.643
R3848 S.n743 S.t2366 3.643
R3849 S.n1349 S.t1099 3.643
R3850 S.n1360 S.n1359 3.643
R3851 S.n1357 S.n1356 3.643
R3852 S.n1352 S.t2348 3.643
R3853 S.n1026 S.t2227 3.643
R3854 S.n1335 S.n1334 3.643
R3855 S.n1338 S.n1337 3.643
R3856 S.n1341 S.t1476 3.643
R3857 S.n2636 S.t1220 3.643
R3858 S.n2648 S.n2647 3.643
R3859 S.n2651 S.n2650 3.643
R3860 S.n2639 S.t64 3.643
R3861 S.n2315 S.t2253 3.643
R3862 S.n2621 S.n2620 3.643
R3863 S.n2624 S.n2623 3.643
R3864 S.n2627 S.t1494 3.643
R3865 S.n3163 S.t2098 3.643
R3866 S.n3175 S.n3174 3.643
R3867 S.n3178 S.n3177 3.643
R3868 S.n3166 S.t108 3.643
R3869 S.n3145 S.t2277 3.643
R3870 S.n3148 S.n3147 3.643
R3871 S.n3151 S.n3150 3.643
R3872 S.n3154 S.t1511 3.643
R3873 S.n3980 S.t2130 3.643
R3874 S.n3992 S.n3991 3.643
R3875 S.n3995 S.n3994 3.643
R3876 S.n3983 S.t145 3.643
R3877 S.n3962 S.t2293 3.643
R3878 S.n3965 S.n3964 3.643
R3879 S.n3968 S.n3967 3.643
R3880 S.n3971 S.t1531 3.643
R3881 S.n4775 S.t2159 3.643
R3882 S.n4787 S.n4786 3.643
R3883 S.n4790 S.n4789 3.643
R3884 S.n4778 S.t179 3.643
R3885 S.n4757 S.t2312 3.643
R3886 S.n4760 S.n4759 3.643
R3887 S.n4763 S.n4762 3.643
R3888 S.n4766 S.t1551 3.643
R3889 S.n5557 S.t2040 3.643
R3890 S.n5569 S.n5568 3.643
R3891 S.n5572 S.n5571 3.643
R3892 S.n5560 S.t5 3.643
R3893 S.n5539 S.t2335 3.643
R3894 S.n5542 S.n5541 3.643
R3895 S.n5545 S.n5544 3.643
R3896 S.n5548 S.t1576 3.643
R3897 S.n6317 S.t2070 3.643
R3898 S.n6329 S.n6328 3.643
R3899 S.n6332 S.n6331 3.643
R3900 S.n6320 S.t70 3.643
R3901 S.n6299 S.t228 3.643
R3902 S.n6302 S.n6301 3.643
R3903 S.n6305 S.n6304 3.643
R3904 S.n6308 S.t1995 3.643
R3905 S.n7064 S.t1598 3.643
R3906 S.n7076 S.n7075 3.643
R3907 S.n7079 S.n7078 3.643
R3908 S.n7067 S.t2176 3.643
R3909 S.n7046 S.t253 3.643
R3910 S.n7049 S.n7048 3.643
R3911 S.n7052 S.n7051 3.643
R3912 S.n7055 S.t2017 3.643
R3913 S.n8075 S.t1623 3.643
R3914 S.n8087 S.n8086 3.643
R3915 S.n8090 S.n8089 3.643
R3916 S.n8078 S.t2205 3.643
R3917 S.n7771 S.t273 3.643
R3918 S.n8060 S.n8059 3.643
R3919 S.n8063 S.n8062 3.643
R3920 S.n8066 S.t2043 3.643
R3921 S.n8787 S.t1437 3.643
R3922 S.n8799 S.n8798 3.643
R3923 S.n8802 S.n8801 3.643
R3924 S.n8790 S.t1958 3.643
R3925 S.n8483 S.t513 3.643
R3926 S.n8772 S.n8771 3.643
R3927 S.n8775 S.n8774 3.643
R3928 S.n8778 S.t651 3.643
R3929 S.n9191 S.t1996 3.643
R3930 S.n9203 S.n9202 3.643
R3931 S.n9206 S.n9205 3.643
R3932 S.n9194 S.t2521 3.643
R3933 S.n9173 S.t975 3.643
R3934 S.n9176 S.n9175 3.643
R3935 S.n9179 S.n9178 3.643
R3936 S.n9182 S.t1238 3.643
R3937 S.n9868 S.t2585 3.643
R3938 S.n9880 S.n9879 3.643
R3939 S.n9883 S.n9882 3.643
R3940 S.n9871 S.t303 3.643
R3941 S.n9850 S.t1524 3.643
R3942 S.n9853 S.n9852 3.643
R3943 S.n9856 S.n9855 3.643
R3944 S.n9859 S.t1834 3.643
R3945 S.n10526 S.t346 3.643
R3946 S.n10538 S.n10537 3.643
R3947 S.n10541 S.n10540 3.643
R3948 S.n10529 S.t893 3.643
R3949 S.n10508 S.t2122 3.643
R3950 S.n10511 S.n10510 3.643
R3951 S.n10514 S.n10513 3.643
R3952 S.n10517 S.t2378 3.643
R3953 S.n11149 S.t960 3.643
R3954 S.n11161 S.n11160 3.643
R3955 S.n11164 S.n11163 3.643
R3956 S.n11152 S.t1478 3.643
R3957 S.n11131 S.t185 3.643
R3958 S.n11134 S.n11133 3.643
R3959 S.n11137 S.n11136 3.643
R3960 S.n11140 S.t471 3.643
R3961 S.n11727 S.t1516 3.643
R3962 S.n11739 S.n11738 3.643
R3963 S.n11742 S.n11741 3.643
R3964 S.n11730 S.t2047 3.643
R3965 S.n12019 S.t737 3.643
R3966 S.n12029 S.n12028 3.643
R3967 S.n12032 S.n12031 3.643
R3968 S.n12022 S.t1063 3.643
R3969 S.n12896 S.t1800 3.643
R3970 S.n12908 S.n12907 3.643
R3971 S.n12911 S.n12910 3.643
R3972 S.n12899 S.t2318 3.643
R3973 S.n12600 S.t232 3.643
R3974 S.n12880 S.n12879 3.643
R3975 S.n12883 S.n12882 3.643
R3976 S.n12886 S.t1376 3.643
R3977 S.n12483 S.t1783 3.643
R3978 S.n1802 S.t139 3.643
R3979 S.n1321 S.t931 3.643
R3980 S.n1329 S.n1328 3.643
R3981 S.n1332 S.n1331 3.643
R3982 S.n1324 S.t1011 3.643
R3983 S.n2659 S.t2250 3.643
R3984 S.n2678 S.n2677 3.643
R3985 S.n2681 S.n2680 3.643
R3986 S.n2656 S.t345 3.643
R3987 S.n12487 S.t911 3.643
R3988 S.n12933 S.t1898 3.643
R3989 S.n12930 S.n12929 3.643
R3990 S.n12927 S.n12926 3.643
R3991 S.n12924 S.t503 3.643
R3992 S.n12919 S.t1067 3.643
R3993 S.n12939 S.n12938 3.643
R3994 S.n12942 S.n12941 3.643
R3995 S.n12916 S.t1555 3.643
R3996 S.n12040 S.t2387 3.643
R3997 S.n12044 S.n12043 3.643
R3998 S.n12047 S.n12046 3.643
R3999 S.n12037 S.t182 3.643
R4000 S.n11750 S.t655 3.643
R4001 S.n11755 S.n11754 3.643
R4002 S.n11758 S.n11757 3.643
R4003 S.n11747 S.t1189 3.643
R4004 S.n11186 S.t1850 3.643
R4005 S.n11183 S.n11182 3.643
R4006 S.n11180 S.n11179 3.643
R4007 S.n11177 S.t2120 3.643
R4008 S.n11172 S.t13 3.643
R4009 S.n11192 S.n11191 3.643
R4010 S.n11195 S.n11194 3.643
R4011 S.n11169 S.t616 3.643
R4012 S.n10563 S.t1255 3.643
R4013 S.n10560 S.n10559 3.643
R4014 S.n10557 S.n10556 3.643
R4015 S.n10554 S.t1522 3.643
R4016 S.n10549 S.t2004 3.643
R4017 S.n10569 S.n10568 3.643
R4018 S.n10572 S.n10571 3.643
R4019 S.n10546 S.t2535 3.643
R4020 S.n9905 S.t663 3.643
R4021 S.n9902 S.n9901 3.643
R4022 S.n9899 S.n9898 3.643
R4023 S.n9896 S.t968 3.643
R4024 S.n9891 S.t1711 3.643
R4025 S.n9911 S.n9910 3.643
R4026 S.n9914 S.n9913 3.643
R4027 S.n9888 S.t1967 3.643
R4028 S.n9228 S.t218 3.643
R4029 S.n9225 S.n9224 3.643
R4030 S.n9222 S.n9221 3.643
R4031 S.n9219 S.t353 3.643
R4032 S.n9214 S.t1145 3.643
R4033 S.n9234 S.n9233 3.643
R4034 S.n9237 S.n9236 3.643
R4035 S.n9211 S.t1643 3.643
R4036 S.n8824 S.t1959 3.643
R4037 S.n8821 S.n8820 3.643
R4038 S.n8818 S.n8817 3.643
R4039 S.n8815 S.t1212 3.643
R4040 S.n8810 S.t787 3.643
R4041 S.n8830 S.n8829 3.643
R4042 S.n8833 S.n8832 3.643
R4043 S.n8807 S.t1369 3.643
R4044 S.n8112 S.t1936 3.643
R4045 S.n8109 S.n8108 3.643
R4046 S.n8106 S.n8105 3.643
R4047 S.n8103 S.t1187 3.643
R4048 S.n8098 S.t758 3.643
R4049 S.n8118 S.n8117 3.643
R4050 S.n8121 S.n8120 3.643
R4051 S.n8095 S.t1346 3.643
R4052 S.n7101 S.t1920 3.643
R4053 S.n7098 S.n7097 3.643
R4054 S.n7095 S.n7094 3.643
R4055 S.n7092 S.t1164 3.643
R4056 S.n7087 S.t735 3.643
R4057 S.n7107 S.n7106 3.643
R4058 S.n7110 S.n7109 3.643
R4059 S.n7084 S.t1312 3.643
R4060 S.n6354 S.t1896 3.643
R4061 S.n6351 S.n6350 3.643
R4062 S.n6348 S.n6347 3.643
R4063 S.n6345 S.t1146 3.643
R4064 S.n6340 S.t1209 3.643
R4065 S.n6360 S.n6359 3.643
R4066 S.n6363 S.n6362 3.643
R4067 S.n6337 S.t1754 3.643
R4068 S.n5594 S.t1477 3.643
R4069 S.n5591 S.n5590 3.643
R4070 S.n5588 S.n5587 3.643
R4071 S.n5585 S.t708 3.643
R4072 S.n5580 S.t1325 3.643
R4073 S.n5600 S.n5599 3.643
R4074 S.n5603 S.n5602 3.643
R4075 S.n5577 S.t1871 3.643
R4076 S.n4812 S.t1454 3.643
R4077 S.n4809 S.n4808 3.643
R4078 S.n4806 S.n4805 3.643
R4079 S.n4803 S.t689 3.643
R4080 S.n4798 S.t1296 3.643
R4081 S.n4818 S.n4817 3.643
R4082 S.n4821 S.n4820 3.643
R4083 S.n4795 S.t1844 3.643
R4084 S.n4020 S.t1438 3.643
R4085 S.n4017 S.n4016 3.643
R4086 S.n4014 S.n4013 3.643
R4087 S.n4011 S.t672 3.643
R4088 S.n4006 S.t1266 3.643
R4089 S.n3998 S.n3997 3.643
R4090 S.n4026 S.n4025 3.643
R4091 S.n4003 S.t1815 3.643
R4092 S.n3498 S.t1421 3.643
R4093 S.n3495 S.n3494 3.643
R4094 S.n3492 S.n3491 3.643
R4095 S.n3191 S.t654 3.643
R4096 S.n3186 S.t1234 3.643
R4097 S.n3504 S.n3503 3.643
R4098 S.n3507 S.n3506 3.643
R4099 S.n3183 S.t1781 3.643
R4100 S.n2673 S.t1394 3.643
R4101 S.n2670 S.n2669 3.643
R4102 S.n2667 S.n2666 3.643
R4103 S.n2664 S.t631 3.643
R4104 S.n1841 S.t158 3.643
R4105 S.n2603 S.t2069 3.643
R4106 S.n2615 S.n2614 3.643
R4107 S.n2618 S.n2617 3.643
R4108 S.n2606 S.t2116 3.643
R4109 S.n3515 S.t241 3.643
R4110 S.n3519 S.n3518 3.643
R4111 S.n3522 S.n3521 3.643
R4112 S.n3512 S.t1507 3.643
R4113 S.n12491 S.t172 3.643
R4114 S.n12677 S.t1038 3.643
R4115 S.n12682 S.n12681 3.643
R4116 S.n12685 S.n12684 3.643
R4117 S.n12674 S.t2149 3.643
R4118 S.n12950 S.t186 3.643
R4119 S.n12954 S.n12953 3.643
R4120 S.n12957 S.n12956 3.643
R4121 S.n12947 S.t693 3.643
R4122 S.n12055 S.t1529 3.643
R4123 S.n12060 S.n12059 3.643
R4124 S.n12063 S.n12062 3.643
R4125 S.n12052 S.t1845 3.643
R4126 S.n11766 S.t2309 3.643
R4127 S.n11770 S.n11769 3.643
R4128 S.n11773 S.n11772 3.643
R4129 S.n11763 S.t313 3.643
R4130 S.n11447 S.t986 3.643
R4131 S.n11452 S.n11451 3.643
R4132 S.n11455 S.n11454 3.643
R4133 S.n11444 S.t1252 3.643
R4134 S.n11203 S.t1723 3.643
R4135 S.n11207 S.n11206 3.643
R4136 S.n11210 S.n11209 3.643
R4137 S.n11200 S.t2272 3.643
R4138 S.n10826 S.t372 3.643
R4139 S.n10831 S.n10830 3.643
R4140 S.n10834 S.n10833 3.643
R4141 S.n10823 S.t661 3.643
R4142 S.n10580 S.t1153 3.643
R4143 S.n10584 S.n10583 3.643
R4144 S.n10587 S.n10586 3.643
R4145 S.n10577 S.t1661 3.643
R4146 S.n10173 S.t2419 3.643
R4147 S.n10178 S.n10177 3.643
R4148 S.n10181 S.n10180 3.643
R4149 S.n10170 S.t31 3.643
R4150 S.n9922 S.t838 3.643
R4151 S.n9926 S.n9925 3.643
R4152 S.n9929 S.n9928 3.643
R4153 S.n9919 S.t1113 3.643
R4154 S.n9497 S.t1126 3.643
R4155 S.n9502 S.n9501 3.643
R4156 S.n9505 S.n9504 3.643
R4157 S.n9494 S.t358 3.643
R4158 S.n9245 S.t2462 3.643
R4159 S.n9249 S.n9248 3.643
R4160 S.n9252 S.n9251 3.643
R4161 S.n9242 S.t525 3.643
R4162 S.n8630 S.t1100 3.643
R4163 S.n8635 S.n8634 3.643
R4164 S.n8638 S.n8637 3.643
R4165 S.n8627 S.t333 3.643
R4166 S.n8841 S.t2438 3.643
R4167 S.n8845 S.n8844 3.643
R4168 S.n8848 S.n8847 3.643
R4169 S.n8838 S.t496 3.643
R4170 S.n7934 S.t1078 3.643
R4171 S.n7939 S.n7938 3.643
R4172 S.n7942 S.n7941 3.643
R4173 S.n7931 S.t312 3.643
R4174 S.n8129 S.t2412 3.643
R4175 S.n8133 S.n8132 3.643
R4176 S.n8136 S.n8135 3.643
R4177 S.n8126 S.t469 3.643
R4178 S.n7381 S.t1060 3.643
R4179 S.n7386 S.n7385 3.643
R4180 S.n7389 S.n7388 3.643
R4181 S.n7378 S.t291 3.643
R4182 S.n7118 S.t2385 3.643
R4183 S.n7122 S.n7121 3.643
R4184 S.n7125 S.n7124 3.643
R4185 S.n7115 S.t435 3.643
R4186 S.n6635 S.t1034 3.643
R4187 S.n6640 S.n6639 3.643
R4188 S.n6643 S.n6642 3.643
R4189 S.n6632 S.t268 3.643
R4190 S.n6371 S.t476 3.643
R4191 S.n6375 S.n6374 3.643
R4192 S.n6378 S.n6377 3.643
R4193 S.n6368 S.t1033 3.643
R4194 S.n5880 S.t615 3.643
R4195 S.n5885 S.n5884 3.643
R4196 S.n5888 S.n5887 3.643
R4197 S.n5877 S.t2365 3.643
R4198 S.n5611 S.t447 3.643
R4199 S.n5615 S.n5614 3.643
R4200 S.n5618 S.n5617 3.643
R4201 S.n5608 S.t1003 3.643
R4202 S.n5099 S.t596 3.643
R4203 S.n5104 S.n5103 3.643
R4204 S.n5107 S.n5106 3.643
R4205 S.n5096 S.t2350 3.643
R4206 S.n4829 S.t412 3.643
R4207 S.n4833 S.n4832 3.643
R4208 S.n4836 S.n4835 3.643
R4209 S.n4826 S.t980 3.643
R4210 S.n4309 S.t575 3.643
R4211 S.n4314 S.n4313 3.643
R4212 S.n4317 S.n4316 3.643
R4213 S.n4306 S.t2329 3.643
R4214 S.n4034 S.t383 3.643
R4215 S.n4038 S.n4037 3.643
R4216 S.n4041 S.n4040 3.643
R4217 S.n4031 S.t948 3.643
R4218 S.n3462 S.t555 3.643
R4219 S.n3466 S.n3465 3.643
R4220 S.n3469 S.n3468 3.643
R4221 S.n3459 S.t2308 3.643
R4222 S.n2724 S.t1855 3.643
R4223 S.n3474 S.t690 3.643
R4224 S.n3486 S.n3485 3.643
R4225 S.n3489 S.n3488 3.643
R4226 S.n3477 S.t692 3.643
R4227 S.n4049 S.t1413 3.643
R4228 S.n4351 S.n4350 3.643
R4229 S.n4354 S.n4353 3.643
R4230 S.n4046 S.t146 3.643
R4231 S.n12495 S.t1835 3.643
R4232 S.n12693 S.t141 3.643
R4233 S.n12698 S.n12697 3.643
R4234 S.n12701 S.n12700 3.643
R4235 S.n12690 S.t1289 3.643
R4236 S.n12965 S.t1853 3.643
R4237 S.n12969 S.n12968 3.643
R4238 S.n12972 S.n12971 3.643
R4239 S.n12962 S.t2353 3.643
R4240 S.n12071 S.t671 3.643
R4241 S.n12076 S.n12075 3.643
R4242 S.n12079 S.n12078 3.643
R4243 S.n12068 S.t983 3.643
R4244 S.n11781 S.t1452 3.643
R4245 S.n11785 S.n11784 3.643
R4246 S.n11788 S.n11787 3.643
R4247 S.n11778 S.t1977 3.643
R4248 S.n11463 S.t66 3.643
R4249 S.n11468 S.n11467 3.643
R4250 S.n11471 S.n11470 3.643
R4251 S.n11460 S.t370 3.643
R4252 S.n11218 S.t851 3.643
R4253 S.n11222 S.n11221 3.643
R4254 S.n11225 S.n11224 3.643
R4255 S.n11215 S.t1416 3.643
R4256 S.n10842 S.t2168 3.643
R4257 S.n10847 S.n10846 3.643
R4258 S.n10850 S.n10849 3.643
R4259 S.n10839 S.t2314 3.643
R4260 S.n10595 S.t277 3.643
R4261 S.n10599 S.n10598 3.643
R4262 S.n10602 S.n10601 3.643
R4263 S.n10592 S.t790 3.643
R4264 S.n10189 S.t270 3.643
R4265 S.n10194 S.n10193 3.643
R4266 S.n10197 S.n10196 3.643
R4267 S.n10186 S.t2037 3.643
R4268 S.n9937 S.t1617 3.643
R4269 S.n9941 S.n9940 3.643
R4270 S.n9944 S.n9943 3.643
R4271 S.n9934 S.t542 3.643
R4272 S.n9513 S.t247 3.643
R4273 S.n9518 S.n9517 3.643
R4274 S.n9521 S.n9520 3.643
R4275 S.n9510 S.t2012 3.643
R4276 S.n9260 S.t1593 3.643
R4277 S.n9264 S.n9263 3.643
R4278 S.n9267 S.n9266 3.643
R4279 S.n9257 S.t2169 3.643
R4280 S.n8646 S.t225 3.643
R4281 S.n8651 S.n8650 3.643
R4282 S.n8654 S.n8653 3.643
R4283 S.n8643 S.t1990 3.643
R4284 S.n8856 S.t1574 3.643
R4285 S.n8860 S.n8859 3.643
R4286 S.n8863 S.n8862 3.643
R4287 S.n8853 S.t2142 3.643
R4288 S.n7950 S.t203 3.643
R4289 S.n7955 S.n7954 3.643
R4290 S.n7958 S.n7957 3.643
R4291 S.n7947 S.t1975 3.643
R4292 S.n8144 S.t1548 3.643
R4293 S.n8148 S.n8147 3.643
R4294 S.n8151 S.n8150 3.643
R4295 S.n8141 S.t2118 3.643
R4296 S.n7397 S.t175 3.643
R4297 S.n7402 S.n7401 3.643
R4298 S.n7405 S.n7404 3.643
R4299 S.n7394 S.t1954 3.643
R4300 S.n7133 S.t1646 3.643
R4301 S.n7137 S.n7136 3.643
R4302 S.n7140 S.n7139 3.643
R4303 S.n7130 S.t2224 3.643
R4304 S.n6651 S.t137 3.643
R4305 S.n6656 S.n6655 3.643
R4306 S.n6659 S.n6658 3.643
R4307 S.n6648 S.t1930 3.643
R4308 S.n6386 S.t2127 3.643
R4309 S.n6390 S.n6389 3.643
R4310 S.n6393 S.n6392 3.643
R4311 S.n6383 S.t136 3.643
R4312 S.n5896 S.t2270 3.643
R4313 S.n5901 S.n5900 3.643
R4314 S.n5904 S.n5903 3.643
R4315 S.n5893 S.t1509 3.643
R4316 S.n5626 S.t2090 3.643
R4317 S.n5630 S.n5629 3.643
R4318 S.n5633 S.n5632 3.643
R4319 S.n5623 S.t99 3.643
R4320 S.n5115 S.t2246 3.643
R4321 S.n5120 S.n5119 3.643
R4322 S.n5123 S.n5122 3.643
R4323 S.n5112 S.t1491 3.643
R4324 S.n4844 S.t2060 3.643
R4325 S.n4848 S.n4847 3.643
R4326 S.n4851 S.n4850 3.643
R4327 S.n4841 S.t54 3.643
R4328 S.n4346 S.t2220 3.643
R4329 S.n4343 S.n4342 3.643
R4330 S.n4340 S.n4339 3.643
R4331 S.n4054 S.t1470 3.643
R4332 S.n3565 S.t1016 3.643
R4333 S.n4322 S.t1881 3.643
R4334 S.n4334 S.n4333 3.643
R4335 S.n4337 S.n4336 3.643
R4336 S.n4325 S.t1852 3.643
R4337 S.n4859 S.t2532 3.643
R4338 S.n5157 S.n5156 3.643
R4339 S.n5160 S.n5159 3.643
R4340 S.n4856 S.t1314 3.643
R4341 S.n12499 S.t969 3.643
R4342 S.n12709 S.t1811 3.643
R4343 S.n12714 S.n12713 3.643
R4344 S.n12717 S.n12716 3.643
R4345 S.n12706 S.t402 3.643
R4346 S.n12980 S.t989 3.643
R4347 S.n12984 S.n12983 3.643
R4348 S.n12987 S.n12986 3.643
R4349 S.n12977 S.t1495 3.643
R4350 S.n12087 S.t2326 3.643
R4351 S.n12092 S.n12091 3.643
R4352 S.n12095 S.n12094 3.643
R4353 S.n12084 S.t58 3.643
R4354 S.n11796 S.t594 3.643
R4355 S.n11800 S.n11799 3.643
R4356 S.n11803 S.n11802 3.643
R4357 S.n11793 S.t1124 3.643
R4358 S.n11479 S.t1894 3.643
R4359 S.n11484 S.n11483 3.643
R4360 S.n11487 S.n11486 3.643
R4361 S.n11476 S.t2021 3.643
R4362 S.n11233 S.t2493 3.643
R4363 S.n11237 S.n11236 3.643
R4364 S.n11240 S.n11239 3.643
R4365 S.n11230 S.t550 3.643
R4366 S.n10858 S.t1956 3.643
R4367 S.n10863 S.n10862 3.643
R4368 S.n10866 S.n10865 3.643
R4369 S.n10855 S.t1206 3.643
R4370 S.n10610 S.t1632 3.643
R4371 S.n10614 S.n10613 3.643
R4372 S.n10617 S.n10616 3.643
R4373 S.n10607 S.t2215 3.643
R4374 S.n10205 S.t1931 3.643
R4375 S.n10210 S.n10209 3.643
R4376 S.n10213 S.n10212 3.643
R4377 S.n10202 S.t1182 3.643
R4378 S.n9952 S.t751 3.643
R4379 S.n9956 S.n9955 3.643
R4380 S.n9959 S.n9958 3.643
R4381 S.n9949 S.t2187 3.643
R4382 S.n9529 S.t1914 3.643
R4383 S.n9534 S.n9533 3.643
R4384 S.n9537 S.n9536 3.643
R4385 S.n9526 S.t1160 3.643
R4386 S.n9275 S.t730 3.643
R4387 S.n9279 S.n9278 3.643
R4388 S.n9282 S.n9281 3.643
R4389 S.n9272 S.t1306 3.643
R4390 S.n8662 S.t1892 3.643
R4391 S.n8667 S.n8666 3.643
R4392 S.n8670 S.n8669 3.643
R4393 S.n8659 S.t1140 3.643
R4394 S.n8871 S.t704 3.643
R4395 S.n8875 S.n8874 3.643
R4396 S.n8878 S.n8877 3.643
R4397 S.n8868 S.t1280 3.643
R4398 S.n7966 S.t1870 3.643
R4399 S.n7971 S.n7970 3.643
R4400 S.n7974 S.n7973 3.643
R4401 S.n7963 S.t1120 3.643
R4402 S.n8159 S.t808 3.643
R4403 S.n8163 S.n8162 3.643
R4404 S.n8166 S.n8165 3.643
R4405 S.n8156 S.t1392 3.643
R4406 S.n7413 S.t1839 3.643
R4407 S.n7418 S.n7417 3.643
R4408 S.n7421 S.n7420 3.643
R4409 S.n7410 S.t1094 3.643
R4410 S.n7148 S.t777 3.643
R4411 S.n7152 S.n7151 3.643
R4412 S.n7155 S.n7154 3.643
R4413 S.n7145 S.t1362 3.643
R4414 S.n6667 S.t1808 3.643
R4415 S.n6672 S.n6671 3.643
R4416 S.n6675 S.n6674 3.643
R4417 S.n6664 S.t1071 3.643
R4418 S.n6401 S.t1261 3.643
R4419 S.n6405 S.n6404 3.643
R4420 S.n6408 S.n6407 3.643
R4421 S.n6398 S.t1806 3.643
R4422 S.n5912 S.t1414 3.643
R4423 S.n5917 S.n5916 3.643
R4424 S.n5920 S.n5919 3.643
R4425 S.n5909 S.t649 3.643
R4426 S.n5641 S.t1228 3.643
R4427 S.n5645 S.n5644 3.643
R4428 S.n5648 S.n5647 3.643
R4429 S.n5638 S.t1776 3.643
R4430 S.n5152 S.t1387 3.643
R4431 S.n5149 S.n5148 3.643
R4432 S.n5146 S.n5145 3.643
R4433 S.n4864 S.t628 3.643
R4434 S.n4397 S.t152 3.643
R4435 S.n5128 S.t511 3.643
R4436 S.n5140 S.n5139 3.643
R4437 S.n5143 S.n5142 3.643
R4438 S.n5131 S.t436 3.643
R4439 S.n5656 S.t1179 3.643
R4440 S.n5954 S.n5953 3.643
R4441 S.n5957 S.n5956 3.643
R4442 S.n5653 S.t2426 3.643
R4443 S.n12503 S.t36 3.643
R4444 S.n12725 S.t944 3.643
R4445 S.n12730 S.n12729 3.643
R4446 S.n12733 S.n12732 3.643
R4447 S.n12722 S.t2051 3.643
R4448 S.n12995 S.t73 3.643
R4449 S.n12999 S.n12998 3.643
R4450 S.n13002 S.n13001 3.643
R4451 S.n12992 S.t632 3.643
R4452 S.n12103 S.t1564 3.643
R4453 S.n12108 S.n12107 3.643
R4454 S.n12111 S.n12110 3.643
R4455 S.n12100 S.t1748 3.643
R4456 S.n11811 S.t2241 3.643
R4457 S.n11815 S.n11814 3.643
R4458 S.n11818 S.n11817 3.643
R4459 S.n11808 S.t245 3.643
R4460 S.n11495 S.t1123 3.643
R4461 S.n11500 S.n11499 3.643
R4462 S.n11503 S.n11502 3.643
R4463 S.n11492 S.t352 3.643
R4464 S.n11248 S.t796 3.643
R4465 S.n11252 S.n11251 3.643
R4466 S.n11255 S.n11254 3.643
R4467 S.n11245 S.t1382 3.643
R4468 S.n10874 S.t1098 3.643
R4469 S.n10879 S.n10878 3.643
R4470 S.n10882 S.n10881 3.643
R4471 S.n10871 S.t328 3.643
R4472 S.n10625 S.t765 3.643
R4473 S.n10629 S.n10628 3.643
R4474 S.n10632 S.n10631 3.643
R4475 S.n10622 S.t1354 3.643
R4476 S.n10221 S.t1073 3.643
R4477 S.n10226 S.n10225 3.643
R4478 S.n10229 S.n10228 3.643
R4479 S.n10218 S.t306 3.643
R4480 S.n9967 S.t2407 3.643
R4481 S.n9971 S.n9970 3.643
R4482 S.n9974 S.n9973 3.643
R4483 S.n9964 S.t1322 3.643
R4484 S.n9545 S.t1054 3.643
R4485 S.n9550 S.n9549 3.643
R4486 S.n9553 S.n9552 3.643
R4487 S.n9542 S.t288 3.643
R4488 S.n9290 S.t2383 3.643
R4489 S.n9294 S.n9293 3.643
R4490 S.n9297 S.n9296 3.643
R4491 S.n9287 S.t424 3.643
R4492 S.n8678 S.t1031 3.643
R4493 S.n8683 S.n8682 3.643
R4494 S.n8686 S.n8685 3.643
R4495 S.n8675 S.t265 3.643
R4496 S.n8886 S.t2486 3.643
R4497 S.n8890 S.n8889 3.643
R4498 S.n8893 S.n8892 3.643
R4499 S.n8883 S.t552 3.643
R4500 S.n7982 S.t1001 3.643
R4501 S.n7987 S.n7986 3.643
R4502 S.n7990 S.n7989 3.643
R4503 S.n7979 S.t243 3.643
R4504 S.n8174 S.t2458 3.643
R4505 S.n8178 S.n8177 3.643
R4506 S.n8181 S.n8180 3.643
R4507 S.n8171 S.t520 3.643
R4508 S.n7429 S.t974 3.643
R4509 S.n7434 S.n7433 3.643
R4510 S.n7437 S.n7436 3.643
R4511 S.n7426 S.t220 3.643
R4512 S.n7163 S.t2429 3.643
R4513 S.n7167 S.n7166 3.643
R4514 S.n7170 S.n7169 3.643
R4515 S.n7160 S.t489 3.643
R4516 S.n6683 S.t942 3.643
R4517 S.n6688 S.n6687 3.643
R4518 S.n6691 S.n6690 3.643
R4519 S.n6680 S.t192 3.643
R4520 S.n6416 S.t378 3.643
R4521 S.n6420 S.n6419 3.643
R4522 S.n6423 S.n6422 3.643
R4523 S.n6413 S.t941 3.643
R4524 S.n5949 S.t549 3.643
R4525 S.n5946 S.n5945 3.643
R4526 S.n5943 S.n5942 3.643
R4527 S.n5661 S.t2305 3.643
R4528 S.n5203 S.t1849 3.643
R4529 S.n5925 S.t1622 3.643
R4530 S.n5937 S.n5936 3.643
R4531 S.n5940 S.n5939 3.643
R4532 S.n5928 S.t1537 3.643
R4533 S.n6431 S.t2328 3.643
R4534 S.n6725 S.n6724 3.643
R4535 S.n6728 S.n6727 3.643
R4536 S.n6428 S.t1101 3.643
R4537 S.n12507 S.t1733 3.643
R4538 S.n12741 S.t193 3.643
R4539 S.n12746 S.n12745 3.643
R4540 S.n12749 S.n12748 3.643
R4541 S.n12738 S.t1191 3.643
R4542 S.n13010 S.t1753 3.643
R4543 S.n13014 S.n13013 3.643
R4544 S.n13017 S.n13016 3.643
R4545 S.n13007 S.t2287 3.643
R4546 S.n12119 S.t266 3.643
R4547 S.n12124 S.n12123 3.643
R4548 S.n12127 S.n12126 3.643
R4549 S.n12116 S.t2034 3.643
R4550 S.n11826 S.t2472 3.643
R4551 S.n11830 S.n11829 3.643
R4552 S.n11833 S.n11832 3.643
R4553 S.n11823 S.t538 3.643
R4554 S.n11511 S.t246 3.643
R4555 S.n11516 S.n11515 3.643
R4556 S.n11519 S.n11518 3.643
R4557 S.n11508 S.t2009 3.643
R4558 S.n11263 S.t2447 3.643
R4559 S.n11267 S.n11266 3.643
R4560 S.n11270 S.n11269 3.643
R4561 S.n11260 S.t507 3.643
R4562 S.n10890 S.t223 3.643
R4563 S.n10895 S.n10894 3.643
R4564 S.n10898 S.n10897 3.643
R4565 S.n10887 S.t1987 3.643
R4566 S.n10640 S.t2418 3.643
R4567 S.n10644 S.n10643 3.643
R4568 S.n10647 S.n10646 3.643
R4569 S.n10637 S.t474 3.643
R4570 S.n10237 S.t196 3.643
R4571 S.n10242 S.n10241 3.643
R4572 S.n10245 S.n10244 3.643
R4573 S.n10234 S.t1969 3.643
R4574 S.n9982 S.t1545 3.643
R4575 S.n9986 S.n9985 3.643
R4576 S.n9989 S.n9988 3.643
R4577 S.n9979 S.t442 3.643
R4578 S.n9561 S.t167 3.643
R4579 S.n9566 S.n9565 3.643
R4580 S.n9569 S.n9568 3.643
R4581 S.n9558 S.t1949 3.643
R4582 S.n9305 S.t1641 3.643
R4583 S.n9309 S.n9308 3.643
R4584 S.n9312 S.n9311 3.643
R4585 S.n9302 S.t2218 3.643
R4586 S.n8694 S.t134 3.643
R4587 S.n8699 S.n8698 3.643
R4588 S.n8702 S.n8701 3.643
R4589 S.n8691 S.t1928 3.643
R4590 S.n8901 S.t1614 3.643
R4591 S.n8905 S.n8904 3.643
R4592 S.n8908 S.n8907 3.643
R4593 S.n8898 S.t2191 3.643
R4594 S.n7998 S.t96 3.643
R4595 S.n8003 S.n8002 3.643
R4596 S.n8006 S.n8005 3.643
R4597 S.n7995 S.t1909 3.643
R4598 S.n8189 S.t1590 3.643
R4599 S.n8193 S.n8192 3.643
R4600 S.n8196 S.n8195 3.643
R4601 S.n8186 S.t2165 3.643
R4602 S.n7445 S.t41 3.643
R4603 S.n7450 S.n7449 3.643
R4604 S.n7453 S.n7452 3.643
R4605 S.n7442 S.t1884 3.643
R4606 S.n7178 S.t1565 3.643
R4607 S.n7182 S.n7181 3.643
R4608 S.n7185 S.n7184 3.643
R4609 S.n7175 S.t2134 3.643
R4610 S.n6720 S.t2581 3.643
R4611 S.n6717 S.n6716 3.643
R4612 S.n6714 S.n6713 3.643
R4613 S.n6436 S.t1861 3.643
R4614 S.n6000 S.t1014 3.643
R4615 S.n6696 S.t2102 3.643
R4616 S.n6708 S.n6707 3.643
R4617 S.n6711 S.n6710 3.643
R4618 S.n6699 S.t1050 3.643
R4619 S.n7193 S.t898 3.643
R4620 S.n7487 S.n7486 3.643
R4621 S.n7490 S.n7489 3.643
R4622 S.n7190 S.t2183 3.643
R4623 S.n12511 S.t859 3.643
R4624 S.n12757 S.t1889 3.643
R4625 S.n12762 S.n12761 3.643
R4626 S.n12765 S.n12764 3.643
R4627 S.n12754 S.t224 3.643
R4628 S.n13025 S.t707 3.643
R4629 S.n13029 S.n13028 3.643
R4630 S.n13032 S.n13031 3.643
R4631 S.n13022 S.t1285 3.643
R4632 S.n12135 S.t1929 3.643
R4633 S.n12140 S.n12139 3.643
R4634 S.n12143 S.n12142 3.643
R4635 S.n12132 S.t1178 3.643
R4636 S.n11841 S.t1602 3.643
R4637 S.n11845 S.n11844 3.643
R4638 S.n11848 S.n11847 3.643
R4639 S.n11838 S.t2179 3.643
R4640 S.n11527 S.t1911 3.643
R4641 S.n11532 S.n11531 3.643
R4642 S.n11535 S.n11534 3.643
R4643 S.n11524 S.t1157 3.643
R4644 S.n11278 S.t1578 3.643
R4645 S.n11282 S.n11281 3.643
R4646 S.n11285 S.n11284 3.643
R4647 S.n11275 S.t2152 3.643
R4648 S.n10906 S.t1888 3.643
R4649 S.n10911 S.n10910 3.643
R4650 S.n10914 S.n10913 3.643
R4651 S.n10903 S.t1137 3.643
R4652 S.n10655 S.t1553 3.643
R4653 S.n10659 S.n10658 3.643
R4654 S.n10662 S.n10661 3.643
R4655 S.n10652 S.t2124 3.643
R4656 S.n10253 S.t1864 3.643
R4657 S.n10258 S.n10257 3.643
R4658 S.n10261 S.n10260 3.643
R4659 S.n10250 S.t1114 3.643
R4660 S.n9997 S.t806 3.643
R4661 S.n10001 S.n10000 3.643
R4662 S.n10004 S.n10003 3.643
R4663 S.n9994 S.t2233 3.643
R4664 S.n9577 S.t1830 3.643
R4665 S.n9582 S.n9581 3.643
R4666 S.n9585 S.n9584 3.643
R4667 S.n9574 S.t1091 3.643
R4668 S.n9320 S.t773 3.643
R4669 S.n9324 S.n9323 3.643
R4670 S.n9327 S.n9326 3.643
R4671 S.n9317 S.t1358 3.643
R4672 S.n8710 S.t1803 3.643
R4673 S.n8715 S.n8714 3.643
R4674 S.n8718 S.n8717 3.643
R4675 S.n8707 S.t1068 3.643
R4676 S.n8916 S.t749 3.643
R4677 S.n8920 S.n8919 3.643
R4678 S.n8923 S.n8922 3.643
R4679 S.n8913 S.t1334 3.643
R4680 S.n8014 S.t1772 3.643
R4681 S.n8019 S.n8018 3.643
R4682 S.n8022 S.n8021 3.643
R4683 S.n8011 S.t1049 3.643
R4684 S.n8204 S.t726 3.643
R4685 S.n8208 S.n8207 3.643
R4686 S.n8211 S.n8210 3.643
R4687 S.n8201 S.t1300 3.643
R4688 S.n7482 S.t1736 3.643
R4689 S.n7479 S.n7478 3.643
R4690 S.n7476 S.n7475 3.643
R4691 S.n7198 S.t1022 3.643
R4692 S.n6771 S.t2204 3.643
R4693 S.n7458 S.t711 3.643
R4694 S.n7470 S.n7469 3.643
R4695 S.n7473 S.n7472 3.643
R4696 S.n7461 S.t2153 3.643
R4697 S.n8219 S.t2042 3.643
R4698 S.n8223 S.n8222 3.643
R4699 S.n8226 S.n8225 3.643
R4700 S.n8216 S.t782 3.643
R4701 S.n12515 S.t1480 3.643
R4702 S.n12773 S.t1027 3.643
R4703 S.n12778 S.n12777 3.643
R4704 S.n12781 S.n12780 3.643
R4705 S.n12770 S.t1891 3.643
R4706 S.n13040 S.t2364 3.643
R4707 S.n13044 S.n13043 3.643
R4708 S.n13047 S.n13046 3.643
R4709 S.n13037 S.t397 3.643
R4710 S.n12151 S.t1070 3.643
R4711 S.n12156 S.n12155 3.643
R4712 S.n12159 S.n12158 3.643
R4713 S.n12148 S.t301 3.643
R4714 S.n11856 S.t738 3.643
R4715 S.n11860 S.n11859 3.643
R4716 S.n11863 S.n11862 3.643
R4717 S.n11853 S.t1318 3.643
R4718 S.n11543 S.t1052 3.643
R4719 S.n11548 S.n11547 3.643
R4720 S.n11551 S.n11550 3.643
R4721 S.n11540 S.t283 3.643
R4722 S.n11293 S.t710 3.643
R4723 S.n11297 S.n11296 3.643
R4724 S.n11300 S.n11299 3.643
R4725 S.n11290 S.t1292 3.643
R4726 S.n10922 S.t1026 3.643
R4727 S.n10927 S.n10926 3.643
R4728 S.n10930 S.n10929 3.643
R4729 S.n10919 S.t259 3.643
R4730 S.n10670 S.t817 3.643
R4731 S.n10674 S.n10673 3.643
R4732 S.n10677 S.n10676 3.643
R4733 S.n10667 S.t1400 3.643
R4734 S.n10269 S.t995 3.643
R4735 S.n10274 S.n10273 3.643
R4736 S.n10277 S.n10276 3.643
R4737 S.n10266 S.t236 3.643
R4738 S.n10012 S.t2455 3.643
R4739 S.n10016 S.n10015 3.643
R4740 S.n10019 S.n10018 3.643
R4741 S.n10009 S.t1371 3.643
R4742 S.n9593 S.t964 3.643
R4743 S.n9598 S.n9597 3.643
R4744 S.n9601 S.n9600 3.643
R4745 S.n9590 S.t213 3.643
R4746 S.n9335 S.t2424 3.643
R4747 S.n9339 S.n9338 3.643
R4748 S.n9342 S.n9341 3.643
R4749 S.n9332 S.t484 3.643
R4750 S.n8726 S.t935 3.643
R4751 S.n8731 S.n8730 3.643
R4752 S.n8734 S.n8733 3.643
R4753 S.n8723 S.t189 3.643
R4754 S.n8931 S.t2401 3.643
R4755 S.n8935 S.n8934 3.643
R4756 S.n8938 S.n8937 3.643
R4757 S.n8928 S.t454 3.643
R4758 S.n8030 S.t900 3.643
R4759 S.n8034 S.n8033 3.643
R4760 S.n8037 S.n8036 3.643
R4761 S.n8027 S.t159 3.643
R4762 S.n7533 S.t1368 3.643
R4763 S.n8042 S.t1907 3.643
R4764 S.n8054 S.n8053 3.643
R4765 S.n8057 S.n8056 3.643
R4766 S.n8045 S.t725 3.643
R4767 S.n8946 S.t674 3.643
R4768 S.n8950 S.n8949 3.643
R4769 S.n8953 S.n8952 3.643
R4770 S.n8943 S.t1963 3.643
R4771 S.n12519 S.t618 3.643
R4772 S.n12789 S.t127 3.643
R4773 S.n12794 S.n12793 3.643
R4774 S.n12797 S.n12796 3.643
R4775 S.n12786 S.t1028 3.643
R4776 S.n13055 S.t1508 3.643
R4777 S.n13059 S.n13058 3.643
R4778 S.n13062 S.n13061 3.643
R4779 S.n13052 S.t2049 3.643
R4780 S.n12167 S.t191 3.643
R4781 S.n12172 S.n12171 3.643
R4782 S.n12175 S.n12174 3.643
R4783 S.n12164 S.t1966 3.643
R4784 S.n11871 S.t2388 3.643
R4785 S.n11875 S.n11874 3.643
R4786 S.n11878 S.n11877 3.643
R4787 S.n11868 S.t440 3.643
R4788 S.n11559 S.t164 3.643
R4789 S.n11564 S.n11563 3.643
R4790 S.n11567 S.n11566 3.643
R4791 S.n11556 S.t1944 3.643
R4792 S.n11308 S.t2496 3.643
R4793 S.n11312 S.n11311 3.643
R4794 S.n11315 S.n11314 3.643
R4795 S.n11305 S.t562 3.643
R4796 S.n10938 S.t123 3.643
R4797 S.n10943 S.n10942 3.643
R4798 S.n10946 S.n10945 3.643
R4799 S.n10935 S.t1925 3.643
R4800 S.n10685 S.t2464 3.643
R4801 S.n10689 S.n10688 3.643
R4802 S.n10692 S.n10691 3.643
R4803 S.n10682 S.t529 3.643
R4804 S.n10285 S.t88 3.643
R4805 S.n10290 S.n10289 3.643
R4806 S.n10293 S.n10292 3.643
R4807 S.n10282 S.t1903 3.643
R4808 S.n10027 S.t1586 3.643
R4809 S.n10031 S.n10030 3.643
R4810 S.n10034 S.n10033 3.643
R4811 S.n10024 S.t498 3.643
R4812 S.n9609 S.t27 3.643
R4813 S.n9614 S.n9613 3.643
R4814 S.n9617 S.n9616 3.643
R4815 S.n9606 S.t1880 3.643
R4816 S.n9350 S.t1559 3.643
R4817 S.n9354 S.n9353 3.643
R4818 S.n9357 S.n9356 3.643
R4819 S.n9347 S.t2131 3.643
R4820 S.n8742 S.t2577 3.643
R4821 S.n8746 S.n8745 3.643
R4822 S.n8749 S.n8748 3.643
R4823 S.n8739 S.t1856 3.643
R4824 S.n8269 S.t524 3.643
R4825 S.n8754 S.t548 3.643
R4826 S.n8766 S.n8765 3.643
R4827 S.n8769 S.n8768 3.643
R4828 S.n8757 S.t1890 3.643
R4829 S.n9365 S.t1860 3.643
R4830 S.n9651 S.n9650 3.643
R4831 S.n9654 S.n9653 3.643
R4832 S.n9362 S.t607 3.643
R4833 S.n12523 S.t2274 3.643
R4834 S.n12805 S.t1798 3.643
R4835 S.n12810 S.n12809 3.643
R4836 S.n12813 S.n12812 3.643
R4837 S.n12802 S.t129 3.643
R4838 S.n13070 S.t648 3.643
R4839 S.n13074 S.n13073 3.643
R4840 S.n13077 S.n13076 3.643
R4841 S.n13067 S.t1190 3.643
R4842 S.n12183 S.t1859 3.643
R4843 S.n12188 S.n12187 3.643
R4844 S.n12191 S.n12190 3.643
R4845 S.n12180 S.t1112 3.643
R4846 S.n11886 S.t1653 3.643
R4847 S.n11890 S.n11889 3.643
R4848 S.n11893 S.n11892 3.643
R4849 S.n11883 S.t2231 3.643
R4850 S.n11575 S.t1827 3.643
R4851 S.n11580 S.n11579 3.643
R4852 S.n11583 S.n11582 3.643
R4853 S.n11572 S.t1087 3.643
R4854 S.n11323 S.t1619 3.643
R4855 S.n11327 S.n11326 3.643
R4856 S.n11330 S.n11329 3.643
R4857 S.n11320 S.t2201 3.643
R4858 S.n10954 S.t1793 3.643
R4859 S.n10959 S.n10958 3.643
R4860 S.n10962 S.n10961 3.643
R4861 S.n10951 S.t1065 3.643
R4862 S.n10700 S.t1594 3.643
R4863 S.n10704 S.n10703 3.643
R4864 S.n10707 S.n10706 3.643
R4865 S.n10697 S.t2171 3.643
R4866 S.n10301 S.t1766 3.643
R4867 S.n10306 S.n10305 3.643
R4868 S.n10309 S.n10308 3.643
R4869 S.n10298 S.t1044 3.643
R4870 S.n10042 S.t721 3.643
R4871 S.n10046 S.n10045 3.643
R4872 S.n10049 S.n10048 3.643
R4873 S.n10039 S.t2144 3.643
R4874 S.n9646 S.t1732 3.643
R4875 S.n9643 S.n9642 3.643
R4876 S.n9640 S.n9639 3.643
R4877 S.n9370 S.t1018 3.643
R4878 S.n8996 S.t2197 3.643
R4879 S.n9622 S.t1659 3.643
R4880 S.n9634 S.n9633 3.643
R4881 S.n9637 S.n9636 3.643
R4882 S.n9625 S.t480 3.643
R4883 S.n10057 S.t485 3.643
R4884 S.n10343 S.n10342 3.643
R4885 S.n10346 S.n10345 3.643
R4886 S.n10054 S.t1130 3.643
R4887 S.n12527 S.t1418 3.643
R4888 S.n12821 S.t928 3.643
R4889 S.n12826 S.n12825 3.643
R4890 S.n12829 S.n12828 3.643
R4891 S.n12818 S.t1799 3.643
R4892 S.n13085 S.t2405 3.643
R4893 S.n13089 S.n13088 3.643
R4894 S.n13092 S.n13091 3.643
R4895 S.n13082 S.t456 3.643
R4896 S.n12199 S.t992 3.643
R4897 S.n12204 S.n12203 3.643
R4898 S.n12207 S.n12206 3.643
R4899 S.n12196 S.t234 3.643
R4900 S.n11901 S.t781 3.643
R4901 S.n11905 S.n11904 3.643
R4902 S.n11908 S.n11907 3.643
R4903 S.n11898 S.t1367 3.643
R4904 S.n11591 S.t959 3.643
R4905 S.n11596 S.n11595 3.643
R4906 S.n11599 S.n11598 3.643
R4907 S.n11588 S.t209 3.643
R4908 S.n11338 S.t752 3.643
R4909 S.n11342 S.n11341 3.643
R4910 S.n11345 S.n11344 3.643
R4911 S.n11335 S.t1344 3.643
R4912 S.n10970 S.t926 3.643
R4913 S.n10975 S.n10974 3.643
R4914 S.n10978 S.n10977 3.643
R4915 S.n10967 S.t184 3.643
R4916 S.n10715 S.t731 3.643
R4917 S.n10719 S.n10718 3.643
R4918 S.n10722 S.n10721 3.643
R4919 S.n10712 S.t1307 3.643
R4920 S.n10338 S.t892 3.643
R4921 S.n10335 S.n10334 3.643
R4922 S.n10332 S.n10331 3.643
R4923 S.n10062 S.t151 3.643
R4924 S.n9697 S.t2212 3.643
R4925 S.n10314 S.t302 3.643
R4926 S.n10326 S.n10325 3.643
R4927 S.n10329 S.n10328 3.643
R4928 S.n10317 S.t1568 3.643
R4929 S.n10730 S.t1017 3.643
R4930 S.n11012 S.n11011 3.643
R4931 S.n11015 S.n11014 3.643
R4932 S.n10727 S.t2281 3.643
R4933 S.n12531 S.t652 3.643
R4934 S.n12837 S.t2569 3.643
R4935 S.n12842 S.n12841 3.643
R4936 S.n12845 S.n12844 3.643
R4937 S.n12834 S.t929 3.643
R4938 S.n13100 S.t1543 3.643
R4939 S.n13104 S.n13103 3.643
R4940 S.n13107 S.n13106 3.643
R4941 S.n13097 S.t2101 3.643
R4942 S.n12215 S.t83 3.643
R4943 S.n12220 S.n12219 3.643
R4944 S.n12223 S.n12222 3.643
R4945 S.n12212 S.t1900 3.643
R4946 S.n11916 S.t2432 3.643
R4947 S.n11920 S.n11919 3.643
R4948 S.n11923 S.n11922 3.643
R4949 S.n11913 S.t495 3.643
R4950 S.n11607 S.t19 3.643
R4951 S.n11612 S.n11611 3.643
R4952 S.n11615 S.n11614 3.643
R4953 S.n11604 S.t1877 3.643
R4954 S.n11353 S.t2408 3.643
R4955 S.n11357 S.n11356 3.643
R4956 S.n11360 S.n11359 3.643
R4957 S.n11350 S.t465 3.643
R4958 S.n11007 S.t2566 3.643
R4959 S.n11004 S.n11003 3.643
R4960 S.n11001 S.n11000 3.643
R4961 S.n10735 S.t1848 3.643
R4962 S.n10389 S.t1377 3.643
R4963 S.n10983 S.t1469 3.643
R4964 S.n10995 S.n10994 3.643
R4965 S.n10998 S.n10997 3.643
R4966 S.n10986 S.t199 3.643
R4967 S.n11368 S.t2155 3.643
R4968 S.n11652 S.n11651 3.643
R4969 S.n11655 S.n11654 3.643
R4970 S.n11365 S.t906 3.643
R4971 S.n12535 S.t2306 3.643
R4972 S.n12853 S.t1693 3.643
R4973 S.n12858 S.n12857 3.643
R4974 S.n12861 S.n12860 3.643
R4975 S.n12850 S.t2572 3.643
R4976 S.n13115 S.t682 3.643
R4977 S.n13119 S.n13118 3.643
R4978 S.n13122 S.n13121 3.643
R4979 S.n13112 S.t1236 3.643
R4980 S.n12231 S.t1762 3.643
R4981 S.n12236 S.n12235 3.643
R4982 S.n12239 S.n12238 3.643
R4983 S.n12228 S.t1041 3.643
R4984 S.n11931 S.t1569 3.643
R4985 S.n11935 S.n11934 3.643
R4986 S.n11938 S.n11937 3.643
R4987 S.n11928 S.t2141 3.643
R4988 S.n11647 S.t1726 3.643
R4989 S.n11644 S.n11643 3.643
R4990 S.n11641 S.n11640 3.643
R4991 S.n11373 S.t1012 3.643
R4992 S.n11048 S.t535 3.643
R4993 S.n11618 S.t71 3.643
R4994 S.n11635 S.n11634 3.643
R4995 S.n11638 S.n11637 3.643
R4996 S.n11621 S.t1335 3.643
R4997 S.n12258 S.t753 3.643
R4998 S.n12267 S.n12266 3.643
R4999 S.n12270 S.n12269 3.643
R5000 S.n12261 S.t2046 3.643
R5001 S.n12539 S.t1450 3.643
R5002 S.n12866 S.t823 3.643
R5003 S.n12874 S.n12873 3.643
R5004 S.n12877 S.n12876 3.643
R5005 S.n12869 S.t1697 3.643
R5006 S.n13129 S.t2341 3.643
R5007 S.n13137 S.n13136 3.643
R5008 S.n13140 S.n13139 3.643
R5009 S.n13132 S.t356 3.643
R5010 S.n11947 S.t885 3.643
R5011 S.n12242 S.n12241 3.643
R5012 S.n12245 S.n12244 3.643
R5013 S.n12248 S.t149 3.643
R5014 S.n12475 S.t2392 3.643
R5015 S.n12657 S.t2336 3.643
R5016 S.n12668 S.n12667 3.643
R5017 S.n12665 S.n12664 3.643
R5018 S.n12660 S.t818 3.643
R5019 S.n13147 S.t427 3.643
R5020 S.n1021 S.t169 3.643
R5021 S.n1023 S.n1022 3.643
R5022 S.n467 S.n465 2.799
R5023 S.n1037 S.n1035 2.799
R5024 S.n2328 S.n2326 2.799
R5025 S.n3202 S.n3200 2.799
R5026 S.n4067 S.n4065 2.799
R5027 S.n4875 S.n4873 2.799
R5028 S.n5674 S.n5672 2.799
R5029 S.n6447 S.n6445 2.799
R5030 S.n7211 S.n7209 2.799
R5031 S.n7782 S.n7780 2.799
R5032 S.n8496 S.n8494 2.799
R5033 S.n9381 S.n9379 2.799
R5034 S.n10075 S.n10073 2.799
R5035 S.n10746 S.n10744 2.799
R5036 S.n11389 S.n11387 2.799
R5037 S.n11960 S.n11958 2.799
R5038 S.n12612 S.n12610 2.799
R5039 S.n106 S.n105 2.645
R5040 S.n461 S.n460 2.645
R5041 S.n1031 S.n1030 2.645
R5042 S.n2322 S.n2321 2.645
R5043 S.n3196 S.n3195 2.645
R5044 S.n4061 S.n4060 2.645
R5045 S.n4869 S.n4868 2.645
R5046 S.n5668 S.n5667 2.645
R5047 S.n6441 S.n6440 2.645
R5048 S.n7205 S.n7204 2.645
R5049 S.n7776 S.n7775 2.645
R5050 S.n8490 S.n8489 2.645
R5051 S.n9375 S.n9374 2.645
R5052 S.n10069 S.n10068 2.645
R5053 S.n10740 S.n10739 2.645
R5054 S.n11383 S.n11382 2.645
R5055 S.n11954 S.n11953 2.645
R5056 S.n11029 S.n11028 0.21
R5057 S.n12314 S.n12311 0.178
R5058 S.n871 S.n870 0.172
R5059 S.n108 S.n104 0.164
R5060 S.n13162 S.n12549 0.141
R5061 S.n2240 S.n2239 0.133
R5062 S.n96 S.n94 0.123
R5063 S.n29 S.n27 0.123
R5064 S.n61 S.n39 0.123
R5065 S.n73 S.n71 0.123
R5066 S.n85 S.n83 0.123
R5067 S.n985 S.n977 0.123
R5068 S.n172 S.n171 0.123
R5069 S.n159 S.n158 0.123
R5070 S.n146 S.n145 0.123
R5071 S.n133 S.n132 0.123
R5072 S.n13177 S.n1809 0.116
R5073 S.n13176 S.n2692 0.111
R5074 S.n13175 S.n3533 0.111
R5075 S.n13174 S.n4365 0.111
R5076 S.n13173 S.n5171 0.111
R5077 S.n13172 S.n5968 0.111
R5078 S.n13171 S.n6739 0.111
R5079 S.n13170 S.n7501 0.111
R5080 S.n13169 S.n8237 0.111
R5081 S.n13168 S.n8964 0.111
R5082 S.n13167 S.n9665 0.111
R5083 S.n13166 S.n10357 0.111
R5084 S.n13165 S.n11026 0.111
R5085 S.n13164 S.n11666 0.111
R5086 S.n12391 S.n12390 0.11
R5087 S.n13162 S.n13161 0.11
R5088 S.n13163 S.n12306 0.11
R5089 S.n11413 S.n11411 0.109
R5090 S.n10792 S.n10790 0.109
R5091 S.n10139 S.n10137 0.109
R5092 S.n9463 S.n9461 0.109
R5093 S.n8596 S.n8594 0.109
R5094 S.n7900 S.n7898 0.109
R5095 S.n7347 S.n7345 0.109
R5096 S.n6601 S.n6599 0.109
R5097 S.n5846 S.n5844 0.109
R5098 S.n5065 S.n5063 0.109
R5099 S.n4275 S.n4273 0.109
R5100 S.n3428 S.n3426 0.109
R5101 S.n2572 S.n2570 0.109
R5102 S.n747 S.n746 0.109
R5103 S.n2611 S.n2608 0.106
R5104 S.n3482 S.n3479 0.106
R5105 S.n4330 S.n4327 0.106
R5106 S.n5136 S.n5133 0.106
R5107 S.n5933 S.n5930 0.106
R5108 S.n6704 S.n6701 0.106
R5109 S.n7466 S.n7463 0.106
R5110 S.n8050 S.n8047 0.106
R5111 S.n8762 S.n8759 0.106
R5112 S.n9630 S.n9627 0.106
R5113 S.n10322 S.n10319 0.106
R5114 S.n10991 S.n10988 0.106
R5115 S.n12007 S.n12002 0.106
R5116 S.n2200 S.n2199 0.097
R5117 S.n3038 S.n3037 0.097
R5118 S.n3850 S.n3849 0.097
R5119 S.n4650 S.n4649 0.097
R5120 S.n5427 S.n5426 0.097
R5121 S.n6192 S.n6191 0.097
R5122 S.n6934 S.n6933 0.097
R5123 S.n7664 S.n7663 0.097
R5124 S.n8371 S.n8370 0.097
R5125 S.n9066 S.n9065 0.097
R5126 S.n9738 S.n9737 0.097
R5127 S.n10398 S.n10397 0.097
R5128 S.n11110 S.n11109 0.097
R5129 S.n1731 S.n1730 0.097
R5130 S.n1759 S.n1758 0.097
R5131 S.n12299 S.n12298 0.095
R5132 S.n12385 S.n12384 0.093
R5133 S.n12606 S.n12605 0.093
R5134 S.n11952 S.n11951 0.093
R5135 S.n12625 S.n12624 0.092
R5136 S.n12648 S.n12647 0.092
R5137 S S.n13178 0.09
R5138 S.n1010 S.n1009 0.087
R5139 S.n12464 S.n12463 0.087
R5140 S.n12383 S.n12382 0.085
R5141 S.n872 S.n869 0.082
R5142 S.n995 S.n992 0.082
R5143 S.n1839 S.n1836 0.082
R5144 S.n2722 S.n2719 0.082
R5145 S.n3563 S.n3560 0.082
R5146 S.n4395 S.n4392 0.082
R5147 S.n5201 S.n5198 0.082
R5148 S.n5998 S.n5995 0.082
R5149 S.n6769 S.n6766 0.082
R5150 S.n7531 S.n7528 0.082
R5151 S.n8267 S.n8264 0.082
R5152 S.n8994 S.n8991 0.082
R5153 S.n9695 S.n9692 0.082
R5154 S.n10387 S.n10384 0.082
R5155 S.n11046 S.n11043 0.082
R5156 S.n12289 S.n12286 0.082
R5157 S.n13159 S.n13156 0.082
R5158 S.n11105 S.n11104 0.08
R5159 S.n10393 S.n10392 0.08
R5160 S.n9733 S.n9732 0.08
R5161 S.n9061 S.n9060 0.08
R5162 S.n8366 S.n8365 0.08
R5163 S.n7659 S.n7658 0.08
R5164 S.n6929 S.n6928 0.08
R5165 S.n6187 S.n6186 0.08
R5166 S.n5422 S.n5421 0.08
R5167 S.n4645 S.n4644 0.08
R5168 S.n3845 S.n3844 0.08
R5169 S.n3033 S.n3032 0.08
R5170 S.n2195 S.n2194 0.08
R5171 S.n1761 S.n1760 0.08
R5172 S.n1733 S.n1732 0.08
R5173 S.n12548 S.n12547 0.079
R5174 S.n1822 S.n1821 0.079
R5175 S.n2705 S.n2704 0.079
R5176 S.n3546 S.n3545 0.079
R5177 S.n4378 S.n4377 0.079
R5178 S.n5184 S.n5183 0.079
R5179 S.n5981 S.n5980 0.079
R5180 S.n6752 S.n6751 0.079
R5181 S.n7514 S.n7513 0.079
R5182 S.n8250 S.n8249 0.079
R5183 S.n8977 S.n8976 0.079
R5184 S.n9678 S.n9677 0.079
R5185 S.n10370 S.n10369 0.079
R5186 S.n1262 S.n1261 0.077
R5187 S.n2542 S.n2541 0.077
R5188 S.n3398 S.n3397 0.077
R5189 S.n4245 S.n4244 0.077
R5190 S.n5035 S.n5034 0.077
R5191 S.n5816 S.n5815 0.077
R5192 S.n6571 S.n6570 0.077
R5193 S.n7317 S.n7316 0.077
R5194 S.n7870 S.n7869 0.077
R5195 S.n8566 S.n8565 0.077
R5196 S.n9433 S.n9432 0.077
R5197 S.n10109 S.n10108 0.077
R5198 S.n10762 S.n10761 0.077
R5199 S.n689 S.n688 0.077
R5200 S.n708 S.n707 0.077
R5201 S.n11394 S.n11393 0.076
R5202 S.n1825 S.n1824 0.075
R5203 S.n2708 S.n2707 0.075
R5204 S.n3549 S.n3548 0.075
R5205 S.n4381 S.n4380 0.075
R5206 S.n5187 S.n5186 0.075
R5207 S.n5984 S.n5983 0.075
R5208 S.n6755 S.n6754 0.075
R5209 S.n7517 S.n7516 0.075
R5210 S.n8253 S.n8252 0.075
R5211 S.n8980 S.n8979 0.075
R5212 S.n9681 S.n9680 0.075
R5213 S.n10373 S.n10372 0.075
R5214 S.n12617 S.n12616 0.074
R5215 S.n10751 S.n10750 0.074
R5216 S.n11965 S.n11964 0.074
R5217 S.n10080 S.n10079 0.074
R5218 S.n9386 S.n9385 0.074
R5219 S.n8501 S.n8500 0.074
R5220 S.n7787 S.n7786 0.074
R5221 S.n7216 S.n7215 0.074
R5222 S.n6452 S.n6451 0.074
R5223 S.n5679 S.n5678 0.074
R5224 S.n4880 S.n4879 0.074
R5225 S.n4072 S.n4071 0.074
R5226 S.n3207 S.n3206 0.074
R5227 S.n2333 S.n2332 0.074
R5228 S.n1042 S.n1041 0.074
R5229 S.n472 S.n471 0.074
R5230 S.n12381 S.n12380 0.073
R5231 S.n12378 S.n12377 0.073
R5232 S.n12374 S.n12373 0.073
R5233 S.n12370 S.n12369 0.073
R5234 S.n12366 S.n12365 0.073
R5235 S.n12362 S.n12361 0.073
R5236 S.n12358 S.n12357 0.073
R5237 S.n12354 S.n12353 0.073
R5238 S.n12350 S.n12349 0.073
R5239 S.n12346 S.n12345 0.073
R5240 S.n12342 S.n12341 0.073
R5241 S.n12338 S.n12337 0.073
R5242 S.n12334 S.n12333 0.073
R5243 S.n12331 S.n12330 0.073
R5244 S.n10400 S.n10399 0.071
R5245 S.n9740 S.n9739 0.071
R5246 S.n9068 S.n9067 0.071
R5247 S.n8373 S.n8372 0.071
R5248 S.n7666 S.n7665 0.071
R5249 S.n6936 S.n6935 0.071
R5250 S.n6194 S.n6193 0.071
R5251 S.n5429 S.n5428 0.071
R5252 S.n4652 S.n4651 0.071
R5253 S.n3852 S.n3851 0.071
R5254 S.n3040 S.n3039 0.071
R5255 S.n2202 S.n2201 0.071
R5256 S.n1727 S.n1726 0.071
R5257 S.n1755 S.n1754 0.071
R5258 S.n12005 S.n12004 0.07
R5259 S.t35 S.n12386 0.068
R5260 S.n942 S.n940 0.067
R5261 S.n942 S.n941 0.067
R5262 S.n205 S.n203 0.067
R5263 S.n205 S.n204 0.067
R5264 S.n906 S.n904 0.067
R5265 S.n906 S.n905 0.067
R5266 S.n936 S.n934 0.067
R5267 S.n936 S.n935 0.067
R5268 S.n9 S.n7 0.067
R5269 S.n9 S.n8 0.067
R5270 S.n192 S.n190 0.067
R5271 S.n192 S.n191 0.067
R5272 S.n20 S.n18 0.067
R5273 S.n20 S.n19 0.067
R5274 S.n180 S.n178 0.067
R5275 S.n180 S.n179 0.067
R5276 S.n32 S.n30 0.067
R5277 S.n32 S.n31 0.067
R5278 S.n167 S.n165 0.067
R5279 S.n167 S.n166 0.067
R5280 S.n64 S.n62 0.067
R5281 S.n64 S.n63 0.067
R5282 S.n154 S.n152 0.067
R5283 S.n154 S.n153 0.067
R5284 S.n76 S.n74 0.067
R5285 S.n76 S.n75 0.067
R5286 S.n141 S.n139 0.067
R5287 S.n141 S.n140 0.067
R5288 S.n88 S.n86 0.067
R5289 S.n88 S.n87 0.067
R5290 S.n128 S.n126 0.067
R5291 S.n128 S.n127 0.067
R5292 S.n92 S.n91 0.067
R5293 S.n92 S.n90 0.067
R5294 S.n872 S.n862 0.067
R5295 S.n872 S.n860 0.067
R5296 S.n1839 S.n1830 0.067
R5297 S.n1839 S.n1829 0.067
R5298 S.n2722 S.n2713 0.067
R5299 S.n2722 S.n2712 0.067
R5300 S.n3563 S.n3554 0.067
R5301 S.n3563 S.n3553 0.067
R5302 S.n4395 S.n4386 0.067
R5303 S.n4395 S.n4385 0.067
R5304 S.n5201 S.n5192 0.067
R5305 S.n5201 S.n5191 0.067
R5306 S.n5998 S.n5989 0.067
R5307 S.n5998 S.n5988 0.067
R5308 S.n6769 S.n6760 0.067
R5309 S.n6769 S.n6759 0.067
R5310 S.n7531 S.n7522 0.067
R5311 S.n7531 S.n7521 0.067
R5312 S.n8267 S.n8258 0.067
R5313 S.n8267 S.n8257 0.067
R5314 S.n8994 S.n8985 0.067
R5315 S.n8994 S.n8984 0.067
R5316 S.n9695 S.n9686 0.067
R5317 S.n9695 S.n9685 0.067
R5318 S.n10387 S.n10378 0.067
R5319 S.n10387 S.n10377 0.067
R5320 S.n11046 S.n11037 0.067
R5321 S.n11046 S.n11036 0.067
R5322 S.n12289 S.n12280 0.067
R5323 S.n13159 S.n13149 0.067
R5324 S.n13159 S.n13150 0.067
R5325 S.n12289 S.n12279 0.067
R5326 S.n121 S.n120 0.066
R5327 S.n901 S.n900 0.066
R5328 S.n873 S.n858 0.065
R5329 S.n937 S.n933 0.063
R5330 S.n12290 S.n12289 0.063
R5331 S.n937 S.n936 0.063
R5332 S.n1785 S.n1784 0.063
R5333 S.n2275 S.n2274 0.063
R5334 S.n2592 S.n2591 0.063
R5335 S.n3110 S.n3109 0.063
R5336 S.n3448 S.n3447 0.063
R5337 S.n3922 S.n3921 0.063
R5338 S.n4295 S.n4294 0.063
R5339 S.n4722 S.n4721 0.063
R5340 S.n5085 S.n5084 0.063
R5341 S.n5499 S.n5498 0.063
R5342 S.n5866 S.n5865 0.063
R5343 S.n6264 S.n6263 0.063
R5344 S.n6621 S.n6620 0.063
R5345 S.n7006 S.n7005 0.063
R5346 S.n7367 S.n7366 0.063
R5347 S.n7736 S.n7735 0.063
R5348 S.n7920 S.n7919 0.063
R5349 S.n8443 S.n8442 0.063
R5350 S.n8616 S.n8615 0.063
R5351 S.n9138 S.n9137 0.063
R5352 S.n9483 S.n9482 0.063
R5353 S.n9810 S.n9809 0.063
R5354 S.n10159 S.n10158 0.063
R5355 S.n10470 S.n10469 0.063
R5356 S.n10812 S.n10811 0.063
R5357 S.n11095 S.n11094 0.063
R5358 S.n11433 S.n11432 0.063
R5359 S.n11692 S.n11691 0.063
R5360 S.n11985 S.n11984 0.063
R5361 S.n823 S.n810 0.063
R5362 S.n729 S.n718 0.063
R5363 S.t320 S.n1019 0.063
R5364 S.n2186 S.n2185 0.063
R5365 S.n2532 S.n2531 0.063
R5366 S.n3024 S.n3023 0.063
R5367 S.n3388 S.n3387 0.063
R5368 S.n3836 S.n3835 0.063
R5369 S.n4235 S.n4234 0.063
R5370 S.n4636 S.n4635 0.063
R5371 S.n5025 S.n5024 0.063
R5372 S.n5413 S.n5412 0.063
R5373 S.n5806 S.n5805 0.063
R5374 S.n6178 S.n6177 0.063
R5375 S.n6561 S.n6560 0.063
R5376 S.n6920 S.n6919 0.063
R5377 S.n7307 S.n7306 0.063
R5378 S.n7650 S.n7649 0.063
R5379 S.n7860 S.n7859 0.063
R5380 S.n8357 S.n8356 0.063
R5381 S.n8556 S.n8555 0.063
R5382 S.n9052 S.n9051 0.063
R5383 S.n9423 S.n9422 0.063
R5384 S.n9724 S.n9723 0.063
R5385 S.n10099 S.n10098 0.063
R5386 S.n1763 S.n1743 0.063
R5387 S.n2241 S.n2228 0.063
R5388 S.n3078 S.n3066 0.063
R5389 S.n3890 S.n3878 0.063
R5390 S.n4690 S.n4678 0.063
R5391 S.n5467 S.n5455 0.063
R5392 S.n6232 S.n6220 0.063
R5393 S.n6974 S.n6962 0.063
R5394 S.n7704 S.n7692 0.063
R5395 S.n8411 S.n8399 0.063
R5396 S.n9106 S.n9094 0.063
R5397 S.n9778 S.n9766 0.063
R5398 S.n10438 S.n10426 0.063
R5399 S.n11063 S.n11051 0.063
R5400 S.n802 S.n788 0.063
R5401 S.n9020 S.n8999 0.063
R5402 S.n8325 S.n8304 0.063
R5403 S.n7618 S.n7597 0.063
R5404 S.n6888 S.n6867 0.063
R5405 S.n6146 S.n6125 0.063
R5406 S.n5381 S.n5360 0.063
R5407 S.n4604 S.n4583 0.063
R5408 S.n3804 S.n3783 0.063
R5409 S.n2992 S.n2971 0.063
R5410 S.n2151 S.n2130 0.063
R5411 S.n1701 S.n1682 0.063
R5412 S.n446 S.n434 0.063
R5413 S.n1673 S.n1672 0.063
R5414 S.n2122 S.n2121 0.063
R5415 S.n2496 S.n2495 0.063
R5416 S.n2963 S.n2962 0.063
R5417 S.n3352 S.n3351 0.063
R5418 S.n3775 S.n3774 0.063
R5419 S.n4199 S.n4198 0.063
R5420 S.n4575 S.n4574 0.063
R5421 S.n4989 S.n4988 0.063
R5422 S.n5352 S.n5351 0.063
R5423 S.n5770 S.n5769 0.063
R5424 S.n6117 S.n6116 0.063
R5425 S.n6525 S.n6524 0.063
R5426 S.n6859 S.n6858 0.063
R5427 S.n7271 S.n7270 0.063
R5428 S.n7589 S.n7588 0.063
R5429 S.n7824 S.n7823 0.063
R5430 S.n8296 S.n8295 0.063
R5431 S.n8520 S.n8519 0.063
R5432 S.n7557 S.n7536 0.063
R5433 S.n6827 S.n6806 0.063
R5434 S.n6085 S.n6064 0.063
R5435 S.n5320 S.n5299 0.063
R5436 S.n4543 S.n4522 0.063
R5437 S.n3743 S.n3722 0.063
R5438 S.n2931 S.n2910 0.063
R5439 S.n2088 S.n2067 0.063
R5440 S.n1643 S.n1623 0.063
R5441 S.n405 S.n393 0.063
R5442 S.n1614 S.n1613 0.063
R5443 S.n2059 S.n2058 0.063
R5444 S.n2460 S.n2459 0.063
R5445 S.n2902 S.n2901 0.063
R5446 S.n3316 S.n3315 0.063
R5447 S.n3714 S.n3713 0.063
R5448 S.n4163 S.n4162 0.063
R5449 S.n4514 S.n4513 0.063
R5450 S.n4953 S.n4952 0.063
R5451 S.n5291 S.n5290 0.063
R5452 S.n5734 S.n5733 0.063
R5453 S.n6056 S.n6055 0.063
R5454 S.n6489 S.n6488 0.063
R5455 S.n6798 S.n6797 0.063
R5456 S.n7235 S.n7234 0.063
R5457 S.n6024 S.n6003 0.063
R5458 S.n5259 S.n5238 0.063
R5459 S.n4482 S.n4461 0.063
R5460 S.n3682 S.n3661 0.063
R5461 S.n2870 S.n2849 0.063
R5462 S.n2025 S.n2004 0.063
R5463 S.n1584 S.n1564 0.063
R5464 S.n364 S.n352 0.063
R5465 S.n1555 S.n1554 0.063
R5466 S.n1996 S.n1995 0.063
R5467 S.n2424 S.n2423 0.063
R5468 S.n2841 S.n2840 0.063
R5469 S.n3280 S.n3279 0.063
R5470 S.n3653 S.n3652 0.063
R5471 S.n4127 S.n4126 0.063
R5472 S.n4453 S.n4452 0.063
R5473 S.n4917 S.n4916 0.063
R5474 S.n5230 S.n5229 0.063
R5475 S.n5698 S.n5697 0.063
R5476 S.n4421 S.n4400 0.063
R5477 S.n3621 S.n3600 0.063
R5478 S.n2809 S.n2788 0.063
R5479 S.n1962 S.n1941 0.063
R5480 S.n1525 S.n1505 0.063
R5481 S.n59 S.n41 0.063
R5482 S.n1496 S.n1495 0.063
R5483 S.n1933 S.n1932 0.063
R5484 S.n2388 S.n2387 0.063
R5485 S.n2780 S.n2779 0.063
R5486 S.n3244 S.n3243 0.063
R5487 S.n3592 S.n3591 0.063
R5488 S.n4091 S.n4090 0.063
R5489 S.n2748 S.n2727 0.063
R5490 S.n1899 S.n1878 0.063
R5491 S.n1469 S.n1446 0.063
R5492 S.n302 S.n290 0.063
R5493 S.n1437 S.n1436 0.063
R5494 S.n1870 S.n1869 0.063
R5495 S.n2352 S.n2351 0.063
R5496 S.n1407 S.n1387 0.063
R5497 S.n261 S.n249 0.063
R5498 S.n851 S.n850 0.063
R5499 S.n943 S.n942 0.062
R5500 S.n193 S.n192 0.062
R5501 S.n181 S.n180 0.062
R5502 S.n168 S.n167 0.062
R5503 S.n155 S.n154 0.062
R5504 S.n142 S.n141 0.062
R5505 S.n129 S.n128 0.062
R5506 S.n917 S.n906 0.061
R5507 S.n10 S.n9 0.06
R5508 S.n21 S.n20 0.06
R5509 S.n33 S.n32 0.06
R5510 S.n65 S.n64 0.06
R5511 S.n77 S.n76 0.06
R5512 S.n89 S.n88 0.06
R5513 S.n93 S.n92 0.06
R5514 S.n12587 S.n12586 0.059
R5515 S.n11701 S.n11700 0.059
R5516 S.n2169 S.n2159 0.059
R5517 S.n206 S.n205 0.059
R5518 S.n13160 S.n13159 0.058
R5519 S.n1811 S.n1810 0.058
R5520 S.n2694 S.n2693 0.058
R5521 S.n3535 S.n3534 0.058
R5522 S.n4367 S.n4366 0.058
R5523 S.n5173 S.n5172 0.058
R5524 S.n5970 S.n5969 0.058
R5525 S.n6741 S.n6740 0.058
R5526 S.n7503 S.n7502 0.058
R5527 S.n8239 S.n8238 0.058
R5528 S.n8966 S.n8965 0.058
R5529 S.n9667 S.n9666 0.058
R5530 S.n10359 S.n10358 0.058
R5531 S.n873 S.n872 0.058
R5532 S.n98 S.n97 0.056
R5533 S.n2 S.n1 0.056
R5534 S.n13 S.n12 0.056
R5535 S.n24 S.n23 0.056
R5536 S.n36 S.n35 0.056
R5537 S.n68 S.n67 0.056
R5538 S.n80 S.n79 0.056
R5539 S.n12546 S.n12545 0.056
R5540 S.n124 S.n102 0.055
R5541 S.n12276 S.n12275 0.055
R5542 S.n885 S.n884 0.055
R5543 S.n1801 S.n1800 0.055
R5544 S.n2684 S.n2683 0.055
R5545 S.n3525 S.n3524 0.055
R5546 S.n4357 S.n4356 0.055
R5547 S.n5163 S.n5162 0.055
R5548 S.n5960 S.n5959 0.055
R5549 S.n6731 S.n6730 0.055
R5550 S.n7493 S.n7492 0.055
R5551 S.n8229 S.n8228 0.055
R5552 S.n8956 S.n8955 0.055
R5553 S.n9657 S.n9656 0.055
R5554 S.n10349 S.n10348 0.055
R5555 S.n11018 S.n11017 0.055
R5556 S.n11658 S.n11657 0.055
R5557 S.n13146 S.n13145 0.055
R5558 S.n474 S.n457 0.054
R5559 S.n12619 S.n12602 0.054
R5560 S.n9389 S.n9372 0.054
R5561 S.n10082 S.n10064 0.054
R5562 S.n10754 S.n10737 0.054
R5563 S.n11396 S.n11375 0.054
R5564 S.n11968 S.n11949 0.054
R5565 S.n7790 S.n7773 0.054
R5566 S.n8503 S.n8485 0.054
R5567 S.n6455 S.n6438 0.054
R5568 S.n7218 S.n7200 0.054
R5569 S.n4883 S.n4866 0.054
R5570 S.n5681 S.n5663 0.054
R5571 S.n3210 S.n3193 0.054
R5572 S.n4074 S.n4056 0.054
R5573 S.n1045 S.n1028 0.054
R5574 S.n2335 S.n2317 0.054
R5575 S.n12315 S.n12314 0.054
R5576 S.n12643 S.n12642 0.054
R5577 S.n12567 S.n12566 0.054
R5578 S.n12012 S.n12011 0.054
R5579 S.n857 S.n856 0.054
R5580 S.n826 S.n825 0.054
R5581 S.n1788 S.n1787 0.054
R5582 S.n12597 S.n12596 0.054
R5583 S.n11988 S.n11987 0.054
R5584 S.n11695 S.n11694 0.054
R5585 S.n11436 S.n11435 0.054
R5586 S.n11098 S.n11097 0.054
R5587 S.n10815 S.n10814 0.054
R5588 S.n10473 S.n10472 0.054
R5589 S.n10162 S.n10161 0.054
R5590 S.n9813 S.n9812 0.054
R5591 S.n9486 S.n9485 0.054
R5592 S.n9141 S.n9140 0.054
R5593 S.n8619 S.n8618 0.054
R5594 S.n8446 S.n8445 0.054
R5595 S.n7923 S.n7922 0.054
R5596 S.n7739 S.n7738 0.054
R5597 S.n7370 S.n7369 0.054
R5598 S.n7009 S.n7008 0.054
R5599 S.n6624 S.n6623 0.054
R5600 S.n6267 S.n6266 0.054
R5601 S.n5869 S.n5868 0.054
R5602 S.n5502 S.n5501 0.054
R5603 S.n5088 S.n5087 0.054
R5604 S.n4725 S.n4724 0.054
R5605 S.n4298 S.n4297 0.054
R5606 S.n3925 S.n3924 0.054
R5607 S.n3451 S.n3450 0.054
R5608 S.n3113 S.n3112 0.054
R5609 S.n2595 S.n2594 0.054
R5610 S.n2278 S.n2277 0.054
R5611 S.n1313 S.n1312 0.054
R5612 S.n732 S.n731 0.054
R5613 S.n429 S.n428 0.054
R5614 S.n1676 S.n1675 0.054
R5615 S.n9170 S.n9169 0.054
R5616 S.n8523 S.n8522 0.054
R5617 S.n8299 S.n8298 0.054
R5618 S.n7827 S.n7826 0.054
R5619 S.n7592 S.n7591 0.054
R5620 S.n7274 S.n7273 0.054
R5621 S.n6862 S.n6861 0.054
R5622 S.n6528 S.n6527 0.054
R5623 S.n6120 S.n6119 0.054
R5624 S.n5773 S.n5772 0.054
R5625 S.n5355 S.n5354 0.054
R5626 S.n4992 S.n4991 0.054
R5627 S.n4578 S.n4577 0.054
R5628 S.n4202 S.n4201 0.054
R5629 S.n3778 S.n3777 0.054
R5630 S.n3355 S.n3354 0.054
R5631 S.n2966 S.n2965 0.054
R5632 S.n2499 S.n2498 0.054
R5633 S.n2125 S.n2124 0.054
R5634 S.n1216 S.n1215 0.054
R5635 S.n449 S.n448 0.054
R5636 S.n9847 S.n9846 0.054
R5637 S.n9407 S.n9406 0.054
R5638 S.n9023 S.n9022 0.054
R5639 S.n8540 S.n8539 0.054
R5640 S.n8328 S.n8327 0.054
R5641 S.n7844 S.n7843 0.054
R5642 S.n7621 S.n7620 0.054
R5643 S.n7291 S.n7290 0.054
R5644 S.n6891 S.n6890 0.054
R5645 S.n6545 S.n6544 0.054
R5646 S.n6149 S.n6148 0.054
R5647 S.n5790 S.n5789 0.054
R5648 S.n5384 S.n5383 0.054
R5649 S.n5009 S.n5008 0.054
R5650 S.n4607 S.n4606 0.054
R5651 S.n4219 S.n4218 0.054
R5652 S.n3807 S.n3806 0.054
R5653 S.n3372 S.n3371 0.054
R5654 S.n2995 S.n2994 0.054
R5655 S.n2516 S.n2515 0.054
R5656 S.n2154 S.n2153 0.054
R5657 S.n1235 S.n1234 0.054
R5658 S.n1255 S.n1254 0.054
R5659 S.n760 S.n759 0.054
R5660 S.n783 S.n782 0.054
R5661 S.n2189 S.n2188 0.054
R5662 S.n3027 S.n3026 0.054
R5663 S.n3839 S.n3838 0.054
R5664 S.n4639 S.n4638 0.054
R5665 S.n5416 S.n5415 0.054
R5666 S.n6181 S.n6180 0.054
R5667 S.n6923 S.n6922 0.054
R5668 S.n7653 S.n7652 0.054
R5669 S.n8360 S.n8359 0.054
R5670 S.n9055 S.n9054 0.054
R5671 S.n9727 S.n9726 0.054
R5672 S.n10505 S.n10504 0.054
R5673 S.n10102 S.n10101 0.054
R5674 S.n9426 S.n9425 0.054
R5675 S.n8559 S.n8558 0.054
R5676 S.n7863 S.n7862 0.054
R5677 S.n7310 S.n7309 0.054
R5678 S.n6564 S.n6563 0.054
R5679 S.n5809 S.n5808 0.054
R5680 S.n5028 S.n5027 0.054
R5681 S.n4238 S.n4237 0.054
R5682 S.n3391 S.n3390 0.054
R5683 S.n2535 S.n2534 0.054
R5684 S.n1738 S.n1737 0.054
R5685 S.n693 S.n692 0.054
R5686 S.n891 S.n890 0.054
R5687 S.n11128 S.n11127 0.054
R5688 S.n10776 S.n10775 0.054
R5689 S.n10421 S.n10420 0.054
R5690 S.n10123 S.n10122 0.054
R5691 S.n9761 S.n9760 0.054
R5692 S.n9447 S.n9446 0.054
R5693 S.n9089 S.n9088 0.054
R5694 S.n8580 S.n8579 0.054
R5695 S.n8394 S.n8393 0.054
R5696 S.n7884 S.n7883 0.054
R5697 S.n7687 S.n7686 0.054
R5698 S.n7331 S.n7330 0.054
R5699 S.n6957 S.n6956 0.054
R5700 S.n6585 S.n6584 0.054
R5701 S.n6215 S.n6214 0.054
R5702 S.n5830 S.n5829 0.054
R5703 S.n5450 S.n5449 0.054
R5704 S.n5049 S.n5048 0.054
R5705 S.n4673 S.n4672 0.054
R5706 S.n4259 S.n4258 0.054
R5707 S.n3873 S.n3872 0.054
R5708 S.n3412 S.n3411 0.054
R5709 S.n3061 S.n3060 0.054
R5710 S.n2556 S.n2555 0.054
R5711 S.n2223 S.n2222 0.054
R5712 S.n1276 S.n1275 0.054
R5713 S.n1766 S.n1765 0.054
R5714 S.n712 S.n711 0.054
R5715 S.n1296 S.n1295 0.054
R5716 S.n2244 S.n2243 0.054
R5717 S.n2576 S.n2575 0.054
R5718 S.n3081 S.n3080 0.054
R5719 S.n3432 S.n3431 0.054
R5720 S.n3893 S.n3892 0.054
R5721 S.n4279 S.n4278 0.054
R5722 S.n4693 S.n4692 0.054
R5723 S.n5069 S.n5068 0.054
R5724 S.n5470 S.n5469 0.054
R5725 S.n5850 S.n5849 0.054
R5726 S.n6235 S.n6234 0.054
R5727 S.n6605 S.n6604 0.054
R5728 S.n6977 S.n6976 0.054
R5729 S.n7351 S.n7350 0.054
R5730 S.n7707 S.n7706 0.054
R5731 S.n7904 S.n7903 0.054
R5732 S.n8414 S.n8413 0.054
R5733 S.n8600 S.n8599 0.054
R5734 S.n9109 S.n9108 0.054
R5735 S.n9467 S.n9466 0.054
R5736 S.n9781 S.n9780 0.054
R5737 S.n10143 S.n10142 0.054
R5738 S.n10441 S.n10440 0.054
R5739 S.n10796 S.n10795 0.054
R5740 S.n11066 S.n11065 0.054
R5741 S.n11417 S.n11416 0.054
R5742 S.n11723 S.n11722 0.054
R5743 S.n805 S.n804 0.054
R5744 S.n1704 S.n1703 0.054
R5745 S.n673 S.n672 0.054
R5746 S.n656 S.n655 0.054
R5747 S.n388 S.n387 0.054
R5748 S.n1617 S.n1616 0.054
R5749 S.n7768 S.n7767 0.054
R5750 S.n7238 S.n7237 0.054
R5751 S.n6801 S.n6800 0.054
R5752 S.n6492 S.n6491 0.054
R5753 S.n6059 S.n6058 0.054
R5754 S.n5737 S.n5736 0.054
R5755 S.n5294 S.n5293 0.054
R5756 S.n4956 S.n4955 0.054
R5757 S.n4517 S.n4516 0.054
R5758 S.n4166 S.n4165 0.054
R5759 S.n3717 S.n3716 0.054
R5760 S.n3319 S.n3318 0.054
R5761 S.n2905 S.n2904 0.054
R5762 S.n2463 S.n2462 0.054
R5763 S.n2062 S.n2061 0.054
R5764 S.n1182 S.n1181 0.054
R5765 S.n408 S.n407 0.054
R5766 S.n8480 S.n8479 0.054
R5767 S.n7808 S.n7807 0.054
R5768 S.n7560 S.n7559 0.054
R5769 S.n7255 S.n7254 0.054
R5770 S.n6830 S.n6829 0.054
R5771 S.n6509 S.n6508 0.054
R5772 S.n6088 S.n6087 0.054
R5773 S.n5754 S.n5753 0.054
R5774 S.n5323 S.n5322 0.054
R5775 S.n4973 S.n4972 0.054
R5776 S.n4546 S.n4545 0.054
R5777 S.n4183 S.n4182 0.054
R5778 S.n3746 S.n3745 0.054
R5779 S.n3336 S.n3335 0.054
R5780 S.n2934 S.n2933 0.054
R5781 S.n2480 S.n2479 0.054
R5782 S.n2091 S.n2090 0.054
R5783 S.n1199 S.n1198 0.054
R5784 S.n1646 S.n1645 0.054
R5785 S.n640 S.n639 0.054
R5786 S.n623 S.n622 0.054
R5787 S.n347 S.n346 0.054
R5788 S.n1558 S.n1557 0.054
R5789 S.n6296 S.n6295 0.054
R5790 S.n5701 S.n5700 0.054
R5791 S.n5233 S.n5232 0.054
R5792 S.n4920 S.n4919 0.054
R5793 S.n4456 S.n4455 0.054
R5794 S.n4130 S.n4129 0.054
R5795 S.n3656 S.n3655 0.054
R5796 S.n3283 S.n3282 0.054
R5797 S.n2844 S.n2843 0.054
R5798 S.n2427 S.n2426 0.054
R5799 S.n1999 S.n1998 0.054
R5800 S.n1148 S.n1147 0.054
R5801 S.n367 S.n366 0.054
R5802 S.n7043 S.n7042 0.054
R5803 S.n6473 S.n6472 0.054
R5804 S.n6027 S.n6026 0.054
R5805 S.n5718 S.n5717 0.054
R5806 S.n5262 S.n5261 0.054
R5807 S.n4937 S.n4936 0.054
R5808 S.n4485 S.n4484 0.054
R5809 S.n4147 S.n4146 0.054
R5810 S.n3685 S.n3684 0.054
R5811 S.n3300 S.n3299 0.054
R5812 S.n2873 S.n2872 0.054
R5813 S.n2444 S.n2443 0.054
R5814 S.n2028 S.n2027 0.054
R5815 S.n1165 S.n1164 0.054
R5816 S.n1587 S.n1586 0.054
R5817 S.n607 S.n606 0.054
R5818 S.n590 S.n589 0.054
R5819 S.n326 S.n325 0.054
R5820 S.n1499 S.n1498 0.054
R5821 S.n4754 S.n4753 0.054
R5822 S.n4094 S.n4093 0.054
R5823 S.n3595 S.n3594 0.054
R5824 S.n3247 S.n3246 0.054
R5825 S.n2783 S.n2782 0.054
R5826 S.n2391 S.n2390 0.054
R5827 S.n1936 S.n1935 0.054
R5828 S.n1114 S.n1113 0.054
R5829 S.n54 S.n53 0.054
R5830 S.n5536 S.n5535 0.054
R5831 S.n4901 S.n4900 0.054
R5832 S.n4424 S.n4423 0.054
R5833 S.n4111 S.n4110 0.054
R5834 S.n3624 S.n3623 0.054
R5835 S.n3264 S.n3263 0.054
R5836 S.n2812 S.n2811 0.054
R5837 S.n2408 S.n2407 0.054
R5838 S.n1965 S.n1964 0.054
R5839 S.n1131 S.n1130 0.054
R5840 S.n1528 S.n1527 0.054
R5841 S.n574 S.n573 0.054
R5842 S.n557 S.n556 0.054
R5843 S.n285 S.n284 0.054
R5844 S.n1440 S.n1439 0.054
R5845 S.n3142 S.n3141 0.054
R5846 S.n2355 S.n2354 0.054
R5847 S.n1873 S.n1872 0.054
R5848 S.n1080 S.n1079 0.054
R5849 S.n305 S.n304 0.054
R5850 S.n3959 S.n3958 0.054
R5851 S.n3228 S.n3227 0.054
R5852 S.n2751 S.n2750 0.054
R5853 S.n2372 S.n2371 0.054
R5854 S.n1902 S.n1901 0.054
R5855 S.n1097 S.n1096 0.054
R5856 S.n1455 S.n1454 0.054
R5857 S.n541 S.n540 0.054
R5858 S.n524 S.n523 0.054
R5859 S.n244 S.n243 0.054
R5860 S.n1381 S.n1380 0.054
R5861 S.n264 S.n263 0.054
R5862 S.n2312 S.n2311 0.054
R5863 S.n1063 S.n1062 0.054
R5864 S.n1410 S.n1409 0.054
R5865 S.n508 S.n507 0.054
R5866 S.n491 S.n490 0.054
R5867 S.n754 S.n753 0.054
R5868 S.n1358 S.n1357 0.054
R5869 S.n1339 S.n1338 0.054
R5870 S.n2652 S.n2651 0.054
R5871 S.n2625 S.n2624 0.054
R5872 S.n3179 S.n3178 0.054
R5873 S.n3152 S.n3151 0.054
R5874 S.n3996 S.n3995 0.054
R5875 S.n3969 S.n3968 0.054
R5876 S.n4791 S.n4790 0.054
R5877 S.n4764 S.n4763 0.054
R5878 S.n5573 S.n5572 0.054
R5879 S.n5546 S.n5545 0.054
R5880 S.n6333 S.n6332 0.054
R5881 S.n6306 S.n6305 0.054
R5882 S.n7080 S.n7079 0.054
R5883 S.n7053 S.n7052 0.054
R5884 S.n8091 S.n8090 0.054
R5885 S.n8064 S.n8063 0.054
R5886 S.n8803 S.n8802 0.054
R5887 S.n8776 S.n8775 0.054
R5888 S.n9207 S.n9206 0.054
R5889 S.n9180 S.n9179 0.054
R5890 S.n9884 S.n9883 0.054
R5891 S.n9857 S.n9856 0.054
R5892 S.n10542 S.n10541 0.054
R5893 S.n10515 S.n10514 0.054
R5894 S.n11165 S.n11164 0.054
R5895 S.n11138 S.n11137 0.054
R5896 S.n11743 S.n11742 0.054
R5897 S.n12033 S.n12032 0.054
R5898 S.n12912 S.n12911 0.054
R5899 S.n12884 S.n12883 0.054
R5900 S.n1333 S.n1332 0.054
R5901 S.n2682 S.n2681 0.054
R5902 S.n12928 S.n12927 0.054
R5903 S.n12943 S.n12942 0.054
R5904 S.n12048 S.n12047 0.054
R5905 S.n11759 S.n11758 0.054
R5906 S.n11181 S.n11180 0.054
R5907 S.n11196 S.n11195 0.054
R5908 S.n10558 S.n10557 0.054
R5909 S.n10573 S.n10572 0.054
R5910 S.n9900 S.n9899 0.054
R5911 S.n9915 S.n9914 0.054
R5912 S.n9223 S.n9222 0.054
R5913 S.n9238 S.n9237 0.054
R5914 S.n8819 S.n8818 0.054
R5915 S.n8834 S.n8833 0.054
R5916 S.n8107 S.n8106 0.054
R5917 S.n8122 S.n8121 0.054
R5918 S.n7096 S.n7095 0.054
R5919 S.n7111 S.n7110 0.054
R5920 S.n6349 S.n6348 0.054
R5921 S.n6364 S.n6363 0.054
R5922 S.n5589 S.n5588 0.054
R5923 S.n5604 S.n5603 0.054
R5924 S.n4807 S.n4806 0.054
R5925 S.n4822 S.n4821 0.054
R5926 S.n4015 S.n4014 0.054
R5927 S.n4027 S.n4026 0.054
R5928 S.n3493 S.n3492 0.054
R5929 S.n3508 S.n3507 0.054
R5930 S.n2668 S.n2667 0.054
R5931 S.n2619 S.n2618 0.054
R5932 S.n3523 S.n3522 0.054
R5933 S.n12686 S.n12685 0.054
R5934 S.n12958 S.n12957 0.054
R5935 S.n12064 S.n12063 0.054
R5936 S.n11774 S.n11773 0.054
R5937 S.n11456 S.n11455 0.054
R5938 S.n11211 S.n11210 0.054
R5939 S.n10835 S.n10834 0.054
R5940 S.n10588 S.n10587 0.054
R5941 S.n10182 S.n10181 0.054
R5942 S.n9930 S.n9929 0.054
R5943 S.n9506 S.n9505 0.054
R5944 S.n9253 S.n9252 0.054
R5945 S.n8639 S.n8638 0.054
R5946 S.n8849 S.n8848 0.054
R5947 S.n7943 S.n7942 0.054
R5948 S.n8137 S.n8136 0.054
R5949 S.n7390 S.n7389 0.054
R5950 S.n7126 S.n7125 0.054
R5951 S.n6644 S.n6643 0.054
R5952 S.n6379 S.n6378 0.054
R5953 S.n5889 S.n5888 0.054
R5954 S.n5619 S.n5618 0.054
R5955 S.n5108 S.n5107 0.054
R5956 S.n4837 S.n4836 0.054
R5957 S.n4318 S.n4317 0.054
R5958 S.n4042 S.n4041 0.054
R5959 S.n3470 S.n3469 0.054
R5960 S.n3490 S.n3489 0.054
R5961 S.n4355 S.n4354 0.054
R5962 S.n12702 S.n12701 0.054
R5963 S.n12973 S.n12972 0.054
R5964 S.n12080 S.n12079 0.054
R5965 S.n11789 S.n11788 0.054
R5966 S.n11472 S.n11471 0.054
R5967 S.n11226 S.n11225 0.054
R5968 S.n10851 S.n10850 0.054
R5969 S.n10603 S.n10602 0.054
R5970 S.n10198 S.n10197 0.054
R5971 S.n9945 S.n9944 0.054
R5972 S.n9522 S.n9521 0.054
R5973 S.n9268 S.n9267 0.054
R5974 S.n8655 S.n8654 0.054
R5975 S.n8864 S.n8863 0.054
R5976 S.n7959 S.n7958 0.054
R5977 S.n8152 S.n8151 0.054
R5978 S.n7406 S.n7405 0.054
R5979 S.n7141 S.n7140 0.054
R5980 S.n6660 S.n6659 0.054
R5981 S.n6394 S.n6393 0.054
R5982 S.n5905 S.n5904 0.054
R5983 S.n5634 S.n5633 0.054
R5984 S.n5124 S.n5123 0.054
R5985 S.n4852 S.n4851 0.054
R5986 S.n4341 S.n4340 0.054
R5987 S.n4338 S.n4337 0.054
R5988 S.n5161 S.n5160 0.054
R5989 S.n12718 S.n12717 0.054
R5990 S.n12988 S.n12987 0.054
R5991 S.n12096 S.n12095 0.054
R5992 S.n11804 S.n11803 0.054
R5993 S.n11488 S.n11487 0.054
R5994 S.n11241 S.n11240 0.054
R5995 S.n10867 S.n10866 0.054
R5996 S.n10618 S.n10617 0.054
R5997 S.n10214 S.n10213 0.054
R5998 S.n9960 S.n9959 0.054
R5999 S.n9538 S.n9537 0.054
R6000 S.n9283 S.n9282 0.054
R6001 S.n8671 S.n8670 0.054
R6002 S.n8879 S.n8878 0.054
R6003 S.n7975 S.n7974 0.054
R6004 S.n8167 S.n8166 0.054
R6005 S.n7422 S.n7421 0.054
R6006 S.n7156 S.n7155 0.054
R6007 S.n6676 S.n6675 0.054
R6008 S.n6409 S.n6408 0.054
R6009 S.n5921 S.n5920 0.054
R6010 S.n5649 S.n5648 0.054
R6011 S.n5147 S.n5146 0.054
R6012 S.n5144 S.n5143 0.054
R6013 S.n5958 S.n5957 0.054
R6014 S.n12734 S.n12733 0.054
R6015 S.n13003 S.n13002 0.054
R6016 S.n12112 S.n12111 0.054
R6017 S.n11819 S.n11818 0.054
R6018 S.n11504 S.n11503 0.054
R6019 S.n11256 S.n11255 0.054
R6020 S.n10883 S.n10882 0.054
R6021 S.n10633 S.n10632 0.054
R6022 S.n10230 S.n10229 0.054
R6023 S.n9975 S.n9974 0.054
R6024 S.n9554 S.n9553 0.054
R6025 S.n9298 S.n9297 0.054
R6026 S.n8687 S.n8686 0.054
R6027 S.n8894 S.n8893 0.054
R6028 S.n7991 S.n7990 0.054
R6029 S.n8182 S.n8181 0.054
R6030 S.n7438 S.n7437 0.054
R6031 S.n7171 S.n7170 0.054
R6032 S.n6692 S.n6691 0.054
R6033 S.n6424 S.n6423 0.054
R6034 S.n5944 S.n5943 0.054
R6035 S.n5941 S.n5940 0.054
R6036 S.n6729 S.n6728 0.054
R6037 S.n12750 S.n12749 0.054
R6038 S.n13018 S.n13017 0.054
R6039 S.n12128 S.n12127 0.054
R6040 S.n11834 S.n11833 0.054
R6041 S.n11520 S.n11519 0.054
R6042 S.n11271 S.n11270 0.054
R6043 S.n10899 S.n10898 0.054
R6044 S.n10648 S.n10647 0.054
R6045 S.n10246 S.n10245 0.054
R6046 S.n9990 S.n9989 0.054
R6047 S.n9570 S.n9569 0.054
R6048 S.n9313 S.n9312 0.054
R6049 S.n8703 S.n8702 0.054
R6050 S.n8909 S.n8908 0.054
R6051 S.n8007 S.n8006 0.054
R6052 S.n8197 S.n8196 0.054
R6053 S.n7454 S.n7453 0.054
R6054 S.n7186 S.n7185 0.054
R6055 S.n6715 S.n6714 0.054
R6056 S.n6712 S.n6711 0.054
R6057 S.n7491 S.n7490 0.054
R6058 S.n12766 S.n12765 0.054
R6059 S.n13033 S.n13032 0.054
R6060 S.n12144 S.n12143 0.054
R6061 S.n11849 S.n11848 0.054
R6062 S.n11536 S.n11535 0.054
R6063 S.n11286 S.n11285 0.054
R6064 S.n10915 S.n10914 0.054
R6065 S.n10663 S.n10662 0.054
R6066 S.n10262 S.n10261 0.054
R6067 S.n10005 S.n10004 0.054
R6068 S.n9586 S.n9585 0.054
R6069 S.n9328 S.n9327 0.054
R6070 S.n8719 S.n8718 0.054
R6071 S.n8924 S.n8923 0.054
R6072 S.n8023 S.n8022 0.054
R6073 S.n8212 S.n8211 0.054
R6074 S.n7477 S.n7476 0.054
R6075 S.n7474 S.n7473 0.054
R6076 S.n8227 S.n8226 0.054
R6077 S.n12782 S.n12781 0.054
R6078 S.n13048 S.n13047 0.054
R6079 S.n12160 S.n12159 0.054
R6080 S.n11864 S.n11863 0.054
R6081 S.n11552 S.n11551 0.054
R6082 S.n11301 S.n11300 0.054
R6083 S.n10931 S.n10930 0.054
R6084 S.n10678 S.n10677 0.054
R6085 S.n10278 S.n10277 0.054
R6086 S.n10020 S.n10019 0.054
R6087 S.n9602 S.n9601 0.054
R6088 S.n9343 S.n9342 0.054
R6089 S.n8735 S.n8734 0.054
R6090 S.n8939 S.n8938 0.054
R6091 S.n8038 S.n8037 0.054
R6092 S.n8058 S.n8057 0.054
R6093 S.n8954 S.n8953 0.054
R6094 S.n12798 S.n12797 0.054
R6095 S.n13063 S.n13062 0.054
R6096 S.n12176 S.n12175 0.054
R6097 S.n11879 S.n11878 0.054
R6098 S.n11568 S.n11567 0.054
R6099 S.n11316 S.n11315 0.054
R6100 S.n10947 S.n10946 0.054
R6101 S.n10693 S.n10692 0.054
R6102 S.n10294 S.n10293 0.054
R6103 S.n10035 S.n10034 0.054
R6104 S.n9618 S.n9617 0.054
R6105 S.n9358 S.n9357 0.054
R6106 S.n8750 S.n8749 0.054
R6107 S.n8770 S.n8769 0.054
R6108 S.n9655 S.n9654 0.054
R6109 S.n12814 S.n12813 0.054
R6110 S.n13078 S.n13077 0.054
R6111 S.n12192 S.n12191 0.054
R6112 S.n11894 S.n11893 0.054
R6113 S.n11584 S.n11583 0.054
R6114 S.n11331 S.n11330 0.054
R6115 S.n10963 S.n10962 0.054
R6116 S.n10708 S.n10707 0.054
R6117 S.n10310 S.n10309 0.054
R6118 S.n10050 S.n10049 0.054
R6119 S.n9641 S.n9640 0.054
R6120 S.n9638 S.n9637 0.054
R6121 S.n10347 S.n10346 0.054
R6122 S.n12830 S.n12829 0.054
R6123 S.n13093 S.n13092 0.054
R6124 S.n12208 S.n12207 0.054
R6125 S.n11909 S.n11908 0.054
R6126 S.n11600 S.n11599 0.054
R6127 S.n11346 S.n11345 0.054
R6128 S.n10979 S.n10978 0.054
R6129 S.n10723 S.n10722 0.054
R6130 S.n10333 S.n10332 0.054
R6131 S.n10330 S.n10329 0.054
R6132 S.n11016 S.n11015 0.054
R6133 S.n12846 S.n12845 0.054
R6134 S.n13108 S.n13107 0.054
R6135 S.n12224 S.n12223 0.054
R6136 S.n11924 S.n11923 0.054
R6137 S.n11616 S.n11615 0.054
R6138 S.n11361 S.n11360 0.054
R6139 S.n11002 S.n11001 0.054
R6140 S.n10999 S.n10998 0.054
R6141 S.n11656 S.n11655 0.054
R6142 S.n12862 S.n12861 0.054
R6143 S.n13123 S.n13122 0.054
R6144 S.n12240 S.n12239 0.054
R6145 S.n11939 S.n11938 0.054
R6146 S.n11642 S.n11641 0.054
R6147 S.n11639 S.n11638 0.054
R6148 S.n12271 S.n12270 0.054
R6149 S.n12878 S.n12877 0.054
R6150 S.n13141 S.n13140 0.054
R6151 S.n12246 S.n12245 0.054
R6152 S.n12666 S.n12665 0.054
R6153 S.t320 S.n1021 0.053
R6154 S.t320 S.n1023 0.052
R6155 S.n470 S.n469 0.052
R6156 S.n1040 S.n1039 0.052
R6157 S.n2331 S.n2330 0.052
R6158 S.n3205 S.n3204 0.052
R6159 S.n4070 S.n4069 0.052
R6160 S.n4878 S.n4877 0.052
R6161 S.n5677 S.n5676 0.052
R6162 S.n6450 S.n6449 0.052
R6163 S.n7214 S.n7213 0.052
R6164 S.n7785 S.n7784 0.052
R6165 S.n8499 S.n8498 0.052
R6166 S.n9384 S.n9383 0.052
R6167 S.n10078 S.n10077 0.052
R6168 S.n10749 S.n10748 0.052
R6169 S.n11392 S.n11391 0.052
R6170 S.n11963 S.n11962 0.052
R6171 S.n12615 S.n12614 0.052
R6172 S.n998 S.n997 0.052
R6173 S.n1821 S.n1820 0.052
R6174 S.n2690 S.n2689 0.052
R6175 S.n2704 S.n2703 0.052
R6176 S.n3531 S.n3530 0.052
R6177 S.n3545 S.n3544 0.052
R6178 S.n4363 S.n4362 0.052
R6179 S.n4377 S.n4376 0.052
R6180 S.n5169 S.n5168 0.052
R6181 S.n5183 S.n5182 0.052
R6182 S.n5966 S.n5965 0.052
R6183 S.n5980 S.n5979 0.052
R6184 S.n6737 S.n6736 0.052
R6185 S.n6751 S.n6750 0.052
R6186 S.n7499 S.n7498 0.052
R6187 S.n7513 S.n7512 0.052
R6188 S.n8235 S.n8234 0.052
R6189 S.n8249 S.n8248 0.052
R6190 S.n8962 S.n8961 0.052
R6191 S.n8976 S.n8975 0.052
R6192 S.n9663 S.n9662 0.052
R6193 S.n9677 S.n9676 0.052
R6194 S.n10355 S.n10354 0.052
R6195 S.n10369 S.n10368 0.052
R6196 S.n11024 S.n11023 0.052
R6197 S.n11664 S.n11663 0.052
R6198 S.n12304 S.n12303 0.052
R6199 S.n12004 S.n12003 0.052
R6200 S.n767 S.n766 0.051
R6201 S.n10497 S.n10495 0.051
R6202 S.n9820 S.n9819 0.051
R6203 S.n9162 S.n9160 0.051
R6204 S.n8453 S.n8452 0.051
R6205 S.n7760 S.n7758 0.051
R6206 S.n7016 S.n7015 0.051
R6207 S.n6288 S.n6286 0.051
R6208 S.n5509 S.n5508 0.051
R6209 S.n4746 S.n4744 0.051
R6210 S.n3932 S.n3931 0.051
R6211 S.n3134 S.n3132 0.051
R6212 S.n2285 S.n2284 0.051
R6213 S.n1376 S.n1374 0.051
R6214 S.n833 S.n832 0.051
R6215 S.n12319 S.n12318 0.051
R6216 S.n12468 S.n12467 0.051
R6217 S.n860 S.n859 0.051
R6218 S.n862 S.n861 0.051
R6219 S.n12591 S.n12590 0.05
R6220 S.n10499 S.n10498 0.05
R6221 S.n11717 S.n11704 0.05
R6222 S.n796 S.n795 0.05
R6223 S.n9838 S.n9835 0.05
R6224 S.n9841 S.n9822 0.05
R6225 S.n9164 S.n9163 0.05
R6226 S.n8469 S.n8468 0.05
R6227 S.n8474 S.n8455 0.05
R6228 S.n7762 S.n7761 0.05
R6229 S.n7032 S.n7031 0.05
R6230 S.n7037 S.n7018 0.05
R6231 S.n6290 S.n6289 0.05
R6232 S.n5527 S.n5524 0.05
R6233 S.n5530 S.n5511 0.05
R6234 S.n4748 S.n4747 0.05
R6235 S.n3948 S.n3947 0.05
R6236 S.n3953 S.n3934 0.05
R6237 S.n3136 S.n3135 0.05
R6238 S.n2301 S.n2300 0.05
R6239 S.n2306 S.n2287 0.05
R6240 S.n1378 S.n1377 0.05
R6241 S.n851 S.n835 0.05
R6242 S.n813 S.n812 0.05
R6243 S.n1265 S.n1264 0.049
R6244 S.n2545 S.n2544 0.049
R6245 S.n3401 S.n3400 0.049
R6246 S.n4248 S.n4247 0.049
R6247 S.n5038 S.n5037 0.049
R6248 S.n5819 S.n5818 0.049
R6249 S.n6574 S.n6573 0.049
R6250 S.n7320 S.n7319 0.049
R6251 S.n7873 S.n7872 0.049
R6252 S.n8569 S.n8568 0.049
R6253 S.n9436 S.n9435 0.049
R6254 S.n10112 S.n10111 0.049
R6255 S.n10765 S.n10764 0.049
R6256 S.n687 S.n686 0.049
R6257 S.n706 S.n705 0.049
R6258 S.n11029 S.n11027 0.049
R6259 S.n11632 S.n11631 0.048
R6260 S.n996 S.n995 0.048
R6261 S.n1840 S.n1839 0.048
R6262 S.n2723 S.n2722 0.048
R6263 S.n3564 S.n3563 0.048
R6264 S.n4396 S.n4395 0.048
R6265 S.n5202 S.n5201 0.048
R6266 S.n5999 S.n5998 0.048
R6267 S.n6770 S.n6769 0.048
R6268 S.n7532 S.n7531 0.048
R6269 S.n8268 S.n8267 0.048
R6270 S.n8995 S.n8994 0.048
R6271 S.n9696 S.n9695 0.048
R6272 S.n10388 S.n10387 0.048
R6273 S.n11047 S.n11046 0.048
R6274 S.n4 S.n3 0.047
R6275 S.n15 S.n14 0.047
R6276 S.n26 S.n25 0.047
R6277 S.n38 S.n37 0.047
R6278 S.n70 S.n69 0.047
R6279 S.n82 S.n81 0.047
R6280 S.n12640 S.n12638 0.047
R6281 S.n12564 S.n12562 0.047
R6282 S.n12009 S.n12000 0.047
R6283 S.n12306 S.n12278 0.047
R6284 S.n851 S.n844 0.047
R6285 S.n823 S.n821 0.047
R6286 S.n1785 S.n1774 0.047
R6287 S.n12591 S.n12576 0.047
R6288 S.n11985 S.n11977 0.047
R6289 S.n11692 S.n11680 0.047
R6290 S.n11433 S.n11425 0.047
R6291 S.n11095 S.n11083 0.047
R6292 S.n10812 S.n10804 0.047
R6293 S.n10470 S.n10458 0.047
R6294 S.n10159 S.n10151 0.047
R6295 S.n9810 S.n9798 0.047
R6296 S.n9483 S.n9475 0.047
R6297 S.n9138 S.n9126 0.047
R6298 S.n8616 S.n8608 0.047
R6299 S.n8443 S.n8431 0.047
R6300 S.n7920 S.n7912 0.047
R6301 S.n7736 S.n7724 0.047
R6302 S.n7367 S.n7359 0.047
R6303 S.n7006 S.n6994 0.047
R6304 S.n6621 S.n6613 0.047
R6305 S.n6264 S.n6252 0.047
R6306 S.n5866 S.n5858 0.047
R6307 S.n5499 S.n5487 0.047
R6308 S.n5085 S.n5077 0.047
R6309 S.n4722 S.n4710 0.047
R6310 S.n4295 S.n4287 0.047
R6311 S.n3922 S.n3910 0.047
R6312 S.n3448 S.n3440 0.047
R6313 S.n3110 S.n3098 0.047
R6314 S.n2592 S.n2584 0.047
R6315 S.n2275 S.n2261 0.047
R6316 S.n1310 S.n1304 0.047
R6317 S.n729 S.n727 0.047
R6318 S.n426 S.n424 0.047
R6319 S.n1673 S.n1663 0.047
R6320 S.n9164 S.n9150 0.047
R6321 S.n8520 S.n8512 0.047
R6322 S.n8296 S.n8284 0.047
R6323 S.n7824 S.n7816 0.047
R6324 S.n7589 S.n7577 0.047
R6325 S.n7271 S.n7263 0.047
R6326 S.n6859 S.n6847 0.047
R6327 S.n6525 S.n6517 0.047
R6328 S.n6117 S.n6105 0.047
R6329 S.n5770 S.n5762 0.047
R6330 S.n5352 S.n5340 0.047
R6331 S.n4989 S.n4981 0.047
R6332 S.n4575 S.n4563 0.047
R6333 S.n4199 S.n4191 0.047
R6334 S.n3775 S.n3763 0.047
R6335 S.n3352 S.n3344 0.047
R6336 S.n2963 S.n2951 0.047
R6337 S.n2496 S.n2488 0.047
R6338 S.n2122 S.n2108 0.047
R6339 S.n1213 S.n1207 0.047
R6340 S.n446 S.n444 0.047
R6341 S.n9841 S.n9832 0.047
R6342 S.n9404 S.n9402 0.047
R6343 S.n9020 S.n9009 0.047
R6344 S.n8537 S.n8535 0.047
R6345 S.n8325 S.n8314 0.047
R6346 S.n7841 S.n7839 0.047
R6347 S.n7618 S.n7607 0.047
R6348 S.n7288 S.n7286 0.047
R6349 S.n6888 S.n6877 0.047
R6350 S.n6542 S.n6540 0.047
R6351 S.n6146 S.n6135 0.047
R6352 S.n5787 S.n5785 0.047
R6353 S.n5381 S.n5370 0.047
R6354 S.n5006 S.n5004 0.047
R6355 S.n4604 S.n4593 0.047
R6356 S.n4216 S.n4214 0.047
R6357 S.n3804 S.n3793 0.047
R6358 S.n3369 S.n3367 0.047
R6359 S.n2992 S.n2981 0.047
R6360 S.n2513 S.n2511 0.047
R6361 S.n2151 S.n2140 0.047
R6362 S.n1232 S.n1228 0.047
R6363 S.n1252 S.n1247 0.047
R6364 S.n765 S.n763 0.047
R6365 S.n780 S.n774 0.047
R6366 S.n2186 S.n2172 0.047
R6367 S.n3024 S.n3012 0.047
R6368 S.n3836 S.n3824 0.047
R6369 S.n4636 S.n4624 0.047
R6370 S.n5413 S.n5401 0.047
R6371 S.n6178 S.n6166 0.047
R6372 S.n6920 S.n6908 0.047
R6373 S.n7650 S.n7638 0.047
R6374 S.n8357 S.n8345 0.047
R6375 S.n9052 S.n9040 0.047
R6376 S.n9724 S.n9712 0.047
R6377 S.n10499 S.n10485 0.047
R6378 S.n10099 S.n10091 0.047
R6379 S.n9423 S.n9415 0.047
R6380 S.n8556 S.n8548 0.047
R6381 S.n7860 S.n7852 0.047
R6382 S.n7307 S.n7299 0.047
R6383 S.n6561 S.n6553 0.047
R6384 S.n5806 S.n5798 0.047
R6385 S.n5025 S.n5017 0.047
R6386 S.n4235 S.n4227 0.047
R6387 S.n3388 S.n3380 0.047
R6388 S.n2532 S.n2524 0.047
R6389 S.n1735 S.n1725 0.047
R6390 S.n690 S.n684 0.047
R6391 S.n901 S.n894 0.047
R6392 S.n11122 S.n11114 0.047
R6393 S.n10773 S.n10768 0.047
R6394 S.n10418 S.n10403 0.047
R6395 S.n10120 S.n10115 0.047
R6396 S.n9758 S.n9743 0.047
R6397 S.n9444 S.n9439 0.047
R6398 S.n9086 S.n9071 0.047
R6399 S.n8577 S.n8572 0.047
R6400 S.n8391 S.n8376 0.047
R6401 S.n7881 S.n7876 0.047
R6402 S.n7684 S.n7669 0.047
R6403 S.n7328 S.n7323 0.047
R6404 S.n6954 S.n6939 0.047
R6405 S.n6582 S.n6577 0.047
R6406 S.n6212 S.n6197 0.047
R6407 S.n5827 S.n5822 0.047
R6408 S.n5447 S.n5432 0.047
R6409 S.n5046 S.n5041 0.047
R6410 S.n4670 S.n4655 0.047
R6411 S.n4256 S.n4251 0.047
R6412 S.n3870 S.n3855 0.047
R6413 S.n3409 S.n3404 0.047
R6414 S.n3058 S.n3043 0.047
R6415 S.n2553 S.n2548 0.047
R6416 S.n2220 S.n2205 0.047
R6417 S.n1273 S.n1268 0.047
R6418 S.n1763 S.n1753 0.047
R6419 S.n709 S.n704 0.047
R6420 S.n1293 S.n1287 0.047
R6421 S.n2241 S.n2238 0.047
R6422 S.n2573 S.n2568 0.047
R6423 S.n3078 S.n3076 0.047
R6424 S.n3429 S.n3424 0.047
R6425 S.n3890 S.n3888 0.047
R6426 S.n4276 S.n4271 0.047
R6427 S.n4690 S.n4688 0.047
R6428 S.n5066 S.n5061 0.047
R6429 S.n5467 S.n5465 0.047
R6430 S.n5847 S.n5842 0.047
R6431 S.n6232 S.n6230 0.047
R6432 S.n6602 S.n6597 0.047
R6433 S.n6974 S.n6972 0.047
R6434 S.n7348 S.n7343 0.047
R6435 S.n7704 S.n7702 0.047
R6436 S.n7901 S.n7896 0.047
R6437 S.n8411 S.n8409 0.047
R6438 S.n8597 S.n8592 0.047
R6439 S.n9106 S.n9104 0.047
R6440 S.n9464 S.n9459 0.047
R6441 S.n9778 S.n9776 0.047
R6442 S.n10140 S.n10135 0.047
R6443 S.n10438 S.n10436 0.047
R6444 S.n10793 S.n10788 0.047
R6445 S.n11063 S.n11061 0.047
R6446 S.n11414 S.n11409 0.047
R6447 S.n11717 S.n11715 0.047
R6448 S.n802 S.n794 0.047
R6449 S.n1701 S.n1691 0.047
R6450 S.n670 S.n668 0.047
R6451 S.n653 S.n651 0.047
R6452 S.n385 S.n383 0.047
R6453 S.n1614 S.n1604 0.047
R6454 S.n7762 S.n7748 0.047
R6455 S.n7235 S.n7227 0.047
R6456 S.n6798 S.n6786 0.047
R6457 S.n6489 S.n6481 0.047
R6458 S.n6056 S.n6044 0.047
R6459 S.n5734 S.n5726 0.047
R6460 S.n5291 S.n5279 0.047
R6461 S.n4953 S.n4945 0.047
R6462 S.n4514 S.n4502 0.047
R6463 S.n4163 S.n4155 0.047
R6464 S.n3714 S.n3702 0.047
R6465 S.n3316 S.n3308 0.047
R6466 S.n2902 S.n2890 0.047
R6467 S.n2460 S.n2452 0.047
R6468 S.n2059 S.n2045 0.047
R6469 S.n1179 S.n1173 0.047
R6470 S.n405 S.n403 0.047
R6471 S.n8474 S.n8465 0.047
R6472 S.n7805 S.n7803 0.047
R6473 S.n7557 S.n7546 0.047
R6474 S.n7252 S.n7250 0.047
R6475 S.n6827 S.n6816 0.047
R6476 S.n6506 S.n6504 0.047
R6477 S.n6085 S.n6074 0.047
R6478 S.n5751 S.n5749 0.047
R6479 S.n5320 S.n5309 0.047
R6480 S.n4970 S.n4968 0.047
R6481 S.n4543 S.n4532 0.047
R6482 S.n4180 S.n4178 0.047
R6483 S.n3743 S.n3732 0.047
R6484 S.n3333 S.n3331 0.047
R6485 S.n2931 S.n2920 0.047
R6486 S.n2477 S.n2475 0.047
R6487 S.n2088 S.n2077 0.047
R6488 S.n1196 S.n1194 0.047
R6489 S.n1643 S.n1632 0.047
R6490 S.n637 S.n635 0.047
R6491 S.n620 S.n618 0.047
R6492 S.n344 S.n342 0.047
R6493 S.n1555 S.n1545 0.047
R6494 S.n6290 S.n6276 0.047
R6495 S.n5698 S.n5690 0.047
R6496 S.n5230 S.n5218 0.047
R6497 S.n4917 S.n4909 0.047
R6498 S.n4453 S.n4441 0.047
R6499 S.n4127 S.n4119 0.047
R6500 S.n3653 S.n3641 0.047
R6501 S.n3280 S.n3272 0.047
R6502 S.n2841 S.n2829 0.047
R6503 S.n2424 S.n2416 0.047
R6504 S.n1996 S.n1982 0.047
R6505 S.n1145 S.n1139 0.047
R6506 S.n364 S.n362 0.047
R6507 S.n7037 S.n7028 0.047
R6508 S.n6470 S.n6468 0.047
R6509 S.n6024 S.n6013 0.047
R6510 S.n5715 S.n5713 0.047
R6511 S.n5259 S.n5248 0.047
R6512 S.n4934 S.n4932 0.047
R6513 S.n4482 S.n4471 0.047
R6514 S.n4144 S.n4142 0.047
R6515 S.n3682 S.n3671 0.047
R6516 S.n3297 S.n3295 0.047
R6517 S.n2870 S.n2859 0.047
R6518 S.n2441 S.n2439 0.047
R6519 S.n2025 S.n2014 0.047
R6520 S.n1162 S.n1160 0.047
R6521 S.n1584 S.n1573 0.047
R6522 S.n604 S.n602 0.047
R6523 S.n587 S.n585 0.047
R6524 S.n323 S.n321 0.047
R6525 S.n1496 S.n1486 0.047
R6526 S.n4748 S.n4734 0.047
R6527 S.n4091 S.n4083 0.047
R6528 S.n3592 S.n3580 0.047
R6529 S.n3244 S.n3236 0.047
R6530 S.n2780 S.n2768 0.047
R6531 S.n2388 S.n2380 0.047
R6532 S.n1933 S.n1919 0.047
R6533 S.n1111 S.n1105 0.047
R6534 S.n59 S.n57 0.047
R6535 S.n5530 S.n5521 0.047
R6536 S.n4898 S.n4896 0.047
R6537 S.n4421 S.n4410 0.047
R6538 S.n4108 S.n4106 0.047
R6539 S.n3621 S.n3610 0.047
R6540 S.n3261 S.n3259 0.047
R6541 S.n2809 S.n2798 0.047
R6542 S.n2405 S.n2403 0.047
R6543 S.n1962 S.n1951 0.047
R6544 S.n1128 S.n1126 0.047
R6545 S.n1525 S.n1514 0.047
R6546 S.n571 S.n569 0.047
R6547 S.n554 S.n552 0.047
R6548 S.n282 S.n280 0.047
R6549 S.n1437 S.n1427 0.047
R6550 S.n3136 S.n3122 0.047
R6551 S.n2352 S.n2344 0.047
R6552 S.n1870 S.n1856 0.047
R6553 S.n1077 S.n1071 0.047
R6554 S.n302 S.n300 0.047
R6555 S.n3953 S.n3944 0.047
R6556 S.n3225 S.n3223 0.047
R6557 S.n2748 S.n2737 0.047
R6558 S.n2369 S.n2367 0.047
R6559 S.n1899 S.n1888 0.047
R6560 S.n1094 S.n1092 0.047
R6561 S.n1469 S.n1458 0.047
R6562 S.n538 S.n536 0.047
R6563 S.n521 S.n519 0.047
R6564 S.n241 S.n239 0.047
R6565 S.n1378 S.n1366 0.047
R6566 S.n261 S.n259 0.047
R6567 S.n2306 S.n2297 0.047
R6568 S.n1060 S.n1058 0.047
R6569 S.n1407 S.n1396 0.047
R6570 S.n505 S.n503 0.047
R6571 S.n488 S.n486 0.047
R6572 S.n880 S.n875 0.047
R6573 S.n748 S.n744 0.047
R6574 S.n1355 S.n1353 0.047
R6575 S.n1346 S.n1342 0.047
R6576 S.n2646 S.n2640 0.047
R6577 S.n2632 S.n2628 0.047
R6578 S.n3173 S.n3167 0.047
R6579 S.n3159 S.n3155 0.047
R6580 S.n3990 S.n3984 0.047
R6581 S.n3976 S.n3972 0.047
R6582 S.n4785 S.n4779 0.047
R6583 S.n4771 S.n4767 0.047
R6584 S.n5567 S.n5561 0.047
R6585 S.n5553 S.n5549 0.047
R6586 S.n6327 S.n6321 0.047
R6587 S.n6313 S.n6309 0.047
R6588 S.n7074 S.n7068 0.047
R6589 S.n7060 S.n7056 0.047
R6590 S.n8085 S.n8079 0.047
R6591 S.n8071 S.n8067 0.047
R6592 S.n8797 S.n8791 0.047
R6593 S.n8783 S.n8779 0.047
R6594 S.n9201 S.n9195 0.047
R6595 S.n9187 S.n9183 0.047
R6596 S.n9878 S.n9872 0.047
R6597 S.n9864 S.n9860 0.047
R6598 S.n10536 S.n10530 0.047
R6599 S.n10522 S.n10518 0.047
R6600 S.n11159 S.n11153 0.047
R6601 S.n11145 S.n11141 0.047
R6602 S.n11737 S.n11731 0.047
R6603 S.n12027 S.n12023 0.047
R6604 S.n12906 S.n12900 0.047
R6605 S.n12891 S.n12887 0.047
R6606 S.n1808 S.n1803 0.047
R6607 S.n1327 S.n1325 0.047
R6608 S.n2676 S.n2657 0.047
R6609 S.n12935 S.n12925 0.047
R6610 S.n12937 S.n12917 0.047
R6611 S.n12042 S.n12038 0.047
R6612 S.n11753 S.n11748 0.047
R6613 S.n11188 S.n11178 0.047
R6614 S.n11190 S.n11170 0.047
R6615 S.n10565 S.n10555 0.047
R6616 S.n10567 S.n10547 0.047
R6617 S.n9907 S.n9897 0.047
R6618 S.n9909 S.n9889 0.047
R6619 S.n9230 S.n9220 0.047
R6620 S.n9232 S.n9212 0.047
R6621 S.n8826 S.n8816 0.047
R6622 S.n8828 S.n8808 0.047
R6623 S.n8114 S.n8104 0.047
R6624 S.n8116 S.n8096 0.047
R6625 S.n7103 S.n7093 0.047
R6626 S.n7105 S.n7085 0.047
R6627 S.n6356 S.n6346 0.047
R6628 S.n6358 S.n6338 0.047
R6629 S.n5596 S.n5586 0.047
R6630 S.n5598 S.n5578 0.047
R6631 S.n4814 S.n4804 0.047
R6632 S.n4816 S.n4796 0.047
R6633 S.n4022 S.n4012 0.047
R6634 S.n4024 S.n4004 0.047
R6635 S.n3500 S.n3192 0.047
R6636 S.n3502 S.n3184 0.047
R6637 S.n2675 S.n2665 0.047
R6638 S.n2692 S.n1842 0.047
R6639 S.n2613 S.n2607 0.047
R6640 S.n3517 S.n3513 0.047
R6641 S.n12680 S.n12675 0.047
R6642 S.n12952 S.n12948 0.047
R6643 S.n12058 S.n12053 0.047
R6644 S.n11768 S.n11764 0.047
R6645 S.n11450 S.n11445 0.047
R6646 S.n11205 S.n11201 0.047
R6647 S.n10829 S.n10824 0.047
R6648 S.n10582 S.n10578 0.047
R6649 S.n10176 S.n10171 0.047
R6650 S.n9924 S.n9920 0.047
R6651 S.n9500 S.n9495 0.047
R6652 S.n9247 S.n9243 0.047
R6653 S.n8633 S.n8628 0.047
R6654 S.n8843 S.n8839 0.047
R6655 S.n7937 S.n7932 0.047
R6656 S.n8131 S.n8127 0.047
R6657 S.n7384 S.n7379 0.047
R6658 S.n7120 S.n7116 0.047
R6659 S.n6638 S.n6633 0.047
R6660 S.n6373 S.n6369 0.047
R6661 S.n5883 S.n5878 0.047
R6662 S.n5613 S.n5609 0.047
R6663 S.n5102 S.n5097 0.047
R6664 S.n4831 S.n4827 0.047
R6665 S.n4312 S.n4307 0.047
R6666 S.n4036 S.n4032 0.047
R6667 S.n3464 S.n3460 0.047
R6668 S.n3533 S.n2725 0.047
R6669 S.n3484 S.n3478 0.047
R6670 S.n4349 S.n4047 0.047
R6671 S.n12696 S.n12691 0.047
R6672 S.n12967 S.n12963 0.047
R6673 S.n12074 S.n12069 0.047
R6674 S.n11783 S.n11779 0.047
R6675 S.n11466 S.n11461 0.047
R6676 S.n11220 S.n11216 0.047
R6677 S.n10845 S.n10840 0.047
R6678 S.n10597 S.n10593 0.047
R6679 S.n10192 S.n10187 0.047
R6680 S.n9939 S.n9935 0.047
R6681 S.n9516 S.n9511 0.047
R6682 S.n9262 S.n9258 0.047
R6683 S.n8649 S.n8644 0.047
R6684 S.n8858 S.n8854 0.047
R6685 S.n7953 S.n7948 0.047
R6686 S.n8146 S.n8142 0.047
R6687 S.n7400 S.n7395 0.047
R6688 S.n7135 S.n7131 0.047
R6689 S.n6654 S.n6649 0.047
R6690 S.n6388 S.n6384 0.047
R6691 S.n5899 S.n5894 0.047
R6692 S.n5628 S.n5624 0.047
R6693 S.n5118 S.n5113 0.047
R6694 S.n4846 S.n4842 0.047
R6695 S.n4348 S.n4055 0.047
R6696 S.n4365 S.n3566 0.047
R6697 S.n4332 S.n4326 0.047
R6698 S.n5155 S.n4857 0.047
R6699 S.n12712 S.n12707 0.047
R6700 S.n12982 S.n12978 0.047
R6701 S.n12090 S.n12085 0.047
R6702 S.n11798 S.n11794 0.047
R6703 S.n11482 S.n11477 0.047
R6704 S.n11235 S.n11231 0.047
R6705 S.n10861 S.n10856 0.047
R6706 S.n10612 S.n10608 0.047
R6707 S.n10208 S.n10203 0.047
R6708 S.n9954 S.n9950 0.047
R6709 S.n9532 S.n9527 0.047
R6710 S.n9277 S.n9273 0.047
R6711 S.n8665 S.n8660 0.047
R6712 S.n8873 S.n8869 0.047
R6713 S.n7969 S.n7964 0.047
R6714 S.n8161 S.n8157 0.047
R6715 S.n7416 S.n7411 0.047
R6716 S.n7150 S.n7146 0.047
R6717 S.n6670 S.n6665 0.047
R6718 S.n6403 S.n6399 0.047
R6719 S.n5915 S.n5910 0.047
R6720 S.n5643 S.n5639 0.047
R6721 S.n5154 S.n4865 0.047
R6722 S.n5171 S.n4398 0.047
R6723 S.n5138 S.n5132 0.047
R6724 S.n5952 S.n5654 0.047
R6725 S.n12728 S.n12723 0.047
R6726 S.n12997 S.n12993 0.047
R6727 S.n12106 S.n12101 0.047
R6728 S.n11813 S.n11809 0.047
R6729 S.n11498 S.n11493 0.047
R6730 S.n11250 S.n11246 0.047
R6731 S.n10877 S.n10872 0.047
R6732 S.n10627 S.n10623 0.047
R6733 S.n10224 S.n10219 0.047
R6734 S.n9969 S.n9965 0.047
R6735 S.n9548 S.n9543 0.047
R6736 S.n9292 S.n9288 0.047
R6737 S.n8681 S.n8676 0.047
R6738 S.n8888 S.n8884 0.047
R6739 S.n7985 S.n7980 0.047
R6740 S.n8176 S.n8172 0.047
R6741 S.n7432 S.n7427 0.047
R6742 S.n7165 S.n7161 0.047
R6743 S.n6686 S.n6681 0.047
R6744 S.n6418 S.n6414 0.047
R6745 S.n5951 S.n5662 0.047
R6746 S.n5968 S.n5204 0.047
R6747 S.n5935 S.n5929 0.047
R6748 S.n6723 S.n6429 0.047
R6749 S.n12744 S.n12739 0.047
R6750 S.n13012 S.n13008 0.047
R6751 S.n12122 S.n12117 0.047
R6752 S.n11828 S.n11824 0.047
R6753 S.n11514 S.n11509 0.047
R6754 S.n11265 S.n11261 0.047
R6755 S.n10893 S.n10888 0.047
R6756 S.n10642 S.n10638 0.047
R6757 S.n10240 S.n10235 0.047
R6758 S.n9984 S.n9980 0.047
R6759 S.n9564 S.n9559 0.047
R6760 S.n9307 S.n9303 0.047
R6761 S.n8697 S.n8692 0.047
R6762 S.n8903 S.n8899 0.047
R6763 S.n8001 S.n7996 0.047
R6764 S.n8191 S.n8187 0.047
R6765 S.n7448 S.n7443 0.047
R6766 S.n7180 S.n7176 0.047
R6767 S.n6722 S.n6437 0.047
R6768 S.n6739 S.n6001 0.047
R6769 S.n6706 S.n6700 0.047
R6770 S.n7485 S.n7191 0.047
R6771 S.n12760 S.n12755 0.047
R6772 S.n13027 S.n13023 0.047
R6773 S.n12138 S.n12133 0.047
R6774 S.n11843 S.n11839 0.047
R6775 S.n11530 S.n11525 0.047
R6776 S.n11280 S.n11276 0.047
R6777 S.n10909 S.n10904 0.047
R6778 S.n10657 S.n10653 0.047
R6779 S.n10256 S.n10251 0.047
R6780 S.n9999 S.n9995 0.047
R6781 S.n9580 S.n9575 0.047
R6782 S.n9322 S.n9318 0.047
R6783 S.n8713 S.n8708 0.047
R6784 S.n8918 S.n8914 0.047
R6785 S.n8017 S.n8012 0.047
R6786 S.n8206 S.n8202 0.047
R6787 S.n7484 S.n7199 0.047
R6788 S.n7501 S.n6772 0.047
R6789 S.n7468 S.n7462 0.047
R6790 S.n8221 S.n8217 0.047
R6791 S.n12776 S.n12771 0.047
R6792 S.n13042 S.n13038 0.047
R6793 S.n12154 S.n12149 0.047
R6794 S.n11858 S.n11854 0.047
R6795 S.n11546 S.n11541 0.047
R6796 S.n11295 S.n11291 0.047
R6797 S.n10925 S.n10920 0.047
R6798 S.n10672 S.n10668 0.047
R6799 S.n10272 S.n10267 0.047
R6800 S.n10014 S.n10010 0.047
R6801 S.n9596 S.n9591 0.047
R6802 S.n9337 S.n9333 0.047
R6803 S.n8729 S.n8724 0.047
R6804 S.n8933 S.n8929 0.047
R6805 S.n8032 S.n8028 0.047
R6806 S.n8237 S.n7534 0.047
R6807 S.n8052 S.n8046 0.047
R6808 S.n8948 S.n8944 0.047
R6809 S.n12792 S.n12787 0.047
R6810 S.n13057 S.n13053 0.047
R6811 S.n12170 S.n12165 0.047
R6812 S.n11873 S.n11869 0.047
R6813 S.n11562 S.n11557 0.047
R6814 S.n11310 S.n11306 0.047
R6815 S.n10941 S.n10936 0.047
R6816 S.n10687 S.n10683 0.047
R6817 S.n10288 S.n10283 0.047
R6818 S.n10029 S.n10025 0.047
R6819 S.n9612 S.n9607 0.047
R6820 S.n9352 S.n9348 0.047
R6821 S.n8744 S.n8740 0.047
R6822 S.n8964 S.n8270 0.047
R6823 S.n8764 S.n8758 0.047
R6824 S.n9649 S.n9363 0.047
R6825 S.n12808 S.n12803 0.047
R6826 S.n13072 S.n13068 0.047
R6827 S.n12186 S.n12181 0.047
R6828 S.n11888 S.n11884 0.047
R6829 S.n11578 S.n11573 0.047
R6830 S.n11325 S.n11321 0.047
R6831 S.n10957 S.n10952 0.047
R6832 S.n10702 S.n10698 0.047
R6833 S.n10304 S.n10299 0.047
R6834 S.n10044 S.n10040 0.047
R6835 S.n9648 S.n9371 0.047
R6836 S.n9665 S.n8997 0.047
R6837 S.n9632 S.n9626 0.047
R6838 S.n10341 S.n10055 0.047
R6839 S.n12824 S.n12819 0.047
R6840 S.n13087 S.n13083 0.047
R6841 S.n12202 S.n12197 0.047
R6842 S.n11903 S.n11899 0.047
R6843 S.n11594 S.n11589 0.047
R6844 S.n11340 S.n11336 0.047
R6845 S.n10973 S.n10968 0.047
R6846 S.n10717 S.n10713 0.047
R6847 S.n10340 S.n10063 0.047
R6848 S.n10357 S.n9698 0.047
R6849 S.n10324 S.n10318 0.047
R6850 S.n11010 S.n10728 0.047
R6851 S.n12840 S.n12835 0.047
R6852 S.n13102 S.n13098 0.047
R6853 S.n12218 S.n12213 0.047
R6854 S.n11918 S.n11914 0.047
R6855 S.n11610 S.n11605 0.047
R6856 S.n11355 S.n11351 0.047
R6857 S.n11009 S.n10736 0.047
R6858 S.n11026 S.n10390 0.047
R6859 S.n10993 S.n10987 0.047
R6860 S.n11650 S.n11366 0.047
R6861 S.n12856 S.n12851 0.047
R6862 S.n13117 S.n13113 0.047
R6863 S.n12234 S.n12229 0.047
R6864 S.n11933 S.n11929 0.047
R6865 S.n11649 S.n11374 0.047
R6866 S.n11666 S.n11049 0.047
R6867 S.n11633 S.n11622 0.047
R6868 S.n12265 S.n12262 0.047
R6869 S.n12872 S.n12870 0.047
R6870 S.n13135 S.n13133 0.047
R6871 S.n12251 S.n12249 0.047
R6872 S.n12663 S.n12661 0.047
R6873 S.n13161 S.n13148 0.047
R6874 S.n1007 S.n1002 0.047
R6875 S.n9708 S.n9707 0.047
R6876 S.n9036 S.n9035 0.047
R6877 S.n8341 S.n8340 0.047
R6878 S.n7634 S.n7633 0.047
R6879 S.n6904 S.n6903 0.047
R6880 S.n6162 S.n6161 0.047
R6881 S.n5397 S.n5396 0.047
R6882 S.n4620 S.n4619 0.047
R6883 S.n3820 S.n3819 0.047
R6884 S.n3008 S.n3007 0.047
R6885 S.n2168 S.n2167 0.047
R6886 S.n925 S.n924 0.046
R6887 S.t28 S.n207 0.046
R6888 S.t28 S.n197 0.046
R6889 S.t28 S.n185 0.046
R6890 S.t28 S.n173 0.046
R6891 S.t28 S.n160 0.046
R6892 S.t28 S.n147 0.046
R6893 S.t28 S.n134 0.046
R6894 S.n1355 S.n1346 0.046
R6895 S.n2676 S.n2675 0.046
R6896 S.n4349 S.n4348 0.045
R6897 S.n5155 S.n5154 0.045
R6898 S.n5952 S.n5951 0.045
R6899 S.n6723 S.n6722 0.045
R6900 S.n7485 S.n7484 0.045
R6901 S.n9649 S.n9648 0.045
R6902 S.n10341 S.n10340 0.045
R6903 S.n11010 S.n11009 0.045
R6904 S.n11650 S.n11649 0.045
R6905 S.n214 S.n212 0.045
R6906 S.n12264 S.n12263 0.045
R6907 S.n12327 S.n12326 0.045
R6908 S.n12466 S.n12465 0.045
R6909 S.n222 S.n221 0.045
R6910 S.n1716 S.n1708 0.045
R6911 S.n2217 S.n2209 0.045
R6912 S.n3055 S.n3047 0.045
R6913 S.n3867 S.n3859 0.045
R6914 S.n4667 S.n4659 0.045
R6915 S.n5444 S.n5436 0.045
R6916 S.n6209 S.n6201 0.045
R6917 S.n6951 S.n6943 0.045
R6918 S.n7681 S.n7673 0.045
R6919 S.n8388 S.n8380 0.045
R6920 S.n9083 S.n9075 0.045
R6921 S.n9755 S.n9747 0.045
R6922 S.n10415 S.n10407 0.045
R6923 S.n1813 S.n1812 0.045
R6924 S.n2696 S.n2695 0.045
R6925 S.n3537 S.n3536 0.045
R6926 S.n4369 S.n4368 0.045
R6927 S.n5175 S.n5174 0.045
R6928 S.n5972 S.n5971 0.045
R6929 S.n6743 S.n6742 0.045
R6930 S.n7505 S.n7504 0.045
R6931 S.n8241 S.n8240 0.045
R6932 S.n8968 S.n8967 0.045
R6933 S.n9669 S.n9668 0.045
R6934 S.n10361 S.n10360 0.045
R6935 S.n12317 S.n12316 0.045
R6936 S.n12265 S.n12251 0.044
R6937 S.n917 S.n916 0.044
R6938 S.n2646 S.n2633 0.044
R6939 S.n3173 S.n3160 0.044
R6940 S.n3990 S.n3977 0.044
R6941 S.n4785 S.n4772 0.044
R6942 S.n5567 S.n5554 0.044
R6943 S.n6327 S.n6314 0.044
R6944 S.n7074 S.n7061 0.044
R6945 S.n8085 S.n8072 0.044
R6946 S.n8797 S.n8784 0.044
R6947 S.n9201 S.n9188 0.044
R6948 S.n9878 S.n9865 0.044
R6949 S.n10536 S.n10523 0.044
R6950 S.n11159 S.n11146 0.044
R6951 S.n11737 S.n11724 0.044
R6952 S.n12906 S.n12893 0.044
R6953 S.n3502 S.n3501 0.044
R6954 S.n4024 S.n4023 0.044
R6955 S.n4816 S.n4815 0.044
R6956 S.n5598 S.n5597 0.044
R6957 S.n6358 S.n6357 0.044
R6958 S.n7105 S.n7104 0.044
R6959 S.n8116 S.n8115 0.044
R6960 S.n8828 S.n8827 0.044
R6961 S.n9232 S.n9231 0.044
R6962 S.n9909 S.n9908 0.044
R6963 S.n10567 S.n10566 0.044
R6964 S.n11190 S.n11189 0.044
R6965 S.n11753 S.n11752 0.044
R6966 S.n12937 S.n12936 0.044
R6967 S.n12391 S.n12389 0.044
R6968 S.n437 S.n436 0.044
R6969 S.n396 S.n395 0.044
R6970 S.n355 S.n354 0.044
R6971 S.n44 S.n43 0.044
R6972 S.n293 S.n292 0.044
R6973 S.n252 S.n251 0.044
R6974 S.n12590 S.n12589 0.043
R6975 S.n11704 S.n11703 0.043
R6976 S.n1669 S.n1668 0.043
R6977 S.n1610 S.n1609 0.043
R6978 S.n1551 S.n1550 0.043
R6979 S.n1492 S.n1491 0.043
R6980 S.n1016 S.n1015 0.043
R6981 S.n929 S.n928 0.043
R6982 S.n1684 S.n1683 0.042
R6983 S.n2132 S.n2131 0.042
R6984 S.n2973 S.n2972 0.042
R6985 S.n3785 S.n3784 0.042
R6986 S.n4585 S.n4584 0.042
R6987 S.n5362 S.n5361 0.042
R6988 S.n6127 S.n6126 0.042
R6989 S.n6869 S.n6868 0.042
R6990 S.n7599 S.n7598 0.042
R6991 S.n8306 S.n8305 0.042
R6992 S.n9001 S.n9000 0.042
R6993 S.n1625 S.n1624 0.042
R6994 S.n2069 S.n2068 0.042
R6995 S.n2912 S.n2911 0.042
R6996 S.n3724 S.n3723 0.042
R6997 S.n4524 S.n4523 0.042
R6998 S.n5301 S.n5300 0.042
R6999 S.n6066 S.n6065 0.042
R7000 S.n6808 S.n6807 0.042
R7001 S.n7538 S.n7537 0.042
R7002 S.n1566 S.n1565 0.042
R7003 S.n2006 S.n2005 0.042
R7004 S.n2851 S.n2850 0.042
R7005 S.n3663 S.n3662 0.042
R7006 S.n4463 S.n4462 0.042
R7007 S.n5240 S.n5239 0.042
R7008 S.n6005 S.n6004 0.042
R7009 S.n1507 S.n1506 0.042
R7010 S.n1943 S.n1942 0.042
R7011 S.n2790 S.n2789 0.042
R7012 S.n3602 S.n3601 0.042
R7013 S.n4402 S.n4401 0.042
R7014 S.n1448 S.n1447 0.042
R7015 S.n1880 S.n1879 0.042
R7016 S.n2729 S.n2728 0.042
R7017 S.n1389 S.n1388 0.042
R7018 S.n11688 S.n11685 0.042
R7019 S.n11091 S.n11088 0.042
R7020 S.n10466 S.n10463 0.042
R7021 S.n9806 S.n9803 0.042
R7022 S.n9134 S.n9131 0.042
R7023 S.n8439 S.n8436 0.042
R7024 S.n7732 S.n7729 0.042
R7025 S.n7002 S.n6999 0.042
R7026 S.n6260 S.n6257 0.042
R7027 S.n5495 S.n5492 0.042
R7028 S.n4718 S.n4715 0.042
R7029 S.n3918 S.n3915 0.042
R7030 S.n3106 S.n3103 0.042
R7031 S.n2271 S.n2266 0.042
R7032 S.n1781 S.n1779 0.042
R7033 S.n720 S.n719 0.042
R7034 S.n8292 S.n8289 0.042
R7035 S.n7585 S.n7582 0.042
R7036 S.n6855 S.n6852 0.042
R7037 S.n6113 S.n6110 0.042
R7038 S.n5348 S.n5345 0.042
R7039 S.n4571 S.n4568 0.042
R7040 S.n3771 S.n3768 0.042
R7041 S.n2959 S.n2956 0.042
R7042 S.n2118 S.n2113 0.042
R7043 S.n9720 S.n9717 0.042
R7044 S.n9048 S.n9045 0.042
R7045 S.n8353 S.n8350 0.042
R7046 S.n7646 S.n7643 0.042
R7047 S.n6916 S.n6913 0.042
R7048 S.n6174 S.n6171 0.042
R7049 S.n5409 S.n5406 0.042
R7050 S.n4632 S.n4629 0.042
R7051 S.n3832 S.n3829 0.042
R7052 S.n3020 S.n3017 0.042
R7053 S.n2182 S.n2177 0.042
R7054 S.n6794 S.n6791 0.042
R7055 S.n6052 S.n6049 0.042
R7056 S.n5287 S.n5284 0.042
R7057 S.n4510 S.n4507 0.042
R7058 S.n3710 S.n3707 0.042
R7059 S.n2898 S.n2895 0.042
R7060 S.n2055 S.n2050 0.042
R7061 S.n5226 S.n5223 0.042
R7062 S.n4449 S.n4446 0.042
R7063 S.n3649 S.n3646 0.042
R7064 S.n2837 S.n2834 0.042
R7065 S.n1992 S.n1987 0.042
R7066 S.n3588 S.n3585 0.042
R7067 S.n2776 S.n2773 0.042
R7068 S.n1929 S.n1924 0.042
R7069 S.n1866 S.n1861 0.042
R7070 S.n96 S.n95 0.042
R7071 S.n6 S.n5 0.042
R7072 S.n903 S.n902 0.042
R7073 S.n17 S.n16 0.042
R7074 S.n29 S.n28 0.042
R7075 S.n61 S.n60 0.042
R7076 S.n73 S.n72 0.042
R7077 S.n85 S.n84 0.042
R7078 S.n11053 S.n11052 0.042
R7079 S.n10428 S.n10427 0.042
R7080 S.n9768 S.n9767 0.042
R7081 S.n9096 S.n9095 0.042
R7082 S.n8401 S.n8400 0.042
R7083 S.n7694 S.n7693 0.042
R7084 S.n6964 S.n6963 0.042
R7085 S.n6222 S.n6221 0.042
R7086 S.n5457 S.n5456 0.042
R7087 S.n4680 S.n4679 0.042
R7088 S.n3880 S.n3879 0.042
R7089 S.n3068 S.n3067 0.042
R7090 S.n2230 S.n2229 0.042
R7091 S.n1745 S.n1744 0.042
R7092 S.n12608 S.n12607 0.042
R7093 S.n933 S.n932 0.041
R7094 S.n10482 S.n10481 0.041
R7095 S.n100 S.n99 0.041
R7096 S.n877 S.n876 0.041
R7097 S.n122 S.n108 0.04
R7098 S.n847 S.n846 0.04
R7099 S.n470 S.n461 0.04
R7100 S.n1040 S.n1031 0.04
R7101 S.n2331 S.n2322 0.04
R7102 S.n3205 S.n3196 0.04
R7103 S.n4070 S.n4061 0.04
R7104 S.n4878 S.n4869 0.04
R7105 S.n5677 S.n5668 0.04
R7106 S.n6450 S.n6441 0.04
R7107 S.n7214 S.n7205 0.04
R7108 S.n7785 S.n7776 0.04
R7109 S.n8499 S.n8490 0.04
R7110 S.n9384 S.n9375 0.04
R7111 S.n10078 S.n10069 0.04
R7112 S.n10749 S.n10740 0.04
R7113 S.n11392 S.n11383 0.04
R7114 S.n11963 S.n11954 0.04
R7115 S.n12420 S.n12419 0.04
R7116 S.n12418 S.n12417 0.04
R7117 S.n12416 S.n12415 0.04
R7118 S.n12414 S.n12413 0.04
R7119 S.n12412 S.n12411 0.04
R7120 S.n12410 S.n12409 0.04
R7121 S.n12408 S.n12407 0.04
R7122 S.n12406 S.n12405 0.04
R7123 S.n12404 S.n12403 0.04
R7124 S.n12402 S.n12401 0.04
R7125 S.n12400 S.n12399 0.04
R7126 S.n12398 S.n12397 0.04
R7127 S.n12396 S.n12395 0.04
R7128 S.n12394 S.n12393 0.04
R7129 S.n12377 S.n12376 0.039
R7130 S.n12373 S.n12372 0.039
R7131 S.n12369 S.n12368 0.039
R7132 S.n12365 S.n12364 0.039
R7133 S.n12361 S.n12360 0.039
R7134 S.n12357 S.n12356 0.039
R7135 S.n12353 S.n12352 0.039
R7136 S.n12349 S.n12348 0.039
R7137 S.n12345 S.n12344 0.039
R7138 S.n12341 S.n12340 0.039
R7139 S.n12337 S.n12336 0.039
R7140 S.n12333 S.n12332 0.039
R7141 S.n12330 S.n12329 0.039
R7142 S.n107 S.n106 0.039
R7143 S.n12295 S.n12294 0.039
R7144 S.n1814 S.n1813 0.039
R7145 S.n1819 S.n1818 0.039
R7146 S.n2697 S.n2696 0.039
R7147 S.n2702 S.n2701 0.039
R7148 S.n3538 S.n3537 0.039
R7149 S.n3543 S.n3542 0.039
R7150 S.n4370 S.n4369 0.039
R7151 S.n4375 S.n4374 0.039
R7152 S.n5176 S.n5175 0.039
R7153 S.n5181 S.n5180 0.039
R7154 S.n5973 S.n5972 0.039
R7155 S.n5978 S.n5977 0.039
R7156 S.n6744 S.n6743 0.039
R7157 S.n6749 S.n6748 0.039
R7158 S.n7506 S.n7505 0.039
R7159 S.n7511 S.n7510 0.039
R7160 S.n8242 S.n8241 0.039
R7161 S.n8247 S.n8246 0.039
R7162 S.n8969 S.n8968 0.039
R7163 S.n8974 S.n8973 0.039
R7164 S.n9670 S.n9669 0.039
R7165 S.n9675 S.n9674 0.039
R7166 S.n10362 S.n10361 0.039
R7167 S.n10367 S.n10366 0.039
R7168 S.n12321 S.n12320 0.039
R7169 S.n12470 S.n12469 0.039
R7170 S.n469 S.n462 0.039
R7171 S.n1039 S.n1032 0.039
R7172 S.n2330 S.n2323 0.039
R7173 S.n3204 S.n3197 0.039
R7174 S.n4069 S.n4062 0.039
R7175 S.n4877 S.n4870 0.039
R7176 S.n5676 S.n5669 0.039
R7177 S.n6449 S.n6442 0.039
R7178 S.n7213 S.n7206 0.039
R7179 S.n7784 S.n7777 0.039
R7180 S.n8498 S.n8491 0.039
R7181 S.n9383 S.n9376 0.039
R7182 S.n10077 S.n10070 0.039
R7183 S.n10748 S.n10741 0.039
R7184 S.n11391 S.n11384 0.039
R7185 S.n11962 S.n11955 0.039
R7186 S.n12606 S.n12604 0.038
R7187 S.n11952 S.n11950 0.038
R7188 S.n11676 S.n11675 0.038
R7189 S.n11079 S.n11078 0.038
R7190 S.n10454 S.n10453 0.038
R7191 S.n9794 S.n9793 0.038
R7192 S.n9122 S.n9121 0.038
R7193 S.n8427 S.n8426 0.038
R7194 S.n7720 S.n7719 0.038
R7195 S.n6990 S.n6989 0.038
R7196 S.n6248 S.n6247 0.038
R7197 S.n5483 S.n5482 0.038
R7198 S.n4706 S.n4705 0.038
R7199 S.n3906 S.n3905 0.038
R7200 S.n3094 S.n3093 0.038
R7201 S.n2257 S.n2256 0.038
R7202 S.n8280 S.n8279 0.038
R7203 S.n7573 S.n7572 0.038
R7204 S.n6843 S.n6842 0.038
R7205 S.n6101 S.n6100 0.038
R7206 S.n5336 S.n5335 0.038
R7207 S.n4559 S.n4558 0.038
R7208 S.n3759 S.n3758 0.038
R7209 S.n2947 S.n2946 0.038
R7210 S.n2104 S.n2103 0.038
R7211 S.n1659 S.n1658 0.038
R7212 S.n9018 S.n9013 0.038
R7213 S.n8323 S.n8318 0.038
R7214 S.n7616 S.n7611 0.038
R7215 S.n6886 S.n6881 0.038
R7216 S.n6144 S.n6139 0.038
R7217 S.n5379 S.n5374 0.038
R7218 S.n4602 S.n4597 0.038
R7219 S.n3802 S.n3797 0.038
R7220 S.n2990 S.n2985 0.038
R7221 S.n2149 S.n2144 0.038
R7222 S.n1699 S.n1695 0.038
R7223 S.n6782 S.n6781 0.038
R7224 S.n6040 S.n6039 0.038
R7225 S.n5275 S.n5274 0.038
R7226 S.n4498 S.n4497 0.038
R7227 S.n3698 S.n3697 0.038
R7228 S.n2886 S.n2885 0.038
R7229 S.n2041 S.n2040 0.038
R7230 S.n1600 S.n1599 0.038
R7231 S.n7555 S.n7550 0.038
R7232 S.n6825 S.n6820 0.038
R7233 S.n6083 S.n6078 0.038
R7234 S.n5318 S.n5313 0.038
R7235 S.n4541 S.n4536 0.038
R7236 S.n3741 S.n3736 0.038
R7237 S.n2929 S.n2924 0.038
R7238 S.n2086 S.n2081 0.038
R7239 S.n1641 S.n1636 0.038
R7240 S.n5214 S.n5213 0.038
R7241 S.n4437 S.n4436 0.038
R7242 S.n3637 S.n3636 0.038
R7243 S.n2825 S.n2824 0.038
R7244 S.n1978 S.n1977 0.038
R7245 S.n1541 S.n1540 0.038
R7246 S.n6022 S.n6017 0.038
R7247 S.n5257 S.n5252 0.038
R7248 S.n4480 S.n4475 0.038
R7249 S.n3680 S.n3675 0.038
R7250 S.n2868 S.n2863 0.038
R7251 S.n2023 S.n2018 0.038
R7252 S.n1582 S.n1577 0.038
R7253 S.n3576 S.n3575 0.038
R7254 S.n2764 S.n2763 0.038
R7255 S.n1915 S.n1914 0.038
R7256 S.n1482 S.n1481 0.038
R7257 S.n4419 S.n4414 0.038
R7258 S.n3619 S.n3614 0.038
R7259 S.n2807 S.n2802 0.038
R7260 S.n1960 S.n1955 0.038
R7261 S.n1523 S.n1518 0.038
R7262 S.n1852 S.n1851 0.038
R7263 S.n1423 S.n1422 0.038
R7264 S.n2746 S.n2741 0.038
R7265 S.n1897 S.n1892 0.038
R7266 S.n1467 S.n1462 0.038
R7267 S.n1405 S.n1400 0.038
R7268 S.n11121 S.n11119 0.037
R7269 S.n12295 S.n12292 0.037
R7270 S.n12294 S.n12293 0.037
R7271 S.n2220 S.n2202 0.037
R7272 S.n3058 S.n3040 0.037
R7273 S.n3870 S.n3852 0.037
R7274 S.n4670 S.n4652 0.037
R7275 S.n5447 S.n5429 0.037
R7276 S.n6212 S.n6194 0.037
R7277 S.n6954 S.n6936 0.037
R7278 S.n7684 S.n7666 0.037
R7279 S.n8391 S.n8373 0.037
R7280 S.n9086 S.n9068 0.037
R7281 S.n9758 S.n9740 0.037
R7282 S.n10418 S.n10400 0.037
R7283 S.n11122 S.n11111 0.037
R7284 S.n1763 S.n1755 0.037
R7285 S.n1735 S.n1727 0.037
R7286 S.n1819 S.n1816 0.037
R7287 S.n1818 S.n1817 0.037
R7288 S.n2702 S.n2699 0.037
R7289 S.n2701 S.n2700 0.037
R7290 S.n3543 S.n3540 0.037
R7291 S.n3542 S.n3541 0.037
R7292 S.n4375 S.n4372 0.037
R7293 S.n4374 S.n4373 0.037
R7294 S.n5181 S.n5178 0.037
R7295 S.n5180 S.n5179 0.037
R7296 S.n5978 S.n5975 0.037
R7297 S.n5977 S.n5976 0.037
R7298 S.n6749 S.n6746 0.037
R7299 S.n6748 S.n6747 0.037
R7300 S.n7511 S.n7508 0.037
R7301 S.n7510 S.n7509 0.037
R7302 S.n8247 S.n8244 0.037
R7303 S.n8246 S.n8245 0.037
R7304 S.n8974 S.n8971 0.037
R7305 S.n8973 S.n8972 0.037
R7306 S.n9675 S.n9672 0.037
R7307 S.n9674 S.n9673 0.037
R7308 S.n10367 S.n10364 0.037
R7309 S.n10366 S.n10365 0.037
R7310 S.n13126 S.n13125 0.037
R7311 S.n12255 S.n12254 0.037
R7312 S.n880 S.n877 0.036
R7313 S.n1292 S.n1291 0.036
R7314 S.n2561 S.n2560 0.036
R7315 S.n3417 S.n3416 0.036
R7316 S.n4264 S.n4263 0.036
R7317 S.n5054 S.n5053 0.036
R7318 S.n5835 S.n5834 0.036
R7319 S.n6590 S.n6589 0.036
R7320 S.n7336 S.n7335 0.036
R7321 S.n7889 S.n7888 0.036
R7322 S.n8585 S.n8584 0.036
R7323 S.n9452 S.n9451 0.036
R7324 S.n10128 S.n10127 0.036
R7325 S.n10781 S.n10780 0.036
R7326 S.n11402 S.n11401 0.036
R7327 S.n9395 S.n9394 0.035
R7328 S.n8528 S.n8527 0.035
R7329 S.n7832 S.n7831 0.035
R7330 S.n7279 S.n7278 0.035
R7331 S.n6533 S.n6532 0.035
R7332 S.n5778 S.n5777 0.035
R7333 S.n4997 S.n4996 0.035
R7334 S.n4207 S.n4206 0.035
R7335 S.n3360 S.n3359 0.035
R7336 S.n2504 S.n2503 0.035
R7337 S.n1221 S.n1220 0.035
R7338 S.n7796 S.n7795 0.035
R7339 S.n7243 S.n7242 0.035
R7340 S.n6497 S.n6496 0.035
R7341 S.n5742 S.n5741 0.035
R7342 S.n4961 S.n4960 0.035
R7343 S.n4171 S.n4170 0.035
R7344 S.n3324 S.n3323 0.035
R7345 S.n2468 S.n2467 0.035
R7346 S.n1187 S.n1186 0.035
R7347 S.n6461 S.n6460 0.035
R7348 S.n5706 S.n5705 0.035
R7349 S.n4925 S.n4924 0.035
R7350 S.n4135 S.n4134 0.035
R7351 S.n3288 S.n3287 0.035
R7352 S.n2432 S.n2431 0.035
R7353 S.n1153 S.n1152 0.035
R7354 S.n4889 S.n4888 0.035
R7355 S.n4099 S.n4098 0.035
R7356 S.n3252 S.n3251 0.035
R7357 S.n2396 S.n2395 0.035
R7358 S.n1119 S.n1118 0.035
R7359 S.n3216 S.n3215 0.035
R7360 S.n2360 S.n2359 0.035
R7361 S.n1085 S.n1084 0.035
R7362 S.n1051 S.n1050 0.035
R7363 S.n12555 S.n12554 0.035
R7364 S.n478 S.n477 0.035
R7365 S.n12623 S.n12622 0.035
R7366 S.n9393 S.n9392 0.035
R7367 S.n10086 S.n10085 0.035
R7368 S.n10758 S.n10757 0.035
R7369 S.n11400 S.n11399 0.035
R7370 S.n11972 S.n11971 0.035
R7371 S.n7794 S.n7793 0.035
R7372 S.n8507 S.n8506 0.035
R7373 S.n6459 S.n6458 0.035
R7374 S.n7222 S.n7221 0.035
R7375 S.n4887 S.n4886 0.035
R7376 S.n5685 S.n5684 0.035
R7377 S.n3214 S.n3213 0.035
R7378 S.n4078 S.n4077 0.035
R7379 S.n1049 S.n1048 0.035
R7380 S.n2339 S.n2338 0.035
R7381 S.n12296 S.n12295 0.035
R7382 S.n11676 S.n11671 0.035
R7383 S.n11079 S.n11074 0.035
R7384 S.n10454 S.n10449 0.035
R7385 S.n9794 S.n9789 0.035
R7386 S.n9122 S.n9117 0.035
R7387 S.n8427 S.n8422 0.035
R7388 S.n7720 S.n7715 0.035
R7389 S.n6990 S.n6985 0.035
R7390 S.n6248 S.n6243 0.035
R7391 S.n5483 S.n5478 0.035
R7392 S.n4706 S.n4701 0.035
R7393 S.n3906 S.n3901 0.035
R7394 S.n3094 S.n3089 0.035
R7395 S.n2257 S.n2252 0.035
R7396 S.n8280 S.n8275 0.035
R7397 S.n7573 S.n7568 0.035
R7398 S.n6843 S.n6838 0.035
R7399 S.n6101 S.n6096 0.035
R7400 S.n5336 S.n5331 0.035
R7401 S.n4559 S.n4554 0.035
R7402 S.n3759 S.n3754 0.035
R7403 S.n2947 S.n2942 0.035
R7404 S.n2104 S.n2099 0.035
R7405 S.n1659 S.n1654 0.035
R7406 S.n10499 S.n10482 0.035
R7407 S.n1699 S.n1698 0.035
R7408 S.n2149 S.n2148 0.035
R7409 S.n2990 S.n2989 0.035
R7410 S.n3802 S.n3801 0.035
R7411 S.n4602 S.n4601 0.035
R7412 S.n5379 S.n5378 0.035
R7413 S.n6144 S.n6143 0.035
R7414 S.n6886 S.n6885 0.035
R7415 S.n7616 S.n7615 0.035
R7416 S.n8323 S.n8322 0.035
R7417 S.n9018 S.n9017 0.035
R7418 S.n6782 S.n6777 0.035
R7419 S.n6040 S.n6035 0.035
R7420 S.n5275 S.n5270 0.035
R7421 S.n4498 S.n4493 0.035
R7422 S.n3698 S.n3693 0.035
R7423 S.n2886 S.n2881 0.035
R7424 S.n2041 S.n2036 0.035
R7425 S.n1600 S.n1595 0.035
R7426 S.n1641 S.n1640 0.035
R7427 S.n2086 S.n2085 0.035
R7428 S.n2929 S.n2928 0.035
R7429 S.n3741 S.n3740 0.035
R7430 S.n4541 S.n4540 0.035
R7431 S.n5318 S.n5317 0.035
R7432 S.n6083 S.n6082 0.035
R7433 S.n6825 S.n6824 0.035
R7434 S.n7555 S.n7554 0.035
R7435 S.n5214 S.n5209 0.035
R7436 S.n4437 S.n4432 0.035
R7437 S.n3637 S.n3632 0.035
R7438 S.n2825 S.n2820 0.035
R7439 S.n1978 S.n1973 0.035
R7440 S.n1541 S.n1536 0.035
R7441 S.n1582 S.n1581 0.035
R7442 S.n2023 S.n2022 0.035
R7443 S.n2868 S.n2867 0.035
R7444 S.n3680 S.n3679 0.035
R7445 S.n4480 S.n4479 0.035
R7446 S.n5257 S.n5256 0.035
R7447 S.n6022 S.n6021 0.035
R7448 S.n3576 S.n3571 0.035
R7449 S.n2764 S.n2759 0.035
R7450 S.n1915 S.n1910 0.035
R7451 S.n1482 S.n1477 0.035
R7452 S.n1523 S.n1522 0.035
R7453 S.n1960 S.n1959 0.035
R7454 S.n2807 S.n2806 0.035
R7455 S.n3619 S.n3618 0.035
R7456 S.n4419 S.n4418 0.035
R7457 S.n1852 S.n1847 0.035
R7458 S.n1423 S.n1418 0.035
R7459 S.n1467 S.n1466 0.035
R7460 S.n1897 S.n1896 0.035
R7461 S.n2746 S.n2745 0.035
R7462 S.n1405 S.n1404 0.035
R7463 S.n1812 S.n1811 0.035
R7464 S.n1822 S.n1819 0.035
R7465 S.n2695 S.n2694 0.035
R7466 S.n2705 S.n2702 0.035
R7467 S.n3536 S.n3535 0.035
R7468 S.n3546 S.n3543 0.035
R7469 S.n4368 S.n4367 0.035
R7470 S.n4378 S.n4375 0.035
R7471 S.n5174 S.n5173 0.035
R7472 S.n5184 S.n5181 0.035
R7473 S.n5971 S.n5970 0.035
R7474 S.n5981 S.n5978 0.035
R7475 S.n6742 S.n6741 0.035
R7476 S.n6752 S.n6749 0.035
R7477 S.n7504 S.n7503 0.035
R7478 S.n7514 S.n7511 0.035
R7479 S.n8240 S.n8239 0.035
R7480 S.n8250 S.n8247 0.035
R7481 S.n8967 S.n8966 0.035
R7482 S.n8977 S.n8974 0.035
R7483 S.n9668 S.n9667 0.035
R7484 S.n9678 S.n9675 0.035
R7485 S.n10360 S.n10359 0.035
R7486 S.n10370 S.n10367 0.035
R7487 S.t35 S.n12540 0.035
R7488 S.t28 S.n949 0.035
R7489 S.t28 S.n945 0.035
R7490 S.t28 S.n195 0.035
R7491 S.t28 S.n973 0.035
R7492 S.t28 S.n209 0.035
R7493 S.t28 S.n220 0.035
R7494 S.t28 S.n927 0.035
R7495 S.t28 S.n183 0.035
R7496 S.t28 S.n969 0.035
R7497 S.t28 S.n170 0.035
R7498 S.t28 S.n965 0.035
R7499 S.t28 S.n157 0.035
R7500 S.t28 S.n961 0.035
R7501 S.t28 S.n144 0.035
R7502 S.t28 S.n957 0.035
R7503 S.t28 S.n131 0.035
R7504 S.t28 S.n953 0.035
R7505 S.t35 S.n12480 0.035
R7506 S.t35 S.n12484 0.035
R7507 S.t35 S.n12488 0.035
R7508 S.t35 S.n12492 0.035
R7509 S.t35 S.n12496 0.035
R7510 S.t35 S.n12500 0.035
R7511 S.t35 S.n12504 0.035
R7512 S.t35 S.n12508 0.035
R7513 S.t35 S.n12512 0.035
R7514 S.t35 S.n12516 0.035
R7515 S.t35 S.n12520 0.035
R7516 S.t35 S.n12524 0.035
R7517 S.t35 S.n12528 0.035
R7518 S.t35 S.n12532 0.035
R7519 S.t35 S.n12536 0.035
R7520 S.t35 S.n12476 0.035
R7521 S.n12388 S.n12387 0.035
R7522 S.n11034 S.n11033 0.034
R7523 S.n206 S.n202 0.034
R7524 S.n199 S.n198 0.034
R7525 S.n187 S.n186 0.034
R7526 S.n175 S.n174 0.034
R7527 S.n162 S.n161 0.034
R7528 S.n149 S.n148 0.034
R7529 S.n136 S.n135 0.034
R7530 S.n12891 S.n12888 0.034
R7531 S.n12906 S.n12902 0.034
R7532 S.n12027 S.n12024 0.034
R7533 S.n11737 S.n11733 0.034
R7534 S.n11145 S.n11142 0.034
R7535 S.n11159 S.n11155 0.034
R7536 S.n10522 S.n10519 0.034
R7537 S.n10536 S.n10532 0.034
R7538 S.n9864 S.n9861 0.034
R7539 S.n9878 S.n9874 0.034
R7540 S.n9187 S.n9184 0.034
R7541 S.n9201 S.n9197 0.034
R7542 S.n8783 S.n8780 0.034
R7543 S.n8797 S.n8793 0.034
R7544 S.n8071 S.n8068 0.034
R7545 S.n8085 S.n8081 0.034
R7546 S.n7060 S.n7057 0.034
R7547 S.n7074 S.n7070 0.034
R7548 S.n6313 S.n6310 0.034
R7549 S.n6327 S.n6323 0.034
R7550 S.n5553 S.n5550 0.034
R7551 S.n5567 S.n5563 0.034
R7552 S.n4771 S.n4768 0.034
R7553 S.n4785 S.n4781 0.034
R7554 S.n3976 S.n3973 0.034
R7555 S.n3990 S.n3986 0.034
R7556 S.n3159 S.n3156 0.034
R7557 S.n3173 S.n3169 0.034
R7558 S.n2632 S.n2629 0.034
R7559 S.n2646 S.n2642 0.034
R7560 S.n1346 S.n1343 0.034
R7561 S.n1808 S.n986 0.034
R7562 S.n2692 S.n2691 0.034
R7563 S.n3533 S.n3532 0.034
R7564 S.n4365 S.n4364 0.034
R7565 S.n5171 S.n5170 0.034
R7566 S.n5968 S.n5967 0.034
R7567 S.n6739 S.n6738 0.034
R7568 S.n7501 S.n7500 0.034
R7569 S.n8237 S.n8236 0.034
R7570 S.n8964 S.n8963 0.034
R7571 S.n9665 S.n9664 0.034
R7572 S.n10357 S.n10356 0.034
R7573 S.n11026 S.n11025 0.034
R7574 S.n11666 S.n11665 0.034
R7575 S.n12306 S.n12305 0.034
R7576 S.n468 S.n463 0.034
R7577 S.n1038 S.n1033 0.034
R7578 S.n2329 S.n2324 0.034
R7579 S.n3203 S.n3198 0.034
R7580 S.n4068 S.n4063 0.034
R7581 S.n4876 S.n4871 0.034
R7582 S.n5675 S.n5670 0.034
R7583 S.n6448 S.n6443 0.034
R7584 S.n7212 S.n7207 0.034
R7585 S.n7783 S.n7778 0.034
R7586 S.n8497 S.n8492 0.034
R7587 S.n9382 S.n9377 0.034
R7588 S.n10076 S.n10071 0.034
R7589 S.n10747 S.n10742 0.034
R7590 S.n11390 S.n11385 0.034
R7591 S.n11961 S.n11956 0.034
R7592 S.n12310 S.n12307 0.034
R7593 S.n10751 S.n10738 0.034
R7594 S.n10080 S.n10067 0.034
R7595 S.n9386 S.n9373 0.034
R7596 S.n8501 S.n8488 0.034
R7597 S.n7787 S.n7774 0.034
R7598 S.n7216 S.n7203 0.034
R7599 S.n6452 S.n6439 0.034
R7600 S.n5679 S.n5666 0.034
R7601 S.n4880 S.n4867 0.034
R7602 S.n4072 S.n4059 0.034
R7603 S.n3207 S.n3194 0.034
R7604 S.n2333 S.n2320 0.034
R7605 S.n1042 S.n1029 0.034
R7606 S.n472 S.n459 0.034
R7607 S.t35 S.n12543 0.034
R7608 S.t28 S.n952 0.034
R7609 S.t28 S.n944 0.034
R7610 S.t28 S.n194 0.034
R7611 S.t28 S.n976 0.034
R7612 S.t28 S.n208 0.034
R7613 S.t28 S.n219 0.034
R7614 S.t28 S.n926 0.034
R7615 S.t28 S.n182 0.034
R7616 S.t28 S.n972 0.034
R7617 S.t28 S.n169 0.034
R7618 S.t28 S.n968 0.034
R7619 S.t28 S.n156 0.034
R7620 S.t28 S.n964 0.034
R7621 S.t28 S.n143 0.034
R7622 S.t28 S.n960 0.034
R7623 S.t28 S.n130 0.034
R7624 S.t28 S.n956 0.034
R7625 S.t35 S.n12483 0.034
R7626 S.t35 S.n12487 0.034
R7627 S.t35 S.n12491 0.034
R7628 S.t35 S.n12495 0.034
R7629 S.t35 S.n12499 0.034
R7630 S.t35 S.n12503 0.034
R7631 S.t35 S.n12507 0.034
R7632 S.t35 S.n12511 0.034
R7633 S.t35 S.n12515 0.034
R7634 S.t35 S.n12519 0.034
R7635 S.t35 S.n12523 0.034
R7636 S.t35 S.n12527 0.034
R7637 S.t35 S.n12531 0.034
R7638 S.t35 S.n12535 0.034
R7639 S.t35 S.n12539 0.034
R7640 S.t35 S.n12475 0.034
R7641 S.n122 S.n121 0.033
R7642 S.n1251 S.n1250 0.033
R7643 S.n12617 S.n12606 0.032
R7644 S.n11965 S.n11952 0.032
R7645 S.n11377 S.n11376 0.032
R7646 S.n1371 S.n1370 0.031
R7647 S.t430 S.n478 0.031
R7648 S.t14 S.n12623 0.031
R7649 S.t26 S.n9393 0.031
R7650 S.t16 S.n10086 0.031
R7651 S.t122 S.n10758 0.031
R7652 S.t18 S.n11400 0.031
R7653 S.t2 S.n11972 0.031
R7654 S.t22 S.n7794 0.031
R7655 S.t0 S.n8507 0.031
R7656 S.t8 S.n6459 0.031
R7657 S.t40 S.n7222 0.031
R7658 S.t81 S.n4887 0.031
R7659 S.t460 S.n5685 0.031
R7660 S.t444 S.n3214 0.031
R7661 S.t51 S.n4078 0.031
R7662 S.t142 S.n1049 0.031
R7663 S.t55 S.n2339 0.031
R7664 S.n11671 S.n11670 0.031
R7665 S.n11074 S.n11073 0.031
R7666 S.n10449 S.n10448 0.031
R7667 S.n9789 S.n9788 0.031
R7668 S.n9117 S.n9116 0.031
R7669 S.n8422 S.n8421 0.031
R7670 S.n7715 S.n7714 0.031
R7671 S.n6985 S.n6984 0.031
R7672 S.n6243 S.n6242 0.031
R7673 S.n5478 S.n5477 0.031
R7674 S.n4701 S.n4700 0.031
R7675 S.n3901 S.n3900 0.031
R7676 S.n3089 S.n3088 0.031
R7677 S.n2252 S.n2251 0.031
R7678 S.n8275 S.n8274 0.031
R7679 S.n7568 S.n7567 0.031
R7680 S.n6838 S.n6837 0.031
R7681 S.n6096 S.n6095 0.031
R7682 S.n5331 S.n5330 0.031
R7683 S.n4554 S.n4553 0.031
R7684 S.n3754 S.n3753 0.031
R7685 S.n2942 S.n2941 0.031
R7686 S.n2099 S.n2098 0.031
R7687 S.n1654 S.n1653 0.031
R7688 S.n1698 S.n1697 0.031
R7689 S.n2148 S.n2147 0.031
R7690 S.n2989 S.n2988 0.031
R7691 S.n3801 S.n3800 0.031
R7692 S.n4601 S.n4600 0.031
R7693 S.n5378 S.n5377 0.031
R7694 S.n6143 S.n6142 0.031
R7695 S.n6885 S.n6884 0.031
R7696 S.n7615 S.n7614 0.031
R7697 S.n8322 S.n8321 0.031
R7698 S.n9017 S.n9016 0.031
R7699 S.n6777 S.n6776 0.031
R7700 S.n6035 S.n6034 0.031
R7701 S.n5270 S.n5269 0.031
R7702 S.n4493 S.n4492 0.031
R7703 S.n3693 S.n3692 0.031
R7704 S.n2881 S.n2880 0.031
R7705 S.n2036 S.n2035 0.031
R7706 S.n1595 S.n1594 0.031
R7707 S.n1640 S.n1639 0.031
R7708 S.n2085 S.n2084 0.031
R7709 S.n2928 S.n2927 0.031
R7710 S.n3740 S.n3739 0.031
R7711 S.n4540 S.n4539 0.031
R7712 S.n5317 S.n5316 0.031
R7713 S.n6082 S.n6081 0.031
R7714 S.n6824 S.n6823 0.031
R7715 S.n7554 S.n7553 0.031
R7716 S.n5209 S.n5208 0.031
R7717 S.n4432 S.n4431 0.031
R7718 S.n3632 S.n3631 0.031
R7719 S.n2820 S.n2819 0.031
R7720 S.n1973 S.n1972 0.031
R7721 S.n1536 S.n1535 0.031
R7722 S.n1581 S.n1580 0.031
R7723 S.n2022 S.n2021 0.031
R7724 S.n2867 S.n2866 0.031
R7725 S.n3679 S.n3678 0.031
R7726 S.n4479 S.n4478 0.031
R7727 S.n5256 S.n5255 0.031
R7728 S.n6021 S.n6020 0.031
R7729 S.n3571 S.n3570 0.031
R7730 S.n2759 S.n2758 0.031
R7731 S.n1910 S.n1909 0.031
R7732 S.n1477 S.n1476 0.031
R7733 S.n1522 S.n1521 0.031
R7734 S.n1959 S.n1958 0.031
R7735 S.n2806 S.n2805 0.031
R7736 S.n3618 S.n3617 0.031
R7737 S.n4418 S.n4417 0.031
R7738 S.n1847 S.n1846 0.031
R7739 S.n1418 S.n1417 0.031
R7740 S.n1466 S.n1465 0.031
R7741 S.n1896 S.n1895 0.031
R7742 S.n2745 S.n2744 0.031
R7743 S.n1404 S.n1403 0.031
R7744 S.n979 S.n978 0.031
R7745 S.n980 S.n979 0.031
R7746 S.n981 S.n980 0.031
R7747 S.n982 S.n981 0.031
R7748 S.n983 S.n982 0.031
R7749 S.n984 S.n983 0.031
R7750 S.n985 S.n984 0.031
R7751 S.n879 S.n878 0.031
R7752 S.n13178 S.n13177 0.031
R7753 S.n13177 S.n13176 0.031
R7754 S.n13176 S.n13175 0.031
R7755 S.n13175 S.n13174 0.031
R7756 S.n13174 S.n13173 0.031
R7757 S.n13173 S.n13172 0.031
R7758 S.n13172 S.n13171 0.031
R7759 S.n13171 S.n13170 0.031
R7760 S.n13170 S.n13169 0.031
R7761 S.n13169 S.n13168 0.031
R7762 S.n13168 S.n13167 0.031
R7763 S.n13167 S.n13166 0.031
R7764 S.n13166 S.n13165 0.031
R7765 S.n13165 S.n13164 0.031
R7766 S.n13164 S.n13163 0.031
R7767 S.n13163 S.n13162 0.031
R7768 S.n12904 S.n12903 0.031
R7769 S.n11735 S.n11734 0.031
R7770 S.n11157 S.n11156 0.031
R7771 S.n10534 S.n10533 0.031
R7772 S.n9876 S.n9875 0.031
R7773 S.n9199 S.n9198 0.031
R7774 S.n8795 S.n8794 0.031
R7775 S.n8083 S.n8082 0.031
R7776 S.n7072 S.n7071 0.031
R7777 S.n6325 S.n6324 0.031
R7778 S.n5565 S.n5564 0.031
R7779 S.n4783 S.n4782 0.031
R7780 S.n3988 S.n3987 0.031
R7781 S.n3171 S.n3170 0.031
R7782 S.n2644 S.n2643 0.031
R7783 S.n8472 S.n8471 0.031
R7784 S.n7035 S.n7034 0.031
R7785 S.n3951 S.n3950 0.031
R7786 S.n2304 S.n2303 0.031
R7787 S.n9824 S.n9823 0.03
R7788 S.n8457 S.n8456 0.03
R7789 S.n7020 S.n7019 0.03
R7790 S.n5513 S.n5512 0.03
R7791 S.n3936 S.n3935 0.03
R7792 S.n2289 S.n2288 0.03
R7793 S.n10412 S.n10411 0.03
R7794 S.n9752 S.n9751 0.03
R7795 S.n9080 S.n9079 0.03
R7796 S.n8385 S.n8384 0.03
R7797 S.n7678 S.n7677 0.03
R7798 S.n6948 S.n6947 0.03
R7799 S.n6206 S.n6205 0.03
R7800 S.n5441 S.n5440 0.03
R7801 S.n4664 S.n4663 0.03
R7802 S.n3864 S.n3863 0.03
R7803 S.n3052 S.n3051 0.03
R7804 S.n2214 S.n2213 0.03
R7805 S.n1713 S.n1712 0.03
R7806 S.n911 S.n910 0.03
R7807 S.n837 S.n836 0.03
R7808 S.n9157 S.n9154 0.029
R7809 S.n10492 S.n10489 0.029
R7810 S.n7755 S.n7752 0.029
R7811 S.n6283 S.n6280 0.029
R7812 S.n4741 S.n4738 0.029
R7813 S.n3129 S.n3126 0.029
R7814 S.n1781 S.n1780 0.029
R7815 S.n2271 S.n2270 0.029
R7816 S.n3106 S.n3105 0.029
R7817 S.n3918 S.n3917 0.029
R7818 S.n4718 S.n4717 0.029
R7819 S.n5495 S.n5494 0.029
R7820 S.n6260 S.n6259 0.029
R7821 S.n7002 S.n7001 0.029
R7822 S.n7732 S.n7731 0.029
R7823 S.n8439 S.n8438 0.029
R7824 S.n9134 S.n9133 0.029
R7825 S.n9806 S.n9805 0.029
R7826 S.n10466 S.n10465 0.029
R7827 S.n11091 S.n11090 0.029
R7828 S.n11688 S.n11687 0.029
R7829 S.n2182 S.n2181 0.029
R7830 S.n3020 S.n3019 0.029
R7831 S.n3832 S.n3831 0.029
R7832 S.n4632 S.n4631 0.029
R7833 S.n5409 S.n5408 0.029
R7834 S.n6174 S.n6173 0.029
R7835 S.n6916 S.n6915 0.029
R7836 S.n7646 S.n7645 0.029
R7837 S.n8353 S.n8352 0.029
R7838 S.n9048 S.n9047 0.029
R7839 S.n9720 S.n9719 0.029
R7840 S.n2118 S.n2117 0.029
R7841 S.n2959 S.n2958 0.029
R7842 S.n3771 S.n3770 0.029
R7843 S.n4571 S.n4570 0.029
R7844 S.n5348 S.n5347 0.029
R7845 S.n6113 S.n6112 0.029
R7846 S.n6855 S.n6854 0.029
R7847 S.n7585 S.n7584 0.029
R7848 S.n8292 S.n8291 0.029
R7849 S.n2055 S.n2054 0.029
R7850 S.n2898 S.n2897 0.029
R7851 S.n3710 S.n3709 0.029
R7852 S.n4510 S.n4509 0.029
R7853 S.n5287 S.n5286 0.029
R7854 S.n6052 S.n6051 0.029
R7855 S.n6794 S.n6793 0.029
R7856 S.n1992 S.n1991 0.029
R7857 S.n2837 S.n2836 0.029
R7858 S.n3649 S.n3648 0.029
R7859 S.n4449 S.n4448 0.029
R7860 S.n5226 S.n5225 0.029
R7861 S.n1929 S.n1928 0.029
R7862 S.n2776 S.n2775 0.029
R7863 S.n3588 S.n3587 0.029
R7864 S.n1866 S.n1865 0.029
R7865 S.n3009 S.n3008 0.029
R7866 S.n3821 S.n3820 0.029
R7867 S.n4621 S.n4620 0.029
R7868 S.n5398 S.n5397 0.029
R7869 S.n6163 S.n6162 0.029
R7870 S.n6905 S.n6904 0.029
R7871 S.n7635 S.n7634 0.029
R7872 S.n8342 S.n8341 0.029
R7873 S.n9037 S.n9036 0.029
R7874 S.n9709 S.n9708 0.029
R7875 S.n10411 S.n10410 0.029
R7876 S.n9751 S.n9750 0.029
R7877 S.n9079 S.n9078 0.029
R7878 S.n8384 S.n8383 0.029
R7879 S.n7677 S.n7676 0.029
R7880 S.n6947 S.n6946 0.029
R7881 S.n6205 S.n6204 0.029
R7882 S.n5440 S.n5439 0.029
R7883 S.n4663 S.n4662 0.029
R7884 S.n3863 S.n3862 0.029
R7885 S.n3051 S.n3050 0.029
R7886 S.n2213 S.n2212 0.029
R7887 S.n1712 S.n1711 0.029
R7888 S.n910 S.n909 0.029
R7889 S.n11671 S.n11668 0.028
R7890 S.n11074 S.n11071 0.028
R7891 S.n10449 S.n10446 0.028
R7892 S.n9789 S.n9786 0.028
R7893 S.n9117 S.n9114 0.028
R7894 S.n8422 S.n8419 0.028
R7895 S.n7715 S.n7712 0.028
R7896 S.n6985 S.n6982 0.028
R7897 S.n6243 S.n6240 0.028
R7898 S.n5478 S.n5475 0.028
R7899 S.n4701 S.n4698 0.028
R7900 S.n3901 S.n3898 0.028
R7901 S.n3089 S.n3086 0.028
R7902 S.n2252 S.n2249 0.028
R7903 S.n8275 S.n8272 0.028
R7904 S.n7568 S.n7565 0.028
R7905 S.n6838 S.n6835 0.028
R7906 S.n6096 S.n6093 0.028
R7907 S.n5331 S.n5328 0.028
R7908 S.n4554 S.n4551 0.028
R7909 S.n3754 S.n3751 0.028
R7910 S.n2942 S.n2939 0.028
R7911 S.n2099 S.n2096 0.028
R7912 S.n1654 S.n1651 0.028
R7913 S.n2148 S.n2145 0.028
R7914 S.n2989 S.n2986 0.028
R7915 S.n3801 S.n3798 0.028
R7916 S.n4601 S.n4598 0.028
R7917 S.n5378 S.n5375 0.028
R7918 S.n6143 S.n6140 0.028
R7919 S.n6885 S.n6882 0.028
R7920 S.n7615 S.n7612 0.028
R7921 S.n8322 S.n8319 0.028
R7922 S.n9017 S.n9014 0.028
R7923 S.n6777 S.n6774 0.028
R7924 S.n6035 S.n6032 0.028
R7925 S.n5270 S.n5267 0.028
R7926 S.n4493 S.n4490 0.028
R7927 S.n3693 S.n3690 0.028
R7928 S.n2881 S.n2878 0.028
R7929 S.n2036 S.n2033 0.028
R7930 S.n1595 S.n1592 0.028
R7931 S.n1640 S.n1637 0.028
R7932 S.n2085 S.n2082 0.028
R7933 S.n2928 S.n2925 0.028
R7934 S.n3740 S.n3737 0.028
R7935 S.n4540 S.n4537 0.028
R7936 S.n5317 S.n5314 0.028
R7937 S.n6082 S.n6079 0.028
R7938 S.n6824 S.n6821 0.028
R7939 S.n7554 S.n7551 0.028
R7940 S.n5209 S.n5206 0.028
R7941 S.n4432 S.n4429 0.028
R7942 S.n3632 S.n3629 0.028
R7943 S.n2820 S.n2817 0.028
R7944 S.n1973 S.n1970 0.028
R7945 S.n1536 S.n1533 0.028
R7946 S.n1581 S.n1578 0.028
R7947 S.n2022 S.n2019 0.028
R7948 S.n2867 S.n2864 0.028
R7949 S.n3679 S.n3676 0.028
R7950 S.n4479 S.n4476 0.028
R7951 S.n5256 S.n5253 0.028
R7952 S.n6021 S.n6018 0.028
R7953 S.n3571 S.n3568 0.028
R7954 S.n2759 S.n2756 0.028
R7955 S.n1910 S.n1907 0.028
R7956 S.n1477 S.n1474 0.028
R7957 S.n1522 S.n1519 0.028
R7958 S.n1959 S.n1956 0.028
R7959 S.n2806 S.n2803 0.028
R7960 S.n3618 S.n3615 0.028
R7961 S.n4418 S.n4415 0.028
R7962 S.n1847 S.n1844 0.028
R7963 S.n1418 S.n1415 0.028
R7964 S.n1466 S.n1463 0.028
R7965 S.n1896 S.n1893 0.028
R7966 S.n2745 S.n2742 0.028
R7967 S.n1404 S.n1401 0.028
R7968 S.n2198 S.n2197 0.028
R7969 S.n2200 S.n2198 0.028
R7970 S.n3036 S.n3035 0.028
R7971 S.n3038 S.n3036 0.028
R7972 S.n3848 S.n3847 0.028
R7973 S.n3850 S.n3848 0.028
R7974 S.n4648 S.n4647 0.028
R7975 S.n4650 S.n4648 0.028
R7976 S.n5425 S.n5424 0.028
R7977 S.n5427 S.n5425 0.028
R7978 S.n6190 S.n6189 0.028
R7979 S.n6192 S.n6190 0.028
R7980 S.n6932 S.n6931 0.028
R7981 S.n6934 S.n6932 0.028
R7982 S.n7662 S.n7661 0.028
R7983 S.n7664 S.n7662 0.028
R7984 S.n8369 S.n8368 0.028
R7985 S.n8371 S.n8369 0.028
R7986 S.n9064 S.n9063 0.028
R7987 S.n9066 S.n9064 0.028
R7988 S.n9736 S.n9735 0.028
R7989 S.n9738 S.n9736 0.028
R7990 S.n10396 S.n10395 0.028
R7991 S.n10398 S.n10396 0.028
R7992 S.n11108 S.n11107 0.028
R7993 S.n11110 S.n11108 0.028
R7994 S.n1729 S.n1728 0.028
R7995 S.n1731 S.n1729 0.028
R7996 S.n1757 S.n1756 0.028
R7997 S.n1759 S.n1757 0.028
R7998 S.n12584 S.n12583 0.028
R7999 S.n10492 S.n10491 0.028
R8000 S.n9157 S.n9156 0.028
R8001 S.n7755 S.n7754 0.028
R8002 S.n6283 S.n6282 0.028
R8003 S.n4741 S.n4740 0.028
R8004 S.n3129 S.n3128 0.028
R8005 S.n2169 S.n2168 0.028
R8006 S.n869 S.n864 0.028
R8007 S.n992 S.n988 0.028
R8008 S.n1836 S.n1832 0.028
R8009 S.n2719 S.n2715 0.028
R8010 S.n3560 S.n3556 0.028
R8011 S.n4392 S.n4388 0.028
R8012 S.n5198 S.n5194 0.028
R8013 S.n5995 S.n5991 0.028
R8014 S.n6766 S.n6762 0.028
R8015 S.n7528 S.n7524 0.028
R8016 S.n8264 S.n8260 0.028
R8017 S.n8991 S.n8987 0.028
R8018 S.n9692 S.n9688 0.028
R8019 S.n10384 S.n10380 0.028
R8020 S.n11043 S.n11039 0.028
R8021 S.n12286 S.n12282 0.028
R8022 S.n13156 S.n13152 0.028
R8023 S.n13126 S.n13124 0.027
R8024 S.n12255 S.n12253 0.027
R8025 S.n12893 S.n12892 0.027
R8026 S.n901 S.n896 0.027
R8027 S.n798 S.n797 0.027
R8028 S.n9837 S.n9836 0.027
R8029 S.n8471 S.n8470 0.027
R8030 S.n7034 S.n7033 0.027
R8031 S.n5526 S.n5525 0.027
R8032 S.n3950 S.n3949 0.027
R8033 S.n2303 S.n2302 0.027
R8034 S.n1808 S.n1807 0.027
R8035 S.n2642 S.n2641 0.027
R8036 S.n3169 S.n3168 0.027
R8037 S.n3986 S.n3985 0.027
R8038 S.n4781 S.n4780 0.027
R8039 S.n5563 S.n5562 0.027
R8040 S.n6323 S.n6322 0.027
R8041 S.n7070 S.n7069 0.027
R8042 S.n8081 S.n8080 0.027
R8043 S.n8793 S.n8792 0.027
R8044 S.n9197 S.n9196 0.027
R8045 S.n9874 S.n9873 0.027
R8046 S.n10532 S.n10531 0.027
R8047 S.n11155 S.n11154 0.027
R8048 S.n11733 S.n11732 0.027
R8049 S.n12902 S.n12901 0.027
R8050 S.n1230 S.n1229 0.027
R8051 S.n1785 S.n1782 0.026
R8052 S.n1310 S.n1309 0.026
R8053 S.n2275 S.n2272 0.026
R8054 S.n2592 S.n2589 0.026
R8055 S.n3110 S.n3107 0.026
R8056 S.n3448 S.n3445 0.026
R8057 S.n3922 S.n3919 0.026
R8058 S.n4295 S.n4292 0.026
R8059 S.n4722 S.n4719 0.026
R8060 S.n5085 S.n5082 0.026
R8061 S.n5499 S.n5496 0.026
R8062 S.n5866 S.n5863 0.026
R8063 S.n6264 S.n6261 0.026
R8064 S.n6621 S.n6618 0.026
R8065 S.n7006 S.n7003 0.026
R8066 S.n7367 S.n7364 0.026
R8067 S.n7736 S.n7733 0.026
R8068 S.n7920 S.n7917 0.026
R8069 S.n8443 S.n8440 0.026
R8070 S.n8616 S.n8613 0.026
R8071 S.n9138 S.n9135 0.026
R8072 S.n9483 S.n9480 0.026
R8073 S.n9810 S.n9807 0.026
R8074 S.n10159 S.n10156 0.026
R8075 S.n10470 S.n10467 0.026
R8076 S.n10812 S.n10809 0.026
R8077 S.n11095 S.n11092 0.026
R8078 S.n11433 S.n11430 0.026
R8079 S.n11692 S.n11689 0.026
R8080 S.n11985 S.n11982 0.026
R8081 S.n12591 S.n12585 0.026
R8082 S.n729 S.n721 0.026
R8083 S.t320 S.n1017 0.026
R8084 S.n1252 S.n1240 0.026
R8085 S.n2186 S.n2183 0.026
R8086 S.n2532 S.n2529 0.026
R8087 S.n3024 S.n3021 0.026
R8088 S.n3388 S.n3385 0.026
R8089 S.n3836 S.n3833 0.026
R8090 S.n4235 S.n4232 0.026
R8091 S.n4636 S.n4633 0.026
R8092 S.n5025 S.n5022 0.026
R8093 S.n5413 S.n5410 0.026
R8094 S.n5806 S.n5803 0.026
R8095 S.n6178 S.n6175 0.026
R8096 S.n6561 S.n6558 0.026
R8097 S.n6920 S.n6917 0.026
R8098 S.n7307 S.n7304 0.026
R8099 S.n7650 S.n7647 0.026
R8100 S.n7860 S.n7857 0.026
R8101 S.n8357 S.n8354 0.026
R8102 S.n8556 S.n8553 0.026
R8103 S.n9052 S.n9049 0.026
R8104 S.n9423 S.n9420 0.026
R8105 S.n9724 S.n9721 0.026
R8106 S.n10099 S.n10096 0.026
R8107 S.n10499 S.n10493 0.026
R8108 S.n1262 S.n1260 0.026
R8109 S.n2542 S.n2540 0.026
R8110 S.n3398 S.n3396 0.026
R8111 S.n4245 S.n4243 0.026
R8112 S.n5035 S.n5033 0.026
R8113 S.n5816 S.n5814 0.026
R8114 S.n6571 S.n6569 0.026
R8115 S.n7317 S.n7315 0.026
R8116 S.n7870 S.n7868 0.026
R8117 S.n8566 S.n8564 0.026
R8118 S.n9433 S.n9431 0.026
R8119 S.n10109 S.n10107 0.026
R8120 S.n10762 S.n10760 0.026
R8121 S.n11413 S.n11412 0.026
R8122 S.n10792 S.n10791 0.026
R8123 S.n10139 S.n10138 0.026
R8124 S.n9463 S.n9462 0.026
R8125 S.n8596 S.n8595 0.026
R8126 S.n7900 S.n7899 0.026
R8127 S.n7347 S.n7346 0.026
R8128 S.n6601 S.n6600 0.026
R8129 S.n5846 S.n5845 0.026
R8130 S.n5065 S.n5064 0.026
R8131 S.n4275 S.n4274 0.026
R8132 S.n3428 S.n3427 0.026
R8133 S.n2572 S.n2571 0.026
R8134 S.n1282 S.n1281 0.026
R8135 S.n1763 S.n1746 0.026
R8136 S.n2241 S.n2231 0.026
R8137 S.n3078 S.n3069 0.026
R8138 S.n3890 S.n3881 0.026
R8139 S.n4690 S.n4681 0.026
R8140 S.n5467 S.n5458 0.026
R8141 S.n6232 S.n6223 0.026
R8142 S.n6974 S.n6965 0.026
R8143 S.n7704 S.n7695 0.026
R8144 S.n8411 S.n8402 0.026
R8145 S.n9106 S.n9097 0.026
R8146 S.n9778 S.n9769 0.026
R8147 S.n10438 S.n10429 0.026
R8148 S.n11063 S.n11054 0.026
R8149 S.n11717 S.n11708 0.026
R8150 S.n9841 S.n9825 0.026
R8151 S.n9020 S.n9002 0.026
R8152 S.n8325 S.n8307 0.026
R8153 S.n7618 S.n7600 0.026
R8154 S.n6888 S.n6870 0.026
R8155 S.n6146 S.n6128 0.026
R8156 S.n5381 S.n5363 0.026
R8157 S.n4604 S.n4586 0.026
R8158 S.n3804 S.n3786 0.026
R8159 S.n2992 S.n2974 0.026
R8160 S.n2151 S.n2133 0.026
R8161 S.n1701 S.n1685 0.026
R8162 S.n1673 S.n1670 0.026
R8163 S.n1213 S.n1212 0.026
R8164 S.n2122 S.n2119 0.026
R8165 S.n2496 S.n2493 0.026
R8166 S.n2963 S.n2960 0.026
R8167 S.n3352 S.n3349 0.026
R8168 S.n3775 S.n3772 0.026
R8169 S.n4199 S.n4196 0.026
R8170 S.n4575 S.n4572 0.026
R8171 S.n4989 S.n4986 0.026
R8172 S.n5352 S.n5349 0.026
R8173 S.n5770 S.n5767 0.026
R8174 S.n6117 S.n6114 0.026
R8175 S.n6525 S.n6522 0.026
R8176 S.n6859 S.n6856 0.026
R8177 S.n7271 S.n7268 0.026
R8178 S.n7589 S.n7586 0.026
R8179 S.n7824 S.n7821 0.026
R8180 S.n8296 S.n8293 0.026
R8181 S.n8520 S.n8517 0.026
R8182 S.n9164 S.n9158 0.026
R8183 S.n8474 S.n8458 0.026
R8184 S.n7557 S.n7539 0.026
R8185 S.n6827 S.n6809 0.026
R8186 S.n6085 S.n6067 0.026
R8187 S.n5320 S.n5302 0.026
R8188 S.n4543 S.n4525 0.026
R8189 S.n3743 S.n3725 0.026
R8190 S.n2931 S.n2913 0.026
R8191 S.n2088 S.n2070 0.026
R8192 S.n1643 S.n1626 0.026
R8193 S.n1614 S.n1611 0.026
R8194 S.n1179 S.n1178 0.026
R8195 S.n2059 S.n2056 0.026
R8196 S.n2460 S.n2457 0.026
R8197 S.n2902 S.n2899 0.026
R8198 S.n3316 S.n3313 0.026
R8199 S.n3714 S.n3711 0.026
R8200 S.n4163 S.n4160 0.026
R8201 S.n4514 S.n4511 0.026
R8202 S.n4953 S.n4950 0.026
R8203 S.n5291 S.n5288 0.026
R8204 S.n5734 S.n5731 0.026
R8205 S.n6056 S.n6053 0.026
R8206 S.n6489 S.n6486 0.026
R8207 S.n6798 S.n6795 0.026
R8208 S.n7235 S.n7232 0.026
R8209 S.n7762 S.n7756 0.026
R8210 S.n7037 S.n7021 0.026
R8211 S.n6024 S.n6006 0.026
R8212 S.n5259 S.n5241 0.026
R8213 S.n4482 S.n4464 0.026
R8214 S.n3682 S.n3664 0.026
R8215 S.n2870 S.n2852 0.026
R8216 S.n2025 S.n2007 0.026
R8217 S.n1584 S.n1567 0.026
R8218 S.n1555 S.n1552 0.026
R8219 S.n1145 S.n1144 0.026
R8220 S.n1996 S.n1993 0.026
R8221 S.n2424 S.n2421 0.026
R8222 S.n2841 S.n2838 0.026
R8223 S.n3280 S.n3277 0.026
R8224 S.n3653 S.n3650 0.026
R8225 S.n4127 S.n4124 0.026
R8226 S.n4453 S.n4450 0.026
R8227 S.n4917 S.n4914 0.026
R8228 S.n5230 S.n5227 0.026
R8229 S.n5698 S.n5695 0.026
R8230 S.n6290 S.n6284 0.026
R8231 S.n5530 S.n5514 0.026
R8232 S.n4421 S.n4403 0.026
R8233 S.n3621 S.n3603 0.026
R8234 S.n2809 S.n2791 0.026
R8235 S.n1962 S.n1944 0.026
R8236 S.n1525 S.n1508 0.026
R8237 S.n1496 S.n1493 0.026
R8238 S.n1111 S.n1110 0.026
R8239 S.n1933 S.n1930 0.026
R8240 S.n2388 S.n2385 0.026
R8241 S.n2780 S.n2777 0.026
R8242 S.n3244 S.n3241 0.026
R8243 S.n3592 S.n3589 0.026
R8244 S.n4091 S.n4088 0.026
R8245 S.n4748 S.n4742 0.026
R8246 S.n3953 S.n3937 0.026
R8247 S.n2748 S.n2730 0.026
R8248 S.n1899 S.n1881 0.026
R8249 S.n1469 S.n1449 0.026
R8250 S.n1437 S.n1432 0.026
R8251 S.n1077 S.n1076 0.026
R8252 S.n1870 S.n1867 0.026
R8253 S.n2352 S.n2349 0.026
R8254 S.n3136 S.n3130 0.026
R8255 S.n2306 S.n2290 0.026
R8256 S.n1407 S.n1390 0.026
R8257 S.n1378 S.n1372 0.026
R8258 S.n851 S.n848 0.026
R8259 S.n851 S.n838 0.026
R8260 S.n12009 S.n11993 0.026
R8261 S.n12654 S.n12653 0.026
R8262 S.n780 S.n779 0.026
R8263 S.n12631 S.n12630 0.026
R8264 S.t28 S.n100 0.025
R8265 S.t28 S.n4 0.025
R8266 S.t28 S.n15 0.025
R8267 S.t28 S.n26 0.025
R8268 S.t28 S.n38 0.025
R8269 S.t28 S.n70 0.025
R8270 S.t28 S.n82 0.025
R8271 S.n920 S.n919 0.024
R8272 S.n994 S.n993 0.024
R8273 S.n1838 S.n1837 0.024
R8274 S.n2721 S.n2720 0.024
R8275 S.n3562 S.n3561 0.024
R8276 S.n4394 S.n4393 0.024
R8277 S.n5200 S.n5199 0.024
R8278 S.n5997 S.n5996 0.024
R8279 S.n6768 S.n6767 0.024
R8280 S.n7530 S.n7529 0.024
R8281 S.n8266 S.n8265 0.024
R8282 S.n8993 S.n8992 0.024
R8283 S.n9694 S.n9693 0.024
R8284 S.n10386 S.n10385 0.024
R8285 S.n11045 S.n11044 0.024
R8286 S.n12288 S.n12287 0.024
R8287 S.n13158 S.n13157 0.024
R8288 S.n12313 S.n12312 0.024
R8289 S.n9708 S.n9703 0.024
R8290 S.n9036 S.n9031 0.024
R8291 S.n8341 S.n8336 0.024
R8292 S.n7634 S.n7629 0.024
R8293 S.n6904 S.n6899 0.024
R8294 S.n6162 S.n6157 0.024
R8295 S.n5397 S.n5392 0.024
R8296 S.n4620 S.n4615 0.024
R8297 S.n3820 S.n3815 0.024
R8298 S.n3008 S.n3003 0.024
R8299 S.n2168 S.n2163 0.024
R8300 S.n2220 S.n2196 0.024
R8301 S.n3058 S.n3034 0.024
R8302 S.n3870 S.n3846 0.024
R8303 S.n4670 S.n4646 0.024
R8304 S.n5447 S.n5423 0.024
R8305 S.n6212 S.n6188 0.024
R8306 S.n6954 S.n6930 0.024
R8307 S.n7684 S.n7660 0.024
R8308 S.n8391 S.n8367 0.024
R8309 S.n9086 S.n9062 0.024
R8310 S.n9758 S.n9734 0.024
R8311 S.n10418 S.n10394 0.024
R8312 S.n11122 S.n11106 0.024
R8313 S.n1763 S.n1762 0.024
R8314 S.n1735 S.n1734 0.024
R8315 S.n1007 S.n1006 0.024
R8316 S.n1807 S.n1806 0.024
R8317 S.n919 S.n918 0.024
R8318 S.n12002 S.n12001 0.023
R8319 S.n12304 S.n12291 0.023
R8320 S.n12474 S.n12466 0.023
R8321 S.n416 S.n415 0.023
R8322 S.n776 S.n775 0.023
R8323 S.n778 S.n776 0.023
R8324 S.n1734 S.n1733 0.023
R8325 S.t28 S.n920 0.023
R8326 S.n11378 S.n11377 0.023
R8327 S.n11106 S.n11105 0.023
R8328 S.n10394 S.n10393 0.023
R8329 S.n9734 S.n9733 0.023
R8330 S.n9062 S.n9061 0.023
R8331 S.n8367 S.n8366 0.023
R8332 S.n7660 S.n7659 0.023
R8333 S.n6930 S.n6929 0.023
R8334 S.n6188 S.n6187 0.023
R8335 S.n5423 S.n5422 0.023
R8336 S.n4646 S.n4645 0.023
R8337 S.n3846 S.n3845 0.023
R8338 S.n3034 S.n3033 0.023
R8339 S.n2196 S.n2195 0.023
R8340 S.n2220 S.n2200 0.023
R8341 S.n3058 S.n3038 0.023
R8342 S.n3870 S.n3850 0.023
R8343 S.n4670 S.n4650 0.023
R8344 S.n5447 S.n5427 0.023
R8345 S.n6212 S.n6192 0.023
R8346 S.n6954 S.n6934 0.023
R8347 S.n7684 S.n7664 0.023
R8348 S.n8391 S.n8371 0.023
R8349 S.n9086 S.n9066 0.023
R8350 S.n9758 S.n9738 0.023
R8351 S.n10418 S.n10398 0.023
R8352 S.n11122 S.n11110 0.023
R8353 S.n687 S.n685 0.023
R8354 S.n1762 S.n1761 0.023
R8355 S.n799 S.n798 0.023
R8356 S.n1763 S.n1759 0.023
R8357 S.n1735 S.n1731 0.023
R8358 S.n9838 S.n9837 0.023
R8359 S.n417 S.n413 0.023
R8360 S.n375 S.n374 0.023
R8361 S.n376 S.n372 0.023
R8362 S.n334 S.n333 0.023
R8363 S.n335 S.n331 0.023
R8364 S.n313 S.n312 0.023
R8365 S.n5527 S.n5526 0.023
R8366 S.n314 S.n310 0.023
R8367 S.n272 S.n271 0.023
R8368 S.n273 S.n269 0.023
R8369 S.n231 S.n230 0.023
R8370 S.n232 S.n228 0.023
R8371 S.n998 S.n996 0.023
R8372 S.n1805 S.n1804 0.023
R8373 S.n2690 S.n2688 0.023
R8374 S.n1816 S.n1815 0.023
R8375 S.n3531 S.n3529 0.023
R8376 S.n2699 S.n2698 0.023
R8377 S.n4363 S.n4361 0.023
R8378 S.n3540 S.n3539 0.023
R8379 S.n5169 S.n5167 0.023
R8380 S.n4372 S.n4371 0.023
R8381 S.n5966 S.n5964 0.023
R8382 S.n5178 S.n5177 0.023
R8383 S.n6737 S.n6735 0.023
R8384 S.n5975 S.n5974 0.023
R8385 S.n7499 S.n7497 0.023
R8386 S.n6746 S.n6745 0.023
R8387 S.n8235 S.n8233 0.023
R8388 S.n7508 S.n7507 0.023
R8389 S.n8962 S.n8960 0.023
R8390 S.n8244 S.n8243 0.023
R8391 S.n9663 S.n9661 0.023
R8392 S.n8971 S.n8970 0.023
R8393 S.n10355 S.n10353 0.023
R8394 S.n9672 S.n9671 0.023
R8395 S.n11024 S.n11022 0.023
R8396 S.n10364 S.n10363 0.023
R8397 S.n11664 S.n11662 0.023
R8398 S.n12325 S.n12317 0.023
R8399 S.n9703 S.n9700 0.023
R8400 S.n9031 S.n9028 0.023
R8401 S.n8336 S.n8333 0.023
R8402 S.n7629 S.n7626 0.023
R8403 S.n6899 S.n6896 0.023
R8404 S.n6157 S.n6155 0.023
R8405 S.n5392 S.n5389 0.023
R8406 S.n4615 S.n4612 0.023
R8407 S.n3815 S.n3812 0.023
R8408 S.n3003 S.n3001 0.023
R8409 S.n2163 S.n2161 0.023
R8410 S.n1006 S.n1003 0.023
R8411 S.n1012 S.n1011 0.023
R8412 S.n12589 S.n12588 0.022
R8413 S.n1011 S.n1010 0.022
R8414 S.n10413 S.n10409 0.022
R8415 S.n9753 S.n9749 0.022
R8416 S.n9081 S.n9077 0.022
R8417 S.n8386 S.n8382 0.022
R8418 S.n7679 S.n7675 0.022
R8419 S.n6949 S.n6945 0.022
R8420 S.n6207 S.n6203 0.022
R8421 S.n5442 S.n5438 0.022
R8422 S.n4665 S.n4661 0.022
R8423 S.n3865 S.n3861 0.022
R8424 S.n3053 S.n3049 0.022
R8425 S.n2215 S.n2211 0.022
R8426 S.n1714 S.n1710 0.022
R8427 S.n912 S.n908 0.022
R8428 S.n11703 S.n11702 0.022
R8429 S.n1825 S.n1823 0.022
R8430 S.n2708 S.n2706 0.022
R8431 S.n3549 S.n3547 0.022
R8432 S.n4381 S.n4379 0.022
R8433 S.n5187 S.n5185 0.022
R8434 S.n5984 S.n5982 0.022
R8435 S.n6755 S.n6753 0.022
R8436 S.n7517 S.n7515 0.022
R8437 S.n8253 S.n8251 0.022
R8438 S.n8980 S.n8978 0.022
R8439 S.n9681 S.n9679 0.022
R8440 S.n10373 S.n10371 0.022
R8441 S.n10497 S.n10496 0.022
R8442 S.n9820 S.n9818 0.022
R8443 S.n9162 S.n9161 0.022
R8444 S.n8453 S.n8451 0.022
R8445 S.n7760 S.n7759 0.022
R8446 S.n7016 S.n7014 0.022
R8447 S.n6288 S.n6287 0.022
R8448 S.n5509 S.n5507 0.022
R8449 S.n4746 S.n4745 0.022
R8450 S.n3932 S.n3930 0.022
R8451 S.n3134 S.n3133 0.022
R8452 S.n2285 S.n2283 0.022
R8453 S.n1376 S.n1375 0.022
R8454 S.n833 S.n831 0.022
R8455 S.n11707 S.n11706 0.022
R8456 S.n12584 S.n12581 0.021
R8457 S.n1779 S.n1778 0.021
R8458 S.n2270 S.n2269 0.021
R8459 S.n2266 S.n2265 0.021
R8460 S.n3105 S.n3104 0.021
R8461 S.n3103 S.n3102 0.021
R8462 S.n3917 S.n3916 0.021
R8463 S.n3915 S.n3914 0.021
R8464 S.n4717 S.n4716 0.021
R8465 S.n4715 S.n4714 0.021
R8466 S.n5494 S.n5493 0.021
R8467 S.n5492 S.n5491 0.021
R8468 S.n6259 S.n6258 0.021
R8469 S.n6257 S.n6256 0.021
R8470 S.n7001 S.n7000 0.021
R8471 S.n6999 S.n6998 0.021
R8472 S.n7731 S.n7730 0.021
R8473 S.n7729 S.n7728 0.021
R8474 S.n8438 S.n8437 0.021
R8475 S.n8436 S.n8435 0.021
R8476 S.n9133 S.n9132 0.021
R8477 S.n9131 S.n9130 0.021
R8478 S.n9805 S.n9804 0.021
R8479 S.n9803 S.n9802 0.021
R8480 S.n10465 S.n10464 0.021
R8481 S.n10463 S.n10462 0.021
R8482 S.n11090 S.n11089 0.021
R8483 S.n11088 S.n11087 0.021
R8484 S.n11687 S.n11686 0.021
R8485 S.n11685 S.n11684 0.021
R8486 S.n12583 S.n12582 0.021
R8487 S.n812 S.n811 0.021
R8488 S.n1015 S.n1014 0.021
R8489 S.n2181 S.n2180 0.021
R8490 S.n2177 S.n2176 0.021
R8491 S.n3019 S.n3018 0.021
R8492 S.n3017 S.n3016 0.021
R8493 S.n3831 S.n3830 0.021
R8494 S.n3829 S.n3828 0.021
R8495 S.n4631 S.n4630 0.021
R8496 S.n4629 S.n4628 0.021
R8497 S.n5408 S.n5407 0.021
R8498 S.n5406 S.n5405 0.021
R8499 S.n6173 S.n6172 0.021
R8500 S.n6171 S.n6170 0.021
R8501 S.n6915 S.n6914 0.021
R8502 S.n6913 S.n6912 0.021
R8503 S.n7645 S.n7644 0.021
R8504 S.n7643 S.n7642 0.021
R8505 S.n8352 S.n8351 0.021
R8506 S.n8350 S.n8349 0.021
R8507 S.n9047 S.n9046 0.021
R8508 S.n9045 S.n9044 0.021
R8509 S.n9719 S.n9718 0.021
R8510 S.n9717 S.n9716 0.021
R8511 S.n10491 S.n10490 0.021
R8512 S.n1668 S.n1667 0.021
R8513 S.n2117 S.n2116 0.021
R8514 S.n2113 S.n2112 0.021
R8515 S.n2958 S.n2957 0.021
R8516 S.n2956 S.n2955 0.021
R8517 S.n3770 S.n3769 0.021
R8518 S.n3768 S.n3767 0.021
R8519 S.n4570 S.n4569 0.021
R8520 S.n4568 S.n4567 0.021
R8521 S.n5347 S.n5346 0.021
R8522 S.n5345 S.n5344 0.021
R8523 S.n6112 S.n6111 0.021
R8524 S.n6110 S.n6109 0.021
R8525 S.n6854 S.n6853 0.021
R8526 S.n6852 S.n6851 0.021
R8527 S.n7584 S.n7583 0.021
R8528 S.n7582 S.n7581 0.021
R8529 S.n8291 S.n8290 0.021
R8530 S.n8289 S.n8288 0.021
R8531 S.n9156 S.n9155 0.021
R8532 S.n1609 S.n1608 0.021
R8533 S.n2054 S.n2053 0.021
R8534 S.n2050 S.n2049 0.021
R8535 S.n2897 S.n2896 0.021
R8536 S.n2895 S.n2894 0.021
R8537 S.n3709 S.n3708 0.021
R8538 S.n3707 S.n3706 0.021
R8539 S.n4509 S.n4508 0.021
R8540 S.n4507 S.n4506 0.021
R8541 S.n5286 S.n5285 0.021
R8542 S.n5284 S.n5283 0.021
R8543 S.n6051 S.n6050 0.021
R8544 S.n6049 S.n6048 0.021
R8545 S.n6793 S.n6792 0.021
R8546 S.n6791 S.n6790 0.021
R8547 S.n7754 S.n7753 0.021
R8548 S.n1550 S.n1549 0.021
R8549 S.n1991 S.n1990 0.021
R8550 S.n1987 S.n1986 0.021
R8551 S.n2836 S.n2835 0.021
R8552 S.n2834 S.n2833 0.021
R8553 S.n3648 S.n3647 0.021
R8554 S.n3646 S.n3645 0.021
R8555 S.n4448 S.n4447 0.021
R8556 S.n4446 S.n4445 0.021
R8557 S.n5225 S.n5224 0.021
R8558 S.n5223 S.n5222 0.021
R8559 S.n6282 S.n6281 0.021
R8560 S.n1491 S.n1490 0.021
R8561 S.n1928 S.n1927 0.021
R8562 S.n1924 S.n1923 0.021
R8563 S.n2775 S.n2774 0.021
R8564 S.n2773 S.n2772 0.021
R8565 S.n3587 S.n3586 0.021
R8566 S.n3585 S.n3584 0.021
R8567 S.n4740 S.n4739 0.021
R8568 S.n1435 S.n1434 0.021
R8569 S.n1865 S.n1864 0.021
R8570 S.n1861 S.n1860 0.021
R8571 S.n3128 S.n3127 0.021
R8572 S.n11381 S.n11380 0.021
R8573 S.n11670 S.n11669 0.021
R8574 S.n11073 S.n11072 0.021
R8575 S.n10448 S.n10447 0.021
R8576 S.n9788 S.n9787 0.021
R8577 S.n9116 S.n9115 0.021
R8578 S.n8421 S.n8420 0.021
R8579 S.n7714 S.n7713 0.021
R8580 S.n6984 S.n6983 0.021
R8581 S.n6242 S.n6241 0.021
R8582 S.n5477 S.n5476 0.021
R8583 S.n4700 S.n4699 0.021
R8584 S.n3900 S.n3899 0.021
R8585 S.n3088 S.n3087 0.021
R8586 S.n2251 S.n2250 0.021
R8587 S.n810 S.n809 0.021
R8588 S.n8274 S.n8273 0.021
R8589 S.n7567 S.n7566 0.021
R8590 S.n6837 S.n6836 0.021
R8591 S.n6095 S.n6094 0.021
R8592 S.n5330 S.n5329 0.021
R8593 S.n4553 S.n4552 0.021
R8594 S.n3753 S.n3752 0.021
R8595 S.n2941 S.n2940 0.021
R8596 S.n2098 S.n2097 0.021
R8597 S.n1653 S.n1652 0.021
R8598 S.n10498 S.n10497 0.021
R8599 S.n11121 S.n11120 0.021
R8600 S.n1697 S.n1696 0.021
R8601 S.n2147 S.n2146 0.021
R8602 S.n2988 S.n2987 0.021
R8603 S.n3800 S.n3799 0.021
R8604 S.n4600 S.n4599 0.021
R8605 S.n5377 S.n5376 0.021
R8606 S.n6142 S.n6141 0.021
R8607 S.n6884 S.n6883 0.021
R8608 S.n7614 S.n7613 0.021
R8609 S.n8321 S.n8320 0.021
R8610 S.n9016 S.n9015 0.021
R8611 S.n9822 S.n9820 0.021
R8612 S.n434 S.n433 0.021
R8613 S.n9163 S.n9162 0.021
R8614 S.n6776 S.n6775 0.021
R8615 S.n6034 S.n6033 0.021
R8616 S.n5269 S.n5268 0.021
R8617 S.n4492 S.n4491 0.021
R8618 S.n3692 S.n3691 0.021
R8619 S.n2880 S.n2879 0.021
R8620 S.n2035 S.n2034 0.021
R8621 S.n1594 S.n1593 0.021
R8622 S.n1639 S.n1638 0.021
R8623 S.n2084 S.n2083 0.021
R8624 S.n2927 S.n2926 0.021
R8625 S.n3739 S.n3738 0.021
R8626 S.n4539 S.n4538 0.021
R8627 S.n5316 S.n5315 0.021
R8628 S.n6081 S.n6080 0.021
R8629 S.n6823 S.n6822 0.021
R8630 S.n7553 S.n7552 0.021
R8631 S.n8455 S.n8453 0.021
R8632 S.n393 S.n392 0.021
R8633 S.n7761 S.n7760 0.021
R8634 S.n5208 S.n5207 0.021
R8635 S.n4431 S.n4430 0.021
R8636 S.n3631 S.n3630 0.021
R8637 S.n2819 S.n2818 0.021
R8638 S.n1972 S.n1971 0.021
R8639 S.n1535 S.n1534 0.021
R8640 S.n1580 S.n1579 0.021
R8641 S.n2021 S.n2020 0.021
R8642 S.n2866 S.n2865 0.021
R8643 S.n3678 S.n3677 0.021
R8644 S.n4478 S.n4477 0.021
R8645 S.n5255 S.n5254 0.021
R8646 S.n6020 S.n6019 0.021
R8647 S.n7018 S.n7016 0.021
R8648 S.n352 S.n351 0.021
R8649 S.n6289 S.n6288 0.021
R8650 S.n3570 S.n3569 0.021
R8651 S.n2758 S.n2757 0.021
R8652 S.n1909 S.n1908 0.021
R8653 S.n1476 S.n1475 0.021
R8654 S.n1521 S.n1520 0.021
R8655 S.n1958 S.n1957 0.021
R8656 S.n2805 S.n2804 0.021
R8657 S.n3617 S.n3616 0.021
R8658 S.n4417 S.n4416 0.021
R8659 S.n5511 S.n5509 0.021
R8660 S.n41 S.n40 0.021
R8661 S.n4747 S.n4746 0.021
R8662 S.n1846 S.n1845 0.021
R8663 S.n1417 S.n1416 0.021
R8664 S.n1465 S.n1464 0.021
R8665 S.n1895 S.n1894 0.021
R8666 S.n2744 S.n2743 0.021
R8667 S.n3934 S.n3932 0.021
R8668 S.n290 S.n289 0.021
R8669 S.n3135 S.n3134 0.021
R8670 S.n1403 S.n1402 0.021
R8671 S.n2287 S.n2285 0.021
R8672 S.n249 S.n248 0.021
R8673 S.n1377 S.n1376 0.021
R8674 S.n835 S.n833 0.021
R8675 S.n12385 S.n12383 0.021
R8676 S.n11030 S.n11029 0.021
R8677 S.n12324 S.n12321 0.02
R8678 S.n12473 S.n12470 0.02
R8679 S.n932 S.n931 0.02
R8680 S.n436 S.n435 0.02
R8681 S.n395 S.n394 0.02
R8682 S.n354 S.n353 0.02
R8683 S.n43 S.n42 0.02
R8684 S.n292 S.n291 0.02
R8685 S.n251 S.n250 0.02
R8686 S.n846 S.n845 0.02
R8687 S.n12554 S.n12553 0.02
R8688 S.n12590 S.n12587 0.02
R8689 S.n9703 S.n9702 0.02
R8690 S.n9031 S.n9030 0.02
R8691 S.n8336 S.n8335 0.02
R8692 S.n7629 S.n7628 0.02
R8693 S.n6899 S.n6898 0.02
R8694 S.n6157 S.n6156 0.02
R8695 S.n5392 S.n5391 0.02
R8696 S.n4615 S.n4614 0.02
R8697 S.n3815 S.n3814 0.02
R8698 S.n3003 S.n3002 0.02
R8699 S.n2163 S.n2162 0.02
R8700 S.n10498 S.n10494 0.02
R8701 S.n11704 S.n11701 0.02
R8702 S.n1006 S.n1005 0.02
R8703 S.n9822 S.n9821 0.02
R8704 S.n9163 S.n9159 0.02
R8705 S.n8455 S.n8454 0.02
R8706 S.n7761 S.n7757 0.02
R8707 S.n7018 S.n7017 0.02
R8708 S.n6289 S.n6285 0.02
R8709 S.n5511 S.n5510 0.02
R8710 S.n4747 S.n4743 0.02
R8711 S.n3934 S.n3933 0.02
R8712 S.n3135 S.n3131 0.02
R8713 S.n2287 S.n2286 0.02
R8714 S.n1377 S.n1373 0.02
R8715 S.n835 S.n834 0.02
R8716 S.n924 S.n923 0.02
R8717 S.t28 S.n214 0.019
R8718 S.n1265 S.n1263 0.019
R8719 S.n2545 S.n2543 0.019
R8720 S.n3401 S.n3399 0.019
R8721 S.n4248 S.n4246 0.019
R8722 S.n5038 S.n5036 0.019
R8723 S.n5819 S.n5817 0.019
R8724 S.n6574 S.n6572 0.019
R8725 S.n7320 S.n7318 0.019
R8726 S.n7873 S.n7871 0.019
R8727 S.n8569 S.n8567 0.019
R8728 S.n9436 S.n9434 0.019
R8729 S.n10112 S.n10110 0.019
R8730 S.n10765 S.n10763 0.019
R8731 S.n223 S.n222 0.019
R8732 S.n1284 S.n1283 0.019
R8733 S.n10417 S.n10416 0.019
R8734 S.n9757 S.n9756 0.019
R8735 S.n9085 S.n9084 0.019
R8736 S.n8390 S.n8389 0.019
R8737 S.n7683 S.n7682 0.019
R8738 S.n6953 S.n6952 0.019
R8739 S.n6211 S.n6210 0.019
R8740 S.n5446 S.n5445 0.019
R8741 S.n4669 S.n4668 0.019
R8742 S.n3869 S.n3868 0.019
R8743 S.n3057 S.n3056 0.019
R8744 S.n2219 S.n2218 0.019
R8745 S.n1718 S.n1717 0.019
R8746 S.n11944 S.n11943 0.019
R8747 S.n898 S.n897 0.018
R8748 S.n869 S.n868 0.018
R8749 S.n992 S.n991 0.018
R8750 S.n1836 S.n1835 0.018
R8751 S.n2719 S.n2718 0.018
R8752 S.n3560 S.n3559 0.018
R8753 S.n4392 S.n4391 0.018
R8754 S.n5198 S.n5197 0.018
R8755 S.n5995 S.n5994 0.018
R8756 S.n6766 S.n6765 0.018
R8757 S.n7528 S.n7527 0.018
R8758 S.n8264 S.n8263 0.018
R8759 S.n8991 S.n8990 0.018
R8760 S.n9692 S.n9691 0.018
R8761 S.n10384 S.n10383 0.018
R8762 S.n11043 S.n11042 0.018
R8763 S.n12286 S.n12285 0.018
R8764 S.n13156 S.n13155 0.018
R8765 S.n214 S.n213 0.018
R8766 S.n413 S.n412 0.018
R8767 S.n372 S.n371 0.018
R8768 S.n331 S.n330 0.018
R8769 S.n310 S.n309 0.018
R8770 S.n269 S.n268 0.018
R8771 S.n228 S.n227 0.018
R8772 S S.n985 0.018
R8773 S.n11629 S.n11628 0.018
R8774 S.n218 S.n217 0.018
R8775 S.n1005 S.n1004 0.018
R8776 S.n9702 S.n9701 0.018
R8777 S.n9030 S.n9029 0.018
R8778 S.n8335 S.n8334 0.018
R8779 S.n7628 S.n7627 0.018
R8780 S.n6898 S.n6897 0.018
R8781 S.n5391 S.n5390 0.018
R8782 S.n4614 S.n4613 0.018
R8783 S.n3814 S.n3813 0.018
R8784 S.n11626 S.n11625 0.017
R8785 S.n12628 S.n12627 0.017
R8786 S.n12651 S.n12650 0.017
R8787 S.n11633 S.n11630 0.017
R8788 S.n12301 S.n12300 0.017
R8789 S.n12300 S.n12299 0.017
R8790 S.n1828 S.n1827 0.017
R8791 S.n2711 S.n2710 0.017
R8792 S.n3552 S.n3551 0.017
R8793 S.n4384 S.n4383 0.017
R8794 S.n5190 S.n5189 0.017
R8795 S.n5987 S.n5986 0.017
R8796 S.n6758 S.n6757 0.017
R8797 S.n7520 S.n7519 0.017
R8798 S.n8256 S.n8255 0.017
R8799 S.n8983 S.n8982 0.017
R8800 S.n9684 S.n9683 0.017
R8801 S.n10376 S.n10375 0.017
R8802 S.t320 S.n1012 0.016
R8803 S.n1252 S.n1248 0.016
R8804 S.n9841 S.n9833 0.016
R8805 S.n8474 S.n8466 0.016
R8806 S.n7037 S.n7029 0.016
R8807 S.n5530 S.n5522 0.016
R8808 S.n3953 S.n3945 0.016
R8809 S.n2306 S.n2298 0.016
R8810 S.n1826 S.n1825 0.016
R8811 S.n2709 S.n2708 0.016
R8812 S.n3550 S.n3549 0.016
R8813 S.n4382 S.n4381 0.016
R8814 S.n5188 S.n5187 0.016
R8815 S.n5985 S.n5984 0.016
R8816 S.n6756 S.n6755 0.016
R8817 S.n7518 S.n7517 0.016
R8818 S.n8254 S.n8253 0.016
R8819 S.n8981 S.n8980 0.016
R8820 S.n9682 S.n9681 0.016
R8821 S.n10374 S.n10373 0.016
R8822 S.n6155 S.n6154 0.015
R8823 S.n3001 S.n3000 0.015
R8824 S.n2161 S.n2160 0.015
R8825 S.n12253 S.n12252 0.015
R8826 S.t320 S.n1008 0.015
R8827 S.n12581 S.n12580 0.015
R8828 S.n10415 S.n10414 0.015
R8829 S.n10414 S.n10413 0.015
R8830 S.n10413 S.n10412 0.015
R8831 S.n9755 S.n9754 0.015
R8832 S.n9754 S.n9753 0.015
R8833 S.n9753 S.n9752 0.015
R8834 S.n9083 S.n9082 0.015
R8835 S.n9082 S.n9081 0.015
R8836 S.n9081 S.n9080 0.015
R8837 S.n8388 S.n8387 0.015
R8838 S.n8387 S.n8386 0.015
R8839 S.n8386 S.n8385 0.015
R8840 S.n7681 S.n7680 0.015
R8841 S.n7680 S.n7679 0.015
R8842 S.n7679 S.n7678 0.015
R8843 S.n6951 S.n6950 0.015
R8844 S.n6950 S.n6949 0.015
R8845 S.n6949 S.n6948 0.015
R8846 S.n6209 S.n6208 0.015
R8847 S.n6208 S.n6207 0.015
R8848 S.n6207 S.n6206 0.015
R8849 S.n5444 S.n5443 0.015
R8850 S.n5443 S.n5442 0.015
R8851 S.n5442 S.n5441 0.015
R8852 S.n4667 S.n4666 0.015
R8853 S.n4666 S.n4665 0.015
R8854 S.n4665 S.n4664 0.015
R8855 S.n3867 S.n3866 0.015
R8856 S.n3866 S.n3865 0.015
R8857 S.n3865 S.n3864 0.015
R8858 S.n3055 S.n3054 0.015
R8859 S.n3054 S.n3053 0.015
R8860 S.n3053 S.n3052 0.015
R8861 S.n2217 S.n2216 0.015
R8862 S.n2216 S.n2215 0.015
R8863 S.n2215 S.n2214 0.015
R8864 S.n1716 S.n1715 0.015
R8865 S.n1715 S.n1714 0.015
R8866 S.n1714 S.n1713 0.015
R8867 S.n913 S.n912 0.015
R8868 S.n912 S.n911 0.015
R8869 S.n11706 S.n11705 0.015
R8870 S.n801 S.n800 0.015
R8871 S.t35 S.n12388 0.015
R8872 S.n2692 S.n1840 0.015
R8873 S.n3533 S.n2723 0.015
R8874 S.n4365 S.n3564 0.015
R8875 S.n5171 S.n4396 0.015
R8876 S.n5968 S.n5202 0.015
R8877 S.n6739 S.n5999 0.015
R8878 S.n7501 S.n6770 0.015
R8879 S.n8237 S.n7532 0.015
R8880 S.n8964 S.n8268 0.015
R8881 S.n9665 S.n8995 0.015
R8882 S.n10357 S.n9696 0.015
R8883 S.n11026 S.n10388 0.015
R8884 S.n11942 S.n11941 0.015
R8885 S.n11941 S.n11940 0.015
R8886 S.n11628 S.n11627 0.015
R8887 S.n11666 S.n11047 0.015
R8888 S.n11673 S.n11672 0.015
R8889 S.n11076 S.n11075 0.015
R8890 S.n10451 S.n10450 0.015
R8891 S.n9791 S.n9790 0.015
R8892 S.n9119 S.n9118 0.015
R8893 S.n8424 S.n8423 0.015
R8894 S.n7717 S.n7716 0.015
R8895 S.n6987 S.n6986 0.015
R8896 S.n6245 S.n6244 0.015
R8897 S.n5480 S.n5479 0.015
R8898 S.n4703 S.n4702 0.015
R8899 S.n3903 S.n3902 0.015
R8900 S.n3091 S.n3090 0.015
R8901 S.n2254 S.n2253 0.015
R8902 S.n8277 S.n8276 0.015
R8903 S.n7570 S.n7569 0.015
R8904 S.n6840 S.n6839 0.015
R8905 S.n6098 S.n6097 0.015
R8906 S.n5333 S.n5332 0.015
R8907 S.n4556 S.n4555 0.015
R8908 S.n3756 S.n3755 0.015
R8909 S.n2944 S.n2943 0.015
R8910 S.n2101 S.n2100 0.015
R8911 S.n1656 S.n1655 0.015
R8912 S.n9011 S.n9010 0.015
R8913 S.n8316 S.n8315 0.015
R8914 S.n7609 S.n7608 0.015
R8915 S.n6879 S.n6878 0.015
R8916 S.n6137 S.n6136 0.015
R8917 S.n5372 S.n5371 0.015
R8918 S.n4595 S.n4594 0.015
R8919 S.n3795 S.n3794 0.015
R8920 S.n2983 S.n2982 0.015
R8921 S.n2142 S.n2141 0.015
R8922 S.n1693 S.n1692 0.015
R8923 S.n6779 S.n6778 0.015
R8924 S.n6037 S.n6036 0.015
R8925 S.n5272 S.n5271 0.015
R8926 S.n4495 S.n4494 0.015
R8927 S.n3695 S.n3694 0.015
R8928 S.n2883 S.n2882 0.015
R8929 S.n2038 S.n2037 0.015
R8930 S.n1597 S.n1596 0.015
R8931 S.n7548 S.n7547 0.015
R8932 S.n6818 S.n6817 0.015
R8933 S.n6076 S.n6075 0.015
R8934 S.n5311 S.n5310 0.015
R8935 S.n4534 S.n4533 0.015
R8936 S.n3734 S.n3733 0.015
R8937 S.n2922 S.n2921 0.015
R8938 S.n2079 S.n2078 0.015
R8939 S.n1634 S.n1633 0.015
R8940 S.n5211 S.n5210 0.015
R8941 S.n4434 S.n4433 0.015
R8942 S.n3634 S.n3633 0.015
R8943 S.n2822 S.n2821 0.015
R8944 S.n1975 S.n1974 0.015
R8945 S.n1538 S.n1537 0.015
R8946 S.n6015 S.n6014 0.015
R8947 S.n5250 S.n5249 0.015
R8948 S.n4473 S.n4472 0.015
R8949 S.n3673 S.n3672 0.015
R8950 S.n2861 S.n2860 0.015
R8951 S.n2016 S.n2015 0.015
R8952 S.n1575 S.n1574 0.015
R8953 S.n3573 S.n3572 0.015
R8954 S.n2761 S.n2760 0.015
R8955 S.n1912 S.n1911 0.015
R8956 S.n1479 S.n1478 0.015
R8957 S.n4412 S.n4411 0.015
R8958 S.n3612 S.n3611 0.015
R8959 S.n2800 S.n2799 0.015
R8960 S.n1953 S.n1952 0.015
R8961 S.n1516 S.n1515 0.015
R8962 S.n1849 S.n1848 0.015
R8963 S.n1420 S.n1419 0.015
R8964 S.n2739 S.n2738 0.015
R8965 S.n1890 S.n1889 0.015
R8966 S.n1460 S.n1459 0.015
R8967 S.n1398 S.n1397 0.015
R8968 S.n916 S.n915 0.014
R8969 S.n11033 S.n11031 0.014
R8970 S.n1660 S.n1659 0.014
R8971 S.n2150 S.n2149 0.014
R8972 S.n2991 S.n2990 0.014
R8973 S.n3803 S.n3802 0.014
R8974 S.n4603 S.n4602 0.014
R8975 S.n5380 S.n5379 0.014
R8976 S.n6145 S.n6144 0.014
R8977 S.n6887 S.n6886 0.014
R8978 S.n7617 S.n7616 0.014
R8979 S.n8324 S.n8323 0.014
R8980 S.n9019 S.n9018 0.014
R8981 S.n1601 S.n1600 0.014
R8982 S.n2087 S.n2086 0.014
R8983 S.n2930 S.n2929 0.014
R8984 S.n3742 S.n3741 0.014
R8985 S.n4542 S.n4541 0.014
R8986 S.n5319 S.n5318 0.014
R8987 S.n6084 S.n6083 0.014
R8988 S.n6826 S.n6825 0.014
R8989 S.n7556 S.n7555 0.014
R8990 S.n1542 S.n1541 0.014
R8991 S.n2024 S.n2023 0.014
R8992 S.n2869 S.n2868 0.014
R8993 S.n3681 S.n3680 0.014
R8994 S.n4481 S.n4480 0.014
R8995 S.n5258 S.n5257 0.014
R8996 S.n6023 S.n6022 0.014
R8997 S.n1483 S.n1482 0.014
R8998 S.n1961 S.n1960 0.014
R8999 S.n2808 S.n2807 0.014
R9000 S.n3620 S.n3619 0.014
R9001 S.n4420 S.n4419 0.014
R9002 S.n1424 S.n1423 0.014
R9003 S.n1898 S.n1897 0.014
R9004 S.n2747 S.n2746 0.014
R9005 S.n13135 S.n13126 0.014
R9006 S.n12265 S.n12255 0.014
R9007 S.n1008 S.n1007 0.014
R9008 S.n1231 S.n1230 0.014
R9009 S.n2612 S.n2611 0.014
R9010 S.n3483 S.n3482 0.014
R9011 S.n4331 S.n4330 0.014
R9012 S.n5137 S.n5136 0.014
R9013 S.n5934 S.n5933 0.014
R9014 S.n6705 S.n6704 0.014
R9015 S.n7467 S.n7466 0.014
R9016 S.n8051 S.n8050 0.014
R9017 S.n8763 S.n8762 0.014
R9018 S.n9631 S.n9630 0.014
R9019 S.n10323 S.n10322 0.014
R9020 S.n10992 S.n10991 0.014
R9021 S.n12008 S.n12007 0.014
R9022 S.n11677 S.n11676 0.013
R9023 S.n11080 S.n11079 0.013
R9024 S.n10455 S.n10454 0.013
R9025 S.n9795 S.n9794 0.013
R9026 S.n9123 S.n9122 0.013
R9027 S.n8428 S.n8427 0.013
R9028 S.n7721 S.n7720 0.013
R9029 S.n6991 S.n6990 0.013
R9030 S.n6249 S.n6248 0.013
R9031 S.n5484 S.n5483 0.013
R9032 S.n4707 S.n4706 0.013
R9033 S.n3907 S.n3906 0.013
R9034 S.n3095 S.n3094 0.013
R9035 S.n2258 S.n2257 0.013
R9036 S.n8281 S.n8280 0.013
R9037 S.n7574 S.n7573 0.013
R9038 S.n6844 S.n6843 0.013
R9039 S.n6102 S.n6101 0.013
R9040 S.n5337 S.n5336 0.013
R9041 S.n4560 S.n4559 0.013
R9042 S.n3760 S.n3759 0.013
R9043 S.n2948 S.n2947 0.013
R9044 S.n2105 S.n2104 0.013
R9045 S.n1700 S.n1699 0.013
R9046 S.n6783 S.n6782 0.013
R9047 S.n6041 S.n6040 0.013
R9048 S.n5276 S.n5275 0.013
R9049 S.n4499 S.n4498 0.013
R9050 S.n3699 S.n3698 0.013
R9051 S.n2887 S.n2886 0.013
R9052 S.n2042 S.n2041 0.013
R9053 S.n1642 S.n1641 0.013
R9054 S.n5215 S.n5214 0.013
R9055 S.n4438 S.n4437 0.013
R9056 S.n3638 S.n3637 0.013
R9057 S.n2826 S.n2825 0.013
R9058 S.n1979 S.n1978 0.013
R9059 S.n1583 S.n1582 0.013
R9060 S.n3577 S.n3576 0.013
R9061 S.n2765 S.n2764 0.013
R9062 S.n1916 S.n1915 0.013
R9063 S.n1524 S.n1523 0.013
R9064 S.n1853 S.n1852 0.013
R9065 S.n1468 S.n1467 0.013
R9066 S.n1406 S.n1405 0.013
R9067 S.n11119 S.n11118 0.013
R9068 S.n2611 S.n2610 0.013
R9069 S.n3482 S.n3481 0.013
R9070 S.n4330 S.n4329 0.013
R9071 S.n5136 S.n5135 0.013
R9072 S.n5933 S.n5932 0.013
R9073 S.n6704 S.n6703 0.013
R9074 S.n7466 S.n7465 0.013
R9075 S.n8050 S.n8049 0.013
R9076 S.n8762 S.n8761 0.013
R9077 S.n9630 S.n9629 0.013
R9078 S.n10322 S.n10321 0.013
R9079 S.n10991 S.n10990 0.013
R9080 S.n12007 S.n12006 0.013
R9081 S.t28 S.n0 0.012
R9082 S.t28 S.n11 0.012
R9083 S.t28 S.n22 0.012
R9084 S.t28 S.n34 0.012
R9085 S.t28 S.n66 0.012
R9086 S.t28 S.n78 0.012
R9087 S.t28 S.n101 0.012
R9088 S.n11047 S.n11035 0.012
R9089 S.n12297 S.n12296 0.012
R9090 S.n11674 S.n11673 0.012
R9091 S.n11077 S.n11076 0.012
R9092 S.n10452 S.n10451 0.012
R9093 S.n9792 S.n9791 0.012
R9094 S.n9120 S.n9119 0.012
R9095 S.n8425 S.n8424 0.012
R9096 S.n7718 S.n7717 0.012
R9097 S.n6988 S.n6987 0.012
R9098 S.n6246 S.n6245 0.012
R9099 S.n5481 S.n5480 0.012
R9100 S.n4704 S.n4703 0.012
R9101 S.n3904 S.n3903 0.012
R9102 S.n3092 S.n3091 0.012
R9103 S.n2255 S.n2254 0.012
R9104 S.n823 S.n814 0.012
R9105 S.n8278 S.n8277 0.012
R9106 S.n7571 S.n7570 0.012
R9107 S.n6841 S.n6840 0.012
R9108 S.n6099 S.n6098 0.012
R9109 S.n5334 S.n5333 0.012
R9110 S.n4557 S.n4556 0.012
R9111 S.n3757 S.n3756 0.012
R9112 S.n2945 S.n2944 0.012
R9113 S.n2102 S.n2101 0.012
R9114 S.n1657 S.n1656 0.012
R9115 S.n9012 S.n9011 0.012
R9116 S.n8317 S.n8316 0.012
R9117 S.n7610 S.n7609 0.012
R9118 S.n6880 S.n6879 0.012
R9119 S.n6138 S.n6137 0.012
R9120 S.n5373 S.n5372 0.012
R9121 S.n4596 S.n4595 0.012
R9122 S.n3796 S.n3795 0.012
R9123 S.n2984 S.n2983 0.012
R9124 S.n2143 S.n2142 0.012
R9125 S.n1001 S.n1000 0.012
R9126 S.n9706 S.n9705 0.012
R9127 S.n9034 S.n9033 0.012
R9128 S.n8339 S.n8338 0.012
R9129 S.n7632 S.n7631 0.012
R9130 S.n6902 S.n6901 0.012
R9131 S.n6160 S.n6159 0.012
R9132 S.n5395 S.n5394 0.012
R9133 S.n4618 S.n4617 0.012
R9134 S.n3818 S.n3817 0.012
R9135 S.n3006 S.n3005 0.012
R9136 S.n2166 S.n2165 0.012
R9137 S.n1694 S.n1693 0.012
R9138 S.n446 S.n438 0.012
R9139 S.n6780 S.n6779 0.012
R9140 S.n6038 S.n6037 0.012
R9141 S.n5273 S.n5272 0.012
R9142 S.n4496 S.n4495 0.012
R9143 S.n3696 S.n3695 0.012
R9144 S.n2884 S.n2883 0.012
R9145 S.n2039 S.n2038 0.012
R9146 S.n1598 S.n1597 0.012
R9147 S.n7549 S.n7548 0.012
R9148 S.n6819 S.n6818 0.012
R9149 S.n6077 S.n6076 0.012
R9150 S.n5312 S.n5311 0.012
R9151 S.n4535 S.n4534 0.012
R9152 S.n3735 S.n3734 0.012
R9153 S.n2923 S.n2922 0.012
R9154 S.n2080 S.n2079 0.012
R9155 S.n1635 S.n1634 0.012
R9156 S.n405 S.n397 0.012
R9157 S.n5212 S.n5211 0.012
R9158 S.n4435 S.n4434 0.012
R9159 S.n3635 S.n3634 0.012
R9160 S.n2823 S.n2822 0.012
R9161 S.n1976 S.n1975 0.012
R9162 S.n1539 S.n1538 0.012
R9163 S.n6016 S.n6015 0.012
R9164 S.n5251 S.n5250 0.012
R9165 S.n4474 S.n4473 0.012
R9166 S.n3674 S.n3673 0.012
R9167 S.n2862 S.n2861 0.012
R9168 S.n2017 S.n2016 0.012
R9169 S.n1576 S.n1575 0.012
R9170 S.n364 S.n356 0.012
R9171 S.n3574 S.n3573 0.012
R9172 S.n2762 S.n2761 0.012
R9173 S.n1913 S.n1912 0.012
R9174 S.n1480 S.n1479 0.012
R9175 S.n4413 S.n4412 0.012
R9176 S.n3613 S.n3612 0.012
R9177 S.n2801 S.n2800 0.012
R9178 S.n1954 S.n1953 0.012
R9179 S.n1517 S.n1516 0.012
R9180 S.n59 S.n45 0.012
R9181 S.n1850 S.n1849 0.012
R9182 S.n1421 S.n1420 0.012
R9183 S.n2740 S.n2739 0.012
R9184 S.n1891 S.n1890 0.012
R9185 S.n1461 S.n1460 0.012
R9186 S.n302 S.n294 0.012
R9187 S.n1399 S.n1398 0.012
R9188 S.n261 S.n253 0.012
R9189 S.n2610 S.n2609 0.012
R9190 S.n1823 S.n1822 0.012
R9191 S.n3481 S.n3480 0.012
R9192 S.n2706 S.n2705 0.012
R9193 S.n4329 S.n4328 0.012
R9194 S.n3547 S.n3546 0.012
R9195 S.n5135 S.n5134 0.012
R9196 S.n4379 S.n4378 0.012
R9197 S.n5932 S.n5931 0.012
R9198 S.n5185 S.n5184 0.012
R9199 S.n6703 S.n6702 0.012
R9200 S.n5982 S.n5981 0.012
R9201 S.n7465 S.n7464 0.012
R9202 S.n6753 S.n6752 0.012
R9203 S.n8049 S.n8048 0.012
R9204 S.n7515 S.n7514 0.012
R9205 S.n8761 S.n8760 0.012
R9206 S.n8251 S.n8250 0.012
R9207 S.n9629 S.n9628 0.012
R9208 S.n8978 S.n8977 0.012
R9209 S.n10321 S.n10320 0.012
R9210 S.n9679 S.n9678 0.012
R9211 S.n10990 S.n10989 0.012
R9212 S.n10371 S.n10370 0.012
R9213 S.n12320 S.n12319 0.012
R9214 S.n12469 S.n12468 0.012
R9215 S.n12006 S.n12005 0.012
R9216 S.n12640 S.n12631 0.011
R9217 S.n12663 S.n12654 0.011
R9218 S.n11633 S.n11626 0.01
R9219 S.n661 S.n660 0.01
R9220 S.n628 S.n627 0.01
R9221 S.n595 S.n594 0.01
R9222 S.n562 S.n561 0.01
R9223 S.n529 S.n528 0.01
R9224 S.n496 S.n495 0.01
R9225 S.n10480 S.n10479 0.01
R9226 S.n780 S.n778 0.01
R9227 S.n1273 S.n1265 0.01
R9228 S.n2553 S.n2545 0.01
R9229 S.n3409 S.n3401 0.01
R9230 S.n4256 S.n4248 0.01
R9231 S.n5046 S.n5038 0.01
R9232 S.n5827 S.n5819 0.01
R9233 S.n6582 S.n6574 0.01
R9234 S.n7328 S.n7320 0.01
R9235 S.n7881 S.n7873 0.01
R9236 S.n8577 S.n8569 0.01
R9237 S.n9444 S.n9436 0.01
R9238 S.n10120 S.n10112 0.01
R9239 S.n10773 S.n10765 0.01
R9240 S.n690 S.n687 0.01
R9241 S.n11414 S.n11410 0.01
R9242 S.n10793 S.n10789 0.01
R9243 S.n10140 S.n10136 0.01
R9244 S.n9464 S.n9460 0.01
R9245 S.n8597 S.n8593 0.01
R9246 S.n7901 S.n7897 0.01
R9247 S.n7348 S.n7344 0.01
R9248 S.n6602 S.n6598 0.01
R9249 S.n5847 S.n5843 0.01
R9250 S.n5066 S.n5062 0.01
R9251 S.n4276 S.n4272 0.01
R9252 S.n3429 S.n3425 0.01
R9253 S.n2573 S.n2569 0.01
R9254 S.n1293 S.n1284 0.01
R9255 S.n709 S.n706 0.01
R9256 S.n417 S.n416 0.01
R9257 S.n376 S.n375 0.01
R9258 S.n335 S.n334 0.01
R9259 S.n314 S.n313 0.01
R9260 S.n273 S.n272 0.01
R9261 S.n232 S.n231 0.01
R9262 S.n748 S.n745 0.01
R9263 S.n1808 S.n1805 0.01
R9264 S.n1808 S.n998 0.01
R9265 S.n2692 S.n2690 0.01
R9266 S.n3533 S.n3531 0.01
R9267 S.n4365 S.n4363 0.01
R9268 S.n5171 S.n5169 0.01
R9269 S.n5968 S.n5966 0.01
R9270 S.n6739 S.n6737 0.01
R9271 S.n7501 S.n7499 0.01
R9272 S.n8237 S.n8235 0.01
R9273 S.n8964 S.n8962 0.01
R9274 S.n9665 S.n9663 0.01
R9275 S.n10357 S.n10355 0.01
R9276 S.n11026 S.n11024 0.01
R9277 S.n11666 S.n11664 0.01
R9278 S.n12640 S.n12628 0.01
R9279 S.n12663 S.n12651 0.01
R9280 S.n12306 S.n12304 0.01
R9281 S.n438 S.n437 0.01
R9282 S.n397 S.n396 0.01
R9283 S.n356 S.n355 0.01
R9284 S.n45 S.n44 0.01
R9285 S.n294 S.n293 0.01
R9286 S.n253 S.n252 0.01
R9287 S.n12299 S.n12297 0.01
R9288 S.n1251 S.n1249 0.01
R9289 S.n415 S.n414 0.01
R9290 S.n374 S.n373 0.01
R9291 S.n333 S.n332 0.01
R9292 S.n312 S.n311 0.01
R9293 S.n271 S.n270 0.01
R9294 S.n230 S.n229 0.01
R9295 S.n11395 S.n11381 0.01
R9296 S.n10081 S.n10066 0.01
R9297 S.n8502 S.n8487 0.01
R9298 S.n7217 S.n7202 0.01
R9299 S.n5680 S.n5665 0.01
R9300 S.n4073 S.n4058 0.01
R9301 S.n2334 S.n2319 0.01
R9302 S.n13161 S.n12550 0.009
R9303 S.n12302 S.n12301 0.009
R9304 S.n11122 S.n11121 0.009
R9305 S.t35 S.n12385 0.009
R9306 S.n12306 S.n12290 0.009
R9307 S.n12627 S.n12626 0.008
R9308 S.n12650 S.n12649 0.008
R9309 S.n12324 S.n12323 0.008
R9310 S.n12473 S.n12472 0.008
R9311 S.n11675 S.n11674 0.008
R9312 S.n11078 S.n11077 0.008
R9313 S.n10453 S.n10452 0.008
R9314 S.n9793 S.n9792 0.008
R9315 S.n9121 S.n9120 0.008
R9316 S.n8426 S.n8425 0.008
R9317 S.n7719 S.n7718 0.008
R9318 S.n6989 S.n6988 0.008
R9319 S.n6247 S.n6246 0.008
R9320 S.n5482 S.n5481 0.008
R9321 S.n4705 S.n4704 0.008
R9322 S.n3905 S.n3904 0.008
R9323 S.n3093 S.n3092 0.008
R9324 S.n2256 S.n2255 0.008
R9325 S.n8279 S.n8278 0.008
R9326 S.n7572 S.n7571 0.008
R9327 S.n6842 S.n6841 0.008
R9328 S.n6100 S.n6099 0.008
R9329 S.n5335 S.n5334 0.008
R9330 S.n4558 S.n4557 0.008
R9331 S.n3758 S.n3757 0.008
R9332 S.n2946 S.n2945 0.008
R9333 S.n2103 S.n2102 0.008
R9334 S.n1658 S.n1657 0.008
R9335 S.n9013 S.n9012 0.008
R9336 S.n8318 S.n8317 0.008
R9337 S.n7611 S.n7610 0.008
R9338 S.n6881 S.n6880 0.008
R9339 S.n6139 S.n6138 0.008
R9340 S.n5374 S.n5373 0.008
R9341 S.n4597 S.n4596 0.008
R9342 S.n3797 S.n3796 0.008
R9343 S.n2985 S.n2984 0.008
R9344 S.n2144 S.n2143 0.008
R9345 S.n1695 S.n1694 0.008
R9346 S.n6781 S.n6780 0.008
R9347 S.n6039 S.n6038 0.008
R9348 S.n5274 S.n5273 0.008
R9349 S.n4497 S.n4496 0.008
R9350 S.n3697 S.n3696 0.008
R9351 S.n2885 S.n2884 0.008
R9352 S.n2040 S.n2039 0.008
R9353 S.n1599 S.n1598 0.008
R9354 S.n7550 S.n7549 0.008
R9355 S.n6820 S.n6819 0.008
R9356 S.n6078 S.n6077 0.008
R9357 S.n5313 S.n5312 0.008
R9358 S.n4536 S.n4535 0.008
R9359 S.n3736 S.n3735 0.008
R9360 S.n2924 S.n2923 0.008
R9361 S.n2081 S.n2080 0.008
R9362 S.n1636 S.n1635 0.008
R9363 S.n5213 S.n5212 0.008
R9364 S.n4436 S.n4435 0.008
R9365 S.n3636 S.n3635 0.008
R9366 S.n2824 S.n2823 0.008
R9367 S.n1977 S.n1976 0.008
R9368 S.n1540 S.n1539 0.008
R9369 S.n6017 S.n6016 0.008
R9370 S.n5252 S.n5251 0.008
R9371 S.n4475 S.n4474 0.008
R9372 S.n3675 S.n3674 0.008
R9373 S.n2863 S.n2862 0.008
R9374 S.n2018 S.n2017 0.008
R9375 S.n1577 S.n1576 0.008
R9376 S.n3575 S.n3574 0.008
R9377 S.n2763 S.n2762 0.008
R9378 S.n1914 S.n1913 0.008
R9379 S.n1481 S.n1480 0.008
R9380 S.n4414 S.n4413 0.008
R9381 S.n3614 S.n3613 0.008
R9382 S.n2802 S.n2801 0.008
R9383 S.n1955 S.n1954 0.008
R9384 S.n1518 S.n1517 0.008
R9385 S.n1851 S.n1850 0.008
R9386 S.n1422 S.n1421 0.008
R9387 S.n2741 S.n2740 0.008
R9388 S.n1892 S.n1891 0.008
R9389 S.n1462 S.n1461 0.008
R9390 S.n1400 S.n1399 0.008
R9391 S.n1784 S.n1783 0.008
R9392 S.n2268 S.n2267 0.008
R9393 S.n2274 S.n2273 0.008
R9394 S.n2591 S.n2590 0.008
R9395 S.n3109 S.n3108 0.008
R9396 S.n3447 S.n3446 0.008
R9397 S.n3921 S.n3920 0.008
R9398 S.n4294 S.n4293 0.008
R9399 S.n4721 S.n4720 0.008
R9400 S.n5084 S.n5083 0.008
R9401 S.n5498 S.n5497 0.008
R9402 S.n5865 S.n5864 0.008
R9403 S.n6263 S.n6262 0.008
R9404 S.n6620 S.n6619 0.008
R9405 S.n7005 S.n7004 0.008
R9406 S.n7366 S.n7365 0.008
R9407 S.n7735 S.n7734 0.008
R9408 S.n7919 S.n7918 0.008
R9409 S.n8442 S.n8441 0.008
R9410 S.n8615 S.n8614 0.008
R9411 S.n9137 S.n9136 0.008
R9412 S.n9482 S.n9481 0.008
R9413 S.n9809 S.n9808 0.008
R9414 S.n10158 S.n10157 0.008
R9415 S.n10469 S.n10468 0.008
R9416 S.n10811 S.n10810 0.008
R9417 S.n11094 S.n11093 0.008
R9418 S.n11432 S.n11431 0.008
R9419 S.n11691 S.n11690 0.008
R9420 S.n11984 S.n11983 0.008
R9421 S.n718 S.n717 0.008
R9422 S.n1019 S.n1018 0.008
R9423 S.n2179 S.n2178 0.008
R9424 S.n2185 S.n2184 0.008
R9425 S.n2531 S.n2530 0.008
R9426 S.n3023 S.n3022 0.008
R9427 S.n3387 S.n3386 0.008
R9428 S.n3835 S.n3834 0.008
R9429 S.n4234 S.n4233 0.008
R9430 S.n4635 S.n4634 0.008
R9431 S.n5024 S.n5023 0.008
R9432 S.n5412 S.n5411 0.008
R9433 S.n5805 S.n5804 0.008
R9434 S.n6177 S.n6176 0.008
R9435 S.n6560 S.n6559 0.008
R9436 S.n6919 S.n6918 0.008
R9437 S.n7306 S.n7305 0.008
R9438 S.n7649 S.n7648 0.008
R9439 S.n7859 S.n7858 0.008
R9440 S.n8356 S.n8355 0.008
R9441 S.n8555 S.n8554 0.008
R9442 S.n9051 S.n9050 0.008
R9443 S.n9422 S.n9421 0.008
R9444 S.n9723 S.n9722 0.008
R9445 S.n10098 S.n10097 0.008
R9446 S.n1273 S.n1262 0.008
R9447 S.n2553 S.n2542 0.008
R9448 S.n3409 S.n3398 0.008
R9449 S.n4256 S.n4245 0.008
R9450 S.n5046 S.n5035 0.008
R9451 S.n5827 S.n5816 0.008
R9452 S.n6582 S.n6571 0.008
R9453 S.n7328 S.n7317 0.008
R9454 S.n7881 S.n7870 0.008
R9455 S.n8577 S.n8566 0.008
R9456 S.n9444 S.n9433 0.008
R9457 S.n10120 S.n10109 0.008
R9458 S.n10773 S.n10762 0.008
R9459 S.n690 S.n689 0.008
R9460 S.n11414 S.n11413 0.008
R9461 S.n10793 S.n10792 0.008
R9462 S.n10140 S.n10139 0.008
R9463 S.n9464 S.n9463 0.008
R9464 S.n8597 S.n8596 0.008
R9465 S.n7901 S.n7900 0.008
R9466 S.n7348 S.n7347 0.008
R9467 S.n6602 S.n6601 0.008
R9468 S.n5847 S.n5846 0.008
R9469 S.n5066 S.n5065 0.008
R9470 S.n4276 S.n4275 0.008
R9471 S.n3429 S.n3428 0.008
R9472 S.n2573 S.n2572 0.008
R9473 S.n1293 S.n1282 0.008
R9474 S.n1743 S.n1742 0.008
R9475 S.n2228 S.n2227 0.008
R9476 S.n3066 S.n3065 0.008
R9477 S.n3878 S.n3877 0.008
R9478 S.n4678 S.n4677 0.008
R9479 S.n5455 S.n5454 0.008
R9480 S.n6220 S.n6219 0.008
R9481 S.n6962 S.n6961 0.008
R9482 S.n7692 S.n7691 0.008
R9483 S.n8399 S.n8398 0.008
R9484 S.n9094 S.n9093 0.008
R9485 S.n9766 S.n9765 0.008
R9486 S.n10426 S.n10425 0.008
R9487 S.n11051 S.n11050 0.008
R9488 S.n788 S.n787 0.008
R9489 S.n800 S.n796 0.008
R9490 S.n800 S.n799 0.008
R9491 S.n709 S.n708 0.008
R9492 S.n9840 S.n9838 0.008
R9493 S.n8999 S.n8998 0.008
R9494 S.n8304 S.n8303 0.008
R9495 S.n7597 S.n7596 0.008
R9496 S.n6867 S.n6866 0.008
R9497 S.n6125 S.n6124 0.008
R9498 S.n5360 S.n5359 0.008
R9499 S.n4583 S.n4582 0.008
R9500 S.n3783 S.n3782 0.008
R9501 S.n2971 S.n2970 0.008
R9502 S.n2130 S.n2129 0.008
R9503 S.n1682 S.n1681 0.008
R9504 S.n1672 S.n1671 0.008
R9505 S.n2115 S.n2114 0.008
R9506 S.n2121 S.n2120 0.008
R9507 S.n2495 S.n2494 0.008
R9508 S.n2962 S.n2961 0.008
R9509 S.n3351 S.n3350 0.008
R9510 S.n3774 S.n3773 0.008
R9511 S.n4198 S.n4197 0.008
R9512 S.n4574 S.n4573 0.008
R9513 S.n4988 S.n4987 0.008
R9514 S.n5351 S.n5350 0.008
R9515 S.n5769 S.n5768 0.008
R9516 S.n6116 S.n6115 0.008
R9517 S.n6524 S.n6523 0.008
R9518 S.n6858 S.n6857 0.008
R9519 S.n7270 S.n7269 0.008
R9520 S.n7588 S.n7587 0.008
R9521 S.n7823 S.n7822 0.008
R9522 S.n8295 S.n8294 0.008
R9523 S.n8519 S.n8518 0.008
R9524 S.n8473 S.n8469 0.008
R9525 S.n7536 S.n7535 0.008
R9526 S.n6806 S.n6805 0.008
R9527 S.n6064 S.n6063 0.008
R9528 S.n5299 S.n5298 0.008
R9529 S.n4522 S.n4521 0.008
R9530 S.n3722 S.n3721 0.008
R9531 S.n2910 S.n2909 0.008
R9532 S.n2067 S.n2066 0.008
R9533 S.n1623 S.n1622 0.008
R9534 S.n1613 S.n1612 0.008
R9535 S.n2052 S.n2051 0.008
R9536 S.n2058 S.n2057 0.008
R9537 S.n2459 S.n2458 0.008
R9538 S.n2901 S.n2900 0.008
R9539 S.n3315 S.n3314 0.008
R9540 S.n3713 S.n3712 0.008
R9541 S.n4162 S.n4161 0.008
R9542 S.n4513 S.n4512 0.008
R9543 S.n4952 S.n4951 0.008
R9544 S.n5290 S.n5289 0.008
R9545 S.n5733 S.n5732 0.008
R9546 S.n6055 S.n6054 0.008
R9547 S.n6488 S.n6487 0.008
R9548 S.n6797 S.n6796 0.008
R9549 S.n7234 S.n7233 0.008
R9550 S.n7036 S.n7032 0.008
R9551 S.n6003 S.n6002 0.008
R9552 S.n5238 S.n5237 0.008
R9553 S.n4461 S.n4460 0.008
R9554 S.n3661 S.n3660 0.008
R9555 S.n2849 S.n2848 0.008
R9556 S.n2004 S.n2003 0.008
R9557 S.n1564 S.n1563 0.008
R9558 S.n1554 S.n1553 0.008
R9559 S.n1989 S.n1988 0.008
R9560 S.n1995 S.n1994 0.008
R9561 S.n2423 S.n2422 0.008
R9562 S.n2840 S.n2839 0.008
R9563 S.n3279 S.n3278 0.008
R9564 S.n3652 S.n3651 0.008
R9565 S.n4126 S.n4125 0.008
R9566 S.n4452 S.n4451 0.008
R9567 S.n4916 S.n4915 0.008
R9568 S.n5229 S.n5228 0.008
R9569 S.n5697 S.n5696 0.008
R9570 S.n5529 S.n5527 0.008
R9571 S.n4400 S.n4399 0.008
R9572 S.n3600 S.n3599 0.008
R9573 S.n2788 S.n2787 0.008
R9574 S.n1941 S.n1940 0.008
R9575 S.n1505 S.n1504 0.008
R9576 S.n1495 S.n1494 0.008
R9577 S.n1926 S.n1925 0.008
R9578 S.n1932 S.n1931 0.008
R9579 S.n2387 S.n2386 0.008
R9580 S.n2779 S.n2778 0.008
R9581 S.n3243 S.n3242 0.008
R9582 S.n3591 S.n3590 0.008
R9583 S.n4090 S.n4089 0.008
R9584 S.n3952 S.n3948 0.008
R9585 S.n2727 S.n2726 0.008
R9586 S.n1878 S.n1877 0.008
R9587 S.n1446 S.n1445 0.008
R9588 S.n1436 S.n1433 0.008
R9589 S.n1863 S.n1862 0.008
R9590 S.n1869 S.n1868 0.008
R9591 S.n2351 S.n2350 0.008
R9592 S.n2305 S.n2301 0.008
R9593 S.n1387 S.n1386 0.008
R9594 S.n850 S.n849 0.008
R9595 S.n748 S.n747 0.008
R9596 S.n880 S.n879 0.008
R9597 S.n11633 S.n11632 0.008
R9598 S.n12552 S.n12551 0.008
R9599 S.n900 S.n899 0.008
R9600 S.n900 S.n898 0.007
R9601 S.t28 S.n206 0.007
R9602 S.t28 S.n199 0.007
R9603 S.t28 S.n187 0.007
R9604 S.t28 S.n175 0.007
R9605 S.t28 S.n162 0.007
R9606 S.t28 S.n149 0.007
R9607 S.t28 S.n136 0.007
R9608 S.n915 S.n914 0.007
R9609 S.n11625 S.n11624 0.007
R9610 S.t35 S.n12379 0.006
R9611 S.t35 S.n12375 0.006
R9612 S.t35 S.n12371 0.006
R9613 S.t35 S.n12367 0.006
R9614 S.t35 S.n12363 0.006
R9615 S.t35 S.n12359 0.006
R9616 S.t35 S.n12355 0.006
R9617 S.t35 S.n12351 0.006
R9618 S.t35 S.n12347 0.006
R9619 S.t35 S.n12343 0.006
R9620 S.t35 S.n12339 0.006
R9621 S.t35 S.n12335 0.006
R9622 S.t35 S.n12328 0.006
R9623 S.n2269 S.n2268 0.006
R9624 S.n2180 S.n2179 0.006
R9625 S.n2116 S.n2115 0.006
R9626 S.n2053 S.n2052 0.006
R9627 S.n1990 S.n1989 0.006
R9628 S.n1927 S.n1926 0.006
R9629 S.n1436 S.n1435 0.006
R9630 S.n1864 S.n1863 0.006
R9631 S.n12553 S.n12552 0.006
R9632 S.n12325 S.n12324 0.006
R9633 S.n12474 S.n12473 0.006
R9634 S.n426 S.n417 0.006
R9635 S.n385 S.n376 0.006
R9636 S.n344 S.n335 0.006
R9637 S.n323 S.n314 0.006
R9638 S.n282 S.n273 0.006
R9639 S.n241 S.n232 0.006
R9640 S.n780 S.n767 0.005
R9641 S.n1002 S.n1001 0.005
R9642 S.n9707 S.n9706 0.005
R9643 S.n9035 S.n9034 0.005
R9644 S.n8340 S.n8339 0.005
R9645 S.n7633 S.n7632 0.005
R9646 S.n6903 S.n6902 0.005
R9647 S.n6161 S.n6160 0.005
R9648 S.n5396 S.n5395 0.005
R9649 S.n4619 S.n4618 0.005
R9650 S.n3819 S.n3818 0.005
R9651 S.n3007 S.n3006 0.005
R9652 S.n2167 S.n2166 0.005
R9653 S.t28 S.n211 0.005
R9654 S.n9835 S.n9834 0.005
R9655 S.n8468 S.n8467 0.005
R9656 S.n7031 S.n7030 0.005
R9657 S.n5524 S.n5523 0.005
R9658 S.n3947 S.n3946 0.005
R9659 S.n2300 S.n2299 0.005
R9660 S.n12323 S.n12322 0.005
R9661 S.n12472 S.n12471 0.005
R9662 S.t28 S.n917 0.005
R9663 S.n12638 S.n12637 0.004
R9664 S.n12562 S.n12561 0.004
R9665 S.n12000 S.n11999 0.004
R9666 S.n12278 S.n12277 0.004
R9667 S.n844 S.n843 0.004
R9668 S.n821 S.n820 0.004
R9669 S.n1774 S.n1773 0.004
R9670 S.n12576 S.n12575 0.004
R9671 S.n11977 S.n11976 0.004
R9672 S.n11680 S.n11679 0.004
R9673 S.n11425 S.n11424 0.004
R9674 S.n11083 S.n11082 0.004
R9675 S.n10804 S.n10803 0.004
R9676 S.n10458 S.n10457 0.004
R9677 S.n10151 S.n10150 0.004
R9678 S.n9798 S.n9797 0.004
R9679 S.n9475 S.n9474 0.004
R9680 S.n9126 S.n9125 0.004
R9681 S.n8608 S.n8607 0.004
R9682 S.n8431 S.n8430 0.004
R9683 S.n7912 S.n7911 0.004
R9684 S.n7724 S.n7723 0.004
R9685 S.n7359 S.n7358 0.004
R9686 S.n6994 S.n6993 0.004
R9687 S.n6613 S.n6612 0.004
R9688 S.n6252 S.n6251 0.004
R9689 S.n5858 S.n5857 0.004
R9690 S.n5487 S.n5486 0.004
R9691 S.n5077 S.n5076 0.004
R9692 S.n4710 S.n4709 0.004
R9693 S.n4287 S.n4286 0.004
R9694 S.n3910 S.n3909 0.004
R9695 S.n3440 S.n3439 0.004
R9696 S.n3098 S.n3097 0.004
R9697 S.n2584 S.n2583 0.004
R9698 S.n2261 S.n2260 0.004
R9699 S.n1304 S.n1303 0.004
R9700 S.n727 S.n726 0.004
R9701 S.n424 S.n423 0.004
R9702 S.n1663 S.n1662 0.004
R9703 S.n9150 S.n9149 0.004
R9704 S.n8512 S.n8511 0.004
R9705 S.n8284 S.n8283 0.004
R9706 S.n7816 S.n7815 0.004
R9707 S.n7577 S.n7576 0.004
R9708 S.n7263 S.n7262 0.004
R9709 S.n6847 S.n6846 0.004
R9710 S.n6517 S.n6516 0.004
R9711 S.n6105 S.n6104 0.004
R9712 S.n5762 S.n5761 0.004
R9713 S.n5340 S.n5339 0.004
R9714 S.n4981 S.n4980 0.004
R9715 S.n4563 S.n4562 0.004
R9716 S.n4191 S.n4190 0.004
R9717 S.n3763 S.n3762 0.004
R9718 S.n3344 S.n3343 0.004
R9719 S.n2951 S.n2950 0.004
R9720 S.n2488 S.n2487 0.004
R9721 S.n2108 S.n2107 0.004
R9722 S.n1207 S.n1206 0.004
R9723 S.n444 S.n443 0.004
R9724 S.n9832 S.n9831 0.004
R9725 S.n9402 S.n9401 0.004
R9726 S.n9009 S.n9008 0.004
R9727 S.n8535 S.n8534 0.004
R9728 S.n8314 S.n8313 0.004
R9729 S.n7839 S.n7838 0.004
R9730 S.n7607 S.n7606 0.004
R9731 S.n7286 S.n7285 0.004
R9732 S.n6877 S.n6876 0.004
R9733 S.n6540 S.n6539 0.004
R9734 S.n6135 S.n6134 0.004
R9735 S.n5785 S.n5784 0.004
R9736 S.n5370 S.n5369 0.004
R9737 S.n5004 S.n5003 0.004
R9738 S.n4593 S.n4592 0.004
R9739 S.n4214 S.n4213 0.004
R9740 S.n3793 S.n3792 0.004
R9741 S.n3367 S.n3366 0.004
R9742 S.n2981 S.n2980 0.004
R9743 S.n2511 S.n2510 0.004
R9744 S.n2140 S.n2139 0.004
R9745 S.n1228 S.n1227 0.004
R9746 S.n1247 S.n1246 0.004
R9747 S.n763 S.n762 0.004
R9748 S.n774 S.n773 0.004
R9749 S.n2172 S.n2171 0.004
R9750 S.n3012 S.n3011 0.004
R9751 S.n3824 S.n3823 0.004
R9752 S.n4624 S.n4623 0.004
R9753 S.n5401 S.n5400 0.004
R9754 S.n6166 S.n6165 0.004
R9755 S.n6908 S.n6907 0.004
R9756 S.n7638 S.n7637 0.004
R9757 S.n8345 S.n8344 0.004
R9758 S.n9040 S.n9039 0.004
R9759 S.n9712 S.n9711 0.004
R9760 S.n10485 S.n10484 0.004
R9761 S.n10091 S.n10090 0.004
R9762 S.n9415 S.n9414 0.004
R9763 S.n8548 S.n8547 0.004
R9764 S.n7852 S.n7851 0.004
R9765 S.n7299 S.n7298 0.004
R9766 S.n6553 S.n6552 0.004
R9767 S.n5798 S.n5797 0.004
R9768 S.n5017 S.n5016 0.004
R9769 S.n4227 S.n4226 0.004
R9770 S.n3380 S.n3379 0.004
R9771 S.n2524 S.n2523 0.004
R9772 S.n1725 S.n1724 0.004
R9773 S.n684 S.n683 0.004
R9774 S.n894 S.n893 0.004
R9775 S.n11114 S.n11113 0.004
R9776 S.n10768 S.n10767 0.004
R9777 S.n10403 S.n10402 0.004
R9778 S.n10115 S.n10114 0.004
R9779 S.n9743 S.n9742 0.004
R9780 S.n9439 S.n9438 0.004
R9781 S.n9071 S.n9070 0.004
R9782 S.n8572 S.n8571 0.004
R9783 S.n8376 S.n8375 0.004
R9784 S.n7876 S.n7875 0.004
R9785 S.n7669 S.n7668 0.004
R9786 S.n7323 S.n7322 0.004
R9787 S.n6939 S.n6938 0.004
R9788 S.n6577 S.n6576 0.004
R9789 S.n6197 S.n6196 0.004
R9790 S.n5822 S.n5821 0.004
R9791 S.n5432 S.n5431 0.004
R9792 S.n5041 S.n5040 0.004
R9793 S.n4655 S.n4654 0.004
R9794 S.n4251 S.n4250 0.004
R9795 S.n3855 S.n3854 0.004
R9796 S.n3404 S.n3403 0.004
R9797 S.n3043 S.n3042 0.004
R9798 S.n2548 S.n2547 0.004
R9799 S.n2205 S.n2204 0.004
R9800 S.n1268 S.n1267 0.004
R9801 S.n1753 S.n1752 0.004
R9802 S.n704 S.n703 0.004
R9803 S.n1287 S.n1286 0.004
R9804 S.n2238 S.n2237 0.004
R9805 S.n2568 S.n2567 0.004
R9806 S.n3076 S.n3075 0.004
R9807 S.n3424 S.n3423 0.004
R9808 S.n3888 S.n3887 0.004
R9809 S.n4271 S.n4270 0.004
R9810 S.n4688 S.n4687 0.004
R9811 S.n5061 S.n5060 0.004
R9812 S.n5465 S.n5464 0.004
R9813 S.n5842 S.n5841 0.004
R9814 S.n6230 S.n6229 0.004
R9815 S.n6597 S.n6596 0.004
R9816 S.n6972 S.n6971 0.004
R9817 S.n7343 S.n7342 0.004
R9818 S.n7702 S.n7701 0.004
R9819 S.n7896 S.n7895 0.004
R9820 S.n8409 S.n8408 0.004
R9821 S.n8592 S.n8591 0.004
R9822 S.n9104 S.n9103 0.004
R9823 S.n9459 S.n9458 0.004
R9824 S.n9776 S.n9775 0.004
R9825 S.n10135 S.n10134 0.004
R9826 S.n10436 S.n10435 0.004
R9827 S.n10788 S.n10787 0.004
R9828 S.n11061 S.n11060 0.004
R9829 S.n11409 S.n11408 0.004
R9830 S.n11715 S.n11714 0.004
R9831 S.n794 S.n793 0.004
R9832 S.n1691 S.n1690 0.004
R9833 S.n668 S.n667 0.004
R9834 S.n651 S.n650 0.004
R9835 S.n383 S.n382 0.004
R9836 S.n1604 S.n1603 0.004
R9837 S.n7748 S.n7747 0.004
R9838 S.n7227 S.n7226 0.004
R9839 S.n6786 S.n6785 0.004
R9840 S.n6481 S.n6480 0.004
R9841 S.n6044 S.n6043 0.004
R9842 S.n5726 S.n5725 0.004
R9843 S.n5279 S.n5278 0.004
R9844 S.n4945 S.n4944 0.004
R9845 S.n4502 S.n4501 0.004
R9846 S.n4155 S.n4154 0.004
R9847 S.n3702 S.n3701 0.004
R9848 S.n3308 S.n3307 0.004
R9849 S.n2890 S.n2889 0.004
R9850 S.n2452 S.n2451 0.004
R9851 S.n2045 S.n2044 0.004
R9852 S.n1173 S.n1172 0.004
R9853 S.n403 S.n402 0.004
R9854 S.n8465 S.n8464 0.004
R9855 S.n7803 S.n7802 0.004
R9856 S.n7546 S.n7545 0.004
R9857 S.n7250 S.n7249 0.004
R9858 S.n6816 S.n6815 0.004
R9859 S.n6504 S.n6503 0.004
R9860 S.n6074 S.n6073 0.004
R9861 S.n5749 S.n5748 0.004
R9862 S.n5309 S.n5308 0.004
R9863 S.n4968 S.n4967 0.004
R9864 S.n4532 S.n4531 0.004
R9865 S.n4178 S.n4177 0.004
R9866 S.n3732 S.n3731 0.004
R9867 S.n3331 S.n3330 0.004
R9868 S.n2920 S.n2919 0.004
R9869 S.n2475 S.n2474 0.004
R9870 S.n2077 S.n2076 0.004
R9871 S.n1194 S.n1193 0.004
R9872 S.n1632 S.n1631 0.004
R9873 S.n635 S.n634 0.004
R9874 S.n618 S.n617 0.004
R9875 S.n342 S.n341 0.004
R9876 S.n1545 S.n1544 0.004
R9877 S.n6276 S.n6275 0.004
R9878 S.n5690 S.n5689 0.004
R9879 S.n5218 S.n5217 0.004
R9880 S.n4909 S.n4908 0.004
R9881 S.n4441 S.n4440 0.004
R9882 S.n4119 S.n4118 0.004
R9883 S.n3641 S.n3640 0.004
R9884 S.n3272 S.n3271 0.004
R9885 S.n2829 S.n2828 0.004
R9886 S.n2416 S.n2415 0.004
R9887 S.n1982 S.n1981 0.004
R9888 S.n1139 S.n1138 0.004
R9889 S.n362 S.n361 0.004
R9890 S.n7028 S.n7027 0.004
R9891 S.n6468 S.n6467 0.004
R9892 S.n6013 S.n6012 0.004
R9893 S.n5713 S.n5712 0.004
R9894 S.n5248 S.n5247 0.004
R9895 S.n4932 S.n4931 0.004
R9896 S.n4471 S.n4470 0.004
R9897 S.n4142 S.n4141 0.004
R9898 S.n3671 S.n3670 0.004
R9899 S.n3295 S.n3294 0.004
R9900 S.n2859 S.n2858 0.004
R9901 S.n2439 S.n2438 0.004
R9902 S.n2014 S.n2013 0.004
R9903 S.n1160 S.n1159 0.004
R9904 S.n1573 S.n1572 0.004
R9905 S.n602 S.n601 0.004
R9906 S.n585 S.n584 0.004
R9907 S.n321 S.n320 0.004
R9908 S.n1486 S.n1485 0.004
R9909 S.n4734 S.n4733 0.004
R9910 S.n4083 S.n4082 0.004
R9911 S.n3580 S.n3579 0.004
R9912 S.n3236 S.n3235 0.004
R9913 S.n2768 S.n2767 0.004
R9914 S.n2380 S.n2379 0.004
R9915 S.n1919 S.n1918 0.004
R9916 S.n1105 S.n1104 0.004
R9917 S.n57 S.n56 0.004
R9918 S.n5521 S.n5520 0.004
R9919 S.n4896 S.n4895 0.004
R9920 S.n4410 S.n4409 0.004
R9921 S.n4106 S.n4105 0.004
R9922 S.n3610 S.n3609 0.004
R9923 S.n3259 S.n3258 0.004
R9924 S.n2798 S.n2797 0.004
R9925 S.n2403 S.n2402 0.004
R9926 S.n1951 S.n1950 0.004
R9927 S.n1126 S.n1125 0.004
R9928 S.n1514 S.n1513 0.004
R9929 S.n569 S.n568 0.004
R9930 S.n552 S.n551 0.004
R9931 S.n280 S.n279 0.004
R9932 S.n1427 S.n1426 0.004
R9933 S.n3122 S.n3121 0.004
R9934 S.n2344 S.n2343 0.004
R9935 S.n1856 S.n1855 0.004
R9936 S.n1071 S.n1070 0.004
R9937 S.n300 S.n299 0.004
R9938 S.n3944 S.n3943 0.004
R9939 S.n3223 S.n3222 0.004
R9940 S.n2737 S.n2736 0.004
R9941 S.n2367 S.n2366 0.004
R9942 S.n1888 S.n1887 0.004
R9943 S.n1092 S.n1091 0.004
R9944 S.n1458 S.n1457 0.004
R9945 S.n536 S.n535 0.004
R9946 S.n519 S.n518 0.004
R9947 S.n239 S.n238 0.004
R9948 S.n1366 S.n1365 0.004
R9949 S.n259 S.n258 0.004
R9950 S.n2297 S.n2296 0.004
R9951 S.n1058 S.n1057 0.004
R9952 S.n1396 S.n1395 0.004
R9953 S.n503 S.n502 0.004
R9954 S.n486 S.n485 0.004
R9955 S.n875 S.n874 0.004
R9956 S.n744 S.n743 0.004
R9957 S.n1353 S.n1352 0.004
R9958 S.n1342 S.n1341 0.004
R9959 S.n2640 S.n2639 0.004
R9960 S.n2628 S.n2627 0.004
R9961 S.n3167 S.n3166 0.004
R9962 S.n3155 S.n3154 0.004
R9963 S.n3984 S.n3983 0.004
R9964 S.n3972 S.n3971 0.004
R9965 S.n4779 S.n4778 0.004
R9966 S.n4767 S.n4766 0.004
R9967 S.n5561 S.n5560 0.004
R9968 S.n5549 S.n5548 0.004
R9969 S.n6321 S.n6320 0.004
R9970 S.n6309 S.n6308 0.004
R9971 S.n7068 S.n7067 0.004
R9972 S.n7056 S.n7055 0.004
R9973 S.n8079 S.n8078 0.004
R9974 S.n8067 S.n8066 0.004
R9975 S.n8791 S.n8790 0.004
R9976 S.n8779 S.n8778 0.004
R9977 S.n9195 S.n9194 0.004
R9978 S.n9183 S.n9182 0.004
R9979 S.n9872 S.n9871 0.004
R9980 S.n9860 S.n9859 0.004
R9981 S.n10530 S.n10529 0.004
R9982 S.n10518 S.n10517 0.004
R9983 S.n11153 S.n11152 0.004
R9984 S.n11141 S.n11140 0.004
R9985 S.n11731 S.n11730 0.004
R9986 S.n12023 S.n12022 0.004
R9987 S.n12900 S.n12899 0.004
R9988 S.n12887 S.n12886 0.004
R9989 S.n1803 S.n1802 0.004
R9990 S.n1325 S.n1324 0.004
R9991 S.n2657 S.n2656 0.004
R9992 S.n12925 S.n12924 0.004
R9993 S.n12917 S.n12916 0.004
R9994 S.n12038 S.n12037 0.004
R9995 S.n11748 S.n11747 0.004
R9996 S.n11178 S.n11177 0.004
R9997 S.n11170 S.n11169 0.004
R9998 S.n10555 S.n10554 0.004
R9999 S.n10547 S.n10546 0.004
R10000 S.n9897 S.n9896 0.004
R10001 S.n9889 S.n9888 0.004
R10002 S.n9220 S.n9219 0.004
R10003 S.n9212 S.n9211 0.004
R10004 S.n8816 S.n8815 0.004
R10005 S.n8808 S.n8807 0.004
R10006 S.n8104 S.n8103 0.004
R10007 S.n8096 S.n8095 0.004
R10008 S.n7093 S.n7092 0.004
R10009 S.n7085 S.n7084 0.004
R10010 S.n6346 S.n6345 0.004
R10011 S.n6338 S.n6337 0.004
R10012 S.n5586 S.n5585 0.004
R10013 S.n5578 S.n5577 0.004
R10014 S.n4804 S.n4803 0.004
R10015 S.n4796 S.n4795 0.004
R10016 S.n4012 S.n4011 0.004
R10017 S.n4004 S.n4003 0.004
R10018 S.n3192 S.n3191 0.004
R10019 S.n3184 S.n3183 0.004
R10020 S.n2665 S.n2664 0.004
R10021 S.n1842 S.n1841 0.004
R10022 S.n2607 S.n2606 0.004
R10023 S.n3513 S.n3512 0.004
R10024 S.n12675 S.n12674 0.004
R10025 S.n12948 S.n12947 0.004
R10026 S.n12053 S.n12052 0.004
R10027 S.n11764 S.n11763 0.004
R10028 S.n11445 S.n11444 0.004
R10029 S.n11201 S.n11200 0.004
R10030 S.n10824 S.n10823 0.004
R10031 S.n10578 S.n10577 0.004
R10032 S.n10171 S.n10170 0.004
R10033 S.n9920 S.n9919 0.004
R10034 S.n9495 S.n9494 0.004
R10035 S.n9243 S.n9242 0.004
R10036 S.n8628 S.n8627 0.004
R10037 S.n8839 S.n8838 0.004
R10038 S.n7932 S.n7931 0.004
R10039 S.n8127 S.n8126 0.004
R10040 S.n7379 S.n7378 0.004
R10041 S.n7116 S.n7115 0.004
R10042 S.n6633 S.n6632 0.004
R10043 S.n6369 S.n6368 0.004
R10044 S.n5878 S.n5877 0.004
R10045 S.n5609 S.n5608 0.004
R10046 S.n5097 S.n5096 0.004
R10047 S.n4827 S.n4826 0.004
R10048 S.n4307 S.n4306 0.004
R10049 S.n4032 S.n4031 0.004
R10050 S.n3460 S.n3459 0.004
R10051 S.n2725 S.n2724 0.004
R10052 S.n3478 S.n3477 0.004
R10053 S.n4047 S.n4046 0.004
R10054 S.n12691 S.n12690 0.004
R10055 S.n12963 S.n12962 0.004
R10056 S.n12069 S.n12068 0.004
R10057 S.n11779 S.n11778 0.004
R10058 S.n11461 S.n11460 0.004
R10059 S.n11216 S.n11215 0.004
R10060 S.n10840 S.n10839 0.004
R10061 S.n10593 S.n10592 0.004
R10062 S.n10187 S.n10186 0.004
R10063 S.n9935 S.n9934 0.004
R10064 S.n9511 S.n9510 0.004
R10065 S.n9258 S.n9257 0.004
R10066 S.n8644 S.n8643 0.004
R10067 S.n8854 S.n8853 0.004
R10068 S.n7948 S.n7947 0.004
R10069 S.n8142 S.n8141 0.004
R10070 S.n7395 S.n7394 0.004
R10071 S.n7131 S.n7130 0.004
R10072 S.n6649 S.n6648 0.004
R10073 S.n6384 S.n6383 0.004
R10074 S.n5894 S.n5893 0.004
R10075 S.n5624 S.n5623 0.004
R10076 S.n5113 S.n5112 0.004
R10077 S.n4842 S.n4841 0.004
R10078 S.n4055 S.n4054 0.004
R10079 S.n3566 S.n3565 0.004
R10080 S.n4326 S.n4325 0.004
R10081 S.n4857 S.n4856 0.004
R10082 S.n12707 S.n12706 0.004
R10083 S.n12978 S.n12977 0.004
R10084 S.n12085 S.n12084 0.004
R10085 S.n11794 S.n11793 0.004
R10086 S.n11477 S.n11476 0.004
R10087 S.n11231 S.n11230 0.004
R10088 S.n10856 S.n10855 0.004
R10089 S.n10608 S.n10607 0.004
R10090 S.n10203 S.n10202 0.004
R10091 S.n9950 S.n9949 0.004
R10092 S.n9527 S.n9526 0.004
R10093 S.n9273 S.n9272 0.004
R10094 S.n8660 S.n8659 0.004
R10095 S.n8869 S.n8868 0.004
R10096 S.n7964 S.n7963 0.004
R10097 S.n8157 S.n8156 0.004
R10098 S.n7411 S.n7410 0.004
R10099 S.n7146 S.n7145 0.004
R10100 S.n6665 S.n6664 0.004
R10101 S.n6399 S.n6398 0.004
R10102 S.n5910 S.n5909 0.004
R10103 S.n5639 S.n5638 0.004
R10104 S.n4865 S.n4864 0.004
R10105 S.n4398 S.n4397 0.004
R10106 S.n5132 S.n5131 0.004
R10107 S.n5654 S.n5653 0.004
R10108 S.n12723 S.n12722 0.004
R10109 S.n12993 S.n12992 0.004
R10110 S.n12101 S.n12100 0.004
R10111 S.n11809 S.n11808 0.004
R10112 S.n11493 S.n11492 0.004
R10113 S.n11246 S.n11245 0.004
R10114 S.n10872 S.n10871 0.004
R10115 S.n10623 S.n10622 0.004
R10116 S.n10219 S.n10218 0.004
R10117 S.n9965 S.n9964 0.004
R10118 S.n9543 S.n9542 0.004
R10119 S.n9288 S.n9287 0.004
R10120 S.n8676 S.n8675 0.004
R10121 S.n8884 S.n8883 0.004
R10122 S.n7980 S.n7979 0.004
R10123 S.n8172 S.n8171 0.004
R10124 S.n7427 S.n7426 0.004
R10125 S.n7161 S.n7160 0.004
R10126 S.n6681 S.n6680 0.004
R10127 S.n6414 S.n6413 0.004
R10128 S.n5662 S.n5661 0.004
R10129 S.n5204 S.n5203 0.004
R10130 S.n5929 S.n5928 0.004
R10131 S.n6429 S.n6428 0.004
R10132 S.n12739 S.n12738 0.004
R10133 S.n13008 S.n13007 0.004
R10134 S.n12117 S.n12116 0.004
R10135 S.n11824 S.n11823 0.004
R10136 S.n11509 S.n11508 0.004
R10137 S.n11261 S.n11260 0.004
R10138 S.n10888 S.n10887 0.004
R10139 S.n10638 S.n10637 0.004
R10140 S.n10235 S.n10234 0.004
R10141 S.n9980 S.n9979 0.004
R10142 S.n9559 S.n9558 0.004
R10143 S.n9303 S.n9302 0.004
R10144 S.n8692 S.n8691 0.004
R10145 S.n8899 S.n8898 0.004
R10146 S.n7996 S.n7995 0.004
R10147 S.n8187 S.n8186 0.004
R10148 S.n7443 S.n7442 0.004
R10149 S.n7176 S.n7175 0.004
R10150 S.n6437 S.n6436 0.004
R10151 S.n6001 S.n6000 0.004
R10152 S.n6700 S.n6699 0.004
R10153 S.n7191 S.n7190 0.004
R10154 S.n12755 S.n12754 0.004
R10155 S.n13023 S.n13022 0.004
R10156 S.n12133 S.n12132 0.004
R10157 S.n11839 S.n11838 0.004
R10158 S.n11525 S.n11524 0.004
R10159 S.n11276 S.n11275 0.004
R10160 S.n10904 S.n10903 0.004
R10161 S.n10653 S.n10652 0.004
R10162 S.n10251 S.n10250 0.004
R10163 S.n9995 S.n9994 0.004
R10164 S.n9575 S.n9574 0.004
R10165 S.n9318 S.n9317 0.004
R10166 S.n8708 S.n8707 0.004
R10167 S.n8914 S.n8913 0.004
R10168 S.n8012 S.n8011 0.004
R10169 S.n8202 S.n8201 0.004
R10170 S.n7199 S.n7198 0.004
R10171 S.n6772 S.n6771 0.004
R10172 S.n7462 S.n7461 0.004
R10173 S.n8217 S.n8216 0.004
R10174 S.n12771 S.n12770 0.004
R10175 S.n13038 S.n13037 0.004
R10176 S.n12149 S.n12148 0.004
R10177 S.n11854 S.n11853 0.004
R10178 S.n11541 S.n11540 0.004
R10179 S.n11291 S.n11290 0.004
R10180 S.n10920 S.n10919 0.004
R10181 S.n10668 S.n10667 0.004
R10182 S.n10267 S.n10266 0.004
R10183 S.n10010 S.n10009 0.004
R10184 S.n9591 S.n9590 0.004
R10185 S.n9333 S.n9332 0.004
R10186 S.n8724 S.n8723 0.004
R10187 S.n8929 S.n8928 0.004
R10188 S.n8028 S.n8027 0.004
R10189 S.n7534 S.n7533 0.004
R10190 S.n8046 S.n8045 0.004
R10191 S.n8944 S.n8943 0.004
R10192 S.n12787 S.n12786 0.004
R10193 S.n13053 S.n13052 0.004
R10194 S.n12165 S.n12164 0.004
R10195 S.n11869 S.n11868 0.004
R10196 S.n11557 S.n11556 0.004
R10197 S.n11306 S.n11305 0.004
R10198 S.n10936 S.n10935 0.004
R10199 S.n10683 S.n10682 0.004
R10200 S.n10283 S.n10282 0.004
R10201 S.n10025 S.n10024 0.004
R10202 S.n9607 S.n9606 0.004
R10203 S.n9348 S.n9347 0.004
R10204 S.n8740 S.n8739 0.004
R10205 S.n8270 S.n8269 0.004
R10206 S.n8758 S.n8757 0.004
R10207 S.n9363 S.n9362 0.004
R10208 S.n12803 S.n12802 0.004
R10209 S.n13068 S.n13067 0.004
R10210 S.n12181 S.n12180 0.004
R10211 S.n11884 S.n11883 0.004
R10212 S.n11573 S.n11572 0.004
R10213 S.n11321 S.n11320 0.004
R10214 S.n10952 S.n10951 0.004
R10215 S.n10698 S.n10697 0.004
R10216 S.n10299 S.n10298 0.004
R10217 S.n10040 S.n10039 0.004
R10218 S.n9371 S.n9370 0.004
R10219 S.n8997 S.n8996 0.004
R10220 S.n9626 S.n9625 0.004
R10221 S.n10055 S.n10054 0.004
R10222 S.n12819 S.n12818 0.004
R10223 S.n13083 S.n13082 0.004
R10224 S.n12197 S.n12196 0.004
R10225 S.n11899 S.n11898 0.004
R10226 S.n11589 S.n11588 0.004
R10227 S.n11336 S.n11335 0.004
R10228 S.n10968 S.n10967 0.004
R10229 S.n10713 S.n10712 0.004
R10230 S.n10063 S.n10062 0.004
R10231 S.n9698 S.n9697 0.004
R10232 S.n10318 S.n10317 0.004
R10233 S.n10728 S.n10727 0.004
R10234 S.n12835 S.n12834 0.004
R10235 S.n13098 S.n13097 0.004
R10236 S.n12213 S.n12212 0.004
R10237 S.n11914 S.n11913 0.004
R10238 S.n11605 S.n11604 0.004
R10239 S.n11351 S.n11350 0.004
R10240 S.n10736 S.n10735 0.004
R10241 S.n10390 S.n10389 0.004
R10242 S.n10987 S.n10986 0.004
R10243 S.n11366 S.n11365 0.004
R10244 S.n12851 S.n12850 0.004
R10245 S.n13113 S.n13112 0.004
R10246 S.n12229 S.n12228 0.004
R10247 S.n11929 S.n11928 0.004
R10248 S.n11374 S.n11373 0.004
R10249 S.n11049 S.n11048 0.004
R10250 S.n11622 S.n11621 0.004
R10251 S.n12262 S.n12261 0.004
R10252 S.n12870 S.n12869 0.004
R10253 S.n13133 S.n13132 0.004
R10254 S.n12249 S.n12248 0.004
R10255 S.n12661 S.n12660 0.004
R10256 S.n13148 S.n13147 0.004
R10257 S.t28 S.n218 0.004
R10258 S.n823 S.n822 0.004
R10259 S.n446 S.n445 0.004
R10260 S.n426 S.n425 0.004
R10261 S.n405 S.n404 0.004
R10262 S.n385 S.n384 0.004
R10263 S.n364 S.n363 0.004
R10264 S.n344 S.n343 0.004
R10265 S.n59 S.n58 0.004
R10266 S.n323 S.n322 0.004
R10267 S.n302 S.n301 0.004
R10268 S.n282 S.n281 0.004
R10269 S.n261 S.n260 0.004
R10270 S.n241 S.n240 0.004
R10271 S.t28 S.n925 0.004
R10272 S.n473 S.n458 0.004
R10273 S.n10753 S.n10752 0.004
R10274 S.n10409 S.n10408 0.004
R10275 S.n9749 S.n9748 0.004
R10276 S.n9077 S.n9076 0.004
R10277 S.n8382 S.n8381 0.004
R10278 S.n7675 S.n7674 0.004
R10279 S.n6945 S.n6944 0.004
R10280 S.n6203 S.n6202 0.004
R10281 S.n5438 S.n5437 0.004
R10282 S.n4661 S.n4660 0.004
R10283 S.n3861 S.n3860 0.004
R10284 S.n3049 S.n3048 0.004
R10285 S.n2211 S.n2210 0.004
R10286 S.n1710 S.n1709 0.004
R10287 S.n908 S.n907 0.004
R10288 S.n12618 S.n12617 0.004
R10289 S.n10753 S.n10751 0.004
R10290 S.n709 S.n697 0.004
R10291 S.n1293 S.n1292 0.004
R10292 S.n2573 S.n2561 0.004
R10293 S.n3429 S.n3417 0.004
R10294 S.n4276 S.n4264 0.004
R10295 S.n5066 S.n5054 0.004
R10296 S.n5847 S.n5835 0.004
R10297 S.n6602 S.n6590 0.004
R10298 S.n7348 S.n7336 0.004
R10299 S.n7901 S.n7889 0.004
R10300 S.n8597 S.n8585 0.004
R10301 S.n9464 S.n9452 0.004
R10302 S.n10140 S.n10128 0.004
R10303 S.n10793 S.n10781 0.004
R10304 S.n11414 S.n11402 0.004
R10305 S.n11967 S.n11965 0.004
R10306 S.n10081 S.n10080 0.004
R10307 S.n670 S.n661 0.004
R10308 S.n9388 S.n9386 0.004
R10309 S.n8502 S.n8501 0.004
R10310 S.n637 S.n628 0.004
R10311 S.n7789 S.n7787 0.004
R10312 S.n7217 S.n7216 0.004
R10313 S.n604 S.n595 0.004
R10314 S.n6454 S.n6452 0.004
R10315 S.n5680 S.n5679 0.004
R10316 S.n571 S.n562 0.004
R10317 S.n4882 S.n4880 0.004
R10318 S.n4073 S.n4072 0.004
R10319 S.n538 S.n529 0.004
R10320 S.n3209 S.n3207 0.004
R10321 S.n2334 S.n2333 0.004
R10322 S.n505 S.n496 0.004
R10323 S.n1044 S.n1042 0.004
R10324 S.n473 S.n472 0.004
R10325 S.n1000 S.n999 0.004
R10326 S.n9705 S.n9704 0.004
R10327 S.n9033 S.n9032 0.004
R10328 S.n8338 S.n8337 0.004
R10329 S.n7631 S.n7630 0.004
R10330 S.n6901 S.n6900 0.004
R10331 S.n6159 S.n6158 0.004
R10332 S.n5394 S.n5393 0.004
R10333 S.n4617 S.n4616 0.004
R10334 S.n3817 S.n3816 0.004
R10335 S.n3005 S.n3004 0.004
R10336 S.n2165 S.n2164 0.004
R10337 S.n11395 S.n11378 0.004
R10338 S.n10417 S.n10415 0.004
R10339 S.n9757 S.n9755 0.004
R10340 S.n9085 S.n9083 0.004
R10341 S.n8390 S.n8388 0.004
R10342 S.n7683 S.n7681 0.004
R10343 S.n6953 S.n6951 0.004
R10344 S.n6211 S.n6209 0.004
R10345 S.n5446 S.n5444 0.004
R10346 S.n4669 S.n4667 0.004
R10347 S.n3869 S.n3867 0.004
R10348 S.n3057 S.n3055 0.004
R10349 S.n2219 S.n2217 0.004
R10350 S.n1718 S.n1716 0.004
R10351 S.n1252 S.n1251 0.004
R10352 S.n9841 S.n9840 0.004
R10353 S.n10081 S.n10065 0.004
R10354 S.n8474 S.n8473 0.004
R10355 S.n8502 S.n8486 0.004
R10356 S.n7037 S.n7036 0.004
R10357 S.n7217 S.n7201 0.004
R10358 S.n5530 S.n5529 0.004
R10359 S.n5680 S.n5664 0.004
R10360 S.n3953 S.n3952 0.004
R10361 S.n4073 S.n4057 0.004
R10362 S.n2306 S.n2305 0.004
R10363 S.n2334 S.n2318 0.004
R10364 S.n1828 S.n1814 0.004
R10365 S.n2692 S.n1828 0.004
R10366 S.n2711 S.n2697 0.004
R10367 S.n3533 S.n2711 0.004
R10368 S.n3552 S.n3538 0.004
R10369 S.n4365 S.n3552 0.004
R10370 S.n4384 S.n4370 0.004
R10371 S.n5171 S.n4384 0.004
R10372 S.n5190 S.n5176 0.004
R10373 S.n5968 S.n5190 0.004
R10374 S.n5987 S.n5973 0.004
R10375 S.n6739 S.n5987 0.004
R10376 S.n6758 S.n6744 0.004
R10377 S.n7501 S.n6758 0.004
R10378 S.n7520 S.n7506 0.004
R10379 S.n8237 S.n7520 0.004
R10380 S.n8256 S.n8242 0.004
R10381 S.n8964 S.n8256 0.004
R10382 S.n8983 S.n8969 0.004
R10383 S.n9665 S.n8983 0.004
R10384 S.n9684 S.n9670 0.004
R10385 S.n10357 S.n9684 0.004
R10386 S.n10376 S.n10362 0.004
R10387 S.n11026 S.n10376 0.004
R10388 S.n11944 S.n11942 0.004
R10389 S.n11035 S.n11034 0.004
R10390 S.n11666 S.n11030 0.004
R10391 S.t35 S.n12381 0.004
R10392 S.t35 S.n12378 0.004
R10393 S.t35 S.n12374 0.004
R10394 S.t35 S.n12370 0.004
R10395 S.t35 S.n12366 0.004
R10396 S.t35 S.n12362 0.004
R10397 S.t35 S.n12358 0.004
R10398 S.t35 S.n12354 0.004
R10399 S.t35 S.n12350 0.004
R10400 S.t35 S.n12346 0.004
R10401 S.t35 S.n12342 0.004
R10402 S.t35 S.n12338 0.004
R10403 S.t35 S.n12334 0.004
R10404 S.t35 S.n12331 0.004
R10405 S.t430 S.n476 0.004
R10406 S.t28 S.n951 0.004
R10407 S.t28 S.n948 0.004
R10408 S.t14 S.n12621 0.004
R10409 S.t28 S.n201 0.004
R10410 S.t26 S.n9391 0.004
R10411 S.t28 S.n975 0.004
R10412 S.t16 S.n10084 0.004
R10413 S.t28 S.n216 0.004
R10414 S.t122 S.n10756 0.004
R10415 S.t28 S.n922 0.004
R10416 S.t18 S.n11398 0.004
R10417 S.t2 S.n11970 0.004
R10418 S.t28 S.n939 0.004
R10419 S.t28 S.n189 0.004
R10420 S.t22 S.n7792 0.004
R10421 S.t28 S.n971 0.004
R10422 S.t0 S.n8505 0.004
R10423 S.t28 S.n177 0.004
R10424 S.t8 S.n6457 0.004
R10425 S.t28 S.n967 0.004
R10426 S.t40 S.n7220 0.004
R10427 S.t28 S.n164 0.004
R10428 S.t81 S.n4885 0.004
R10429 S.t28 S.n963 0.004
R10430 S.t460 S.n5683 0.004
R10431 S.t28 S.n151 0.004
R10432 S.t444 S.n3212 0.004
R10433 S.t28 S.n959 0.004
R10434 S.t51 S.n4076 0.004
R10435 S.t28 S.n138 0.004
R10436 S.t142 S.n1047 0.004
R10437 S.t28 S.n955 0.004
R10438 S.t55 S.n2337 0.004
R10439 S.t28 S.n125 0.004
R10440 S.t35 S.n12542 0.004
R10441 S.t35 S.n12544 0.004
R10442 S.t35 S.n12482 0.004
R10443 S.t35 S.n12486 0.004
R10444 S.t35 S.n12490 0.004
R10445 S.t35 S.n12494 0.004
R10446 S.t35 S.n12498 0.004
R10447 S.t35 S.n12502 0.004
R10448 S.t35 S.n12506 0.004
R10449 S.t35 S.n12510 0.004
R10450 S.t35 S.n12514 0.004
R10451 S.t35 S.n12518 0.004
R10452 S.t35 S.n12522 0.004
R10453 S.t35 S.n12526 0.004
R10454 S.t35 S.n12530 0.004
R10455 S.t35 S.n12534 0.004
R10456 S.t35 S.n12538 0.004
R10457 S.t35 S.n12478 0.004
R10458 S.t28 S.n946 0.004
R10459 S.t35 S.n12391 0.004
R10460 S.t28 S.n10 0.004
R10461 S.t28 S.n21 0.004
R10462 S.t28 S.n33 0.004
R10463 S.t28 S.n65 0.004
R10464 S.t28 S.n77 0.004
R10465 S.t28 S.n89 0.004
R10466 S.t28 S.n93 0.004
R10467 S.n765 S.n764 0.004
R10468 S.t28 S.n943 0.004
R10469 S.t28 S.n193 0.004
R10470 S.t28 S.n181 0.004
R10471 S.t28 S.n168 0.004
R10472 S.t28 S.n155 0.004
R10473 S.t28 S.n142 0.004
R10474 S.t28 S.n129 0.004
R10475 S.n11967 S.n11966 0.004
R10476 S.n10099 S.n10088 0.004
R10477 S.n9423 S.n9412 0.004
R10478 S.n8556 S.n8545 0.004
R10479 S.n7860 S.n7849 0.004
R10480 S.n7307 S.n7296 0.004
R10481 S.n6561 S.n6550 0.004
R10482 S.n5806 S.n5795 0.004
R10483 S.n5025 S.n5014 0.004
R10484 S.n4235 S.n4224 0.004
R10485 S.n3388 S.n3377 0.004
R10486 S.n2532 S.n2521 0.004
R10487 S.n12646 S.n12645 0.003
R10488 S.n12570 S.n12569 0.003
R10489 S.n12015 S.n12014 0.003
R10490 S.n12274 S.n12273 0.003
R10491 S.n854 S.n853 0.003
R10492 S.n829 S.n828 0.003
R10493 S.n1791 S.n1790 0.003
R10494 S.n12594 S.n12593 0.003
R10495 S.n11991 S.n11990 0.003
R10496 S.n11698 S.n11697 0.003
R10497 S.n11439 S.n11438 0.003
R10498 S.n11101 S.n11100 0.003
R10499 S.n10818 S.n10817 0.003
R10500 S.n10476 S.n10475 0.003
R10501 S.n10165 S.n10164 0.003
R10502 S.n9816 S.n9815 0.003
R10503 S.n9489 S.n9488 0.003
R10504 S.n9144 S.n9143 0.003
R10505 S.n8622 S.n8621 0.003
R10506 S.n8449 S.n8448 0.003
R10507 S.n7926 S.n7925 0.003
R10508 S.n7742 S.n7741 0.003
R10509 S.n7373 S.n7372 0.003
R10510 S.n7012 S.n7011 0.003
R10511 S.n6627 S.n6626 0.003
R10512 S.n6270 S.n6269 0.003
R10513 S.n5872 S.n5871 0.003
R10514 S.n5505 S.n5504 0.003
R10515 S.n5091 S.n5090 0.003
R10516 S.n4728 S.n4727 0.003
R10517 S.n4301 S.n4300 0.003
R10518 S.n3928 S.n3927 0.003
R10519 S.n3454 S.n3453 0.003
R10520 S.n3116 S.n3115 0.003
R10521 S.n2598 S.n2597 0.003
R10522 S.n2281 S.n2280 0.003
R10523 S.n1316 S.n1315 0.003
R10524 S.n735 S.n734 0.003
R10525 S.n432 S.n431 0.003
R10526 S.n1679 S.n1678 0.003
R10527 S.n9167 S.n9166 0.003
R10528 S.n8526 S.n8525 0.003
R10529 S.n8302 S.n8301 0.003
R10530 S.n7830 S.n7829 0.003
R10531 S.n7595 S.n7594 0.003
R10532 S.n7277 S.n7276 0.003
R10533 S.n6865 S.n6864 0.003
R10534 S.n6531 S.n6530 0.003
R10535 S.n6123 S.n6122 0.003
R10536 S.n5776 S.n5775 0.003
R10537 S.n5358 S.n5357 0.003
R10538 S.n4995 S.n4994 0.003
R10539 S.n4581 S.n4580 0.003
R10540 S.n4205 S.n4204 0.003
R10541 S.n3781 S.n3780 0.003
R10542 S.n3358 S.n3357 0.003
R10543 S.n2969 S.n2968 0.003
R10544 S.n2502 S.n2501 0.003
R10545 S.n2128 S.n2127 0.003
R10546 S.n1219 S.n1218 0.003
R10547 S.n452 S.n451 0.003
R10548 S.n9844 S.n9843 0.003
R10549 S.n9410 S.n9409 0.003
R10550 S.n9026 S.n9025 0.003
R10551 S.n8543 S.n8542 0.003
R10552 S.n8331 S.n8330 0.003
R10553 S.n7847 S.n7846 0.003
R10554 S.n7624 S.n7623 0.003
R10555 S.n7294 S.n7293 0.003
R10556 S.n6894 S.n6893 0.003
R10557 S.n6548 S.n6547 0.003
R10558 S.n6152 S.n6151 0.003
R10559 S.n5793 S.n5792 0.003
R10560 S.n5387 S.n5386 0.003
R10561 S.n5012 S.n5011 0.003
R10562 S.n4610 S.n4609 0.003
R10563 S.n4222 S.n4221 0.003
R10564 S.n3810 S.n3809 0.003
R10565 S.n3375 S.n3374 0.003
R10566 S.n2998 S.n2997 0.003
R10567 S.n2519 S.n2518 0.003
R10568 S.n2157 S.n2156 0.003
R10569 S.n1238 S.n1237 0.003
R10570 S.n1258 S.n1257 0.003
R10571 S.n757 S.n756 0.003
R10572 S.n786 S.n785 0.003
R10573 S.n2192 S.n2191 0.003
R10574 S.n3030 S.n3029 0.003
R10575 S.n3842 S.n3841 0.003
R10576 S.n4642 S.n4641 0.003
R10577 S.n5419 S.n5418 0.003
R10578 S.n6184 S.n6183 0.003
R10579 S.n6926 S.n6925 0.003
R10580 S.n7656 S.n7655 0.003
R10581 S.n8363 S.n8362 0.003
R10582 S.n9058 S.n9057 0.003
R10583 S.n9730 S.n9729 0.003
R10584 S.n10502 S.n10501 0.003
R10585 S.n10105 S.n10104 0.003
R10586 S.n9429 S.n9428 0.003
R10587 S.n8562 S.n8561 0.003
R10588 S.n7866 S.n7865 0.003
R10589 S.n7313 S.n7312 0.003
R10590 S.n6567 S.n6566 0.003
R10591 S.n5812 S.n5811 0.003
R10592 S.n5031 S.n5030 0.003
R10593 S.n4241 S.n4240 0.003
R10594 S.n3394 S.n3393 0.003
R10595 S.n2538 S.n2537 0.003
R10596 S.n1741 S.n1740 0.003
R10597 S.n696 S.n695 0.003
R10598 S.n888 S.n887 0.003
R10599 S.n11125 S.n11124 0.003
R10600 S.n10779 S.n10778 0.003
R10601 S.n10424 S.n10423 0.003
R10602 S.n10126 S.n10125 0.003
R10603 S.n9764 S.n9763 0.003
R10604 S.n9450 S.n9449 0.003
R10605 S.n9092 S.n9091 0.003
R10606 S.n8583 S.n8582 0.003
R10607 S.n8397 S.n8396 0.003
R10608 S.n7887 S.n7886 0.003
R10609 S.n7690 S.n7689 0.003
R10610 S.n7334 S.n7333 0.003
R10611 S.n6960 S.n6959 0.003
R10612 S.n6588 S.n6587 0.003
R10613 S.n6218 S.n6217 0.003
R10614 S.n5833 S.n5832 0.003
R10615 S.n5453 S.n5452 0.003
R10616 S.n5052 S.n5051 0.003
R10617 S.n4676 S.n4675 0.003
R10618 S.n4262 S.n4261 0.003
R10619 S.n3876 S.n3875 0.003
R10620 S.n3415 S.n3414 0.003
R10621 S.n3064 S.n3063 0.003
R10622 S.n2559 S.n2558 0.003
R10623 S.n2226 S.n2225 0.003
R10624 S.n1279 S.n1278 0.003
R10625 S.n1769 S.n1768 0.003
R10626 S.n715 S.n714 0.003
R10627 S.n1299 S.n1298 0.003
R10628 S.n2247 S.n2246 0.003
R10629 S.n2579 S.n2578 0.003
R10630 S.n3084 S.n3083 0.003
R10631 S.n3435 S.n3434 0.003
R10632 S.n3896 S.n3895 0.003
R10633 S.n4282 S.n4281 0.003
R10634 S.n4696 S.n4695 0.003
R10635 S.n5072 S.n5071 0.003
R10636 S.n5473 S.n5472 0.003
R10637 S.n5853 S.n5852 0.003
R10638 S.n6238 S.n6237 0.003
R10639 S.n6608 S.n6607 0.003
R10640 S.n6980 S.n6979 0.003
R10641 S.n7354 S.n7353 0.003
R10642 S.n7710 S.n7709 0.003
R10643 S.n7907 S.n7906 0.003
R10644 S.n8417 S.n8416 0.003
R10645 S.n8603 S.n8602 0.003
R10646 S.n9112 S.n9111 0.003
R10647 S.n9470 S.n9469 0.003
R10648 S.n9784 S.n9783 0.003
R10649 S.n10146 S.n10145 0.003
R10650 S.n10444 S.n10443 0.003
R10651 S.n10799 S.n10798 0.003
R10652 S.n11069 S.n11068 0.003
R10653 S.n11420 S.n11419 0.003
R10654 S.n11720 S.n11719 0.003
R10655 S.n808 S.n807 0.003
R10656 S.n1707 S.n1706 0.003
R10657 S.n676 S.n675 0.003
R10658 S.n659 S.n658 0.003
R10659 S.n391 S.n390 0.003
R10660 S.n1620 S.n1619 0.003
R10661 S.n7765 S.n7764 0.003
R10662 S.n7241 S.n7240 0.003
R10663 S.n6804 S.n6803 0.003
R10664 S.n6495 S.n6494 0.003
R10665 S.n6062 S.n6061 0.003
R10666 S.n5740 S.n5739 0.003
R10667 S.n5297 S.n5296 0.003
R10668 S.n4959 S.n4958 0.003
R10669 S.n4520 S.n4519 0.003
R10670 S.n4169 S.n4168 0.003
R10671 S.n3720 S.n3719 0.003
R10672 S.n3322 S.n3321 0.003
R10673 S.n2908 S.n2907 0.003
R10674 S.n2466 S.n2465 0.003
R10675 S.n2065 S.n2064 0.003
R10676 S.n1185 S.n1184 0.003
R10677 S.n411 S.n410 0.003
R10678 S.n8477 S.n8476 0.003
R10679 S.n7811 S.n7810 0.003
R10680 S.n7563 S.n7562 0.003
R10681 S.n7258 S.n7257 0.003
R10682 S.n6833 S.n6832 0.003
R10683 S.n6512 S.n6511 0.003
R10684 S.n6091 S.n6090 0.003
R10685 S.n5757 S.n5756 0.003
R10686 S.n5326 S.n5325 0.003
R10687 S.n4976 S.n4975 0.003
R10688 S.n4549 S.n4548 0.003
R10689 S.n4186 S.n4185 0.003
R10690 S.n3749 S.n3748 0.003
R10691 S.n3339 S.n3338 0.003
R10692 S.n2937 S.n2936 0.003
R10693 S.n2483 S.n2482 0.003
R10694 S.n2094 S.n2093 0.003
R10695 S.n1202 S.n1201 0.003
R10696 S.n1649 S.n1648 0.003
R10697 S.n643 S.n642 0.003
R10698 S.n626 S.n625 0.003
R10699 S.n350 S.n349 0.003
R10700 S.n1561 S.n1560 0.003
R10701 S.n6293 S.n6292 0.003
R10702 S.n5704 S.n5703 0.003
R10703 S.n5236 S.n5235 0.003
R10704 S.n4923 S.n4922 0.003
R10705 S.n4459 S.n4458 0.003
R10706 S.n4133 S.n4132 0.003
R10707 S.n3659 S.n3658 0.003
R10708 S.n3286 S.n3285 0.003
R10709 S.n2847 S.n2846 0.003
R10710 S.n2430 S.n2429 0.003
R10711 S.n2002 S.n2001 0.003
R10712 S.n1151 S.n1150 0.003
R10713 S.n370 S.n369 0.003
R10714 S.n7040 S.n7039 0.003
R10715 S.n6476 S.n6475 0.003
R10716 S.n6030 S.n6029 0.003
R10717 S.n5721 S.n5720 0.003
R10718 S.n5265 S.n5264 0.003
R10719 S.n4940 S.n4939 0.003
R10720 S.n4488 S.n4487 0.003
R10721 S.n4150 S.n4149 0.003
R10722 S.n3688 S.n3687 0.003
R10723 S.n3303 S.n3302 0.003
R10724 S.n2876 S.n2875 0.003
R10725 S.n2447 S.n2446 0.003
R10726 S.n2031 S.n2030 0.003
R10727 S.n1168 S.n1167 0.003
R10728 S.n1590 S.n1589 0.003
R10729 S.n610 S.n609 0.003
R10730 S.n593 S.n592 0.003
R10731 S.n329 S.n328 0.003
R10732 S.n1502 S.n1501 0.003
R10733 S.n4751 S.n4750 0.003
R10734 S.n4097 S.n4096 0.003
R10735 S.n3598 S.n3597 0.003
R10736 S.n3250 S.n3249 0.003
R10737 S.n2786 S.n2785 0.003
R10738 S.n2394 S.n2393 0.003
R10739 S.n1939 S.n1938 0.003
R10740 S.n1117 S.n1116 0.003
R10741 S.n51 S.n50 0.003
R10742 S.n5533 S.n5532 0.003
R10743 S.n4904 S.n4903 0.003
R10744 S.n4427 S.n4426 0.003
R10745 S.n4114 S.n4113 0.003
R10746 S.n3627 S.n3626 0.003
R10747 S.n3267 S.n3266 0.003
R10748 S.n2815 S.n2814 0.003
R10749 S.n2411 S.n2410 0.003
R10750 S.n1968 S.n1967 0.003
R10751 S.n1134 S.n1133 0.003
R10752 S.n1531 S.n1530 0.003
R10753 S.n577 S.n576 0.003
R10754 S.n560 S.n559 0.003
R10755 S.n288 S.n287 0.003
R10756 S.n1443 S.n1442 0.003
R10757 S.n3139 S.n3138 0.003
R10758 S.n2358 S.n2357 0.003
R10759 S.n1876 S.n1875 0.003
R10760 S.n1083 S.n1082 0.003
R10761 S.n308 S.n307 0.003
R10762 S.n3956 S.n3955 0.003
R10763 S.n3231 S.n3230 0.003
R10764 S.n2754 S.n2753 0.003
R10765 S.n2375 S.n2374 0.003
R10766 S.n1905 S.n1904 0.003
R10767 S.n1100 S.n1099 0.003
R10768 S.n1472 S.n1471 0.003
R10769 S.n544 S.n543 0.003
R10770 S.n527 S.n526 0.003
R10771 S.n247 S.n246 0.003
R10772 S.n1384 S.n1383 0.003
R10773 S.n267 S.n266 0.003
R10774 S.n2309 S.n2308 0.003
R10775 S.n1066 S.n1065 0.003
R10776 S.n1413 S.n1412 0.003
R10777 S.n511 S.n510 0.003
R10778 S.n494 S.n493 0.003
R10779 S.n883 S.n882 0.003
R10780 S.n751 S.n750 0.003
R10781 S.n1361 S.n1360 0.003
R10782 S.n1336 S.n1335 0.003
R10783 S.n2649 S.n2648 0.003
R10784 S.n2622 S.n2621 0.003
R10785 S.n3176 S.n3175 0.003
R10786 S.n3149 S.n3148 0.003
R10787 S.n3993 S.n3992 0.003
R10788 S.n3966 S.n3965 0.003
R10789 S.n4788 S.n4787 0.003
R10790 S.n4761 S.n4760 0.003
R10791 S.n5570 S.n5569 0.003
R10792 S.n5543 S.n5542 0.003
R10793 S.n6330 S.n6329 0.003
R10794 S.n6303 S.n6302 0.003
R10795 S.n7077 S.n7076 0.003
R10796 S.n7050 S.n7049 0.003
R10797 S.n8088 S.n8087 0.003
R10798 S.n8061 S.n8060 0.003
R10799 S.n8800 S.n8799 0.003
R10800 S.n8773 S.n8772 0.003
R10801 S.n9204 S.n9203 0.003
R10802 S.n9177 S.n9176 0.003
R10803 S.n9881 S.n9880 0.003
R10804 S.n9854 S.n9853 0.003
R10805 S.n10539 S.n10538 0.003
R10806 S.n10512 S.n10511 0.003
R10807 S.n11162 S.n11161 0.003
R10808 S.n11135 S.n11134 0.003
R10809 S.n11740 S.n11739 0.003
R10810 S.n12030 S.n12029 0.003
R10811 S.n12909 S.n12908 0.003
R10812 S.n12881 S.n12880 0.003
R10813 S.n1799 S.n1798 0.003
R10814 S.n1330 S.n1329 0.003
R10815 S.n2679 S.n2678 0.003
R10816 S.n12931 S.n12930 0.003
R10817 S.n12940 S.n12939 0.003
R10818 S.n12045 S.n12044 0.003
R10819 S.n11756 S.n11755 0.003
R10820 S.n11184 S.n11183 0.003
R10821 S.n11193 S.n11192 0.003
R10822 S.n10561 S.n10560 0.003
R10823 S.n10570 S.n10569 0.003
R10824 S.n9903 S.n9902 0.003
R10825 S.n9912 S.n9911 0.003
R10826 S.n9226 S.n9225 0.003
R10827 S.n9235 S.n9234 0.003
R10828 S.n8822 S.n8821 0.003
R10829 S.n8831 S.n8830 0.003
R10830 S.n8110 S.n8109 0.003
R10831 S.n8119 S.n8118 0.003
R10832 S.n7099 S.n7098 0.003
R10833 S.n7108 S.n7107 0.003
R10834 S.n6352 S.n6351 0.003
R10835 S.n6361 S.n6360 0.003
R10836 S.n5592 S.n5591 0.003
R10837 S.n5601 S.n5600 0.003
R10838 S.n4810 S.n4809 0.003
R10839 S.n4819 S.n4818 0.003
R10840 S.n4018 S.n4017 0.003
R10841 S.n3999 S.n3998 0.003
R10842 S.n3496 S.n3495 0.003
R10843 S.n3505 S.n3504 0.003
R10844 S.n2671 S.n2670 0.003
R10845 S.n2687 S.n2686 0.003
R10846 S.n2616 S.n2615 0.003
R10847 S.n3520 S.n3519 0.003
R10848 S.n12683 S.n12682 0.003
R10849 S.n12955 S.n12954 0.003
R10850 S.n12061 S.n12060 0.003
R10851 S.n11771 S.n11770 0.003
R10852 S.n11453 S.n11452 0.003
R10853 S.n11208 S.n11207 0.003
R10854 S.n10832 S.n10831 0.003
R10855 S.n10585 S.n10584 0.003
R10856 S.n10179 S.n10178 0.003
R10857 S.n9927 S.n9926 0.003
R10858 S.n9503 S.n9502 0.003
R10859 S.n9250 S.n9249 0.003
R10860 S.n8636 S.n8635 0.003
R10861 S.n8846 S.n8845 0.003
R10862 S.n7940 S.n7939 0.003
R10863 S.n8134 S.n8133 0.003
R10864 S.n7387 S.n7386 0.003
R10865 S.n7123 S.n7122 0.003
R10866 S.n6641 S.n6640 0.003
R10867 S.n6376 S.n6375 0.003
R10868 S.n5886 S.n5885 0.003
R10869 S.n5616 S.n5615 0.003
R10870 S.n5105 S.n5104 0.003
R10871 S.n4834 S.n4833 0.003
R10872 S.n4315 S.n4314 0.003
R10873 S.n4039 S.n4038 0.003
R10874 S.n3467 S.n3466 0.003
R10875 S.n3528 S.n3527 0.003
R10876 S.n3487 S.n3486 0.003
R10877 S.n4352 S.n4351 0.003
R10878 S.n12699 S.n12698 0.003
R10879 S.n12970 S.n12969 0.003
R10880 S.n12077 S.n12076 0.003
R10881 S.n11786 S.n11785 0.003
R10882 S.n11469 S.n11468 0.003
R10883 S.n11223 S.n11222 0.003
R10884 S.n10848 S.n10847 0.003
R10885 S.n10600 S.n10599 0.003
R10886 S.n10195 S.n10194 0.003
R10887 S.n9942 S.n9941 0.003
R10888 S.n9519 S.n9518 0.003
R10889 S.n9265 S.n9264 0.003
R10890 S.n8652 S.n8651 0.003
R10891 S.n8861 S.n8860 0.003
R10892 S.n7956 S.n7955 0.003
R10893 S.n8149 S.n8148 0.003
R10894 S.n7403 S.n7402 0.003
R10895 S.n7138 S.n7137 0.003
R10896 S.n6657 S.n6656 0.003
R10897 S.n6391 S.n6390 0.003
R10898 S.n5902 S.n5901 0.003
R10899 S.n5631 S.n5630 0.003
R10900 S.n5121 S.n5120 0.003
R10901 S.n4849 S.n4848 0.003
R10902 S.n4344 S.n4343 0.003
R10903 S.n4360 S.n4359 0.003
R10904 S.n4335 S.n4334 0.003
R10905 S.n5158 S.n5157 0.003
R10906 S.n12715 S.n12714 0.003
R10907 S.n12985 S.n12984 0.003
R10908 S.n12093 S.n12092 0.003
R10909 S.n11801 S.n11800 0.003
R10910 S.n11485 S.n11484 0.003
R10911 S.n11238 S.n11237 0.003
R10912 S.n10864 S.n10863 0.003
R10913 S.n10615 S.n10614 0.003
R10914 S.n10211 S.n10210 0.003
R10915 S.n9957 S.n9956 0.003
R10916 S.n9535 S.n9534 0.003
R10917 S.n9280 S.n9279 0.003
R10918 S.n8668 S.n8667 0.003
R10919 S.n8876 S.n8875 0.003
R10920 S.n7972 S.n7971 0.003
R10921 S.n8164 S.n8163 0.003
R10922 S.n7419 S.n7418 0.003
R10923 S.n7153 S.n7152 0.003
R10924 S.n6673 S.n6672 0.003
R10925 S.n6406 S.n6405 0.003
R10926 S.n5918 S.n5917 0.003
R10927 S.n5646 S.n5645 0.003
R10928 S.n5150 S.n5149 0.003
R10929 S.n5166 S.n5165 0.003
R10930 S.n5141 S.n5140 0.003
R10931 S.n5955 S.n5954 0.003
R10932 S.n12731 S.n12730 0.003
R10933 S.n13000 S.n12999 0.003
R10934 S.n12109 S.n12108 0.003
R10935 S.n11816 S.n11815 0.003
R10936 S.n11501 S.n11500 0.003
R10937 S.n11253 S.n11252 0.003
R10938 S.n10880 S.n10879 0.003
R10939 S.n10630 S.n10629 0.003
R10940 S.n10227 S.n10226 0.003
R10941 S.n9972 S.n9971 0.003
R10942 S.n9551 S.n9550 0.003
R10943 S.n9295 S.n9294 0.003
R10944 S.n8684 S.n8683 0.003
R10945 S.n8891 S.n8890 0.003
R10946 S.n7988 S.n7987 0.003
R10947 S.n8179 S.n8178 0.003
R10948 S.n7435 S.n7434 0.003
R10949 S.n7168 S.n7167 0.003
R10950 S.n6689 S.n6688 0.003
R10951 S.n6421 S.n6420 0.003
R10952 S.n5947 S.n5946 0.003
R10953 S.n5963 S.n5962 0.003
R10954 S.n5938 S.n5937 0.003
R10955 S.n6726 S.n6725 0.003
R10956 S.n12747 S.n12746 0.003
R10957 S.n13015 S.n13014 0.003
R10958 S.n12125 S.n12124 0.003
R10959 S.n11831 S.n11830 0.003
R10960 S.n11517 S.n11516 0.003
R10961 S.n11268 S.n11267 0.003
R10962 S.n10896 S.n10895 0.003
R10963 S.n10645 S.n10644 0.003
R10964 S.n10243 S.n10242 0.003
R10965 S.n9987 S.n9986 0.003
R10966 S.n9567 S.n9566 0.003
R10967 S.n9310 S.n9309 0.003
R10968 S.n8700 S.n8699 0.003
R10969 S.n8906 S.n8905 0.003
R10970 S.n8004 S.n8003 0.003
R10971 S.n8194 S.n8193 0.003
R10972 S.n7451 S.n7450 0.003
R10973 S.n7183 S.n7182 0.003
R10974 S.n6718 S.n6717 0.003
R10975 S.n6734 S.n6733 0.003
R10976 S.n6709 S.n6708 0.003
R10977 S.n7488 S.n7487 0.003
R10978 S.n12763 S.n12762 0.003
R10979 S.n13030 S.n13029 0.003
R10980 S.n12141 S.n12140 0.003
R10981 S.n11846 S.n11845 0.003
R10982 S.n11533 S.n11532 0.003
R10983 S.n11283 S.n11282 0.003
R10984 S.n10912 S.n10911 0.003
R10985 S.n10660 S.n10659 0.003
R10986 S.n10259 S.n10258 0.003
R10987 S.n10002 S.n10001 0.003
R10988 S.n9583 S.n9582 0.003
R10989 S.n9325 S.n9324 0.003
R10990 S.n8716 S.n8715 0.003
R10991 S.n8921 S.n8920 0.003
R10992 S.n8020 S.n8019 0.003
R10993 S.n8209 S.n8208 0.003
R10994 S.n7480 S.n7479 0.003
R10995 S.n7496 S.n7495 0.003
R10996 S.n7471 S.n7470 0.003
R10997 S.n8224 S.n8223 0.003
R10998 S.n12779 S.n12778 0.003
R10999 S.n13045 S.n13044 0.003
R11000 S.n12157 S.n12156 0.003
R11001 S.n11861 S.n11860 0.003
R11002 S.n11549 S.n11548 0.003
R11003 S.n11298 S.n11297 0.003
R11004 S.n10928 S.n10927 0.003
R11005 S.n10675 S.n10674 0.003
R11006 S.n10275 S.n10274 0.003
R11007 S.n10017 S.n10016 0.003
R11008 S.n9599 S.n9598 0.003
R11009 S.n9340 S.n9339 0.003
R11010 S.n8732 S.n8731 0.003
R11011 S.n8936 S.n8935 0.003
R11012 S.n8035 S.n8034 0.003
R11013 S.n8232 S.n8231 0.003
R11014 S.n8055 S.n8054 0.003
R11015 S.n8951 S.n8950 0.003
R11016 S.n12795 S.n12794 0.003
R11017 S.n13060 S.n13059 0.003
R11018 S.n12173 S.n12172 0.003
R11019 S.n11876 S.n11875 0.003
R11020 S.n11565 S.n11564 0.003
R11021 S.n11313 S.n11312 0.003
R11022 S.n10944 S.n10943 0.003
R11023 S.n10690 S.n10689 0.003
R11024 S.n10291 S.n10290 0.003
R11025 S.n10032 S.n10031 0.003
R11026 S.n9615 S.n9614 0.003
R11027 S.n9355 S.n9354 0.003
R11028 S.n8747 S.n8746 0.003
R11029 S.n8959 S.n8958 0.003
R11030 S.n8767 S.n8766 0.003
R11031 S.n9652 S.n9651 0.003
R11032 S.n12811 S.n12810 0.003
R11033 S.n13075 S.n13074 0.003
R11034 S.n12189 S.n12188 0.003
R11035 S.n11891 S.n11890 0.003
R11036 S.n11581 S.n11580 0.003
R11037 S.n11328 S.n11327 0.003
R11038 S.n10960 S.n10959 0.003
R11039 S.n10705 S.n10704 0.003
R11040 S.n10307 S.n10306 0.003
R11041 S.n10047 S.n10046 0.003
R11042 S.n9644 S.n9643 0.003
R11043 S.n9660 S.n9659 0.003
R11044 S.n9635 S.n9634 0.003
R11045 S.n10344 S.n10343 0.003
R11046 S.n12827 S.n12826 0.003
R11047 S.n13090 S.n13089 0.003
R11048 S.n12205 S.n12204 0.003
R11049 S.n11906 S.n11905 0.003
R11050 S.n11597 S.n11596 0.003
R11051 S.n11343 S.n11342 0.003
R11052 S.n10976 S.n10975 0.003
R11053 S.n10720 S.n10719 0.003
R11054 S.n10336 S.n10335 0.003
R11055 S.n10352 S.n10351 0.003
R11056 S.n10327 S.n10326 0.003
R11057 S.n11013 S.n11012 0.003
R11058 S.n12843 S.n12842 0.003
R11059 S.n13105 S.n13104 0.003
R11060 S.n12221 S.n12220 0.003
R11061 S.n11921 S.n11920 0.003
R11062 S.n11613 S.n11612 0.003
R11063 S.n11358 S.n11357 0.003
R11064 S.n11005 S.n11004 0.003
R11065 S.n11021 S.n11020 0.003
R11066 S.n10996 S.n10995 0.003
R11067 S.n11653 S.n11652 0.003
R11068 S.n12859 S.n12858 0.003
R11069 S.n13120 S.n13119 0.003
R11070 S.n12237 S.n12236 0.003
R11071 S.n11936 S.n11935 0.003
R11072 S.n11645 S.n11644 0.003
R11073 S.n11661 S.n11660 0.003
R11074 S.n11636 S.n11635 0.003
R11075 S.n12268 S.n12267 0.003
R11076 S.n12875 S.n12874 0.003
R11077 S.n13138 S.n13137 0.003
R11078 S.n12243 S.n12242 0.003
R11079 S.n12669 S.n12668 0.003
R11080 S.n13144 S.n13143 0.003
R11081 S.n1232 S.n1231 0.003
R11082 S.n12640 S.n12635 0.003
R11083 S.n12564 S.n12559 0.003
R11084 S.n12009 S.n11997 0.003
R11085 S.n851 S.n841 0.003
R11086 S.n823 S.n818 0.003
R11087 S.n1785 S.n1777 0.003
R11088 S.n12591 S.n12579 0.003
R11089 S.n11985 S.n11980 0.003
R11090 S.n11692 S.n11683 0.003
R11091 S.n11433 S.n11428 0.003
R11092 S.n11095 S.n11086 0.003
R11093 S.n10812 S.n10807 0.003
R11094 S.n10470 S.n10461 0.003
R11095 S.n10159 S.n10154 0.003
R11096 S.n9810 S.n9801 0.003
R11097 S.n9483 S.n9478 0.003
R11098 S.n9138 S.n9129 0.003
R11099 S.n8616 S.n8611 0.003
R11100 S.n8443 S.n8434 0.003
R11101 S.n7920 S.n7915 0.003
R11102 S.n7736 S.n7727 0.003
R11103 S.n7367 S.n7362 0.003
R11104 S.n7006 S.n6997 0.003
R11105 S.n6621 S.n6616 0.003
R11106 S.n6264 S.n6255 0.003
R11107 S.n5866 S.n5861 0.003
R11108 S.n5499 S.n5490 0.003
R11109 S.n5085 S.n5080 0.003
R11110 S.n4722 S.n4713 0.003
R11111 S.n4295 S.n4290 0.003
R11112 S.n3922 S.n3913 0.003
R11113 S.n3448 S.n3443 0.003
R11114 S.n3110 S.n3101 0.003
R11115 S.n2592 S.n2587 0.003
R11116 S.n2275 S.n2264 0.003
R11117 S.n1310 S.n1307 0.003
R11118 S.n729 S.n724 0.003
R11119 S.n426 S.n421 0.003
R11120 S.n1673 S.n1666 0.003
R11121 S.n9164 S.n9153 0.003
R11122 S.n8520 S.n8515 0.003
R11123 S.n8296 S.n8287 0.003
R11124 S.n7824 S.n7819 0.003
R11125 S.n7589 S.n7580 0.003
R11126 S.n7271 S.n7266 0.003
R11127 S.n6859 S.n6850 0.003
R11128 S.n6525 S.n6520 0.003
R11129 S.n6117 S.n6108 0.003
R11130 S.n5770 S.n5765 0.003
R11131 S.n5352 S.n5343 0.003
R11132 S.n4989 S.n4984 0.003
R11133 S.n4575 S.n4566 0.003
R11134 S.n4199 S.n4194 0.003
R11135 S.n3775 S.n3766 0.003
R11136 S.n3352 S.n3347 0.003
R11137 S.n2963 S.n2954 0.003
R11138 S.n2496 S.n2491 0.003
R11139 S.n2122 S.n2111 0.003
R11140 S.n1213 S.n1210 0.003
R11141 S.n446 S.n441 0.003
R11142 S.n9841 S.n9829 0.003
R11143 S.n9404 S.n9399 0.003
R11144 S.n9020 S.n9006 0.003
R11145 S.n8537 S.n8532 0.003
R11146 S.n8325 S.n8311 0.003
R11147 S.n7841 S.n7836 0.003
R11148 S.n7618 S.n7604 0.003
R11149 S.n7288 S.n7283 0.003
R11150 S.n6888 S.n6874 0.003
R11151 S.n6542 S.n6537 0.003
R11152 S.n6146 S.n6132 0.003
R11153 S.n5787 S.n5782 0.003
R11154 S.n5381 S.n5367 0.003
R11155 S.n5006 S.n5001 0.003
R11156 S.n4604 S.n4590 0.003
R11157 S.n4216 S.n4211 0.003
R11158 S.n3804 S.n3790 0.003
R11159 S.n3369 S.n3364 0.003
R11160 S.n2992 S.n2978 0.003
R11161 S.n2513 S.n2508 0.003
R11162 S.n2151 S.n2137 0.003
R11163 S.n1232 S.n1225 0.003
R11164 S.n1252 S.n1244 0.003
R11165 S.n765 S.n456 0.003
R11166 S.n780 S.n771 0.003
R11167 S.n2186 S.n2175 0.003
R11168 S.n3024 S.n3015 0.003
R11169 S.n3836 S.n3827 0.003
R11170 S.n4636 S.n4627 0.003
R11171 S.n5413 S.n5404 0.003
R11172 S.n6178 S.n6169 0.003
R11173 S.n6920 S.n6911 0.003
R11174 S.n7650 S.n7641 0.003
R11175 S.n8357 S.n8348 0.003
R11176 S.n9052 S.n9043 0.003
R11177 S.n9724 S.n9715 0.003
R11178 S.n10499 S.n10488 0.003
R11179 S.n10099 S.n10094 0.003
R11180 S.n9423 S.n9418 0.003
R11181 S.n8556 S.n8551 0.003
R11182 S.n7860 S.n7855 0.003
R11183 S.n7307 S.n7302 0.003
R11184 S.n6561 S.n6556 0.003
R11185 S.n5806 S.n5801 0.003
R11186 S.n5025 S.n5020 0.003
R11187 S.n4235 S.n4230 0.003
R11188 S.n3388 S.n3383 0.003
R11189 S.n2532 S.n2527 0.003
R11190 S.n1735 S.n1722 0.003
R11191 S.n690 S.n681 0.003
R11192 S.n901 S.n226 0.003
R11193 S.n11122 S.n11117 0.003
R11194 S.n10773 S.n10771 0.003
R11195 S.n10418 S.n10406 0.003
R11196 S.n10120 S.n10118 0.003
R11197 S.n9758 S.n9746 0.003
R11198 S.n9444 S.n9442 0.003
R11199 S.n9086 S.n9074 0.003
R11200 S.n8577 S.n8575 0.003
R11201 S.n8391 S.n8379 0.003
R11202 S.n7881 S.n7879 0.003
R11203 S.n7684 S.n7672 0.003
R11204 S.n7328 S.n7326 0.003
R11205 S.n6954 S.n6942 0.003
R11206 S.n6582 S.n6580 0.003
R11207 S.n6212 S.n6200 0.003
R11208 S.n5827 S.n5825 0.003
R11209 S.n5447 S.n5435 0.003
R11210 S.n5046 S.n5044 0.003
R11211 S.n4670 S.n4658 0.003
R11212 S.n4256 S.n4254 0.003
R11213 S.n3870 S.n3858 0.003
R11214 S.n3409 S.n3407 0.003
R11215 S.n3058 S.n3046 0.003
R11216 S.n2553 S.n2551 0.003
R11217 S.n2220 S.n2208 0.003
R11218 S.n1273 S.n1271 0.003
R11219 S.n1763 S.n1750 0.003
R11220 S.n709 S.n701 0.003
R11221 S.n1293 S.n1290 0.003
R11222 S.n2241 S.n2235 0.003
R11223 S.n2573 S.n2565 0.003
R11224 S.n3078 S.n3073 0.003
R11225 S.n3429 S.n3421 0.003
R11226 S.n3890 S.n3885 0.003
R11227 S.n4276 S.n4268 0.003
R11228 S.n4690 S.n4685 0.003
R11229 S.n5066 S.n5058 0.003
R11230 S.n5467 S.n5462 0.003
R11231 S.n5847 S.n5839 0.003
R11232 S.n6232 S.n6227 0.003
R11233 S.n6602 S.n6594 0.003
R11234 S.n6974 S.n6969 0.003
R11235 S.n7348 S.n7340 0.003
R11236 S.n7704 S.n7699 0.003
R11237 S.n7901 S.n7893 0.003
R11238 S.n8411 S.n8406 0.003
R11239 S.n8597 S.n8589 0.003
R11240 S.n9106 S.n9101 0.003
R11241 S.n9464 S.n9456 0.003
R11242 S.n9778 S.n9773 0.003
R11243 S.n10140 S.n10132 0.003
R11244 S.n10438 S.n10433 0.003
R11245 S.n10793 S.n10785 0.003
R11246 S.n11063 S.n11058 0.003
R11247 S.n11414 S.n11406 0.003
R11248 S.n11717 S.n11712 0.003
R11249 S.n802 S.n791 0.003
R11250 S.n1701 S.n1688 0.003
R11251 S.n670 S.n665 0.003
R11252 S.n653 S.n648 0.003
R11253 S.n385 S.n380 0.003
R11254 S.n1614 S.n1607 0.003
R11255 S.n7762 S.n7751 0.003
R11256 S.n7235 S.n7230 0.003
R11257 S.n6798 S.n6789 0.003
R11258 S.n6489 S.n6484 0.003
R11259 S.n6056 S.n6047 0.003
R11260 S.n5734 S.n5729 0.003
R11261 S.n5291 S.n5282 0.003
R11262 S.n4953 S.n4948 0.003
R11263 S.n4514 S.n4505 0.003
R11264 S.n4163 S.n4158 0.003
R11265 S.n3714 S.n3705 0.003
R11266 S.n3316 S.n3311 0.003
R11267 S.n2902 S.n2893 0.003
R11268 S.n2460 S.n2455 0.003
R11269 S.n2059 S.n2048 0.003
R11270 S.n1179 S.n1176 0.003
R11271 S.n405 S.n400 0.003
R11272 S.n8474 S.n8462 0.003
R11273 S.n7805 S.n7800 0.003
R11274 S.n7557 S.n7543 0.003
R11275 S.n7252 S.n7247 0.003
R11276 S.n6827 S.n6813 0.003
R11277 S.n6506 S.n6501 0.003
R11278 S.n6085 S.n6071 0.003
R11279 S.n5751 S.n5746 0.003
R11280 S.n5320 S.n5306 0.003
R11281 S.n4970 S.n4965 0.003
R11282 S.n4543 S.n4529 0.003
R11283 S.n4180 S.n4175 0.003
R11284 S.n3743 S.n3729 0.003
R11285 S.n3333 S.n3328 0.003
R11286 S.n2931 S.n2917 0.003
R11287 S.n2477 S.n2472 0.003
R11288 S.n2088 S.n2074 0.003
R11289 S.n1196 S.n1191 0.003
R11290 S.n1643 S.n1629 0.003
R11291 S.n637 S.n632 0.003
R11292 S.n620 S.n615 0.003
R11293 S.n344 S.n339 0.003
R11294 S.n1555 S.n1548 0.003
R11295 S.n6290 S.n6279 0.003
R11296 S.n5698 S.n5693 0.003
R11297 S.n5230 S.n5221 0.003
R11298 S.n4917 S.n4912 0.003
R11299 S.n4453 S.n4444 0.003
R11300 S.n4127 S.n4122 0.003
R11301 S.n3653 S.n3644 0.003
R11302 S.n3280 S.n3275 0.003
R11303 S.n2841 S.n2832 0.003
R11304 S.n2424 S.n2419 0.003
R11305 S.n1996 S.n1985 0.003
R11306 S.n1145 S.n1142 0.003
R11307 S.n364 S.n359 0.003
R11308 S.n7037 S.n7025 0.003
R11309 S.n6470 S.n6465 0.003
R11310 S.n6024 S.n6010 0.003
R11311 S.n5715 S.n5710 0.003
R11312 S.n5259 S.n5245 0.003
R11313 S.n4934 S.n4929 0.003
R11314 S.n4482 S.n4468 0.003
R11315 S.n4144 S.n4139 0.003
R11316 S.n3682 S.n3668 0.003
R11317 S.n3297 S.n3292 0.003
R11318 S.n2870 S.n2856 0.003
R11319 S.n2441 S.n2436 0.003
R11320 S.n2025 S.n2011 0.003
R11321 S.n1162 S.n1157 0.003
R11322 S.n1584 S.n1570 0.003
R11323 S.n604 S.n599 0.003
R11324 S.n587 S.n582 0.003
R11325 S.n323 S.n318 0.003
R11326 S.n1496 S.n1489 0.003
R11327 S.n4748 S.n4737 0.003
R11328 S.n4091 S.n4086 0.003
R11329 S.n3592 S.n3583 0.003
R11330 S.n3244 S.n3239 0.003
R11331 S.n2780 S.n2771 0.003
R11332 S.n2388 S.n2383 0.003
R11333 S.n1933 S.n1922 0.003
R11334 S.n1111 S.n1108 0.003
R11335 S.n59 S.n48 0.003
R11336 S.n5530 S.n5518 0.003
R11337 S.n4898 S.n4893 0.003
R11338 S.n4421 S.n4407 0.003
R11339 S.n4108 S.n4103 0.003
R11340 S.n3621 S.n3607 0.003
R11341 S.n3261 S.n3256 0.003
R11342 S.n2809 S.n2795 0.003
R11343 S.n2405 S.n2400 0.003
R11344 S.n1962 S.n1948 0.003
R11345 S.n1128 S.n1123 0.003
R11346 S.n1525 S.n1511 0.003
R11347 S.n571 S.n566 0.003
R11348 S.n554 S.n549 0.003
R11349 S.n282 S.n277 0.003
R11350 S.n1437 S.n1430 0.003
R11351 S.n3136 S.n3125 0.003
R11352 S.n2352 S.n2347 0.003
R11353 S.n1870 S.n1859 0.003
R11354 S.n1077 S.n1074 0.003
R11355 S.n302 S.n297 0.003
R11356 S.n3953 S.n3941 0.003
R11357 S.n3225 S.n3220 0.003
R11358 S.n2748 S.n2734 0.003
R11359 S.n2369 S.n2364 0.003
R11360 S.n1899 S.n1885 0.003
R11361 S.n1094 S.n1089 0.003
R11362 S.n1469 S.n1452 0.003
R11363 S.n538 S.n533 0.003
R11364 S.n521 S.n516 0.003
R11365 S.n241 S.n236 0.003
R11366 S.n1378 S.n1369 0.003
R11367 S.n261 S.n256 0.003
R11368 S.n2306 S.n2294 0.003
R11369 S.n1060 S.n1055 0.003
R11370 S.n1407 S.n1393 0.003
R11371 S.n505 S.n500 0.003
R11372 S.n488 S.n483 0.003
R11373 S.n748 S.n741 0.003
R11374 S.n1355 S.n1350 0.003
R11375 S.n1346 S.n1027 0.003
R11376 S.n2646 S.n2637 0.003
R11377 S.n2632 S.n2316 0.003
R11378 S.n3173 S.n3164 0.003
R11379 S.n3159 S.n3146 0.003
R11380 S.n3990 S.n3981 0.003
R11381 S.n3976 S.n3963 0.003
R11382 S.n4785 S.n4776 0.003
R11383 S.n4771 S.n4758 0.003
R11384 S.n5567 S.n5558 0.003
R11385 S.n5553 S.n5540 0.003
R11386 S.n6327 S.n6318 0.003
R11387 S.n6313 S.n6300 0.003
R11388 S.n7074 S.n7065 0.003
R11389 S.n7060 S.n7047 0.003
R11390 S.n8085 S.n8076 0.003
R11391 S.n8071 S.n7772 0.003
R11392 S.n8797 S.n8788 0.003
R11393 S.n8783 S.n8484 0.003
R11394 S.n9201 S.n9192 0.003
R11395 S.n9187 S.n9174 0.003
R11396 S.n9878 S.n9869 0.003
R11397 S.n9864 S.n9851 0.003
R11398 S.n10536 S.n10527 0.003
R11399 S.n10522 S.n10509 0.003
R11400 S.n11159 S.n11150 0.003
R11401 S.n11145 S.n11132 0.003
R11402 S.n11737 S.n11728 0.003
R11403 S.n12027 S.n12020 0.003
R11404 S.n12906 S.n12897 0.003
R11405 S.n12891 S.n12601 0.003
R11406 S.n1327 S.n1322 0.003
R11407 S.n2676 S.n2660 0.003
R11408 S.n12935 S.n12934 0.003
R11409 S.n12937 S.n12920 0.003
R11410 S.n12042 S.n12041 0.003
R11411 S.n11753 S.n11751 0.003
R11412 S.n11188 S.n11187 0.003
R11413 S.n11190 S.n11173 0.003
R11414 S.n10565 S.n10564 0.003
R11415 S.n10567 S.n10550 0.003
R11416 S.n9907 S.n9906 0.003
R11417 S.n9909 S.n9892 0.003
R11418 S.n9230 S.n9229 0.003
R11419 S.n9232 S.n9215 0.003
R11420 S.n8826 S.n8825 0.003
R11421 S.n8828 S.n8811 0.003
R11422 S.n8114 S.n8113 0.003
R11423 S.n8116 S.n8099 0.003
R11424 S.n7103 S.n7102 0.003
R11425 S.n7105 S.n7088 0.003
R11426 S.n6356 S.n6355 0.003
R11427 S.n6358 S.n6341 0.003
R11428 S.n5596 S.n5595 0.003
R11429 S.n5598 S.n5581 0.003
R11430 S.n4814 S.n4813 0.003
R11431 S.n4816 S.n4799 0.003
R11432 S.n4022 S.n4021 0.003
R11433 S.n4024 S.n4007 0.003
R11434 S.n3500 S.n3499 0.003
R11435 S.n3502 S.n3187 0.003
R11436 S.n2675 S.n2674 0.003
R11437 S.n2613 S.n2604 0.003
R11438 S.n3517 S.n3516 0.003
R11439 S.n12680 S.n12678 0.003
R11440 S.n12952 S.n12951 0.003
R11441 S.n12058 S.n12056 0.003
R11442 S.n11768 S.n11767 0.003
R11443 S.n11450 S.n11448 0.003
R11444 S.n11205 S.n11204 0.003
R11445 S.n10829 S.n10827 0.003
R11446 S.n10582 S.n10581 0.003
R11447 S.n10176 S.n10174 0.003
R11448 S.n9924 S.n9923 0.003
R11449 S.n9500 S.n9498 0.003
R11450 S.n9247 S.n9246 0.003
R11451 S.n8633 S.n8631 0.003
R11452 S.n8843 S.n8842 0.003
R11453 S.n7937 S.n7935 0.003
R11454 S.n8131 S.n8130 0.003
R11455 S.n7384 S.n7382 0.003
R11456 S.n7120 S.n7119 0.003
R11457 S.n6638 S.n6636 0.003
R11458 S.n6373 S.n6372 0.003
R11459 S.n5883 S.n5881 0.003
R11460 S.n5613 S.n5612 0.003
R11461 S.n5102 S.n5100 0.003
R11462 S.n4831 S.n4830 0.003
R11463 S.n4312 S.n4310 0.003
R11464 S.n4036 S.n4035 0.003
R11465 S.n3464 S.n3463 0.003
R11466 S.n3484 S.n3475 0.003
R11467 S.n4349 S.n4050 0.003
R11468 S.n12696 S.n12694 0.003
R11469 S.n12967 S.n12966 0.003
R11470 S.n12074 S.n12072 0.003
R11471 S.n11783 S.n11782 0.003
R11472 S.n11466 S.n11464 0.003
R11473 S.n11220 S.n11219 0.003
R11474 S.n10845 S.n10843 0.003
R11475 S.n10597 S.n10596 0.003
R11476 S.n10192 S.n10190 0.003
R11477 S.n9939 S.n9938 0.003
R11478 S.n9516 S.n9514 0.003
R11479 S.n9262 S.n9261 0.003
R11480 S.n8649 S.n8647 0.003
R11481 S.n8858 S.n8857 0.003
R11482 S.n7953 S.n7951 0.003
R11483 S.n8146 S.n8145 0.003
R11484 S.n7400 S.n7398 0.003
R11485 S.n7135 S.n7134 0.003
R11486 S.n6654 S.n6652 0.003
R11487 S.n6388 S.n6387 0.003
R11488 S.n5899 S.n5897 0.003
R11489 S.n5628 S.n5627 0.003
R11490 S.n5118 S.n5116 0.003
R11491 S.n4846 S.n4845 0.003
R11492 S.n4348 S.n4347 0.003
R11493 S.n4332 S.n4323 0.003
R11494 S.n5155 S.n4860 0.003
R11495 S.n12712 S.n12710 0.003
R11496 S.n12982 S.n12981 0.003
R11497 S.n12090 S.n12088 0.003
R11498 S.n11798 S.n11797 0.003
R11499 S.n11482 S.n11480 0.003
R11500 S.n11235 S.n11234 0.003
R11501 S.n10861 S.n10859 0.003
R11502 S.n10612 S.n10611 0.003
R11503 S.n10208 S.n10206 0.003
R11504 S.n9954 S.n9953 0.003
R11505 S.n9532 S.n9530 0.003
R11506 S.n9277 S.n9276 0.003
R11507 S.n8665 S.n8663 0.003
R11508 S.n8873 S.n8872 0.003
R11509 S.n7969 S.n7967 0.003
R11510 S.n8161 S.n8160 0.003
R11511 S.n7416 S.n7414 0.003
R11512 S.n7150 S.n7149 0.003
R11513 S.n6670 S.n6668 0.003
R11514 S.n6403 S.n6402 0.003
R11515 S.n5915 S.n5913 0.003
R11516 S.n5643 S.n5642 0.003
R11517 S.n5154 S.n5153 0.003
R11518 S.n5138 S.n5129 0.003
R11519 S.n5952 S.n5657 0.003
R11520 S.n12728 S.n12726 0.003
R11521 S.n12997 S.n12996 0.003
R11522 S.n12106 S.n12104 0.003
R11523 S.n11813 S.n11812 0.003
R11524 S.n11498 S.n11496 0.003
R11525 S.n11250 S.n11249 0.003
R11526 S.n10877 S.n10875 0.003
R11527 S.n10627 S.n10626 0.003
R11528 S.n10224 S.n10222 0.003
R11529 S.n9969 S.n9968 0.003
R11530 S.n9548 S.n9546 0.003
R11531 S.n9292 S.n9291 0.003
R11532 S.n8681 S.n8679 0.003
R11533 S.n8888 S.n8887 0.003
R11534 S.n7985 S.n7983 0.003
R11535 S.n8176 S.n8175 0.003
R11536 S.n7432 S.n7430 0.003
R11537 S.n7165 S.n7164 0.003
R11538 S.n6686 S.n6684 0.003
R11539 S.n6418 S.n6417 0.003
R11540 S.n5951 S.n5950 0.003
R11541 S.n5935 S.n5926 0.003
R11542 S.n6723 S.n6432 0.003
R11543 S.n12744 S.n12742 0.003
R11544 S.n13012 S.n13011 0.003
R11545 S.n12122 S.n12120 0.003
R11546 S.n11828 S.n11827 0.003
R11547 S.n11514 S.n11512 0.003
R11548 S.n11265 S.n11264 0.003
R11549 S.n10893 S.n10891 0.003
R11550 S.n10642 S.n10641 0.003
R11551 S.n10240 S.n10238 0.003
R11552 S.n9984 S.n9983 0.003
R11553 S.n9564 S.n9562 0.003
R11554 S.n9307 S.n9306 0.003
R11555 S.n8697 S.n8695 0.003
R11556 S.n8903 S.n8902 0.003
R11557 S.n8001 S.n7999 0.003
R11558 S.n8191 S.n8190 0.003
R11559 S.n7448 S.n7446 0.003
R11560 S.n7180 S.n7179 0.003
R11561 S.n6722 S.n6721 0.003
R11562 S.n6706 S.n6697 0.003
R11563 S.n7485 S.n7194 0.003
R11564 S.n12760 S.n12758 0.003
R11565 S.n13027 S.n13026 0.003
R11566 S.n12138 S.n12136 0.003
R11567 S.n11843 S.n11842 0.003
R11568 S.n11530 S.n11528 0.003
R11569 S.n11280 S.n11279 0.003
R11570 S.n10909 S.n10907 0.003
R11571 S.n10657 S.n10656 0.003
R11572 S.n10256 S.n10254 0.003
R11573 S.n9999 S.n9998 0.003
R11574 S.n9580 S.n9578 0.003
R11575 S.n9322 S.n9321 0.003
R11576 S.n8713 S.n8711 0.003
R11577 S.n8918 S.n8917 0.003
R11578 S.n8017 S.n8015 0.003
R11579 S.n8206 S.n8205 0.003
R11580 S.n7484 S.n7483 0.003
R11581 S.n7468 S.n7459 0.003
R11582 S.n8221 S.n8220 0.003
R11583 S.n12776 S.n12774 0.003
R11584 S.n13042 S.n13041 0.003
R11585 S.n12154 S.n12152 0.003
R11586 S.n11858 S.n11857 0.003
R11587 S.n11546 S.n11544 0.003
R11588 S.n11295 S.n11294 0.003
R11589 S.n10925 S.n10923 0.003
R11590 S.n10672 S.n10671 0.003
R11591 S.n10272 S.n10270 0.003
R11592 S.n10014 S.n10013 0.003
R11593 S.n9596 S.n9594 0.003
R11594 S.n9337 S.n9336 0.003
R11595 S.n8729 S.n8727 0.003
R11596 S.n8933 S.n8932 0.003
R11597 S.n8032 S.n8031 0.003
R11598 S.n8052 S.n8043 0.003
R11599 S.n8948 S.n8947 0.003
R11600 S.n12792 S.n12790 0.003
R11601 S.n13057 S.n13056 0.003
R11602 S.n12170 S.n12168 0.003
R11603 S.n11873 S.n11872 0.003
R11604 S.n11562 S.n11560 0.003
R11605 S.n11310 S.n11309 0.003
R11606 S.n10941 S.n10939 0.003
R11607 S.n10687 S.n10686 0.003
R11608 S.n10288 S.n10286 0.003
R11609 S.n10029 S.n10028 0.003
R11610 S.n9612 S.n9610 0.003
R11611 S.n9352 S.n9351 0.003
R11612 S.n8744 S.n8743 0.003
R11613 S.n8764 S.n8755 0.003
R11614 S.n9649 S.n9366 0.003
R11615 S.n12808 S.n12806 0.003
R11616 S.n13072 S.n13071 0.003
R11617 S.n12186 S.n12184 0.003
R11618 S.n11888 S.n11887 0.003
R11619 S.n11578 S.n11576 0.003
R11620 S.n11325 S.n11324 0.003
R11621 S.n10957 S.n10955 0.003
R11622 S.n10702 S.n10701 0.003
R11623 S.n10304 S.n10302 0.003
R11624 S.n10044 S.n10043 0.003
R11625 S.n9648 S.n9647 0.003
R11626 S.n9632 S.n9623 0.003
R11627 S.n10341 S.n10058 0.003
R11628 S.n12824 S.n12822 0.003
R11629 S.n13087 S.n13086 0.003
R11630 S.n12202 S.n12200 0.003
R11631 S.n11903 S.n11902 0.003
R11632 S.n11594 S.n11592 0.003
R11633 S.n11340 S.n11339 0.003
R11634 S.n10973 S.n10971 0.003
R11635 S.n10717 S.n10716 0.003
R11636 S.n10340 S.n10339 0.003
R11637 S.n10324 S.n10315 0.003
R11638 S.n11010 S.n10731 0.003
R11639 S.n12840 S.n12838 0.003
R11640 S.n13102 S.n13101 0.003
R11641 S.n12218 S.n12216 0.003
R11642 S.n11918 S.n11917 0.003
R11643 S.n11610 S.n11608 0.003
R11644 S.n11355 S.n11354 0.003
R11645 S.n11009 S.n11008 0.003
R11646 S.n10993 S.n10984 0.003
R11647 S.n11650 S.n11369 0.003
R11648 S.n12856 S.n12854 0.003
R11649 S.n13117 S.n13116 0.003
R11650 S.n12234 S.n12232 0.003
R11651 S.n11933 S.n11932 0.003
R11652 S.n11649 S.n11648 0.003
R11653 S.n11633 S.n11619 0.003
R11654 S.n12265 S.n12259 0.003
R11655 S.n12872 S.n12867 0.003
R11656 S.n13135 S.n13130 0.003
R11657 S.n12251 S.n11948 0.003
R11658 S.n12663 S.n12658 0.003
R11659 S.n880 S.n873 0.003
R11660 S.n4 S.n2 0.003
R11661 S.n15 S.n13 0.003
R11662 S.n26 S.n24 0.003
R11663 S.n38 S.n36 0.003
R11664 S.n70 S.n68 0.003
R11665 S.n82 S.n80 0.003
R11666 S.n100 S.n98 0.003
R11667 S.n12549 S.n12315 0.003
R11668 S.n12549 S.n12548 0.003
R11669 S.n11395 S.n11394 0.003
R11670 S.n848 S.n847 0.003
R11671 S.n778 S.n777 0.003
R11672 S.n11380 S.n11379 0.003
R11673 S.n10418 S.n10417 0.003
R11674 S.n9758 S.n9757 0.003
R11675 S.n9086 S.n9085 0.003
R11676 S.n8391 S.n8390 0.003
R11677 S.n7684 S.n7683 0.003
R11678 S.n6954 S.n6953 0.003
R11679 S.n6212 S.n6211 0.003
R11680 S.n5447 S.n5446 0.003
R11681 S.n4670 S.n4669 0.003
R11682 S.n3870 S.n3869 0.003
R11683 S.n3058 S.n3057 0.003
R11684 S.n2220 S.n2219 0.003
R11685 S.n1735 S.n1718 0.003
R11686 S.n12251 S.n11944 0.003
R11687 S.t320 S.n1796 0.003
R11688 S.t320 S.n1794 0.003
R11689 S.n12618 S.n12603 0.003
R11690 S.n9388 S.n9387 0.003
R11691 S.n7789 S.n7788 0.003
R11692 S.n6454 S.n6453 0.003
R11693 S.n4882 S.n4881 0.003
R11694 S.n3209 S.n3208 0.003
R11695 S.n1044 S.n1043 0.003
R11696 S.n11708 S.n11707 0.003
R11697 S.n9404 S.n9395 0.003
R11698 S.n8537 S.n8528 0.003
R11699 S.n7841 S.n7832 0.003
R11700 S.n7288 S.n7279 0.003
R11701 S.n6542 S.n6533 0.003
R11702 S.n5787 S.n5778 0.003
R11703 S.n5006 S.n4997 0.003
R11704 S.n4216 S.n4207 0.003
R11705 S.n3369 S.n3360 0.003
R11706 S.n2513 S.n2504 0.003
R11707 S.n1232 S.n1221 0.003
R11708 S.n7805 S.n7796 0.003
R11709 S.n7252 S.n7243 0.003
R11710 S.n6506 S.n6497 0.003
R11711 S.n5751 S.n5742 0.003
R11712 S.n4970 S.n4961 0.003
R11713 S.n4180 S.n4171 0.003
R11714 S.n3333 S.n3324 0.003
R11715 S.n2477 S.n2468 0.003
R11716 S.n1196 S.n1187 0.003
R11717 S.n6470 S.n6461 0.003
R11718 S.n5715 S.n5706 0.003
R11719 S.n4934 S.n4925 0.003
R11720 S.n4144 S.n4135 0.003
R11721 S.n3297 S.n3288 0.003
R11722 S.n2441 S.n2432 0.003
R11723 S.n1162 S.n1153 0.003
R11724 S.n4898 S.n4889 0.003
R11725 S.n4108 S.n4099 0.003
R11726 S.n3261 S.n3252 0.003
R11727 S.n2405 S.n2396 0.003
R11728 S.n1128 S.n1119 0.003
R11729 S.n3225 S.n3216 0.003
R11730 S.n2369 S.n2360 0.003
R11731 S.n1094 S.n1085 0.003
R11732 S.n1060 S.n1051 0.003
R11733 S.n12564 S.n12555 0.003
R11734 S.n13161 S.n13160 0.003
R11735 S.t35 S.n12464 0.003
R11736 S.t35 S.n12327 0.003
R11737 S.n1372 S.n1371 0.003
R11738 S.n814 S.n813 0.003
R11739 S.n914 S.n913 0.003
R11740 S.n670 S.n662 0.002
R11741 S.n1701 S.n1680 0.002
R11742 S.n1232 S.n1222 0.002
R11743 S.n2151 S.n2134 0.002
R11744 S.n2513 S.n2505 0.002
R11745 S.n2992 S.n2975 0.002
R11746 S.n3369 S.n3361 0.002
R11747 S.n3804 S.n3787 0.002
R11748 S.n4216 S.n4208 0.002
R11749 S.n4604 S.n4587 0.002
R11750 S.n5006 S.n4998 0.002
R11751 S.n5381 S.n5364 0.002
R11752 S.n5787 S.n5779 0.002
R11753 S.n6146 S.n6129 0.002
R11754 S.n6542 S.n6534 0.002
R11755 S.n6888 S.n6871 0.002
R11756 S.n7288 S.n7280 0.002
R11757 S.n7618 S.n7601 0.002
R11758 S.n7841 S.n7833 0.002
R11759 S.n8325 S.n8308 0.002
R11760 S.n8537 S.n8529 0.002
R11761 S.n9020 S.n9003 0.002
R11762 S.n9404 S.n9396 0.002
R11763 S.n902 S.n901 0.002
R11764 S.n690 S.n678 0.002
R11765 S.n1735 S.n1719 0.002
R11766 S.n1273 S.n1259 0.002
R11767 S.n2220 S.n2193 0.002
R11768 S.n2553 S.n2539 0.002
R11769 S.n3058 S.n3031 0.002
R11770 S.n3409 S.n3395 0.002
R11771 S.n3870 S.n3843 0.002
R11772 S.n4256 S.n4242 0.002
R11773 S.n4670 S.n4643 0.002
R11774 S.n5046 S.n5032 0.002
R11775 S.n5447 S.n5420 0.002
R11776 S.n5827 S.n5813 0.002
R11777 S.n6212 S.n6185 0.002
R11778 S.n6582 S.n6568 0.002
R11779 S.n6954 S.n6927 0.002
R11780 S.n7328 S.n7314 0.002
R11781 S.n7684 S.n7657 0.002
R11782 S.n7881 S.n7867 0.002
R11783 S.n8391 S.n8364 0.002
R11784 S.n8577 S.n8563 0.002
R11785 S.n9086 S.n9059 0.002
R11786 S.n9444 S.n9430 0.002
R11787 S.n9758 S.n9731 0.002
R11788 S.n10120 S.n10106 0.002
R11789 S.n10418 S.n10391 0.002
R11790 S.n10773 S.n10759 0.002
R11791 S.n11414 S.n11403 0.002
R11792 S.n11063 S.n11055 0.002
R11793 S.n10793 S.n10782 0.002
R11794 S.n10438 S.n10430 0.002
R11795 S.n10140 S.n10129 0.002
R11796 S.n9778 S.n9770 0.002
R11797 S.n9464 S.n9453 0.002
R11798 S.n9106 S.n9098 0.002
R11799 S.n8597 S.n8586 0.002
R11800 S.n8411 S.n8403 0.002
R11801 S.n7901 S.n7890 0.002
R11802 S.n7704 S.n7696 0.002
R11803 S.n7348 S.n7337 0.002
R11804 S.n6974 S.n6966 0.002
R11805 S.n6602 S.n6591 0.002
R11806 S.n6232 S.n6224 0.002
R11807 S.n5847 S.n5836 0.002
R11808 S.n5467 S.n5459 0.002
R11809 S.n5066 S.n5055 0.002
R11810 S.n4690 S.n4682 0.002
R11811 S.n4276 S.n4265 0.002
R11812 S.n3890 S.n3882 0.002
R11813 S.n3429 S.n3418 0.002
R11814 S.n3078 S.n3070 0.002
R11815 S.n2573 S.n2562 0.002
R11816 S.n2241 S.n2232 0.002
R11817 S.n1293 S.n1280 0.002
R11818 S.n1763 S.n1747 0.002
R11819 S.n709 S.n698 0.002
R11820 S.n637 S.n629 0.002
R11821 S.n1643 S.n1621 0.002
R11822 S.n1196 S.n1188 0.002
R11823 S.n2088 S.n2071 0.002
R11824 S.n2477 S.n2469 0.002
R11825 S.n2931 S.n2914 0.002
R11826 S.n3333 S.n3325 0.002
R11827 S.n3743 S.n3726 0.002
R11828 S.n4180 S.n4172 0.002
R11829 S.n4543 S.n4526 0.002
R11830 S.n4970 S.n4962 0.002
R11831 S.n5320 S.n5303 0.002
R11832 S.n5751 S.n5743 0.002
R11833 S.n6085 S.n6068 0.002
R11834 S.n6506 S.n6498 0.002
R11835 S.n6827 S.n6810 0.002
R11836 S.n7252 S.n7244 0.002
R11837 S.n7557 S.n7540 0.002
R11838 S.n7805 S.n7797 0.002
R11839 S.n604 S.n596 0.002
R11840 S.n1584 S.n1562 0.002
R11841 S.n1162 S.n1154 0.002
R11842 S.n2025 S.n2008 0.002
R11843 S.n2441 S.n2433 0.002
R11844 S.n2870 S.n2853 0.002
R11845 S.n3297 S.n3289 0.002
R11846 S.n3682 S.n3665 0.002
R11847 S.n4144 S.n4136 0.002
R11848 S.n4482 S.n4465 0.002
R11849 S.n4934 S.n4926 0.002
R11850 S.n5259 S.n5242 0.002
R11851 S.n5715 S.n5707 0.002
R11852 S.n6024 S.n6007 0.002
R11853 S.n6470 S.n6462 0.002
R11854 S.n60 S.n59 0.002
R11855 S.n571 S.n563 0.002
R11856 S.n1525 S.n1503 0.002
R11857 S.n1128 S.n1120 0.002
R11858 S.n1962 S.n1945 0.002
R11859 S.n2405 S.n2397 0.002
R11860 S.n2809 S.n2792 0.002
R11861 S.n3261 S.n3253 0.002
R11862 S.n3621 S.n3604 0.002
R11863 S.n4108 S.n4100 0.002
R11864 S.n4421 S.n4404 0.002
R11865 S.n4898 S.n4890 0.002
R11866 S.n538 S.n530 0.002
R11867 S.n1469 S.n1444 0.002
R11868 S.n1094 S.n1086 0.002
R11869 S.n1899 S.n1882 0.002
R11870 S.n2369 S.n2361 0.002
R11871 S.n2748 S.n2731 0.002
R11872 S.n3225 S.n3217 0.002
R11873 S.n505 S.n497 0.002
R11874 S.n1407 S.n1385 0.002
R11875 S.n1060 S.n1052 0.002
R11876 S.n12891 S.n12598 0.002
R11877 S.n12906 S.n12894 0.002
R11878 S.n12027 S.n12017 0.002
R11879 S.n11737 S.n11725 0.002
R11880 S.n11145 S.n11129 0.002
R11881 S.n11159 S.n11147 0.002
R11882 S.n10522 S.n10506 0.002
R11883 S.n10536 S.n10524 0.002
R11884 S.n9864 S.n9848 0.002
R11885 S.n9878 S.n9866 0.002
R11886 S.n9187 S.n9171 0.002
R11887 S.n9201 S.n9189 0.002
R11888 S.n8783 S.n8481 0.002
R11889 S.n8797 S.n8785 0.002
R11890 S.n8071 S.n7769 0.002
R11891 S.n8085 S.n8073 0.002
R11892 S.n7060 S.n7044 0.002
R11893 S.n7074 S.n7062 0.002
R11894 S.n6313 S.n6297 0.002
R11895 S.n6327 S.n6315 0.002
R11896 S.n5553 S.n5537 0.002
R11897 S.n5567 S.n5555 0.002
R11898 S.n4771 S.n4755 0.002
R11899 S.n4785 S.n4773 0.002
R11900 S.n3976 S.n3960 0.002
R11901 S.n3990 S.n3978 0.002
R11902 S.n3159 S.n3143 0.002
R11903 S.n3173 S.n3161 0.002
R11904 S.n2632 S.n2313 0.002
R11905 S.n2646 S.n2634 0.002
R11906 S.n1346 S.n1024 0.002
R11907 S.n1355 S.n1347 0.002
R11908 S.n12935 S.n12921 0.002
R11909 S.n12937 S.n12913 0.002
R11910 S.n12042 S.n12034 0.002
R11911 S.n11753 S.n11744 0.002
R11912 S.n11188 S.n11174 0.002
R11913 S.n11190 S.n11166 0.002
R11914 S.n10565 S.n10551 0.002
R11915 S.n10567 S.n10543 0.002
R11916 S.n9907 S.n9893 0.002
R11917 S.n9909 S.n9885 0.002
R11918 S.n9230 S.n9216 0.002
R11919 S.n9232 S.n9208 0.002
R11920 S.n8826 S.n8812 0.002
R11921 S.n8828 S.n8804 0.002
R11922 S.n8114 S.n8100 0.002
R11923 S.n8116 S.n8092 0.002
R11924 S.n7103 S.n7089 0.002
R11925 S.n7105 S.n7081 0.002
R11926 S.n6356 S.n6342 0.002
R11927 S.n6358 S.n6334 0.002
R11928 S.n5596 S.n5582 0.002
R11929 S.n5598 S.n5574 0.002
R11930 S.n4814 S.n4800 0.002
R11931 S.n4816 S.n4792 0.002
R11932 S.n4022 S.n4008 0.002
R11933 S.n4024 S.n4000 0.002
R11934 S.n3500 S.n3188 0.002
R11935 S.n3502 S.n3180 0.002
R11936 S.n2675 S.n2661 0.002
R11937 S.n2676 S.n2653 0.002
R11938 S.n1327 S.n1319 0.002
R11939 S.n12680 S.n12671 0.002
R11940 S.n12952 S.n12944 0.002
R11941 S.n12058 S.n12049 0.002
R11942 S.n11768 S.n11760 0.002
R11943 S.n11450 S.n11441 0.002
R11944 S.n11205 S.n11197 0.002
R11945 S.n10829 S.n10820 0.002
R11946 S.n10582 S.n10574 0.002
R11947 S.n10176 S.n10167 0.002
R11948 S.n9924 S.n9916 0.002
R11949 S.n9500 S.n9491 0.002
R11950 S.n9247 S.n9239 0.002
R11951 S.n8633 S.n8624 0.002
R11952 S.n8843 S.n8835 0.002
R11953 S.n7937 S.n7928 0.002
R11954 S.n8131 S.n8123 0.002
R11955 S.n7384 S.n7375 0.002
R11956 S.n7120 S.n7112 0.002
R11957 S.n6638 S.n6629 0.002
R11958 S.n6373 S.n6365 0.002
R11959 S.n5883 S.n5874 0.002
R11960 S.n5613 S.n5605 0.002
R11961 S.n5102 S.n5093 0.002
R11962 S.n4831 S.n4823 0.002
R11963 S.n4312 S.n4303 0.002
R11964 S.n4036 S.n4028 0.002
R11965 S.n3464 S.n3456 0.002
R11966 S.n3517 S.n3509 0.002
R11967 S.n2613 S.n2601 0.002
R11968 S.n12696 S.n12687 0.002
R11969 S.n12967 S.n12959 0.002
R11970 S.n12074 S.n12065 0.002
R11971 S.n11783 S.n11775 0.002
R11972 S.n11466 S.n11457 0.002
R11973 S.n11220 S.n11212 0.002
R11974 S.n10845 S.n10836 0.002
R11975 S.n10597 S.n10589 0.002
R11976 S.n10192 S.n10183 0.002
R11977 S.n9939 S.n9931 0.002
R11978 S.n9516 S.n9507 0.002
R11979 S.n9262 S.n9254 0.002
R11980 S.n8649 S.n8640 0.002
R11981 S.n8858 S.n8850 0.002
R11982 S.n7953 S.n7944 0.002
R11983 S.n8146 S.n8138 0.002
R11984 S.n7400 S.n7391 0.002
R11985 S.n7135 S.n7127 0.002
R11986 S.n6654 S.n6645 0.002
R11987 S.n6388 S.n6380 0.002
R11988 S.n5899 S.n5890 0.002
R11989 S.n5628 S.n5620 0.002
R11990 S.n5118 S.n5109 0.002
R11991 S.n4846 S.n4838 0.002
R11992 S.n4348 S.n4051 0.002
R11993 S.n4349 S.n4043 0.002
R11994 S.n3484 S.n3472 0.002
R11995 S.n12712 S.n12703 0.002
R11996 S.n12982 S.n12974 0.002
R11997 S.n12090 S.n12081 0.002
R11998 S.n11798 S.n11790 0.002
R11999 S.n11482 S.n11473 0.002
R12000 S.n11235 S.n11227 0.002
R12001 S.n10861 S.n10852 0.002
R12002 S.n10612 S.n10604 0.002
R12003 S.n10208 S.n10199 0.002
R12004 S.n9954 S.n9946 0.002
R12005 S.n9532 S.n9523 0.002
R12006 S.n9277 S.n9269 0.002
R12007 S.n8665 S.n8656 0.002
R12008 S.n8873 S.n8865 0.002
R12009 S.n7969 S.n7960 0.002
R12010 S.n8161 S.n8153 0.002
R12011 S.n7416 S.n7407 0.002
R12012 S.n7150 S.n7142 0.002
R12013 S.n6670 S.n6661 0.002
R12014 S.n6403 S.n6395 0.002
R12015 S.n5915 S.n5906 0.002
R12016 S.n5643 S.n5635 0.002
R12017 S.n5154 S.n4861 0.002
R12018 S.n5155 S.n4853 0.002
R12019 S.n4332 S.n4320 0.002
R12020 S.n12728 S.n12719 0.002
R12021 S.n12997 S.n12989 0.002
R12022 S.n12106 S.n12097 0.002
R12023 S.n11813 S.n11805 0.002
R12024 S.n11498 S.n11489 0.002
R12025 S.n11250 S.n11242 0.002
R12026 S.n10877 S.n10868 0.002
R12027 S.n10627 S.n10619 0.002
R12028 S.n10224 S.n10215 0.002
R12029 S.n9969 S.n9961 0.002
R12030 S.n9548 S.n9539 0.002
R12031 S.n9292 S.n9284 0.002
R12032 S.n8681 S.n8672 0.002
R12033 S.n8888 S.n8880 0.002
R12034 S.n7985 S.n7976 0.002
R12035 S.n8176 S.n8168 0.002
R12036 S.n7432 S.n7423 0.002
R12037 S.n7165 S.n7157 0.002
R12038 S.n6686 S.n6677 0.002
R12039 S.n6418 S.n6410 0.002
R12040 S.n5951 S.n5658 0.002
R12041 S.n5952 S.n5650 0.002
R12042 S.n5138 S.n5126 0.002
R12043 S.n12744 S.n12735 0.002
R12044 S.n13012 S.n13004 0.002
R12045 S.n12122 S.n12113 0.002
R12046 S.n11828 S.n11820 0.002
R12047 S.n11514 S.n11505 0.002
R12048 S.n11265 S.n11257 0.002
R12049 S.n10893 S.n10884 0.002
R12050 S.n10642 S.n10634 0.002
R12051 S.n10240 S.n10231 0.002
R12052 S.n9984 S.n9976 0.002
R12053 S.n9564 S.n9555 0.002
R12054 S.n9307 S.n9299 0.002
R12055 S.n8697 S.n8688 0.002
R12056 S.n8903 S.n8895 0.002
R12057 S.n8001 S.n7992 0.002
R12058 S.n8191 S.n8183 0.002
R12059 S.n7448 S.n7439 0.002
R12060 S.n7180 S.n7172 0.002
R12061 S.n6722 S.n6433 0.002
R12062 S.n6723 S.n6425 0.002
R12063 S.n5935 S.n5923 0.002
R12064 S.n12760 S.n12751 0.002
R12065 S.n13027 S.n13019 0.002
R12066 S.n12138 S.n12129 0.002
R12067 S.n11843 S.n11835 0.002
R12068 S.n11530 S.n11521 0.002
R12069 S.n11280 S.n11272 0.002
R12070 S.n10909 S.n10900 0.002
R12071 S.n10657 S.n10649 0.002
R12072 S.n10256 S.n10247 0.002
R12073 S.n9999 S.n9991 0.002
R12074 S.n9580 S.n9571 0.002
R12075 S.n9322 S.n9314 0.002
R12076 S.n8713 S.n8704 0.002
R12077 S.n8918 S.n8910 0.002
R12078 S.n8017 S.n8008 0.002
R12079 S.n8206 S.n8198 0.002
R12080 S.n7484 S.n7195 0.002
R12081 S.n7485 S.n7187 0.002
R12082 S.n6706 S.n6694 0.002
R12083 S.n12776 S.n12767 0.002
R12084 S.n13042 S.n13034 0.002
R12085 S.n12154 S.n12145 0.002
R12086 S.n11858 S.n11850 0.002
R12087 S.n11546 S.n11537 0.002
R12088 S.n11295 S.n11287 0.002
R12089 S.n10925 S.n10916 0.002
R12090 S.n10672 S.n10664 0.002
R12091 S.n10272 S.n10263 0.002
R12092 S.n10014 S.n10006 0.002
R12093 S.n9596 S.n9587 0.002
R12094 S.n9337 S.n9329 0.002
R12095 S.n8729 S.n8720 0.002
R12096 S.n8933 S.n8925 0.002
R12097 S.n8032 S.n8024 0.002
R12098 S.n8221 S.n8213 0.002
R12099 S.n7468 S.n7456 0.002
R12100 S.n12792 S.n12783 0.002
R12101 S.n13057 S.n13049 0.002
R12102 S.n12170 S.n12161 0.002
R12103 S.n11873 S.n11865 0.002
R12104 S.n11562 S.n11553 0.002
R12105 S.n11310 S.n11302 0.002
R12106 S.n10941 S.n10932 0.002
R12107 S.n10687 S.n10679 0.002
R12108 S.n10288 S.n10279 0.002
R12109 S.n10029 S.n10021 0.002
R12110 S.n9612 S.n9603 0.002
R12111 S.n9352 S.n9344 0.002
R12112 S.n8744 S.n8736 0.002
R12113 S.n8948 S.n8940 0.002
R12114 S.n8052 S.n8040 0.002
R12115 S.n12808 S.n12799 0.002
R12116 S.n13072 S.n13064 0.002
R12117 S.n12186 S.n12177 0.002
R12118 S.n11888 S.n11880 0.002
R12119 S.n11578 S.n11569 0.002
R12120 S.n11325 S.n11317 0.002
R12121 S.n10957 S.n10948 0.002
R12122 S.n10702 S.n10694 0.002
R12123 S.n10304 S.n10295 0.002
R12124 S.n10044 S.n10036 0.002
R12125 S.n9648 S.n9367 0.002
R12126 S.n9649 S.n9359 0.002
R12127 S.n8764 S.n8752 0.002
R12128 S.n12824 S.n12815 0.002
R12129 S.n13087 S.n13079 0.002
R12130 S.n12202 S.n12193 0.002
R12131 S.n11903 S.n11895 0.002
R12132 S.n11594 S.n11585 0.002
R12133 S.n11340 S.n11332 0.002
R12134 S.n10973 S.n10964 0.002
R12135 S.n10717 S.n10709 0.002
R12136 S.n10340 S.n10059 0.002
R12137 S.n10341 S.n10051 0.002
R12138 S.n9632 S.n9620 0.002
R12139 S.n12840 S.n12831 0.002
R12140 S.n13102 S.n13094 0.002
R12141 S.n12218 S.n12209 0.002
R12142 S.n11918 S.n11910 0.002
R12143 S.n11610 S.n11601 0.002
R12144 S.n11355 S.n11347 0.002
R12145 S.n11009 S.n10732 0.002
R12146 S.n11010 S.n10724 0.002
R12147 S.n10324 S.n10312 0.002
R12148 S.n12856 S.n12847 0.002
R12149 S.n13117 S.n13109 0.002
R12150 S.n12234 S.n12225 0.002
R12151 S.n11933 S.n11925 0.002
R12152 S.n11649 S.n11370 0.002
R12153 S.n11650 S.n11362 0.002
R12154 S.n10993 S.n10981 0.002
R12155 S.n12251 S.n11945 0.002
R12156 S.n13135 S.n13127 0.002
R12157 S.n12872 S.n12864 0.002
R12158 S.n11633 S.n11623 0.002
R12159 S.n12265 S.n12256 0.002
R12160 S.n12009 S.n11994 0.002
R12161 S.n12564 S.n12556 0.002
R12162 S.n12640 S.n12632 0.002
R12163 S.n9841 S.n9826 0.002
R12164 S.n11122 S.n11103 0.002
R12165 S.n11717 S.n11709 0.002
R12166 S.n8474 S.n8459 0.002
R12167 S.n7037 S.n7022 0.002
R12168 S.n5530 S.n5515 0.002
R12169 S.n3953 S.n3938 0.002
R12170 S.n2306 S.n2291 0.002
R12171 S.n1827 S.n1826 0.002
R12172 S.n2710 S.n2709 0.002
R12173 S.n3551 S.n3550 0.002
R12174 S.n4383 S.n4382 0.002
R12175 S.n5189 S.n5188 0.002
R12176 S.n5986 S.n5985 0.002
R12177 S.n6757 S.n6756 0.002
R12178 S.n7519 S.n7518 0.002
R12179 S.n8255 S.n8254 0.002
R12180 S.n8982 S.n8981 0.002
R12181 S.n9683 S.n9682 0.002
R12182 S.n10375 S.n10374 0.002
R12183 S.n12626 S.n12625 0.002
R12184 S.n12649 S.n12648 0.002
R12185 S.n12422 S.n12421 0.002
R12186 S.n12425 S.n12424 0.002
R12187 S.n12428 S.n12427 0.002
R12188 S.n12431 S.n12430 0.002
R12189 S.n12434 S.n12433 0.002
R12190 S.n12437 S.n12436 0.002
R12191 S.n12440 S.n12439 0.002
R12192 S.n12443 S.n12442 0.002
R12193 S.n12446 S.n12445 0.002
R12194 S.n12449 S.n12448 0.002
R12195 S.n12452 S.n12451 0.002
R12196 S.n12455 S.n12454 0.002
R12197 S.n12458 S.n12457 0.002
R12198 S.n12461 S.n12460 0.002
R12199 S.t28 S.n937 0.002
R12200 S.n1355 S.n1354 0.002
R12201 S.n838 S.n837 0.002
R12202 S.n12585 S.n12584 0.002
R12203 S.n10493 S.n10492 0.002
R12204 S.n9158 S.n9157 0.002
R12205 S.n7756 S.n7755 0.002
R12206 S.n6284 S.n6283 0.002
R12207 S.n4742 S.n4741 0.002
R12208 S.n3130 S.n3129 0.002
R12209 S.n1785 S.n1771 0.002
R12210 S.n1673 S.n1660 0.002
R12211 S.n2151 S.n2150 0.002
R12212 S.n2513 S.n2512 0.002
R12213 S.n2992 S.n2991 0.002
R12214 S.n3369 S.n3368 0.002
R12215 S.n3804 S.n3803 0.002
R12216 S.n4216 S.n4215 0.002
R12217 S.n4604 S.n4603 0.002
R12218 S.n5006 S.n5005 0.002
R12219 S.n5381 S.n5380 0.002
R12220 S.n5787 S.n5786 0.002
R12221 S.n6146 S.n6145 0.002
R12222 S.n6542 S.n6541 0.002
R12223 S.n6888 S.n6887 0.002
R12224 S.n7288 S.n7287 0.002
R12225 S.n7618 S.n7617 0.002
R12226 S.n7841 S.n7840 0.002
R12227 S.n8325 S.n8324 0.002
R12228 S.n8537 S.n8536 0.002
R12229 S.n9020 S.n9019 0.002
R12230 S.n9404 S.n9403 0.002
R12231 S.n1614 S.n1601 0.002
R12232 S.n1196 S.n1195 0.002
R12233 S.n2088 S.n2087 0.002
R12234 S.n2477 S.n2476 0.002
R12235 S.n2931 S.n2930 0.002
R12236 S.n3333 S.n3332 0.002
R12237 S.n3743 S.n3742 0.002
R12238 S.n4180 S.n4179 0.002
R12239 S.n4543 S.n4542 0.002
R12240 S.n4970 S.n4969 0.002
R12241 S.n5320 S.n5319 0.002
R12242 S.n5751 S.n5750 0.002
R12243 S.n6085 S.n6084 0.002
R12244 S.n6506 S.n6505 0.002
R12245 S.n6827 S.n6826 0.002
R12246 S.n7252 S.n7251 0.002
R12247 S.n7557 S.n7556 0.002
R12248 S.n7805 S.n7804 0.002
R12249 S.n1555 S.n1542 0.002
R12250 S.n1162 S.n1161 0.002
R12251 S.n2025 S.n2024 0.002
R12252 S.n2441 S.n2440 0.002
R12253 S.n2870 S.n2869 0.002
R12254 S.n3297 S.n3296 0.002
R12255 S.n3682 S.n3681 0.002
R12256 S.n4144 S.n4143 0.002
R12257 S.n4482 S.n4481 0.002
R12258 S.n4934 S.n4933 0.002
R12259 S.n5259 S.n5258 0.002
R12260 S.n5715 S.n5714 0.002
R12261 S.n6024 S.n6023 0.002
R12262 S.n6470 S.n6469 0.002
R12263 S.n1496 S.n1483 0.002
R12264 S.n1128 S.n1127 0.002
R12265 S.n1962 S.n1961 0.002
R12266 S.n2405 S.n2404 0.002
R12267 S.n2809 S.n2808 0.002
R12268 S.n3261 S.n3260 0.002
R12269 S.n3621 S.n3620 0.002
R12270 S.n4108 S.n4107 0.002
R12271 S.n4421 S.n4420 0.002
R12272 S.n4898 S.n4897 0.002
R12273 S.n1437 S.n1424 0.002
R12274 S.n1094 S.n1093 0.002
R12275 S.n1899 S.n1898 0.002
R12276 S.n2369 S.n2368 0.002
R12277 S.n2748 S.n2747 0.002
R12278 S.n3225 S.n3224 0.002
R12279 S.n1060 S.n1059 0.002
R12280 S.n2676 S.n2654 0.002
R12281 S.n3517 S.n3510 0.002
R12282 S.n4349 S.n4044 0.002
R12283 S.n5155 S.n4854 0.002
R12284 S.n5952 S.n5651 0.002
R12285 S.n6723 S.n6426 0.002
R12286 S.n7485 S.n7188 0.002
R12287 S.n8221 S.n8214 0.002
R12288 S.n8948 S.n8941 0.002
R12289 S.n9649 S.n9360 0.002
R12290 S.n10341 S.n10052 0.002
R12291 S.n11010 S.n10725 0.002
R12292 S.n11650 S.n11363 0.002
R12293 S.n12251 S.n12250 0.002
R12294 S.n13135 S.n13134 0.002
R12295 S.n12872 S.n12871 0.002
R12296 S.n12663 S.n12662 0.002
R12297 S.n12009 S.n12008 0.002
R12298 S.n12564 S.n12563 0.002
R12299 S.n12640 S.n12639 0.002
R12300 S.n9825 S.n9824 0.002
R12301 S.n8458 S.n8457 0.002
R12302 S.n7021 S.n7020 0.002
R12303 S.n5514 S.n5513 0.002
R12304 S.n3937 S.n3936 0.002
R12305 S.n2290 S.n2289 0.002
R12306 S.n11985 S.n11974 0.002
R12307 S.n11692 S.n11677 0.002
R12308 S.n11433 S.n11422 0.002
R12309 S.n11095 S.n11080 0.002
R12310 S.n10812 S.n10801 0.002
R12311 S.n10470 S.n10455 0.002
R12312 S.n10159 S.n10148 0.002
R12313 S.n9810 S.n9795 0.002
R12314 S.n9483 S.n9472 0.002
R12315 S.n9138 S.n9123 0.002
R12316 S.n8616 S.n8605 0.002
R12317 S.n8443 S.n8428 0.002
R12318 S.n7920 S.n7909 0.002
R12319 S.n7736 S.n7721 0.002
R12320 S.n7367 S.n7356 0.002
R12321 S.n7006 S.n6991 0.002
R12322 S.n6621 S.n6610 0.002
R12323 S.n6264 S.n6249 0.002
R12324 S.n5866 S.n5855 0.002
R12325 S.n5499 S.n5484 0.002
R12326 S.n5085 S.n5074 0.002
R12327 S.n4722 S.n4707 0.002
R12328 S.n4295 S.n4284 0.002
R12329 S.n3922 S.n3907 0.002
R12330 S.n3448 S.n3437 0.002
R12331 S.n3110 S.n3095 0.002
R12332 S.n2592 S.n2581 0.002
R12333 S.n2275 S.n2258 0.002
R12334 S.n1310 S.n1301 0.002
R12335 S.n729 S.n728 0.002
R12336 S.n8520 S.n8509 0.002
R12337 S.n8296 S.n8281 0.002
R12338 S.n7824 S.n7813 0.002
R12339 S.n7589 S.n7574 0.002
R12340 S.n7271 S.n7260 0.002
R12341 S.n6859 S.n6844 0.002
R12342 S.n6525 S.n6514 0.002
R12343 S.n6117 S.n6102 0.002
R12344 S.n5770 S.n5759 0.002
R12345 S.n5352 S.n5337 0.002
R12346 S.n4989 S.n4978 0.002
R12347 S.n4575 S.n4560 0.002
R12348 S.n4199 S.n4188 0.002
R12349 S.n3775 S.n3760 0.002
R12350 S.n3352 S.n3341 0.002
R12351 S.n2963 S.n2948 0.002
R12352 S.n2496 S.n2485 0.002
R12353 S.n2122 S.n2105 0.002
R12354 S.n1213 S.n1204 0.002
R12355 S.n1701 S.n1700 0.002
R12356 S.n670 S.n669 0.002
R12357 S.n653 S.n652 0.002
R12358 S.n7235 S.n7224 0.002
R12359 S.n6798 S.n6783 0.002
R12360 S.n6489 S.n6478 0.002
R12361 S.n6056 S.n6041 0.002
R12362 S.n5734 S.n5723 0.002
R12363 S.n5291 S.n5276 0.002
R12364 S.n4953 S.n4942 0.002
R12365 S.n4514 S.n4499 0.002
R12366 S.n4163 S.n4152 0.002
R12367 S.n3714 S.n3699 0.002
R12368 S.n3316 S.n3305 0.002
R12369 S.n2902 S.n2887 0.002
R12370 S.n2460 S.n2449 0.002
R12371 S.n2059 S.n2042 0.002
R12372 S.n1179 S.n1170 0.002
R12373 S.n1643 S.n1642 0.002
R12374 S.n637 S.n636 0.002
R12375 S.n620 S.n619 0.002
R12376 S.n5698 S.n5687 0.002
R12377 S.n5230 S.n5215 0.002
R12378 S.n4917 S.n4906 0.002
R12379 S.n4453 S.n4438 0.002
R12380 S.n4127 S.n4116 0.002
R12381 S.n3653 S.n3638 0.002
R12382 S.n3280 S.n3269 0.002
R12383 S.n2841 S.n2826 0.002
R12384 S.n2424 S.n2413 0.002
R12385 S.n1996 S.n1979 0.002
R12386 S.n1145 S.n1136 0.002
R12387 S.n1584 S.n1583 0.002
R12388 S.n604 S.n603 0.002
R12389 S.n587 S.n586 0.002
R12390 S.n4091 S.n4080 0.002
R12391 S.n3592 S.n3577 0.002
R12392 S.n3244 S.n3233 0.002
R12393 S.n2780 S.n2765 0.002
R12394 S.n2388 S.n2377 0.002
R12395 S.n1933 S.n1916 0.002
R12396 S.n1111 S.n1102 0.002
R12397 S.n1525 S.n1524 0.002
R12398 S.n571 S.n570 0.002
R12399 S.n554 S.n553 0.002
R12400 S.n2352 S.n2341 0.002
R12401 S.n1870 S.n1853 0.002
R12402 S.n1077 S.n1068 0.002
R12403 S.n1469 S.n1468 0.002
R12404 S.n538 S.n537 0.002
R12405 S.n521 S.n520 0.002
R12406 S.n1407 S.n1406 0.002
R12407 S.n505 S.n504 0.002
R12408 S.n488 S.n487 0.002
R12409 S.n12935 S.n12922 0.002
R12410 S.n12937 S.n12914 0.002
R12411 S.n12042 S.n12035 0.002
R12412 S.n11753 S.n11745 0.002
R12413 S.n11188 S.n11175 0.002
R12414 S.n11190 S.n11167 0.002
R12415 S.n10565 S.n10552 0.002
R12416 S.n10567 S.n10544 0.002
R12417 S.n9907 S.n9894 0.002
R12418 S.n9909 S.n9886 0.002
R12419 S.n9230 S.n9217 0.002
R12420 S.n9232 S.n9209 0.002
R12421 S.n8826 S.n8813 0.002
R12422 S.n8828 S.n8805 0.002
R12423 S.n8114 S.n8101 0.002
R12424 S.n8116 S.n8093 0.002
R12425 S.n7103 S.n7090 0.002
R12426 S.n7105 S.n7082 0.002
R12427 S.n6356 S.n6343 0.002
R12428 S.n6358 S.n6335 0.002
R12429 S.n5596 S.n5583 0.002
R12430 S.n5598 S.n5575 0.002
R12431 S.n4814 S.n4801 0.002
R12432 S.n4816 S.n4793 0.002
R12433 S.n4022 S.n4009 0.002
R12434 S.n4024 S.n4001 0.002
R12435 S.n3500 S.n3189 0.002
R12436 S.n3502 S.n3181 0.002
R12437 S.n2675 S.n2662 0.002
R12438 S.n1327 S.n1326 0.002
R12439 S.n12680 S.n12672 0.002
R12440 S.n12952 S.n12945 0.002
R12441 S.n12058 S.n12050 0.002
R12442 S.n11768 S.n11761 0.002
R12443 S.n11450 S.n11442 0.002
R12444 S.n11205 S.n11198 0.002
R12445 S.n10829 S.n10821 0.002
R12446 S.n10582 S.n10575 0.002
R12447 S.n10176 S.n10168 0.002
R12448 S.n9924 S.n9917 0.002
R12449 S.n9500 S.n9492 0.002
R12450 S.n9247 S.n9240 0.002
R12451 S.n8633 S.n8625 0.002
R12452 S.n8843 S.n8836 0.002
R12453 S.n7937 S.n7929 0.002
R12454 S.n8131 S.n8124 0.002
R12455 S.n7384 S.n7376 0.002
R12456 S.n7120 S.n7113 0.002
R12457 S.n6638 S.n6630 0.002
R12458 S.n6373 S.n6366 0.002
R12459 S.n5883 S.n5875 0.002
R12460 S.n5613 S.n5606 0.002
R12461 S.n5102 S.n5094 0.002
R12462 S.n4831 S.n4824 0.002
R12463 S.n4312 S.n4304 0.002
R12464 S.n4036 S.n4029 0.002
R12465 S.n3464 S.n3457 0.002
R12466 S.n2613 S.n2612 0.002
R12467 S.n12696 S.n12688 0.002
R12468 S.n12967 S.n12960 0.002
R12469 S.n12074 S.n12066 0.002
R12470 S.n11783 S.n11776 0.002
R12471 S.n11466 S.n11458 0.002
R12472 S.n11220 S.n11213 0.002
R12473 S.n10845 S.n10837 0.002
R12474 S.n10597 S.n10590 0.002
R12475 S.n10192 S.n10184 0.002
R12476 S.n9939 S.n9932 0.002
R12477 S.n9516 S.n9508 0.002
R12478 S.n9262 S.n9255 0.002
R12479 S.n8649 S.n8641 0.002
R12480 S.n8858 S.n8851 0.002
R12481 S.n7953 S.n7945 0.002
R12482 S.n8146 S.n8139 0.002
R12483 S.n7400 S.n7392 0.002
R12484 S.n7135 S.n7128 0.002
R12485 S.n6654 S.n6646 0.002
R12486 S.n6388 S.n6381 0.002
R12487 S.n5899 S.n5891 0.002
R12488 S.n5628 S.n5621 0.002
R12489 S.n5118 S.n5110 0.002
R12490 S.n4846 S.n4839 0.002
R12491 S.n4348 S.n4052 0.002
R12492 S.n3484 S.n3483 0.002
R12493 S.n12712 S.n12704 0.002
R12494 S.n12982 S.n12975 0.002
R12495 S.n12090 S.n12082 0.002
R12496 S.n11798 S.n11791 0.002
R12497 S.n11482 S.n11474 0.002
R12498 S.n11235 S.n11228 0.002
R12499 S.n10861 S.n10853 0.002
R12500 S.n10612 S.n10605 0.002
R12501 S.n10208 S.n10200 0.002
R12502 S.n9954 S.n9947 0.002
R12503 S.n9532 S.n9524 0.002
R12504 S.n9277 S.n9270 0.002
R12505 S.n8665 S.n8657 0.002
R12506 S.n8873 S.n8866 0.002
R12507 S.n7969 S.n7961 0.002
R12508 S.n8161 S.n8154 0.002
R12509 S.n7416 S.n7408 0.002
R12510 S.n7150 S.n7143 0.002
R12511 S.n6670 S.n6662 0.002
R12512 S.n6403 S.n6396 0.002
R12513 S.n5915 S.n5907 0.002
R12514 S.n5643 S.n5636 0.002
R12515 S.n5154 S.n4862 0.002
R12516 S.n4332 S.n4331 0.002
R12517 S.n12728 S.n12720 0.002
R12518 S.n12997 S.n12990 0.002
R12519 S.n12106 S.n12098 0.002
R12520 S.n11813 S.n11806 0.002
R12521 S.n11498 S.n11490 0.002
R12522 S.n11250 S.n11243 0.002
R12523 S.n10877 S.n10869 0.002
R12524 S.n10627 S.n10620 0.002
R12525 S.n10224 S.n10216 0.002
R12526 S.n9969 S.n9962 0.002
R12527 S.n9548 S.n9540 0.002
R12528 S.n9292 S.n9285 0.002
R12529 S.n8681 S.n8673 0.002
R12530 S.n8888 S.n8881 0.002
R12531 S.n7985 S.n7977 0.002
R12532 S.n8176 S.n8169 0.002
R12533 S.n7432 S.n7424 0.002
R12534 S.n7165 S.n7158 0.002
R12535 S.n6686 S.n6678 0.002
R12536 S.n6418 S.n6411 0.002
R12537 S.n5951 S.n5659 0.002
R12538 S.n5138 S.n5137 0.002
R12539 S.n12744 S.n12736 0.002
R12540 S.n13012 S.n13005 0.002
R12541 S.n12122 S.n12114 0.002
R12542 S.n11828 S.n11821 0.002
R12543 S.n11514 S.n11506 0.002
R12544 S.n11265 S.n11258 0.002
R12545 S.n10893 S.n10885 0.002
R12546 S.n10642 S.n10635 0.002
R12547 S.n10240 S.n10232 0.002
R12548 S.n9984 S.n9977 0.002
R12549 S.n9564 S.n9556 0.002
R12550 S.n9307 S.n9300 0.002
R12551 S.n8697 S.n8689 0.002
R12552 S.n8903 S.n8896 0.002
R12553 S.n8001 S.n7993 0.002
R12554 S.n8191 S.n8184 0.002
R12555 S.n7448 S.n7440 0.002
R12556 S.n7180 S.n7173 0.002
R12557 S.n6722 S.n6434 0.002
R12558 S.n5935 S.n5934 0.002
R12559 S.n12760 S.n12752 0.002
R12560 S.n13027 S.n13020 0.002
R12561 S.n12138 S.n12130 0.002
R12562 S.n11843 S.n11836 0.002
R12563 S.n11530 S.n11522 0.002
R12564 S.n11280 S.n11273 0.002
R12565 S.n10909 S.n10901 0.002
R12566 S.n10657 S.n10650 0.002
R12567 S.n10256 S.n10248 0.002
R12568 S.n9999 S.n9992 0.002
R12569 S.n9580 S.n9572 0.002
R12570 S.n9322 S.n9315 0.002
R12571 S.n8713 S.n8705 0.002
R12572 S.n8918 S.n8911 0.002
R12573 S.n8017 S.n8009 0.002
R12574 S.n8206 S.n8199 0.002
R12575 S.n7484 S.n7196 0.002
R12576 S.n6706 S.n6705 0.002
R12577 S.n12776 S.n12768 0.002
R12578 S.n13042 S.n13035 0.002
R12579 S.n12154 S.n12146 0.002
R12580 S.n11858 S.n11851 0.002
R12581 S.n11546 S.n11538 0.002
R12582 S.n11295 S.n11288 0.002
R12583 S.n10925 S.n10917 0.002
R12584 S.n10672 S.n10665 0.002
R12585 S.n10272 S.n10264 0.002
R12586 S.n10014 S.n10007 0.002
R12587 S.n9596 S.n9588 0.002
R12588 S.n9337 S.n9330 0.002
R12589 S.n8729 S.n8721 0.002
R12590 S.n8933 S.n8926 0.002
R12591 S.n8032 S.n8025 0.002
R12592 S.n7468 S.n7467 0.002
R12593 S.n12792 S.n12784 0.002
R12594 S.n13057 S.n13050 0.002
R12595 S.n12170 S.n12162 0.002
R12596 S.n11873 S.n11866 0.002
R12597 S.n11562 S.n11554 0.002
R12598 S.n11310 S.n11303 0.002
R12599 S.n10941 S.n10933 0.002
R12600 S.n10687 S.n10680 0.002
R12601 S.n10288 S.n10280 0.002
R12602 S.n10029 S.n10022 0.002
R12603 S.n9612 S.n9604 0.002
R12604 S.n9352 S.n9345 0.002
R12605 S.n8744 S.n8737 0.002
R12606 S.n8052 S.n8051 0.002
R12607 S.n12808 S.n12800 0.002
R12608 S.n13072 S.n13065 0.002
R12609 S.n12186 S.n12178 0.002
R12610 S.n11888 S.n11881 0.002
R12611 S.n11578 S.n11570 0.002
R12612 S.n11325 S.n11318 0.002
R12613 S.n10957 S.n10949 0.002
R12614 S.n10702 S.n10695 0.002
R12615 S.n10304 S.n10296 0.002
R12616 S.n10044 S.n10037 0.002
R12617 S.n9648 S.n9368 0.002
R12618 S.n8764 S.n8763 0.002
R12619 S.n12824 S.n12816 0.002
R12620 S.n13087 S.n13080 0.002
R12621 S.n12202 S.n12194 0.002
R12622 S.n11903 S.n11896 0.002
R12623 S.n11594 S.n11586 0.002
R12624 S.n11340 S.n11333 0.002
R12625 S.n10973 S.n10965 0.002
R12626 S.n10717 S.n10710 0.002
R12627 S.n10340 S.n10060 0.002
R12628 S.n9632 S.n9631 0.002
R12629 S.n12840 S.n12832 0.002
R12630 S.n13102 S.n13095 0.002
R12631 S.n12218 S.n12210 0.002
R12632 S.n11918 S.n11911 0.002
R12633 S.n11610 S.n11602 0.002
R12634 S.n11355 S.n11348 0.002
R12635 S.n11009 S.n10733 0.002
R12636 S.n10324 S.n10323 0.002
R12637 S.n12856 S.n12848 0.002
R12638 S.n13117 S.n13110 0.002
R12639 S.n12234 S.n12226 0.002
R12640 S.n11933 S.n11926 0.002
R12641 S.n11649 S.n11371 0.002
R12642 S.n10993 S.n10992 0.002
R12643 S.n12265 S.n12264 0.002
R12644 S.n901 S.n223 0.002
R12645 S.n802 S.n801 0.002
R12646 S.n11633 S.n11629 0.002
R12647 S.n119 S.n116 0.002
R12648 S.t35 S.n12325 0.002
R12649 S.t35 S.n12474 0.002
R12650 S.n1809 S.n1808 0.002
R12651 S.n12591 S.n12573 0.002
R12652 S.n9164 S.n9147 0.002
R12653 S.n7762 S.n7745 0.002
R12654 S.n6290 S.n6273 0.002
R12655 S.n4748 S.n4731 0.002
R12656 S.n3136 S.n3119 0.002
R12657 S.n1378 S.n1363 0.002
R12658 S.n123 S.n122 0.002
R12659 S.n11717 S.n11716 0.002
R12660 S.n11063 S.n11062 0.002
R12661 S.n10438 S.n10437 0.002
R12662 S.n9778 S.n9777 0.002
R12663 S.n9106 S.n9105 0.002
R12664 S.n8411 S.n8410 0.002
R12665 S.n7704 S.n7703 0.002
R12666 S.n6974 S.n6973 0.002
R12667 S.n6232 S.n6231 0.002
R12668 S.n5467 S.n5466 0.002
R12669 S.n4690 S.n4689 0.002
R12670 S.n3890 S.n3889 0.002
R12671 S.n3078 S.n3077 0.002
R12672 S.n2241 S.n2240 0.002
R12673 S.n2613 S.n2600 0.002
R12674 S.n4312 S.n4311 0.002
R12675 S.n5102 S.n5101 0.002
R12676 S.n5883 S.n5882 0.002
R12677 S.n6638 S.n6637 0.002
R12678 S.n7384 S.n7383 0.002
R12679 S.n7937 S.n7936 0.002
R12680 S.n8633 S.n8632 0.002
R12681 S.n9500 S.n9499 0.002
R12682 S.n10176 S.n10175 0.002
R12683 S.n10829 S.n10828 0.002
R12684 S.n11450 S.n11449 0.002
R12685 S.n12058 S.n12057 0.002
R12686 S.n12680 S.n12679 0.002
R12687 S.n3484 S.n3471 0.002
R12688 S.n5118 S.n5117 0.002
R12689 S.n5899 S.n5898 0.002
R12690 S.n6654 S.n6653 0.002
R12691 S.n7400 S.n7399 0.002
R12692 S.n7953 S.n7952 0.002
R12693 S.n8649 S.n8648 0.002
R12694 S.n9516 S.n9515 0.002
R12695 S.n10192 S.n10191 0.002
R12696 S.n10845 S.n10844 0.002
R12697 S.n11466 S.n11465 0.002
R12698 S.n12074 S.n12073 0.002
R12699 S.n12696 S.n12695 0.002
R12700 S.n4332 S.n4319 0.002
R12701 S.n5915 S.n5914 0.002
R12702 S.n6670 S.n6669 0.002
R12703 S.n7416 S.n7415 0.002
R12704 S.n7969 S.n7968 0.002
R12705 S.n8665 S.n8664 0.002
R12706 S.n9532 S.n9531 0.002
R12707 S.n10208 S.n10207 0.002
R12708 S.n10861 S.n10860 0.002
R12709 S.n11482 S.n11481 0.002
R12710 S.n12090 S.n12089 0.002
R12711 S.n12712 S.n12711 0.002
R12712 S.n5138 S.n5125 0.002
R12713 S.n6686 S.n6685 0.002
R12714 S.n7432 S.n7431 0.002
R12715 S.n7985 S.n7984 0.002
R12716 S.n8681 S.n8680 0.002
R12717 S.n9548 S.n9547 0.002
R12718 S.n10224 S.n10223 0.002
R12719 S.n10877 S.n10876 0.002
R12720 S.n11498 S.n11497 0.002
R12721 S.n12106 S.n12105 0.002
R12722 S.n12728 S.n12727 0.002
R12723 S.n5935 S.n5922 0.002
R12724 S.n7448 S.n7447 0.002
R12725 S.n8001 S.n8000 0.002
R12726 S.n8697 S.n8696 0.002
R12727 S.n9564 S.n9563 0.002
R12728 S.n10240 S.n10239 0.002
R12729 S.n10893 S.n10892 0.002
R12730 S.n11514 S.n11513 0.002
R12731 S.n12122 S.n12121 0.002
R12732 S.n12744 S.n12743 0.002
R12733 S.n6706 S.n6693 0.002
R12734 S.n8017 S.n8016 0.002
R12735 S.n8713 S.n8712 0.002
R12736 S.n9580 S.n9579 0.002
R12737 S.n10256 S.n10255 0.002
R12738 S.n10909 S.n10908 0.002
R12739 S.n11530 S.n11529 0.002
R12740 S.n12138 S.n12137 0.002
R12741 S.n12760 S.n12759 0.002
R12742 S.n7468 S.n7455 0.002
R12743 S.n8729 S.n8728 0.002
R12744 S.n9596 S.n9595 0.002
R12745 S.n10272 S.n10271 0.002
R12746 S.n10925 S.n10924 0.002
R12747 S.n11546 S.n11545 0.002
R12748 S.n12154 S.n12153 0.002
R12749 S.n12776 S.n12775 0.002
R12750 S.n8052 S.n8039 0.002
R12751 S.n9612 S.n9611 0.002
R12752 S.n10288 S.n10287 0.002
R12753 S.n10941 S.n10940 0.002
R12754 S.n11562 S.n11561 0.002
R12755 S.n12170 S.n12169 0.002
R12756 S.n12792 S.n12791 0.002
R12757 S.n8764 S.n8751 0.002
R12758 S.n10304 S.n10303 0.002
R12759 S.n10957 S.n10956 0.002
R12760 S.n11578 S.n11577 0.002
R12761 S.n12186 S.n12185 0.002
R12762 S.n12808 S.n12807 0.002
R12763 S.n9632 S.n9619 0.002
R12764 S.n10973 S.n10972 0.002
R12765 S.n11594 S.n11593 0.002
R12766 S.n12202 S.n12201 0.002
R12767 S.n12824 S.n12823 0.002
R12768 S.n10324 S.n10311 0.002
R12769 S.n11610 S.n11609 0.002
R12770 S.n12218 S.n12217 0.002
R12771 S.n12840 S.n12839 0.002
R12772 S.n10993 S.n10980 0.002
R12773 S.n12234 S.n12233 0.002
R12774 S.n12856 S.n12855 0.002
R12775 S.n12872 S.n12863 0.002
R12776 S.n10773 S.n10772 0.002
R12777 S.n10120 S.n10119 0.002
R12778 S.n9444 S.n9443 0.002
R12779 S.n8577 S.n8576 0.002
R12780 S.n7881 S.n7880 0.002
R12781 S.n7328 S.n7327 0.002
R12782 S.n6582 S.n6581 0.002
R12783 S.n5827 S.n5826 0.002
R12784 S.n5046 S.n5045 0.002
R12785 S.n4256 S.n4255 0.002
R12786 S.n3409 S.n3408 0.002
R12787 S.n2553 S.n2552 0.002
R12788 S.n1273 S.n1272 0.002
R12789 S.n690 S.n677 0.002
R12790 S.n748 S.n737 0.002
R12791 S.n2633 S.n2632 0.002
R12792 S.n3160 S.n3159 0.002
R12793 S.n3977 S.n3976 0.002
R12794 S.n4772 S.n4771 0.002
R12795 S.n5554 S.n5553 0.002
R12796 S.n6314 S.n6313 0.002
R12797 S.n7061 S.n7060 0.002
R12798 S.n8072 S.n8071 0.002
R12799 S.n8784 S.n8783 0.002
R12800 S.n9188 S.n9187 0.002
R12801 S.n9865 S.n9864 0.002
R12802 S.n10523 S.n10522 0.002
R12803 S.n11146 S.n11145 0.002
R12804 S.n12893 S.n12891 0.002
R12805 S.n1327 S.n1318 0.002
R12806 S.n3501 S.n3500 0.002
R12807 S.n4023 S.n4022 0.002
R12808 S.n4815 S.n4814 0.002
R12809 S.n5597 S.n5596 0.002
R12810 S.n6357 S.n6356 0.002
R12811 S.n7104 S.n7103 0.002
R12812 S.n8115 S.n8114 0.002
R12813 S.n8827 S.n8826 0.002
R12814 S.n9231 S.n9230 0.002
R12815 S.n9908 S.n9907 0.002
R12816 S.n10566 S.n10565 0.002
R12817 S.n11189 S.n11188 0.002
R12818 S.n12936 S.n12935 0.002
R12819 S.n12591 S.n12572 0.002
R12820 S.n11985 S.n11973 0.002
R12821 S.n11692 S.n11667 0.002
R12822 S.n11433 S.n11421 0.002
R12823 S.n11095 S.n11070 0.002
R12824 S.n10812 S.n10800 0.002
R12825 S.n10470 S.n10445 0.002
R12826 S.n10159 S.n10147 0.002
R12827 S.n9810 S.n9785 0.002
R12828 S.n9483 S.n9471 0.002
R12829 S.n9138 S.n9113 0.002
R12830 S.n8616 S.n8604 0.002
R12831 S.n8443 S.n8418 0.002
R12832 S.n7920 S.n7908 0.002
R12833 S.n7736 S.n7711 0.002
R12834 S.n7367 S.n7355 0.002
R12835 S.n7006 S.n6981 0.002
R12836 S.n6621 S.n6609 0.002
R12837 S.n6264 S.n6239 0.002
R12838 S.n5866 S.n5854 0.002
R12839 S.n5499 S.n5474 0.002
R12840 S.n5085 S.n5073 0.002
R12841 S.n4722 S.n4697 0.002
R12842 S.n4295 S.n4283 0.002
R12843 S.n3922 S.n3897 0.002
R12844 S.n3448 S.n3436 0.002
R12845 S.n3110 S.n3085 0.002
R12846 S.n2592 S.n2580 0.002
R12847 S.n2275 S.n2248 0.002
R12848 S.n1310 S.n1300 0.002
R12849 S.n1785 S.n1770 0.002
R12850 S.n729 S.n716 0.002
R12851 S.n823 S.n815 0.002
R12852 S.n10499 S.n10478 0.002
R12853 S.n10099 S.n10087 0.002
R12854 S.n9724 S.n9699 0.002
R12855 S.n9423 S.n9411 0.002
R12856 S.n9052 S.n9027 0.002
R12857 S.n8556 S.n8544 0.002
R12858 S.n8357 S.n8332 0.002
R12859 S.n7860 S.n7848 0.002
R12860 S.n7650 S.n7625 0.002
R12861 S.n7307 S.n7295 0.002
R12862 S.n6920 S.n6895 0.002
R12863 S.n6561 S.n6549 0.002
R12864 S.n6178 S.n6153 0.002
R12865 S.n5806 S.n5794 0.002
R12866 S.n5413 S.n5388 0.002
R12867 S.n5025 S.n5013 0.002
R12868 S.n4636 S.n4611 0.002
R12869 S.n4235 S.n4223 0.002
R12870 S.n3836 S.n3811 0.002
R12871 S.n3388 S.n3376 0.002
R12872 S.n3024 S.n2999 0.002
R12873 S.n2532 S.n2520 0.002
R12874 S.n2186 S.n2158 0.002
R12875 S.n1252 S.n1241 0.002
R12876 S.t320 S.n1013 0.002
R12877 S.n780 S.n768 0.002
R12878 S.n765 S.n453 0.002
R12879 S.n9164 S.n9146 0.002
R12880 S.n8520 S.n8508 0.002
R12881 S.n8296 S.n8271 0.002
R12882 S.n7824 S.n7812 0.002
R12883 S.n7589 S.n7564 0.002
R12884 S.n7271 S.n7259 0.002
R12885 S.n6859 S.n6834 0.002
R12886 S.n6525 S.n6513 0.002
R12887 S.n6117 S.n6092 0.002
R12888 S.n5770 S.n5758 0.002
R12889 S.n5352 S.n5327 0.002
R12890 S.n4989 S.n4977 0.002
R12891 S.n4575 S.n4550 0.002
R12892 S.n4199 S.n4187 0.002
R12893 S.n3775 S.n3750 0.002
R12894 S.n3352 S.n3340 0.002
R12895 S.n2963 S.n2938 0.002
R12896 S.n2496 S.n2484 0.002
R12897 S.n2122 S.n2095 0.002
R12898 S.n1213 S.n1203 0.002
R12899 S.n1673 S.n1650 0.002
R12900 S.n653 S.n644 0.002
R12901 S.n426 S.n418 0.002
R12902 S.n7762 S.n7744 0.002
R12903 S.n7235 S.n7223 0.002
R12904 S.n6798 S.n6773 0.002
R12905 S.n6489 S.n6477 0.002
R12906 S.n6056 S.n6031 0.002
R12907 S.n5734 S.n5722 0.002
R12908 S.n5291 S.n5266 0.002
R12909 S.n4953 S.n4941 0.002
R12910 S.n4514 S.n4489 0.002
R12911 S.n4163 S.n4151 0.002
R12912 S.n3714 S.n3689 0.002
R12913 S.n3316 S.n3304 0.002
R12914 S.n2902 S.n2877 0.002
R12915 S.n2460 S.n2448 0.002
R12916 S.n2059 S.n2032 0.002
R12917 S.n1179 S.n1169 0.002
R12918 S.n1614 S.n1591 0.002
R12919 S.n620 S.n611 0.002
R12920 S.n385 S.n377 0.002
R12921 S.n6290 S.n6272 0.002
R12922 S.n5698 S.n5686 0.002
R12923 S.n5230 S.n5205 0.002
R12924 S.n4917 S.n4905 0.002
R12925 S.n4453 S.n4428 0.002
R12926 S.n4127 S.n4115 0.002
R12927 S.n3653 S.n3628 0.002
R12928 S.n3280 S.n3268 0.002
R12929 S.n2841 S.n2816 0.002
R12930 S.n2424 S.n2412 0.002
R12931 S.n1996 S.n1969 0.002
R12932 S.n1145 S.n1135 0.002
R12933 S.n1555 S.n1532 0.002
R12934 S.n587 S.n578 0.002
R12935 S.n344 S.n336 0.002
R12936 S.n4748 S.n4730 0.002
R12937 S.n4091 S.n4079 0.002
R12938 S.n3592 S.n3567 0.002
R12939 S.n3244 S.n3232 0.002
R12940 S.n2780 S.n2755 0.002
R12941 S.n2388 S.n2376 0.002
R12942 S.n1933 S.n1906 0.002
R12943 S.n1111 S.n1101 0.002
R12944 S.n1496 S.n1473 0.002
R12945 S.n554 S.n545 0.002
R12946 S.n323 S.n315 0.002
R12947 S.n3136 S.n3118 0.002
R12948 S.n2352 S.n2340 0.002
R12949 S.n1870 S.n1843 0.002
R12950 S.n1077 S.n1067 0.002
R12951 S.n1437 S.n1414 0.002
R12952 S.n521 S.n512 0.002
R12953 S.n282 S.n274 0.002
R12954 S.n1378 S.n1362 0.002
R12955 S.n488 S.n479 0.002
R12956 S.n241 S.n233 0.002
R12957 S.n12663 S.n12655 0.002
R12958 S.n933 S.n930 0.002
R12959 S.n12463 S.n12423 0.001
R12960 S.n12463 S.n12426 0.001
R12961 S.n12463 S.n12429 0.001
R12962 S.n12463 S.n12432 0.001
R12963 S.n12463 S.n12435 0.001
R12964 S.n12463 S.n12438 0.001
R12965 S.n12463 S.n12441 0.001
R12966 S.n12463 S.n12444 0.001
R12967 S.n12463 S.n12447 0.001
R12968 S.n12463 S.n12450 0.001
R12969 S.n12463 S.n12453 0.001
R12970 S.n12463 S.n12456 0.001
R12971 S.n12463 S.n12459 0.001
R12972 S.n12463 S.n12462 0.001
R12973 S.n1017 S.n1016 0.001
R12974 S.n1670 S.n1669 0.001
R12975 S.n1611 S.n1610 0.001
R12976 S.n1552 S.n1551 0.001
R12977 S.n1493 S.n1492 0.001
R12978 S.n1432 S.n1431 0.001
R12979 S.n12309 S.n12308 0.001
R12980 S.n124 S.n123 0.001
R12981 S.t28 S.n124 0.001
R12982 S.n11054 S.n11053 0.001
R12983 S.n10429 S.n10428 0.001
R12984 S.n9769 S.n9768 0.001
R12985 S.n9097 S.n9096 0.001
R12986 S.n8402 S.n8401 0.001
R12987 S.n7695 S.n7694 0.001
R12988 S.n6965 S.n6964 0.001
R12989 S.n6223 S.n6222 0.001
R12990 S.n5458 S.n5457 0.001
R12991 S.n4681 S.n4680 0.001
R12992 S.n3881 S.n3880 0.001
R12993 S.n3069 S.n3068 0.001
R12994 S.n2231 S.n2230 0.001
R12995 S.n1746 S.n1745 0.001
R12996 S.n11033 S.n11032 0.001
R12997 S.n2186 S.n2169 0.001
R12998 S.n9840 S.n9839 0.001
R12999 S.n8473 S.n8472 0.001
R13000 S.n7036 S.n7035 0.001
R13001 S.n5529 S.n5528 0.001
R13002 S.n3952 S.n3951 0.001
R13003 S.n2305 S.n2304 0.001
R13004 S.n12303 S.n12302 0.001
R13005 S.n1782 S.n1781 0.001
R13006 S.n1309 S.n1308 0.001
R13007 S.n2272 S.n2271 0.001
R13008 S.n2589 S.n2588 0.001
R13009 S.n3107 S.n3106 0.001
R13010 S.n3445 S.n3444 0.001
R13011 S.n3919 S.n3918 0.001
R13012 S.n4292 S.n4291 0.001
R13013 S.n4719 S.n4718 0.001
R13014 S.n5082 S.n5081 0.001
R13015 S.n5496 S.n5495 0.001
R13016 S.n5863 S.n5862 0.001
R13017 S.n6261 S.n6260 0.001
R13018 S.n6618 S.n6617 0.001
R13019 S.n7003 S.n7002 0.001
R13020 S.n7364 S.n7363 0.001
R13021 S.n7733 S.n7732 0.001
R13022 S.n7917 S.n7916 0.001
R13023 S.n8440 S.n8439 0.001
R13024 S.n8613 S.n8612 0.001
R13025 S.n9135 S.n9134 0.001
R13026 S.n9480 S.n9479 0.001
R13027 S.n9807 S.n9806 0.001
R13028 S.n10156 S.n10155 0.001
R13029 S.n10467 S.n10466 0.001
R13030 S.n10809 S.n10808 0.001
R13031 S.n11092 S.n11091 0.001
R13032 S.n11430 S.n11429 0.001
R13033 S.n11689 S.n11688 0.001
R13034 S.n11982 S.n11981 0.001
R13035 S.n721 S.n720 0.001
R13036 S.n1240 S.n1239 0.001
R13037 S.n2183 S.n2182 0.001
R13038 S.n2529 S.n2528 0.001
R13039 S.n3021 S.n3020 0.001
R13040 S.n3385 S.n3384 0.001
R13041 S.n3833 S.n3832 0.001
R13042 S.n4232 S.n4231 0.001
R13043 S.n4633 S.n4632 0.001
R13044 S.n5022 S.n5021 0.001
R13045 S.n5410 S.n5409 0.001
R13046 S.n5803 S.n5802 0.001
R13047 S.n6175 S.n6174 0.001
R13048 S.n6558 S.n6557 0.001
R13049 S.n6917 S.n6916 0.001
R13050 S.n7304 S.n7303 0.001
R13051 S.n7647 S.n7646 0.001
R13052 S.n7857 S.n7856 0.001
R13053 S.n8354 S.n8353 0.001
R13054 S.n8553 S.n8552 0.001
R13055 S.n9049 S.n9048 0.001
R13056 S.n9420 S.n9419 0.001
R13057 S.n9721 S.n9720 0.001
R13058 S.n10096 S.n10095 0.001
R13059 S.n1212 S.n1211 0.001
R13060 S.n2119 S.n2118 0.001
R13061 S.n2493 S.n2492 0.001
R13062 S.n2960 S.n2959 0.001
R13063 S.n3349 S.n3348 0.001
R13064 S.n3772 S.n3771 0.001
R13065 S.n4196 S.n4195 0.001
R13066 S.n4572 S.n4571 0.001
R13067 S.n4986 S.n4985 0.001
R13068 S.n5349 S.n5348 0.001
R13069 S.n5767 S.n5766 0.001
R13070 S.n6114 S.n6113 0.001
R13071 S.n6522 S.n6521 0.001
R13072 S.n6856 S.n6855 0.001
R13073 S.n7268 S.n7267 0.001
R13074 S.n7586 S.n7585 0.001
R13075 S.n7821 S.n7820 0.001
R13076 S.n8293 S.n8292 0.001
R13077 S.n8517 S.n8516 0.001
R13078 S.n1178 S.n1177 0.001
R13079 S.n2056 S.n2055 0.001
R13080 S.n2457 S.n2456 0.001
R13081 S.n2899 S.n2898 0.001
R13082 S.n3313 S.n3312 0.001
R13083 S.n3711 S.n3710 0.001
R13084 S.n4160 S.n4159 0.001
R13085 S.n4511 S.n4510 0.001
R13086 S.n4950 S.n4949 0.001
R13087 S.n5288 S.n5287 0.001
R13088 S.n5731 S.n5730 0.001
R13089 S.n6053 S.n6052 0.001
R13090 S.n6486 S.n6485 0.001
R13091 S.n6795 S.n6794 0.001
R13092 S.n7232 S.n7231 0.001
R13093 S.n1144 S.n1143 0.001
R13094 S.n1993 S.n1992 0.001
R13095 S.n2421 S.n2420 0.001
R13096 S.n2838 S.n2837 0.001
R13097 S.n3277 S.n3276 0.001
R13098 S.n3650 S.n3649 0.001
R13099 S.n4124 S.n4123 0.001
R13100 S.n4450 S.n4449 0.001
R13101 S.n4914 S.n4913 0.001
R13102 S.n5227 S.n5226 0.001
R13103 S.n5695 S.n5694 0.001
R13104 S.n1110 S.n1109 0.001
R13105 S.n1930 S.n1929 0.001
R13106 S.n2385 S.n2384 0.001
R13107 S.n2777 S.n2776 0.001
R13108 S.n3241 S.n3240 0.001
R13109 S.n3589 S.n3588 0.001
R13110 S.n4088 S.n4087 0.001
R13111 S.n1076 S.n1075 0.001
R13112 S.n1867 S.n1866 0.001
R13113 S.n2349 S.n2348 0.001
R13114 S.n12463 S.n12392 0.001
R13115 S.n9002 S.n9001 0.001
R13116 S.n8307 S.n8306 0.001
R13117 S.n7600 S.n7599 0.001
R13118 S.n6870 S.n6869 0.001
R13119 S.n6128 S.n6127 0.001
R13120 S.n5363 S.n5362 0.001
R13121 S.n4586 S.n4585 0.001
R13122 S.n3786 S.n3785 0.001
R13123 S.n2974 S.n2973 0.001
R13124 S.n2133 S.n2132 0.001
R13125 S.n1685 S.n1684 0.001
R13126 S.n7539 S.n7538 0.001
R13127 S.n6809 S.n6808 0.001
R13128 S.n6067 S.n6066 0.001
R13129 S.n5302 S.n5301 0.001
R13130 S.n4525 S.n4524 0.001
R13131 S.n3725 S.n3724 0.001
R13132 S.n2913 S.n2912 0.001
R13133 S.n2070 S.n2069 0.001
R13134 S.n1626 S.n1625 0.001
R13135 S.n6006 S.n6005 0.001
R13136 S.n5241 S.n5240 0.001
R13137 S.n4464 S.n4463 0.001
R13138 S.n3664 S.n3663 0.001
R13139 S.n2852 S.n2851 0.001
R13140 S.n2007 S.n2006 0.001
R13141 S.n1567 S.n1566 0.001
R13142 S.n4403 S.n4402 0.001
R13143 S.n3603 S.n3602 0.001
R13144 S.n2791 S.n2790 0.001
R13145 S.n1944 S.n1943 0.001
R13146 S.n1508 S.n1507 0.001
R13147 S.n2730 S.n2729 0.001
R13148 S.n1881 S.n1880 0.001
R13149 S.n1449 S.n1448 0.001
R13150 S.n1390 S.n1389 0.001
R13151 S.n748 S.n738 0.001
R13152 S.n469 S.n468 0.001
R13153 S.n1039 S.n1038 0.001
R13154 S.n2330 S.n2329 0.001
R13155 S.n3204 S.n3203 0.001
R13156 S.n4069 S.n4068 0.001
R13157 S.n4877 S.n4876 0.001
R13158 S.n5676 S.n5675 0.001
R13159 S.n6449 S.n6448 0.001
R13160 S.n7213 S.n7212 0.001
R13161 S.n7784 S.n7783 0.001
R13162 S.n8498 S.n8497 0.001
R13163 S.n9383 S.n9382 0.001
R13164 S.n10077 S.n10076 0.001
R13165 S.n10748 S.n10747 0.001
R13166 S.n11391 S.n11390 0.001
R13167 S.n11962 S.n11961 0.001
R13168 S.n12311 S.n12310 0.001
R13169 S.t28 S.n96 0.001
R13170 S.t28 S.n6 0.001
R13171 S.t28 S.n210 0.001
R13172 S.t28 S.n903 0.001
R13173 S.t28 S.n17 0.001
R13174 S.t28 S.n29 0.001
R13175 S.t28 S.n61 0.001
R13176 S.t28 S.n73 0.001
R13177 S.t28 S.n85 0.001
R13178 S.n977 S.t28 0.001
R13179 S.t28 S.n929 0.001
R13180 S.t28 S.n196 0.001
R13181 S.t28 S.n184 0.001
R13182 S.t28 S.n172 0.001
R13183 S.t28 S.n159 0.001
R13184 S.t28 S.n146 0.001
R13185 S.t28 S.n133 0.001
R13186 S.n120 S.n119 0.001
R13187 S.n9724 S.n9709 0.001
R13188 S.n9052 S.n9037 0.001
R13189 S.n8357 S.n8342 0.001
R13190 S.n7650 S.n7635 0.001
R13191 S.n6920 S.n6905 0.001
R13192 S.n6178 S.n6163 0.001
R13193 S.n5413 S.n5398 0.001
R13194 S.n4636 S.n4621 0.001
R13195 S.n3836 S.n3821 0.001
R13196 S.n3024 S.n3009 0.001
R13197 S.n12549 S.n12546 0.001
R13198 S.n12619 S.n12618 0.001
R13199 S.n9389 S.n9388 0.001
R13200 S.n10754 S.n10753 0.001
R13201 S.n11396 S.n11395 0.001
R13202 S.n11968 S.n11967 0.001
R13203 S.n10082 S.n10081 0.001
R13204 S.n7790 S.n7789 0.001
R13205 S.n8503 S.n8502 0.001
R13206 S.n6455 S.n6454 0.001
R13207 S.n7218 S.n7217 0.001
R13208 S.n4883 S.n4882 0.001
R13209 S.n5681 S.n5680 0.001
R13210 S.n3210 S.n3209 0.001
R13211 S.n4074 S.n4073 0.001
R13212 S.n1045 S.n1044 0.001
R13213 S.n2335 S.n2334 0.001
R13214 S.n474 S.n473 0.001
R13215 S.n119 S.n118 0.001
R13216 S.n10499 S.n10480 0.001
R13217 S.n12891 S.n12890 0.001
R13218 S.n12906 S.n12905 0.001
R13219 S.n12027 S.n12026 0.001
R13220 S.n11737 S.n11736 0.001
R13221 S.n11145 S.n11144 0.001
R13222 S.n11159 S.n11158 0.001
R13223 S.n10522 S.n10521 0.001
R13224 S.n10536 S.n10535 0.001
R13225 S.n9864 S.n9863 0.001
R13226 S.n9878 S.n9877 0.001
R13227 S.n9187 S.n9186 0.001
R13228 S.n9201 S.n9200 0.001
R13229 S.n8783 S.n8782 0.001
R13230 S.n8797 S.n8796 0.001
R13231 S.n8071 S.n8070 0.001
R13232 S.n8085 S.n8084 0.001
R13233 S.n7060 S.n7059 0.001
R13234 S.n7074 S.n7073 0.001
R13235 S.n6313 S.n6312 0.001
R13236 S.n6327 S.n6326 0.001
R13237 S.n5553 S.n5552 0.001
R13238 S.n5567 S.n5566 0.001
R13239 S.n4771 S.n4770 0.001
R13240 S.n4785 S.n4784 0.001
R13241 S.n3976 S.n3975 0.001
R13242 S.n3990 S.n3989 0.001
R13243 S.n3159 S.n3158 0.001
R13244 S.n3173 S.n3172 0.001
R13245 S.n2632 S.n2631 0.001
R13246 S.n2646 S.n2645 0.001
R13247 S.n1346 S.n1345 0.001
R13248 S.n12630 S.n12629 0.001
R13249 S.n12653 S.n12652 0.001
R13250 S.n467 S.n466 0.001
R13251 S.n1037 S.n1036 0.001
R13252 S.n2328 S.n2327 0.001
R13253 S.n3202 S.n3201 0.001
R13254 S.n4067 S.n4066 0.001
R13255 S.n4875 S.n4874 0.001
R13256 S.n5674 S.n5673 0.001
R13257 S.n6447 S.n6446 0.001
R13258 S.n7211 S.n7210 0.001
R13259 S.n7782 S.n7781 0.001
R13260 S.n8496 S.n8495 0.001
R13261 S.n9381 S.n9380 0.001
R13262 S.n10075 S.n10074 0.001
R13263 S.n10746 S.n10745 0.001
R13264 S.n11389 S.n11388 0.001
R13265 S.n11960 S.n11959 0.001
R13266 S.n12612 S.n12611 0.001
R13267 S.t430 S.n474 0.001
R13268 S.t14 S.n12619 0.001
R13269 S.t26 S.n9389 0.001
R13270 S.t16 S.n10082 0.001
R13271 S.t122 S.n10754 0.001
R13272 S.t18 S.n11396 0.001
R13273 S.t2 S.n11968 0.001
R13274 S.t22 S.n7790 0.001
R13275 S.t0 S.n8503 0.001
R13276 S.t8 S.n6455 0.001
R13277 S.t40 S.n7218 0.001
R13278 S.t81 S.n4883 0.001
R13279 S.t460 S.n5681 0.001
R13280 S.t444 S.n3210 0.001
R13281 S.t51 S.n4074 0.001
R13282 S.t142 S.n1045 0.001
R13283 S.t55 S.n2335 0.001
R13284 S.n12546 S.t35 0.001
R13285 S.n12310 S.n12309 0.001
R13286 S.n468 S.n467 0.001
R13287 S.n1038 S.n1037 0.001
R13288 S.n2329 S.n2328 0.001
R13289 S.n3203 S.n3202 0.001
R13290 S.n4068 S.n4067 0.001
R13291 S.n4876 S.n4875 0.001
R13292 S.n5675 S.n5674 0.001
R13293 S.n6448 S.n6447 0.001
R13294 S.n7212 S.n7211 0.001
R13295 S.n7783 S.n7782 0.001
R13296 S.n8497 S.n8496 0.001
R13297 S.n9382 S.n9381 0.001
R13298 S.n10076 S.n10075 0.001
R13299 S.n10747 S.n10746 0.001
R13300 S.n11390 S.n11389 0.001
R13301 S.n11961 S.n11960 0.001
R13302 S.n12614 S.n12608 0.001
R13303 S.n12463 S.n12420 0.001
R13304 S.n11993 S.n11992 0.001
R13305 S.n766 S.n765 0.001
R13306 S.n653 S.n645 0.001
R13307 S.n620 S.n612 0.001
R13308 S.n587 S.n579 0.001
R13309 S.n554 S.n546 0.001
R13310 S.n521 S.n513 0.001
R13311 S.n488 S.n480 0.001
R13312 S.n868 S.n867 0.001
R13313 S.n991 S.n990 0.001
R13314 S.n1835 S.n1834 0.001
R13315 S.n2718 S.n2717 0.001
R13316 S.n3559 S.n3558 0.001
R13317 S.n4391 S.n4390 0.001
R13318 S.n5197 S.n5196 0.001
R13319 S.n5994 S.n5993 0.001
R13320 S.n6765 S.n6764 0.001
R13321 S.n7527 S.n7526 0.001
R13322 S.n8263 S.n8262 0.001
R13323 S.n8990 S.n8989 0.001
R13324 S.n9691 S.n9690 0.001
R13325 S.n10383 S.n10382 0.001
R13326 S.n11042 S.n11041 0.001
R13327 S.n12285 S.n12284 0.001
R13328 S.n13155 S.n13154 0.001
R13329 S.n896 S.n895 0.001
R13330 S.n119 S.n109 0.001
R13331 S.n119 S.n115 0.001
R13332 S.n119 S.n114 0.001
R13333 S.n119 S.n113 0.001
R13334 S.n119 S.n112 0.001
R13335 S.n119 S.n111 0.001
R13336 S.n119 S.n110 0.001
R13337 S.n12635 S.n12634 0.001
R13338 S.n12559 S.n12558 0.001
R13339 S.n11997 S.n11996 0.001
R13340 S.n841 S.n840 0.001
R13341 S.n818 S.n817 0.001
R13342 S.n1777 S.n1776 0.001
R13343 S.n12579 S.n12578 0.001
R13344 S.n11980 S.n11979 0.001
R13345 S.n11683 S.n11682 0.001
R13346 S.n11428 S.n11427 0.001
R13347 S.n11086 S.n11085 0.001
R13348 S.n10807 S.n10806 0.001
R13349 S.n10461 S.n10460 0.001
R13350 S.n10154 S.n10153 0.001
R13351 S.n9801 S.n9800 0.001
R13352 S.n9478 S.n9477 0.001
R13353 S.n9129 S.n9128 0.001
R13354 S.n8611 S.n8610 0.001
R13355 S.n8434 S.n8433 0.001
R13356 S.n7915 S.n7914 0.001
R13357 S.n7727 S.n7726 0.001
R13358 S.n7362 S.n7361 0.001
R13359 S.n6997 S.n6996 0.001
R13360 S.n6616 S.n6615 0.001
R13361 S.n6255 S.n6254 0.001
R13362 S.n5861 S.n5860 0.001
R13363 S.n5490 S.n5489 0.001
R13364 S.n5080 S.n5079 0.001
R13365 S.n4713 S.n4712 0.001
R13366 S.n4290 S.n4289 0.001
R13367 S.n3913 S.n3912 0.001
R13368 S.n3443 S.n3442 0.001
R13369 S.n3101 S.n3100 0.001
R13370 S.n2587 S.n2586 0.001
R13371 S.n2264 S.n2263 0.001
R13372 S.n1307 S.n1306 0.001
R13373 S.n724 S.n723 0.001
R13374 S.n421 S.n420 0.001
R13375 S.n1666 S.n1665 0.001
R13376 S.n9153 S.n9152 0.001
R13377 S.n8515 S.n8514 0.001
R13378 S.n8287 S.n8286 0.001
R13379 S.n7819 S.n7818 0.001
R13380 S.n7580 S.n7579 0.001
R13381 S.n7266 S.n7265 0.001
R13382 S.n6850 S.n6849 0.001
R13383 S.n6520 S.n6519 0.001
R13384 S.n6108 S.n6107 0.001
R13385 S.n5765 S.n5764 0.001
R13386 S.n5343 S.n5342 0.001
R13387 S.n4984 S.n4983 0.001
R13388 S.n4566 S.n4565 0.001
R13389 S.n4194 S.n4193 0.001
R13390 S.n3766 S.n3765 0.001
R13391 S.n3347 S.n3346 0.001
R13392 S.n2954 S.n2953 0.001
R13393 S.n2491 S.n2490 0.001
R13394 S.n2111 S.n2110 0.001
R13395 S.n1210 S.n1209 0.001
R13396 S.n441 S.n440 0.001
R13397 S.n9829 S.n9828 0.001
R13398 S.n9399 S.n9398 0.001
R13399 S.n9006 S.n9005 0.001
R13400 S.n8532 S.n8531 0.001
R13401 S.n8311 S.n8310 0.001
R13402 S.n7836 S.n7835 0.001
R13403 S.n7604 S.n7603 0.001
R13404 S.n7283 S.n7282 0.001
R13405 S.n6874 S.n6873 0.001
R13406 S.n6537 S.n6536 0.001
R13407 S.n6132 S.n6131 0.001
R13408 S.n5782 S.n5781 0.001
R13409 S.n5367 S.n5366 0.001
R13410 S.n5001 S.n5000 0.001
R13411 S.n4590 S.n4589 0.001
R13412 S.n4211 S.n4210 0.001
R13413 S.n3790 S.n3789 0.001
R13414 S.n3364 S.n3363 0.001
R13415 S.n2978 S.n2977 0.001
R13416 S.n2508 S.n2507 0.001
R13417 S.n2137 S.n2136 0.001
R13418 S.n1225 S.n1224 0.001
R13419 S.n1244 S.n1243 0.001
R13420 S.n456 S.n455 0.001
R13421 S.n771 S.n770 0.001
R13422 S.n2175 S.n2174 0.001
R13423 S.n3015 S.n3014 0.001
R13424 S.n3827 S.n3826 0.001
R13425 S.n4627 S.n4626 0.001
R13426 S.n5404 S.n5403 0.001
R13427 S.n6169 S.n6168 0.001
R13428 S.n6911 S.n6910 0.001
R13429 S.n7641 S.n7640 0.001
R13430 S.n8348 S.n8347 0.001
R13431 S.n9043 S.n9042 0.001
R13432 S.n9715 S.n9714 0.001
R13433 S.n10488 S.n10487 0.001
R13434 S.n10094 S.n10093 0.001
R13435 S.n9418 S.n9417 0.001
R13436 S.n8551 S.n8550 0.001
R13437 S.n7855 S.n7854 0.001
R13438 S.n7302 S.n7301 0.001
R13439 S.n6556 S.n6555 0.001
R13440 S.n5801 S.n5800 0.001
R13441 S.n5020 S.n5019 0.001
R13442 S.n4230 S.n4229 0.001
R13443 S.n3383 S.n3382 0.001
R13444 S.n2527 S.n2526 0.001
R13445 S.n1722 S.n1721 0.001
R13446 S.n681 S.n680 0.001
R13447 S.n226 S.n225 0.001
R13448 S.n11117 S.n11116 0.001
R13449 S.n10771 S.n10770 0.001
R13450 S.n10406 S.n10405 0.001
R13451 S.n10118 S.n10117 0.001
R13452 S.n9746 S.n9745 0.001
R13453 S.n9442 S.n9441 0.001
R13454 S.n9074 S.n9073 0.001
R13455 S.n8575 S.n8574 0.001
R13456 S.n8379 S.n8378 0.001
R13457 S.n7879 S.n7878 0.001
R13458 S.n7672 S.n7671 0.001
R13459 S.n7326 S.n7325 0.001
R13460 S.n6942 S.n6941 0.001
R13461 S.n6580 S.n6579 0.001
R13462 S.n6200 S.n6199 0.001
R13463 S.n5825 S.n5824 0.001
R13464 S.n5435 S.n5434 0.001
R13465 S.n5044 S.n5043 0.001
R13466 S.n4658 S.n4657 0.001
R13467 S.n4254 S.n4253 0.001
R13468 S.n3858 S.n3857 0.001
R13469 S.n3407 S.n3406 0.001
R13470 S.n3046 S.n3045 0.001
R13471 S.n2551 S.n2550 0.001
R13472 S.n2208 S.n2207 0.001
R13473 S.n1271 S.n1270 0.001
R13474 S.n1750 S.n1749 0.001
R13475 S.n701 S.n700 0.001
R13476 S.n1290 S.n1289 0.001
R13477 S.n2235 S.n2234 0.001
R13478 S.n2565 S.n2564 0.001
R13479 S.n3073 S.n3072 0.001
R13480 S.n3421 S.n3420 0.001
R13481 S.n3885 S.n3884 0.001
R13482 S.n4268 S.n4267 0.001
R13483 S.n4685 S.n4684 0.001
R13484 S.n5058 S.n5057 0.001
R13485 S.n5462 S.n5461 0.001
R13486 S.n5839 S.n5838 0.001
R13487 S.n6227 S.n6226 0.001
R13488 S.n6594 S.n6593 0.001
R13489 S.n6969 S.n6968 0.001
R13490 S.n7340 S.n7339 0.001
R13491 S.n7699 S.n7698 0.001
R13492 S.n7893 S.n7892 0.001
R13493 S.n8406 S.n8405 0.001
R13494 S.n8589 S.n8588 0.001
R13495 S.n9101 S.n9100 0.001
R13496 S.n9456 S.n9455 0.001
R13497 S.n9773 S.n9772 0.001
R13498 S.n10132 S.n10131 0.001
R13499 S.n10433 S.n10432 0.001
R13500 S.n10785 S.n10784 0.001
R13501 S.n11058 S.n11057 0.001
R13502 S.n11406 S.n11405 0.001
R13503 S.n11712 S.n11711 0.001
R13504 S.n791 S.n790 0.001
R13505 S.n1688 S.n1687 0.001
R13506 S.n665 S.n664 0.001
R13507 S.n648 S.n647 0.001
R13508 S.n380 S.n379 0.001
R13509 S.n1607 S.n1606 0.001
R13510 S.n7751 S.n7750 0.001
R13511 S.n7230 S.n7229 0.001
R13512 S.n6789 S.n6788 0.001
R13513 S.n6484 S.n6483 0.001
R13514 S.n6047 S.n6046 0.001
R13515 S.n5729 S.n5728 0.001
R13516 S.n5282 S.n5281 0.001
R13517 S.n4948 S.n4947 0.001
R13518 S.n4505 S.n4504 0.001
R13519 S.n4158 S.n4157 0.001
R13520 S.n3705 S.n3704 0.001
R13521 S.n3311 S.n3310 0.001
R13522 S.n2893 S.n2892 0.001
R13523 S.n2455 S.n2454 0.001
R13524 S.n2048 S.n2047 0.001
R13525 S.n1176 S.n1175 0.001
R13526 S.n400 S.n399 0.001
R13527 S.n8462 S.n8461 0.001
R13528 S.n7800 S.n7799 0.001
R13529 S.n7543 S.n7542 0.001
R13530 S.n7247 S.n7246 0.001
R13531 S.n6813 S.n6812 0.001
R13532 S.n6501 S.n6500 0.001
R13533 S.n6071 S.n6070 0.001
R13534 S.n5746 S.n5745 0.001
R13535 S.n5306 S.n5305 0.001
R13536 S.n4965 S.n4964 0.001
R13537 S.n4529 S.n4528 0.001
R13538 S.n4175 S.n4174 0.001
R13539 S.n3729 S.n3728 0.001
R13540 S.n3328 S.n3327 0.001
R13541 S.n2917 S.n2916 0.001
R13542 S.n2472 S.n2471 0.001
R13543 S.n2074 S.n2073 0.001
R13544 S.n1191 S.n1190 0.001
R13545 S.n1629 S.n1628 0.001
R13546 S.n632 S.n631 0.001
R13547 S.n615 S.n614 0.001
R13548 S.n339 S.n338 0.001
R13549 S.n1548 S.n1547 0.001
R13550 S.n6279 S.n6278 0.001
R13551 S.n5693 S.n5692 0.001
R13552 S.n5221 S.n5220 0.001
R13553 S.n4912 S.n4911 0.001
R13554 S.n4444 S.n4443 0.001
R13555 S.n4122 S.n4121 0.001
R13556 S.n3644 S.n3643 0.001
R13557 S.n3275 S.n3274 0.001
R13558 S.n2832 S.n2831 0.001
R13559 S.n2419 S.n2418 0.001
R13560 S.n1985 S.n1984 0.001
R13561 S.n1142 S.n1141 0.001
R13562 S.n359 S.n358 0.001
R13563 S.n7025 S.n7024 0.001
R13564 S.n6465 S.n6464 0.001
R13565 S.n6010 S.n6009 0.001
R13566 S.n5710 S.n5709 0.001
R13567 S.n5245 S.n5244 0.001
R13568 S.n4929 S.n4928 0.001
R13569 S.n4468 S.n4467 0.001
R13570 S.n4139 S.n4138 0.001
R13571 S.n3668 S.n3667 0.001
R13572 S.n3292 S.n3291 0.001
R13573 S.n2856 S.n2855 0.001
R13574 S.n2436 S.n2435 0.001
R13575 S.n2011 S.n2010 0.001
R13576 S.n1157 S.n1156 0.001
R13577 S.n1570 S.n1569 0.001
R13578 S.n599 S.n598 0.001
R13579 S.n582 S.n581 0.001
R13580 S.n318 S.n317 0.001
R13581 S.n1489 S.n1488 0.001
R13582 S.n4737 S.n4736 0.001
R13583 S.n4086 S.n4085 0.001
R13584 S.n3583 S.n3582 0.001
R13585 S.n3239 S.n3238 0.001
R13586 S.n2771 S.n2770 0.001
R13587 S.n2383 S.n2382 0.001
R13588 S.n1922 S.n1921 0.001
R13589 S.n1108 S.n1107 0.001
R13590 S.n48 S.n47 0.001
R13591 S.n5518 S.n5517 0.001
R13592 S.n4893 S.n4892 0.001
R13593 S.n4407 S.n4406 0.001
R13594 S.n4103 S.n4102 0.001
R13595 S.n3607 S.n3606 0.001
R13596 S.n3256 S.n3255 0.001
R13597 S.n2795 S.n2794 0.001
R13598 S.n2400 S.n2399 0.001
R13599 S.n1948 S.n1947 0.001
R13600 S.n1123 S.n1122 0.001
R13601 S.n1511 S.n1510 0.001
R13602 S.n566 S.n565 0.001
R13603 S.n549 S.n548 0.001
R13604 S.n277 S.n276 0.001
R13605 S.n1430 S.n1429 0.001
R13606 S.n3125 S.n3124 0.001
R13607 S.n2347 S.n2346 0.001
R13608 S.n1859 S.n1858 0.001
R13609 S.n1074 S.n1073 0.001
R13610 S.n297 S.n296 0.001
R13611 S.n3941 S.n3940 0.001
R13612 S.n3220 S.n3219 0.001
R13613 S.n2734 S.n2733 0.001
R13614 S.n2364 S.n2363 0.001
R13615 S.n1885 S.n1884 0.001
R13616 S.n1089 S.n1088 0.001
R13617 S.n1452 S.n1451 0.001
R13618 S.n533 S.n532 0.001
R13619 S.n516 S.n515 0.001
R13620 S.n236 S.n235 0.001
R13621 S.n1369 S.n1368 0.001
R13622 S.n256 S.n255 0.001
R13623 S.n2294 S.n2293 0.001
R13624 S.n1055 S.n1054 0.001
R13625 S.n1393 S.n1392 0.001
R13626 S.n500 S.n499 0.001
R13627 S.n483 S.n482 0.001
R13628 S.n741 S.n740 0.001
R13629 S.n1350 S.n1349 0.001
R13630 S.n1027 S.n1026 0.001
R13631 S.n2637 S.n2636 0.001
R13632 S.n2316 S.n2315 0.001
R13633 S.n3164 S.n3163 0.001
R13634 S.n3146 S.n3145 0.001
R13635 S.n3981 S.n3980 0.001
R13636 S.n3963 S.n3962 0.001
R13637 S.n4776 S.n4775 0.001
R13638 S.n4758 S.n4757 0.001
R13639 S.n5558 S.n5557 0.001
R13640 S.n5540 S.n5539 0.001
R13641 S.n6318 S.n6317 0.001
R13642 S.n6300 S.n6299 0.001
R13643 S.n7065 S.n7064 0.001
R13644 S.n7047 S.n7046 0.001
R13645 S.n8076 S.n8075 0.001
R13646 S.n7772 S.n7771 0.001
R13647 S.n8788 S.n8787 0.001
R13648 S.n8484 S.n8483 0.001
R13649 S.n9192 S.n9191 0.001
R13650 S.n9174 S.n9173 0.001
R13651 S.n9869 S.n9868 0.001
R13652 S.n9851 S.n9850 0.001
R13653 S.n10527 S.n10526 0.001
R13654 S.n10509 S.n10508 0.001
R13655 S.n11150 S.n11149 0.001
R13656 S.n11132 S.n11131 0.001
R13657 S.n11728 S.n11727 0.001
R13658 S.n12020 S.n12019 0.001
R13659 S.n12897 S.n12896 0.001
R13660 S.n12601 S.n12600 0.001
R13661 S.n1322 S.n1321 0.001
R13662 S.n2660 S.n2659 0.001
R13663 S.n12934 S.n12933 0.001
R13664 S.n12920 S.n12919 0.001
R13665 S.n12041 S.n12040 0.001
R13666 S.n11751 S.n11750 0.001
R13667 S.n11187 S.n11186 0.001
R13668 S.n11173 S.n11172 0.001
R13669 S.n10564 S.n10563 0.001
R13670 S.n10550 S.n10549 0.001
R13671 S.n9906 S.n9905 0.001
R13672 S.n9892 S.n9891 0.001
R13673 S.n9229 S.n9228 0.001
R13674 S.n9215 S.n9214 0.001
R13675 S.n8825 S.n8824 0.001
R13676 S.n8811 S.n8810 0.001
R13677 S.n8113 S.n8112 0.001
R13678 S.n8099 S.n8098 0.001
R13679 S.n7102 S.n7101 0.001
R13680 S.n7088 S.n7087 0.001
R13681 S.n6355 S.n6354 0.001
R13682 S.n6341 S.n6340 0.001
R13683 S.n5595 S.n5594 0.001
R13684 S.n5581 S.n5580 0.001
R13685 S.n4813 S.n4812 0.001
R13686 S.n4799 S.n4798 0.001
R13687 S.n4021 S.n4020 0.001
R13688 S.n4007 S.n4006 0.001
R13689 S.n3499 S.n3498 0.001
R13690 S.n3187 S.n3186 0.001
R13691 S.n2674 S.n2673 0.001
R13692 S.n2604 S.n2603 0.001
R13693 S.n3516 S.n3515 0.001
R13694 S.n12678 S.n12677 0.001
R13695 S.n12951 S.n12950 0.001
R13696 S.n12056 S.n12055 0.001
R13697 S.n11767 S.n11766 0.001
R13698 S.n11448 S.n11447 0.001
R13699 S.n11204 S.n11203 0.001
R13700 S.n10827 S.n10826 0.001
R13701 S.n10581 S.n10580 0.001
R13702 S.n10174 S.n10173 0.001
R13703 S.n9923 S.n9922 0.001
R13704 S.n9498 S.n9497 0.001
R13705 S.n9246 S.n9245 0.001
R13706 S.n8631 S.n8630 0.001
R13707 S.n8842 S.n8841 0.001
R13708 S.n7935 S.n7934 0.001
R13709 S.n8130 S.n8129 0.001
R13710 S.n7382 S.n7381 0.001
R13711 S.n7119 S.n7118 0.001
R13712 S.n6636 S.n6635 0.001
R13713 S.n6372 S.n6371 0.001
R13714 S.n5881 S.n5880 0.001
R13715 S.n5612 S.n5611 0.001
R13716 S.n5100 S.n5099 0.001
R13717 S.n4830 S.n4829 0.001
R13718 S.n4310 S.n4309 0.001
R13719 S.n4035 S.n4034 0.001
R13720 S.n3463 S.n3462 0.001
R13721 S.n3475 S.n3474 0.001
R13722 S.n4050 S.n4049 0.001
R13723 S.n12694 S.n12693 0.001
R13724 S.n12966 S.n12965 0.001
R13725 S.n12072 S.n12071 0.001
R13726 S.n11782 S.n11781 0.001
R13727 S.n11464 S.n11463 0.001
R13728 S.n11219 S.n11218 0.001
R13729 S.n10843 S.n10842 0.001
R13730 S.n10596 S.n10595 0.001
R13731 S.n10190 S.n10189 0.001
R13732 S.n9938 S.n9937 0.001
R13733 S.n9514 S.n9513 0.001
R13734 S.n9261 S.n9260 0.001
R13735 S.n8647 S.n8646 0.001
R13736 S.n8857 S.n8856 0.001
R13737 S.n7951 S.n7950 0.001
R13738 S.n8145 S.n8144 0.001
R13739 S.n7398 S.n7397 0.001
R13740 S.n7134 S.n7133 0.001
R13741 S.n6652 S.n6651 0.001
R13742 S.n6387 S.n6386 0.001
R13743 S.n5897 S.n5896 0.001
R13744 S.n5627 S.n5626 0.001
R13745 S.n5116 S.n5115 0.001
R13746 S.n4845 S.n4844 0.001
R13747 S.n4347 S.n4346 0.001
R13748 S.n4323 S.n4322 0.001
R13749 S.n4860 S.n4859 0.001
R13750 S.n12710 S.n12709 0.001
R13751 S.n12981 S.n12980 0.001
R13752 S.n12088 S.n12087 0.001
R13753 S.n11797 S.n11796 0.001
R13754 S.n11480 S.n11479 0.001
R13755 S.n11234 S.n11233 0.001
R13756 S.n10859 S.n10858 0.001
R13757 S.n10611 S.n10610 0.001
R13758 S.n10206 S.n10205 0.001
R13759 S.n9953 S.n9952 0.001
R13760 S.n9530 S.n9529 0.001
R13761 S.n9276 S.n9275 0.001
R13762 S.n8663 S.n8662 0.001
R13763 S.n8872 S.n8871 0.001
R13764 S.n7967 S.n7966 0.001
R13765 S.n8160 S.n8159 0.001
R13766 S.n7414 S.n7413 0.001
R13767 S.n7149 S.n7148 0.001
R13768 S.n6668 S.n6667 0.001
R13769 S.n6402 S.n6401 0.001
R13770 S.n5913 S.n5912 0.001
R13771 S.n5642 S.n5641 0.001
R13772 S.n5153 S.n5152 0.001
R13773 S.n5129 S.n5128 0.001
R13774 S.n5657 S.n5656 0.001
R13775 S.n12726 S.n12725 0.001
R13776 S.n12996 S.n12995 0.001
R13777 S.n12104 S.n12103 0.001
R13778 S.n11812 S.n11811 0.001
R13779 S.n11496 S.n11495 0.001
R13780 S.n11249 S.n11248 0.001
R13781 S.n10875 S.n10874 0.001
R13782 S.n10626 S.n10625 0.001
R13783 S.n10222 S.n10221 0.001
R13784 S.n9968 S.n9967 0.001
R13785 S.n9546 S.n9545 0.001
R13786 S.n9291 S.n9290 0.001
R13787 S.n8679 S.n8678 0.001
R13788 S.n8887 S.n8886 0.001
R13789 S.n7983 S.n7982 0.001
R13790 S.n8175 S.n8174 0.001
R13791 S.n7430 S.n7429 0.001
R13792 S.n7164 S.n7163 0.001
R13793 S.n6684 S.n6683 0.001
R13794 S.n6417 S.n6416 0.001
R13795 S.n5950 S.n5949 0.001
R13796 S.n5926 S.n5925 0.001
R13797 S.n6432 S.n6431 0.001
R13798 S.n12742 S.n12741 0.001
R13799 S.n13011 S.n13010 0.001
R13800 S.n12120 S.n12119 0.001
R13801 S.n11827 S.n11826 0.001
R13802 S.n11512 S.n11511 0.001
R13803 S.n11264 S.n11263 0.001
R13804 S.n10891 S.n10890 0.001
R13805 S.n10641 S.n10640 0.001
R13806 S.n10238 S.n10237 0.001
R13807 S.n9983 S.n9982 0.001
R13808 S.n9562 S.n9561 0.001
R13809 S.n9306 S.n9305 0.001
R13810 S.n8695 S.n8694 0.001
R13811 S.n8902 S.n8901 0.001
R13812 S.n7999 S.n7998 0.001
R13813 S.n8190 S.n8189 0.001
R13814 S.n7446 S.n7445 0.001
R13815 S.n7179 S.n7178 0.001
R13816 S.n6721 S.n6720 0.001
R13817 S.n6697 S.n6696 0.001
R13818 S.n7194 S.n7193 0.001
R13819 S.n12758 S.n12757 0.001
R13820 S.n13026 S.n13025 0.001
R13821 S.n12136 S.n12135 0.001
R13822 S.n11842 S.n11841 0.001
R13823 S.n11528 S.n11527 0.001
R13824 S.n11279 S.n11278 0.001
R13825 S.n10907 S.n10906 0.001
R13826 S.n10656 S.n10655 0.001
R13827 S.n10254 S.n10253 0.001
R13828 S.n9998 S.n9997 0.001
R13829 S.n9578 S.n9577 0.001
R13830 S.n9321 S.n9320 0.001
R13831 S.n8711 S.n8710 0.001
R13832 S.n8917 S.n8916 0.001
R13833 S.n8015 S.n8014 0.001
R13834 S.n8205 S.n8204 0.001
R13835 S.n7483 S.n7482 0.001
R13836 S.n7459 S.n7458 0.001
R13837 S.n8220 S.n8219 0.001
R13838 S.n12774 S.n12773 0.001
R13839 S.n13041 S.n13040 0.001
R13840 S.n12152 S.n12151 0.001
R13841 S.n11857 S.n11856 0.001
R13842 S.n11544 S.n11543 0.001
R13843 S.n11294 S.n11293 0.001
R13844 S.n10923 S.n10922 0.001
R13845 S.n10671 S.n10670 0.001
R13846 S.n10270 S.n10269 0.001
R13847 S.n10013 S.n10012 0.001
R13848 S.n9594 S.n9593 0.001
R13849 S.n9336 S.n9335 0.001
R13850 S.n8727 S.n8726 0.001
R13851 S.n8932 S.n8931 0.001
R13852 S.n8031 S.n8030 0.001
R13853 S.n8043 S.n8042 0.001
R13854 S.n8947 S.n8946 0.001
R13855 S.n12790 S.n12789 0.001
R13856 S.n13056 S.n13055 0.001
R13857 S.n12168 S.n12167 0.001
R13858 S.n11872 S.n11871 0.001
R13859 S.n11560 S.n11559 0.001
R13860 S.n11309 S.n11308 0.001
R13861 S.n10939 S.n10938 0.001
R13862 S.n10686 S.n10685 0.001
R13863 S.n10286 S.n10285 0.001
R13864 S.n10028 S.n10027 0.001
R13865 S.n9610 S.n9609 0.001
R13866 S.n9351 S.n9350 0.001
R13867 S.n8743 S.n8742 0.001
R13868 S.n8755 S.n8754 0.001
R13869 S.n9366 S.n9365 0.001
R13870 S.n12806 S.n12805 0.001
R13871 S.n13071 S.n13070 0.001
R13872 S.n12184 S.n12183 0.001
R13873 S.n11887 S.n11886 0.001
R13874 S.n11576 S.n11575 0.001
R13875 S.n11324 S.n11323 0.001
R13876 S.n10955 S.n10954 0.001
R13877 S.n10701 S.n10700 0.001
R13878 S.n10302 S.n10301 0.001
R13879 S.n10043 S.n10042 0.001
R13880 S.n9647 S.n9646 0.001
R13881 S.n9623 S.n9622 0.001
R13882 S.n10058 S.n10057 0.001
R13883 S.n12822 S.n12821 0.001
R13884 S.n13086 S.n13085 0.001
R13885 S.n12200 S.n12199 0.001
R13886 S.n11902 S.n11901 0.001
R13887 S.n11592 S.n11591 0.001
R13888 S.n11339 S.n11338 0.001
R13889 S.n10971 S.n10970 0.001
R13890 S.n10716 S.n10715 0.001
R13891 S.n10339 S.n10338 0.001
R13892 S.n10315 S.n10314 0.001
R13893 S.n10731 S.n10730 0.001
R13894 S.n12838 S.n12837 0.001
R13895 S.n13101 S.n13100 0.001
R13896 S.n12216 S.n12215 0.001
R13897 S.n11917 S.n11916 0.001
R13898 S.n11608 S.n11607 0.001
R13899 S.n11354 S.n11353 0.001
R13900 S.n11008 S.n11007 0.001
R13901 S.n10984 S.n10983 0.001
R13902 S.n11369 S.n11368 0.001
R13903 S.n12854 S.n12853 0.001
R13904 S.n13116 S.n13115 0.001
R13905 S.n12232 S.n12231 0.001
R13906 S.n11932 S.n11931 0.001
R13907 S.n11648 S.n11647 0.001
R13908 S.n11619 S.n11618 0.001
R13909 S.n12259 S.n12258 0.001
R13910 S.n12867 S.n12866 0.001
R13911 S.n13130 S.n13129 0.001
R13912 S.n11948 S.n11947 0.001
R13913 S.n12658 S.n12657 0.001
R13914 S.n12423 S.n12422 0.001
R13915 S.n12426 S.n12425 0.001
R13916 S.n12429 S.n12428 0.001
R13917 S.n12432 S.n12431 0.001
R13918 S.n12435 S.n12434 0.001
R13919 S.n12438 S.n12437 0.001
R13920 S.n12441 S.n12440 0.001
R13921 S.n12444 S.n12443 0.001
R13922 S.n12447 S.n12446 0.001
R13923 S.n12450 S.n12449 0.001
R13924 S.n12453 S.n12452 0.001
R13925 S.n12456 S.n12455 0.001
R13926 S.n12459 S.n12458 0.001
R13927 S.n12462 S.n12461 0.001
R13928 S.n119 S.n117 0.001
R13929 S.n12616 S.n12615 0.001
R13930 S.n11964 S.n11963 0.001
R13931 S.n11393 S.n11392 0.001
R13932 S.n10750 S.n10749 0.001
R13933 S.n10079 S.n10078 0.001
R13934 S.n9385 S.n9384 0.001
R13935 S.n8500 S.n8499 0.001
R13936 S.n7786 S.n7785 0.001
R13937 S.n7215 S.n7214 0.001
R13938 S.n6451 S.n6450 0.001
R13939 S.n5678 S.n5677 0.001
R13940 S.n4879 S.n4878 0.001
R13941 S.n4071 S.n4070 0.001
R13942 S.n3206 S.n3205 0.001
R13943 S.n2332 S.n2331 0.001
R13944 S.n1041 S.n1040 0.001
R13945 S.n471 S.n470 0.001
R13946 S.t14 S.n12646 0.001
R13947 S.t14 S.n12643 0.001
R13948 S.n12643 S.n12640 0.001
R13949 S.t72 S.n12570 0.001
R13950 S.t72 S.n12567 0.001
R13951 S.n12567 S.n12564 0.001
R13952 S.t2 S.n12015 0.001
R13953 S.t2 S.n12012 0.001
R13954 S.n12012 S.n12009 0.001
R13955 S.n12274 S.t44 0.001
R13956 S.n12306 S.n12276 0.001
R13957 S.t116 S.n854 0.001
R13958 S.t116 S.n857 0.001
R13959 S.t116 S.n829 0.001
R13960 S.t116 S.n826 0.001
R13961 S.n826 S.n823 0.001
R13962 S.t320 S.n1791 0.001
R13963 S.t320 S.n1788 0.001
R13964 S.n1788 S.n1785 0.001
R13965 S.t72 S.n12594 0.001
R13966 S.t72 S.n12597 0.001
R13967 S.t2 S.n11991 0.001
R13968 S.t2 S.n11988 0.001
R13969 S.n11988 S.n11985 0.001
R13970 S.t44 S.n11698 0.001
R13971 S.t44 S.n11695 0.001
R13972 S.n11695 S.n11692 0.001
R13973 S.t18 S.n11439 0.001
R13974 S.t18 S.n11436 0.001
R13975 S.n11436 S.n11433 0.001
R13976 S.t12 S.n11101 0.001
R13977 S.t12 S.n11098 0.001
R13978 S.n11098 S.n11095 0.001
R13979 S.t122 S.n10818 0.001
R13980 S.t122 S.n10815 0.001
R13981 S.n10815 S.n10812 0.001
R13982 S.t103 S.n10476 0.001
R13983 S.t103 S.n10473 0.001
R13984 S.n10473 S.n10470 0.001
R13985 S.t16 S.n10165 0.001
R13986 S.t16 S.n10162 0.001
R13987 S.n10162 S.n10159 0.001
R13988 S.t86 S.n9816 0.001
R13989 S.t86 S.n9813 0.001
R13990 S.n9813 S.n9810 0.001
R13991 S.t26 S.n9489 0.001
R13992 S.t26 S.n9486 0.001
R13993 S.n9486 S.n9483 0.001
R13994 S.t24 S.n9144 0.001
R13995 S.t24 S.n9141 0.001
R13996 S.n9141 S.n9138 0.001
R13997 S.t0 S.n8622 0.001
R13998 S.t0 S.n8619 0.001
R13999 S.n8619 S.n8616 0.001
R14000 S.t131 S.n8449 0.001
R14001 S.t131 S.n8446 0.001
R14002 S.n8446 S.n8443 0.001
R14003 S.t22 S.n7926 0.001
R14004 S.t22 S.n7923 0.001
R14005 S.n7923 S.n7920 0.001
R14006 S.t59 S.n7742 0.001
R14007 S.t59 S.n7739 0.001
R14008 S.n7739 S.n7736 0.001
R14009 S.t40 S.n7373 0.001
R14010 S.t40 S.n7370 0.001
R14011 S.n7370 S.n7367 0.001
R14012 S.t37 S.n7012 0.001
R14013 S.t37 S.n7009 0.001
R14014 S.n7009 S.n7006 0.001
R14015 S.t8 S.n6627 0.001
R14016 S.t8 S.n6624 0.001
R14017 S.n6624 S.n6621 0.001
R14018 S.t119 S.n6270 0.001
R14019 S.t119 S.n6267 0.001
R14020 S.n6267 S.n6264 0.001
R14021 S.t460 S.n5872 0.001
R14022 S.t460 S.n5869 0.001
R14023 S.n5869 S.n5866 0.001
R14024 S.t390 S.n5505 0.001
R14025 S.t390 S.n5502 0.001
R14026 S.n5502 S.n5499 0.001
R14027 S.t81 S.n5091 0.001
R14028 S.t81 S.n5088 0.001
R14029 S.n5088 S.n5085 0.001
R14030 S.t360 S.n4728 0.001
R14031 S.t360 S.n4725 0.001
R14032 S.n4725 S.n4722 0.001
R14033 S.t51 S.n4301 0.001
R14034 S.t51 S.n4298 0.001
R14035 S.n4298 S.n4295 0.001
R14036 S.t109 S.n3928 0.001
R14037 S.t109 S.n3925 0.001
R14038 S.n3925 S.n3922 0.001
R14039 S.t444 S.n3454 0.001
R14040 S.t444 S.n3451 0.001
R14041 S.n3451 S.n3448 0.001
R14042 S.t240 S.n3116 0.001
R14043 S.t240 S.n3113 0.001
R14044 S.n3113 S.n3110 0.001
R14045 S.t55 S.n2598 0.001
R14046 S.t55 S.n2595 0.001
R14047 S.n2595 S.n2592 0.001
R14048 S.t200 S.n2281 0.001
R14049 S.t200 S.n2278 0.001
R14050 S.n2278 S.n2275 0.001
R14051 S.t142 S.n1316 0.001
R14052 S.t142 S.n1313 0.001
R14053 S.n1313 S.n1310 0.001
R14054 S.t430 S.n735 0.001
R14055 S.t430 S.n732 0.001
R14056 S.n732 S.n729 0.001
R14057 S.t116 S.n432 0.001
R14058 S.t116 S.n429 0.001
R14059 S.n429 S.n426 0.001
R14060 S.t320 S.n1679 0.001
R14061 S.t320 S.n1676 0.001
R14062 S.n1676 S.n1673 0.001
R14063 S.t24 S.n9167 0.001
R14064 S.t24 S.n9170 0.001
R14065 S.t0 S.n8526 0.001
R14066 S.t0 S.n8523 0.001
R14067 S.n8523 S.n8520 0.001
R14068 S.t131 S.n8302 0.001
R14069 S.t131 S.n8299 0.001
R14070 S.n8299 S.n8296 0.001
R14071 S.t22 S.n7830 0.001
R14072 S.t22 S.n7827 0.001
R14073 S.n7827 S.n7824 0.001
R14074 S.t59 S.n7595 0.001
R14075 S.t59 S.n7592 0.001
R14076 S.n7592 S.n7589 0.001
R14077 S.t40 S.n7277 0.001
R14078 S.t40 S.n7274 0.001
R14079 S.n7274 S.n7271 0.001
R14080 S.t37 S.n6865 0.001
R14081 S.t37 S.n6862 0.001
R14082 S.n6862 S.n6859 0.001
R14083 S.t8 S.n6531 0.001
R14084 S.t8 S.n6528 0.001
R14085 S.n6528 S.n6525 0.001
R14086 S.t119 S.n6123 0.001
R14087 S.t119 S.n6120 0.001
R14088 S.n6120 S.n6117 0.001
R14089 S.t460 S.n5776 0.001
R14090 S.t460 S.n5773 0.001
R14091 S.n5773 S.n5770 0.001
R14092 S.t390 S.n5358 0.001
R14093 S.t390 S.n5355 0.001
R14094 S.n5355 S.n5352 0.001
R14095 S.t81 S.n4995 0.001
R14096 S.t81 S.n4992 0.001
R14097 S.n4992 S.n4989 0.001
R14098 S.t360 S.n4581 0.001
R14099 S.t360 S.n4578 0.001
R14100 S.n4578 S.n4575 0.001
R14101 S.t51 S.n4205 0.001
R14102 S.t51 S.n4202 0.001
R14103 S.n4202 S.n4199 0.001
R14104 S.t109 S.n3781 0.001
R14105 S.t109 S.n3778 0.001
R14106 S.n3778 S.n3775 0.001
R14107 S.t444 S.n3358 0.001
R14108 S.t444 S.n3355 0.001
R14109 S.n3355 S.n3352 0.001
R14110 S.t240 S.n2969 0.001
R14111 S.t240 S.n2966 0.001
R14112 S.n2966 S.n2963 0.001
R14113 S.t55 S.n2502 0.001
R14114 S.t55 S.n2499 0.001
R14115 S.n2499 S.n2496 0.001
R14116 S.t200 S.n2128 0.001
R14117 S.t200 S.n2125 0.001
R14118 S.n2125 S.n2122 0.001
R14119 S.t142 S.n1219 0.001
R14120 S.t142 S.n1216 0.001
R14121 S.n1216 S.n1213 0.001
R14122 S.t116 S.n452 0.001
R14123 S.t116 S.n449 0.001
R14124 S.n449 S.n446 0.001
R14125 S.t86 S.n9844 0.001
R14126 S.t86 S.n9847 0.001
R14127 S.t26 S.n9410 0.001
R14128 S.t26 S.n9407 0.001
R14129 S.n9407 S.n9404 0.001
R14130 S.t24 S.n9026 0.001
R14131 S.t24 S.n9023 0.001
R14132 S.n9023 S.n9020 0.001
R14133 S.t0 S.n8543 0.001
R14134 S.t0 S.n8540 0.001
R14135 S.n8540 S.n8537 0.001
R14136 S.t131 S.n8331 0.001
R14137 S.t131 S.n8328 0.001
R14138 S.n8328 S.n8325 0.001
R14139 S.t22 S.n7847 0.001
R14140 S.t22 S.n7844 0.001
R14141 S.n7844 S.n7841 0.001
R14142 S.t59 S.n7624 0.001
R14143 S.t59 S.n7621 0.001
R14144 S.n7621 S.n7618 0.001
R14145 S.t40 S.n7294 0.001
R14146 S.t40 S.n7291 0.001
R14147 S.n7291 S.n7288 0.001
R14148 S.t37 S.n6894 0.001
R14149 S.t37 S.n6891 0.001
R14150 S.n6891 S.n6888 0.001
R14151 S.t8 S.n6548 0.001
R14152 S.t8 S.n6545 0.001
R14153 S.n6545 S.n6542 0.001
R14154 S.t119 S.n6152 0.001
R14155 S.t119 S.n6149 0.001
R14156 S.n6149 S.n6146 0.001
R14157 S.t460 S.n5793 0.001
R14158 S.t460 S.n5790 0.001
R14159 S.n5790 S.n5787 0.001
R14160 S.t390 S.n5387 0.001
R14161 S.t390 S.n5384 0.001
R14162 S.n5384 S.n5381 0.001
R14163 S.t81 S.n5012 0.001
R14164 S.t81 S.n5009 0.001
R14165 S.n5009 S.n5006 0.001
R14166 S.t360 S.n4610 0.001
R14167 S.t360 S.n4607 0.001
R14168 S.n4607 S.n4604 0.001
R14169 S.t51 S.n4222 0.001
R14170 S.t51 S.n4219 0.001
R14171 S.n4219 S.n4216 0.001
R14172 S.t109 S.n3810 0.001
R14173 S.t109 S.n3807 0.001
R14174 S.n3807 S.n3804 0.001
R14175 S.t444 S.n3375 0.001
R14176 S.t444 S.n3372 0.001
R14177 S.n3372 S.n3369 0.001
R14178 S.t240 S.n2998 0.001
R14179 S.t240 S.n2995 0.001
R14180 S.n2995 S.n2992 0.001
R14181 S.t55 S.n2519 0.001
R14182 S.t55 S.n2516 0.001
R14183 S.n2516 S.n2513 0.001
R14184 S.t200 S.n2157 0.001
R14185 S.t200 S.n2154 0.001
R14186 S.n2154 S.n2151 0.001
R14187 S.t142 S.n1238 0.001
R14188 S.t142 S.n1235 0.001
R14189 S.n1235 S.n1232 0.001
R14190 S.t142 S.n1258 0.001
R14191 S.t142 S.n1255 0.001
R14192 S.n1255 S.n1252 0.001
R14193 S.n757 S.t430 0.001
R14194 S.n765 S.n760 0.001
R14195 S.t116 S.n786 0.001
R14196 S.t116 S.n783 0.001
R14197 S.n783 S.n780 0.001
R14198 S.t200 S.n2192 0.001
R14199 S.t200 S.n2189 0.001
R14200 S.n2189 S.n2186 0.001
R14201 S.t240 S.n3030 0.001
R14202 S.t240 S.n3027 0.001
R14203 S.n3027 S.n3024 0.001
R14204 S.t109 S.n3842 0.001
R14205 S.t109 S.n3839 0.001
R14206 S.n3839 S.n3836 0.001
R14207 S.t360 S.n4642 0.001
R14208 S.t360 S.n4639 0.001
R14209 S.n4639 S.n4636 0.001
R14210 S.t390 S.n5419 0.001
R14211 S.t390 S.n5416 0.001
R14212 S.n5416 S.n5413 0.001
R14213 S.t119 S.n6184 0.001
R14214 S.t119 S.n6181 0.001
R14215 S.n6181 S.n6178 0.001
R14216 S.t37 S.n6926 0.001
R14217 S.t37 S.n6923 0.001
R14218 S.n6923 S.n6920 0.001
R14219 S.t59 S.n7656 0.001
R14220 S.t59 S.n7653 0.001
R14221 S.n7653 S.n7650 0.001
R14222 S.t131 S.n8363 0.001
R14223 S.t131 S.n8360 0.001
R14224 S.n8360 S.n8357 0.001
R14225 S.t24 S.n9058 0.001
R14226 S.t24 S.n9055 0.001
R14227 S.n9055 S.n9052 0.001
R14228 S.t86 S.n9730 0.001
R14229 S.t86 S.n9727 0.001
R14230 S.n9727 S.n9724 0.001
R14231 S.t103 S.n10502 0.001
R14232 S.t103 S.n10505 0.001
R14233 S.t16 S.n10105 0.001
R14234 S.t16 S.n10102 0.001
R14235 S.n10102 S.n10099 0.001
R14236 S.t26 S.n9429 0.001
R14237 S.t26 S.n9426 0.001
R14238 S.n9426 S.n9423 0.001
R14239 S.t0 S.n8562 0.001
R14240 S.t0 S.n8559 0.001
R14241 S.n8559 S.n8556 0.001
R14242 S.t22 S.n7866 0.001
R14243 S.t22 S.n7863 0.001
R14244 S.n7863 S.n7860 0.001
R14245 S.t40 S.n7313 0.001
R14246 S.t40 S.n7310 0.001
R14247 S.n7310 S.n7307 0.001
R14248 S.t8 S.n6567 0.001
R14249 S.t8 S.n6564 0.001
R14250 S.n6564 S.n6561 0.001
R14251 S.t460 S.n5812 0.001
R14252 S.t460 S.n5809 0.001
R14253 S.n5809 S.n5806 0.001
R14254 S.t81 S.n5031 0.001
R14255 S.t81 S.n5028 0.001
R14256 S.n5028 S.n5025 0.001
R14257 S.t51 S.n4241 0.001
R14258 S.t51 S.n4238 0.001
R14259 S.n4238 S.n4235 0.001
R14260 S.t444 S.n3394 0.001
R14261 S.t444 S.n3391 0.001
R14262 S.n3391 S.n3388 0.001
R14263 S.t55 S.n2538 0.001
R14264 S.t55 S.n2535 0.001
R14265 S.n2535 S.n2532 0.001
R14266 S.t320 S.n1741 0.001
R14267 S.t320 S.n1738 0.001
R14268 S.n1738 S.n1735 0.001
R14269 S.t430 S.n696 0.001
R14270 S.t430 S.n693 0.001
R14271 S.n693 S.n690 0.001
R14272 S.n888 S.t116 0.001
R14273 S.n901 S.n891 0.001
R14274 S.t12 S.n11125 0.001
R14275 S.t12 S.n11128 0.001
R14276 S.t122 S.n10779 0.001
R14277 S.t122 S.n10776 0.001
R14278 S.n10776 S.n10773 0.001
R14279 S.t103 S.n10424 0.001
R14280 S.t103 S.n10421 0.001
R14281 S.n10421 S.n10418 0.001
R14282 S.t16 S.n10126 0.001
R14283 S.t16 S.n10123 0.001
R14284 S.n10123 S.n10120 0.001
R14285 S.t86 S.n9764 0.001
R14286 S.t86 S.n9761 0.001
R14287 S.n9761 S.n9758 0.001
R14288 S.t26 S.n9450 0.001
R14289 S.t26 S.n9447 0.001
R14290 S.n9447 S.n9444 0.001
R14291 S.t24 S.n9092 0.001
R14292 S.t24 S.n9089 0.001
R14293 S.n9089 S.n9086 0.001
R14294 S.t0 S.n8583 0.001
R14295 S.t0 S.n8580 0.001
R14296 S.n8580 S.n8577 0.001
R14297 S.t131 S.n8397 0.001
R14298 S.t131 S.n8394 0.001
R14299 S.n8394 S.n8391 0.001
R14300 S.t22 S.n7887 0.001
R14301 S.t22 S.n7884 0.001
R14302 S.n7884 S.n7881 0.001
R14303 S.t59 S.n7690 0.001
R14304 S.t59 S.n7687 0.001
R14305 S.n7687 S.n7684 0.001
R14306 S.t40 S.n7334 0.001
R14307 S.t40 S.n7331 0.001
R14308 S.n7331 S.n7328 0.001
R14309 S.t37 S.n6960 0.001
R14310 S.t37 S.n6957 0.001
R14311 S.n6957 S.n6954 0.001
R14312 S.t8 S.n6588 0.001
R14313 S.t8 S.n6585 0.001
R14314 S.n6585 S.n6582 0.001
R14315 S.t119 S.n6218 0.001
R14316 S.t119 S.n6215 0.001
R14317 S.n6215 S.n6212 0.001
R14318 S.t460 S.n5833 0.001
R14319 S.t460 S.n5830 0.001
R14320 S.n5830 S.n5827 0.001
R14321 S.t390 S.n5453 0.001
R14322 S.t390 S.n5450 0.001
R14323 S.n5450 S.n5447 0.001
R14324 S.t81 S.n5052 0.001
R14325 S.t81 S.n5049 0.001
R14326 S.n5049 S.n5046 0.001
R14327 S.t360 S.n4676 0.001
R14328 S.t360 S.n4673 0.001
R14329 S.n4673 S.n4670 0.001
R14330 S.t51 S.n4262 0.001
R14331 S.t51 S.n4259 0.001
R14332 S.n4259 S.n4256 0.001
R14333 S.t109 S.n3876 0.001
R14334 S.t109 S.n3873 0.001
R14335 S.n3873 S.n3870 0.001
R14336 S.t444 S.n3415 0.001
R14337 S.t444 S.n3412 0.001
R14338 S.n3412 S.n3409 0.001
R14339 S.t240 S.n3064 0.001
R14340 S.t240 S.n3061 0.001
R14341 S.n3061 S.n3058 0.001
R14342 S.t55 S.n2559 0.001
R14343 S.t55 S.n2556 0.001
R14344 S.n2556 S.n2553 0.001
R14345 S.t200 S.n2226 0.001
R14346 S.t200 S.n2223 0.001
R14347 S.n2223 S.n2220 0.001
R14348 S.t142 S.n1279 0.001
R14349 S.t142 S.n1276 0.001
R14350 S.n1276 S.n1273 0.001
R14351 S.t320 S.n1769 0.001
R14352 S.t320 S.n1766 0.001
R14353 S.n1766 S.n1763 0.001
R14354 S.t430 S.n715 0.001
R14355 S.t430 S.n712 0.001
R14356 S.n712 S.n709 0.001
R14357 S.t142 S.n1299 0.001
R14358 S.t142 S.n1296 0.001
R14359 S.n1296 S.n1293 0.001
R14360 S.t200 S.n2247 0.001
R14361 S.t200 S.n2244 0.001
R14362 S.n2244 S.n2241 0.001
R14363 S.t55 S.n2579 0.001
R14364 S.t55 S.n2576 0.001
R14365 S.n2576 S.n2573 0.001
R14366 S.t240 S.n3084 0.001
R14367 S.t240 S.n3081 0.001
R14368 S.n3081 S.n3078 0.001
R14369 S.t444 S.n3435 0.001
R14370 S.t444 S.n3432 0.001
R14371 S.n3432 S.n3429 0.001
R14372 S.t109 S.n3896 0.001
R14373 S.t109 S.n3893 0.001
R14374 S.n3893 S.n3890 0.001
R14375 S.t51 S.n4282 0.001
R14376 S.t51 S.n4279 0.001
R14377 S.n4279 S.n4276 0.001
R14378 S.t360 S.n4696 0.001
R14379 S.t360 S.n4693 0.001
R14380 S.n4693 S.n4690 0.001
R14381 S.t81 S.n5072 0.001
R14382 S.t81 S.n5069 0.001
R14383 S.n5069 S.n5066 0.001
R14384 S.t390 S.n5473 0.001
R14385 S.t390 S.n5470 0.001
R14386 S.n5470 S.n5467 0.001
R14387 S.t460 S.n5853 0.001
R14388 S.t460 S.n5850 0.001
R14389 S.n5850 S.n5847 0.001
R14390 S.t119 S.n6238 0.001
R14391 S.t119 S.n6235 0.001
R14392 S.n6235 S.n6232 0.001
R14393 S.t8 S.n6608 0.001
R14394 S.t8 S.n6605 0.001
R14395 S.n6605 S.n6602 0.001
R14396 S.t37 S.n6980 0.001
R14397 S.t37 S.n6977 0.001
R14398 S.n6977 S.n6974 0.001
R14399 S.t40 S.n7354 0.001
R14400 S.t40 S.n7351 0.001
R14401 S.n7351 S.n7348 0.001
R14402 S.t59 S.n7710 0.001
R14403 S.t59 S.n7707 0.001
R14404 S.n7707 S.n7704 0.001
R14405 S.t22 S.n7907 0.001
R14406 S.t22 S.n7904 0.001
R14407 S.n7904 S.n7901 0.001
R14408 S.t131 S.n8417 0.001
R14409 S.t131 S.n8414 0.001
R14410 S.n8414 S.n8411 0.001
R14411 S.t0 S.n8603 0.001
R14412 S.t0 S.n8600 0.001
R14413 S.n8600 S.n8597 0.001
R14414 S.t24 S.n9112 0.001
R14415 S.t24 S.n9109 0.001
R14416 S.n9109 S.n9106 0.001
R14417 S.t26 S.n9470 0.001
R14418 S.t26 S.n9467 0.001
R14419 S.n9467 S.n9464 0.001
R14420 S.t86 S.n9784 0.001
R14421 S.t86 S.n9781 0.001
R14422 S.n9781 S.n9778 0.001
R14423 S.t16 S.n10146 0.001
R14424 S.t16 S.n10143 0.001
R14425 S.n10143 S.n10140 0.001
R14426 S.t103 S.n10444 0.001
R14427 S.t103 S.n10441 0.001
R14428 S.n10441 S.n10438 0.001
R14429 S.t122 S.n10799 0.001
R14430 S.t122 S.n10796 0.001
R14431 S.n10796 S.n10793 0.001
R14432 S.t12 S.n11069 0.001
R14433 S.t12 S.n11066 0.001
R14434 S.n11066 S.n11063 0.001
R14435 S.t18 S.n11420 0.001
R14436 S.t18 S.n11417 0.001
R14437 S.n11417 S.n11414 0.001
R14438 S.t44 S.n11720 0.001
R14439 S.t44 S.n11723 0.001
R14440 S.t116 S.n808 0.001
R14441 S.t116 S.n805 0.001
R14442 S.n805 S.n802 0.001
R14443 S.t320 S.n1707 0.001
R14444 S.t320 S.n1704 0.001
R14445 S.n1704 S.n1701 0.001
R14446 S.t430 S.n676 0.001
R14447 S.t430 S.n673 0.001
R14448 S.n673 S.n670 0.001
R14449 S.t430 S.n659 0.001
R14450 S.t430 S.n656 0.001
R14451 S.n656 S.n653 0.001
R14452 S.t116 S.n391 0.001
R14453 S.t116 S.n388 0.001
R14454 S.n388 S.n385 0.001
R14455 S.t320 S.n1620 0.001
R14456 S.t320 S.n1617 0.001
R14457 S.n1617 S.n1614 0.001
R14458 S.t59 S.n7765 0.001
R14459 S.t59 S.n7768 0.001
R14460 S.t40 S.n7241 0.001
R14461 S.t40 S.n7238 0.001
R14462 S.n7238 S.n7235 0.001
R14463 S.t37 S.n6804 0.001
R14464 S.t37 S.n6801 0.001
R14465 S.n6801 S.n6798 0.001
R14466 S.t8 S.n6495 0.001
R14467 S.t8 S.n6492 0.001
R14468 S.n6492 S.n6489 0.001
R14469 S.t119 S.n6062 0.001
R14470 S.t119 S.n6059 0.001
R14471 S.n6059 S.n6056 0.001
R14472 S.t460 S.n5740 0.001
R14473 S.t460 S.n5737 0.001
R14474 S.n5737 S.n5734 0.001
R14475 S.t390 S.n5297 0.001
R14476 S.t390 S.n5294 0.001
R14477 S.n5294 S.n5291 0.001
R14478 S.t81 S.n4959 0.001
R14479 S.t81 S.n4956 0.001
R14480 S.n4956 S.n4953 0.001
R14481 S.t360 S.n4520 0.001
R14482 S.t360 S.n4517 0.001
R14483 S.n4517 S.n4514 0.001
R14484 S.t51 S.n4169 0.001
R14485 S.t51 S.n4166 0.001
R14486 S.n4166 S.n4163 0.001
R14487 S.t109 S.n3720 0.001
R14488 S.t109 S.n3717 0.001
R14489 S.n3717 S.n3714 0.001
R14490 S.t444 S.n3322 0.001
R14491 S.t444 S.n3319 0.001
R14492 S.n3319 S.n3316 0.001
R14493 S.t240 S.n2908 0.001
R14494 S.t240 S.n2905 0.001
R14495 S.n2905 S.n2902 0.001
R14496 S.t55 S.n2466 0.001
R14497 S.t55 S.n2463 0.001
R14498 S.n2463 S.n2460 0.001
R14499 S.t200 S.n2065 0.001
R14500 S.t200 S.n2062 0.001
R14501 S.n2062 S.n2059 0.001
R14502 S.t142 S.n1185 0.001
R14503 S.t142 S.n1182 0.001
R14504 S.n1182 S.n1179 0.001
R14505 S.t116 S.n411 0.001
R14506 S.t116 S.n408 0.001
R14507 S.n408 S.n405 0.001
R14508 S.t131 S.n8477 0.001
R14509 S.t131 S.n8480 0.001
R14510 S.t22 S.n7811 0.001
R14511 S.t22 S.n7808 0.001
R14512 S.n7808 S.n7805 0.001
R14513 S.t59 S.n7563 0.001
R14514 S.t59 S.n7560 0.001
R14515 S.n7560 S.n7557 0.001
R14516 S.t40 S.n7258 0.001
R14517 S.t40 S.n7255 0.001
R14518 S.n7255 S.n7252 0.001
R14519 S.t37 S.n6833 0.001
R14520 S.t37 S.n6830 0.001
R14521 S.n6830 S.n6827 0.001
R14522 S.t8 S.n6512 0.001
R14523 S.t8 S.n6509 0.001
R14524 S.n6509 S.n6506 0.001
R14525 S.t119 S.n6091 0.001
R14526 S.t119 S.n6088 0.001
R14527 S.n6088 S.n6085 0.001
R14528 S.t460 S.n5757 0.001
R14529 S.t460 S.n5754 0.001
R14530 S.n5754 S.n5751 0.001
R14531 S.t390 S.n5326 0.001
R14532 S.t390 S.n5323 0.001
R14533 S.n5323 S.n5320 0.001
R14534 S.t81 S.n4976 0.001
R14535 S.t81 S.n4973 0.001
R14536 S.n4973 S.n4970 0.001
R14537 S.t360 S.n4549 0.001
R14538 S.t360 S.n4546 0.001
R14539 S.n4546 S.n4543 0.001
R14540 S.t51 S.n4186 0.001
R14541 S.t51 S.n4183 0.001
R14542 S.n4183 S.n4180 0.001
R14543 S.t109 S.n3749 0.001
R14544 S.t109 S.n3746 0.001
R14545 S.n3746 S.n3743 0.001
R14546 S.t444 S.n3339 0.001
R14547 S.t444 S.n3336 0.001
R14548 S.n3336 S.n3333 0.001
R14549 S.t240 S.n2937 0.001
R14550 S.t240 S.n2934 0.001
R14551 S.n2934 S.n2931 0.001
R14552 S.t55 S.n2483 0.001
R14553 S.t55 S.n2480 0.001
R14554 S.n2480 S.n2477 0.001
R14555 S.t200 S.n2094 0.001
R14556 S.t200 S.n2091 0.001
R14557 S.n2091 S.n2088 0.001
R14558 S.t142 S.n1202 0.001
R14559 S.t142 S.n1199 0.001
R14560 S.n1199 S.n1196 0.001
R14561 S.t320 S.n1649 0.001
R14562 S.t320 S.n1646 0.001
R14563 S.n1646 S.n1643 0.001
R14564 S.t430 S.n643 0.001
R14565 S.t430 S.n640 0.001
R14566 S.n640 S.n637 0.001
R14567 S.t430 S.n626 0.001
R14568 S.t430 S.n623 0.001
R14569 S.n623 S.n620 0.001
R14570 S.t116 S.n350 0.001
R14571 S.t116 S.n347 0.001
R14572 S.n347 S.n344 0.001
R14573 S.t320 S.n1561 0.001
R14574 S.t320 S.n1558 0.001
R14575 S.n1558 S.n1555 0.001
R14576 S.t119 S.n6293 0.001
R14577 S.t119 S.n6296 0.001
R14578 S.t460 S.n5704 0.001
R14579 S.t460 S.n5701 0.001
R14580 S.n5701 S.n5698 0.001
R14581 S.t390 S.n5236 0.001
R14582 S.t390 S.n5233 0.001
R14583 S.n5233 S.n5230 0.001
R14584 S.t81 S.n4923 0.001
R14585 S.t81 S.n4920 0.001
R14586 S.n4920 S.n4917 0.001
R14587 S.t360 S.n4459 0.001
R14588 S.t360 S.n4456 0.001
R14589 S.n4456 S.n4453 0.001
R14590 S.t51 S.n4133 0.001
R14591 S.t51 S.n4130 0.001
R14592 S.n4130 S.n4127 0.001
R14593 S.t109 S.n3659 0.001
R14594 S.t109 S.n3656 0.001
R14595 S.n3656 S.n3653 0.001
R14596 S.t444 S.n3286 0.001
R14597 S.t444 S.n3283 0.001
R14598 S.n3283 S.n3280 0.001
R14599 S.t240 S.n2847 0.001
R14600 S.t240 S.n2844 0.001
R14601 S.n2844 S.n2841 0.001
R14602 S.t55 S.n2430 0.001
R14603 S.t55 S.n2427 0.001
R14604 S.n2427 S.n2424 0.001
R14605 S.t200 S.n2002 0.001
R14606 S.t200 S.n1999 0.001
R14607 S.n1999 S.n1996 0.001
R14608 S.t142 S.n1151 0.001
R14609 S.t142 S.n1148 0.001
R14610 S.n1148 S.n1145 0.001
R14611 S.t116 S.n370 0.001
R14612 S.t116 S.n367 0.001
R14613 S.n367 S.n364 0.001
R14614 S.t37 S.n7040 0.001
R14615 S.t37 S.n7043 0.001
R14616 S.t8 S.n6476 0.001
R14617 S.t8 S.n6473 0.001
R14618 S.n6473 S.n6470 0.001
R14619 S.t119 S.n6030 0.001
R14620 S.t119 S.n6027 0.001
R14621 S.n6027 S.n6024 0.001
R14622 S.t460 S.n5721 0.001
R14623 S.t460 S.n5718 0.001
R14624 S.n5718 S.n5715 0.001
R14625 S.t390 S.n5265 0.001
R14626 S.t390 S.n5262 0.001
R14627 S.n5262 S.n5259 0.001
R14628 S.t81 S.n4940 0.001
R14629 S.t81 S.n4937 0.001
R14630 S.n4937 S.n4934 0.001
R14631 S.t360 S.n4488 0.001
R14632 S.t360 S.n4485 0.001
R14633 S.n4485 S.n4482 0.001
R14634 S.t51 S.n4150 0.001
R14635 S.t51 S.n4147 0.001
R14636 S.n4147 S.n4144 0.001
R14637 S.t109 S.n3688 0.001
R14638 S.t109 S.n3685 0.001
R14639 S.n3685 S.n3682 0.001
R14640 S.t444 S.n3303 0.001
R14641 S.t444 S.n3300 0.001
R14642 S.n3300 S.n3297 0.001
R14643 S.t240 S.n2876 0.001
R14644 S.t240 S.n2873 0.001
R14645 S.n2873 S.n2870 0.001
R14646 S.t55 S.n2447 0.001
R14647 S.t55 S.n2444 0.001
R14648 S.n2444 S.n2441 0.001
R14649 S.t200 S.n2031 0.001
R14650 S.t200 S.n2028 0.001
R14651 S.n2028 S.n2025 0.001
R14652 S.t142 S.n1168 0.001
R14653 S.t142 S.n1165 0.001
R14654 S.n1165 S.n1162 0.001
R14655 S.t320 S.n1590 0.001
R14656 S.t320 S.n1587 0.001
R14657 S.n1587 S.n1584 0.001
R14658 S.t430 S.n610 0.001
R14659 S.t430 S.n607 0.001
R14660 S.n607 S.n604 0.001
R14661 S.t430 S.n593 0.001
R14662 S.t430 S.n590 0.001
R14663 S.n590 S.n587 0.001
R14664 S.t116 S.n329 0.001
R14665 S.t116 S.n326 0.001
R14666 S.n326 S.n323 0.001
R14667 S.t320 S.n1502 0.001
R14668 S.t320 S.n1499 0.001
R14669 S.n1499 S.n1496 0.001
R14670 S.t360 S.n4751 0.001
R14671 S.t360 S.n4754 0.001
R14672 S.t51 S.n4097 0.001
R14673 S.t51 S.n4094 0.001
R14674 S.n4094 S.n4091 0.001
R14675 S.t109 S.n3598 0.001
R14676 S.t109 S.n3595 0.001
R14677 S.n3595 S.n3592 0.001
R14678 S.t444 S.n3250 0.001
R14679 S.t444 S.n3247 0.001
R14680 S.n3247 S.n3244 0.001
R14681 S.t240 S.n2786 0.001
R14682 S.t240 S.n2783 0.001
R14683 S.n2783 S.n2780 0.001
R14684 S.t55 S.n2394 0.001
R14685 S.t55 S.n2391 0.001
R14686 S.n2391 S.n2388 0.001
R14687 S.t200 S.n1939 0.001
R14688 S.t200 S.n1936 0.001
R14689 S.n1936 S.n1933 0.001
R14690 S.t142 S.n1117 0.001
R14691 S.t142 S.n1114 0.001
R14692 S.n1114 S.n1111 0.001
R14693 S.n59 S.n54 0.001
R14694 S.t390 S.n5533 0.001
R14695 S.t390 S.n5536 0.001
R14696 S.t81 S.n4904 0.001
R14697 S.t81 S.n4901 0.001
R14698 S.n4901 S.n4898 0.001
R14699 S.t360 S.n4427 0.001
R14700 S.t360 S.n4424 0.001
R14701 S.n4424 S.n4421 0.001
R14702 S.t51 S.n4114 0.001
R14703 S.t51 S.n4111 0.001
R14704 S.n4111 S.n4108 0.001
R14705 S.t109 S.n3627 0.001
R14706 S.t109 S.n3624 0.001
R14707 S.n3624 S.n3621 0.001
R14708 S.t444 S.n3267 0.001
R14709 S.t444 S.n3264 0.001
R14710 S.n3264 S.n3261 0.001
R14711 S.t240 S.n2815 0.001
R14712 S.t240 S.n2812 0.001
R14713 S.n2812 S.n2809 0.001
R14714 S.t55 S.n2411 0.001
R14715 S.t55 S.n2408 0.001
R14716 S.n2408 S.n2405 0.001
R14717 S.t200 S.n1968 0.001
R14718 S.t200 S.n1965 0.001
R14719 S.n1965 S.n1962 0.001
R14720 S.t142 S.n1134 0.001
R14721 S.t142 S.n1131 0.001
R14722 S.n1131 S.n1128 0.001
R14723 S.t320 S.n1531 0.001
R14724 S.t320 S.n1528 0.001
R14725 S.n1528 S.n1525 0.001
R14726 S.t430 S.n577 0.001
R14727 S.t430 S.n574 0.001
R14728 S.n574 S.n571 0.001
R14729 S.t430 S.n560 0.001
R14730 S.t430 S.n557 0.001
R14731 S.n557 S.n554 0.001
R14732 S.t116 S.n288 0.001
R14733 S.t116 S.n285 0.001
R14734 S.n285 S.n282 0.001
R14735 S.t320 S.n1443 0.001
R14736 S.t320 S.n1440 0.001
R14737 S.n1440 S.n1437 0.001
R14738 S.t240 S.n3139 0.001
R14739 S.t240 S.n3142 0.001
R14740 S.t55 S.n2358 0.001
R14741 S.t55 S.n2355 0.001
R14742 S.n2355 S.n2352 0.001
R14743 S.t200 S.n1876 0.001
R14744 S.t200 S.n1873 0.001
R14745 S.n1873 S.n1870 0.001
R14746 S.t142 S.n1083 0.001
R14747 S.t142 S.n1080 0.001
R14748 S.n1080 S.n1077 0.001
R14749 S.t116 S.n308 0.001
R14750 S.t116 S.n305 0.001
R14751 S.n305 S.n302 0.001
R14752 S.t109 S.n3956 0.001
R14753 S.t109 S.n3959 0.001
R14754 S.t444 S.n3231 0.001
R14755 S.t444 S.n3228 0.001
R14756 S.n3228 S.n3225 0.001
R14757 S.t240 S.n2754 0.001
R14758 S.t240 S.n2751 0.001
R14759 S.n2751 S.n2748 0.001
R14760 S.t55 S.n2375 0.001
R14761 S.t55 S.n2372 0.001
R14762 S.n2372 S.n2369 0.001
R14763 S.t200 S.n1905 0.001
R14764 S.t200 S.n1902 0.001
R14765 S.n1902 S.n1899 0.001
R14766 S.t142 S.n1100 0.001
R14767 S.t142 S.n1097 0.001
R14768 S.n1097 S.n1094 0.001
R14769 S.t320 S.n1472 0.001
R14770 S.n1469 S.n1455 0.001
R14771 S.t430 S.n544 0.001
R14772 S.t430 S.n541 0.001
R14773 S.n541 S.n538 0.001
R14774 S.t430 S.n527 0.001
R14775 S.t430 S.n524 0.001
R14776 S.n524 S.n521 0.001
R14777 S.t116 S.n247 0.001
R14778 S.t116 S.n244 0.001
R14779 S.n244 S.n241 0.001
R14780 S.t320 S.n1384 0.001
R14781 S.t320 S.n1381 0.001
R14782 S.n1381 S.n1378 0.001
R14783 S.t116 S.n267 0.001
R14784 S.t116 S.n264 0.001
R14785 S.n264 S.n261 0.001
R14786 S.t200 S.n2309 0.001
R14787 S.t200 S.n2312 0.001
R14788 S.t142 S.n1066 0.001
R14789 S.t142 S.n1063 0.001
R14790 S.n1063 S.n1060 0.001
R14791 S.t320 S.n1413 0.001
R14792 S.t320 S.n1410 0.001
R14793 S.n1410 S.n1407 0.001
R14794 S.t430 S.n511 0.001
R14795 S.t430 S.n508 0.001
R14796 S.n508 S.n505 0.001
R14797 S.t430 S.n494 0.001
R14798 S.t430 S.n491 0.001
R14799 S.n491 S.n488 0.001
R14800 S.t116 S.n883 0.001
R14801 S.t116 S.n885 0.001
R14802 S.t430 S.n751 0.001
R14803 S.t430 S.n754 0.001
R14804 S.t320 S.n1361 0.001
R14805 S.t320 S.n1358 0.001
R14806 S.n1358 S.n1355 0.001
R14807 S.n1336 S.t142 0.001
R14808 S.n1346 S.n1339 0.001
R14809 S.t200 S.n2649 0.001
R14810 S.t200 S.n2652 0.001
R14811 S.n2622 S.t55 0.001
R14812 S.n2632 S.n2625 0.001
R14813 S.t240 S.n3176 0.001
R14814 S.t240 S.n3179 0.001
R14815 S.n3159 S.n3152 0.001
R14816 S.t109 S.n3993 0.001
R14817 S.t109 S.n3996 0.001
R14818 S.n3976 S.n3969 0.001
R14819 S.t360 S.n4788 0.001
R14820 S.t360 S.n4791 0.001
R14821 S.n4771 S.n4764 0.001
R14822 S.t390 S.n5570 0.001
R14823 S.t390 S.n5573 0.001
R14824 S.n5553 S.n5546 0.001
R14825 S.t119 S.n6330 0.001
R14826 S.t119 S.n6333 0.001
R14827 S.n6313 S.n6306 0.001
R14828 S.t37 S.n7077 0.001
R14829 S.t37 S.n7080 0.001
R14830 S.n7060 S.n7053 0.001
R14831 S.t59 S.n8088 0.001
R14832 S.t59 S.n8091 0.001
R14833 S.n8061 S.t22 0.001
R14834 S.n8071 S.n8064 0.001
R14835 S.t131 S.n8800 0.001
R14836 S.t131 S.n8803 0.001
R14837 S.n8773 S.t0 0.001
R14838 S.n8783 S.n8776 0.001
R14839 S.t24 S.n9204 0.001
R14840 S.t24 S.n9207 0.001
R14841 S.n9187 S.n9180 0.001
R14842 S.t86 S.n9881 0.001
R14843 S.t86 S.n9884 0.001
R14844 S.n9864 S.n9857 0.001
R14845 S.t103 S.n10539 0.001
R14846 S.t103 S.n10542 0.001
R14847 S.n10522 S.n10515 0.001
R14848 S.t12 S.n11162 0.001
R14849 S.t12 S.n11165 0.001
R14850 S.n11145 S.n11138 0.001
R14851 S.t44 S.n11740 0.001
R14852 S.t44 S.n11743 0.001
R14853 S.t2 S.n12030 0.001
R14854 S.t2 S.n12033 0.001
R14855 S.t72 S.n12909 0.001
R14856 S.t72 S.n12912 0.001
R14857 S.n12881 S.t14 0.001
R14858 S.n12891 S.n12884 0.001
R14859 S.n12890 S.n12889 0.001
R14860 S.n12905 S.n12904 0.001
R14861 S.n12026 S.n12025 0.001
R14862 S.n11736 S.n11735 0.001
R14863 S.n11144 S.n11143 0.001
R14864 S.n11158 S.n11157 0.001
R14865 S.n10521 S.n10520 0.001
R14866 S.n10535 S.n10534 0.001
R14867 S.n9863 S.n9862 0.001
R14868 S.n9877 S.n9876 0.001
R14869 S.n9186 S.n9185 0.001
R14870 S.n9200 S.n9199 0.001
R14871 S.n8782 S.n8781 0.001
R14872 S.n8796 S.n8795 0.001
R14873 S.n8070 S.n8069 0.001
R14874 S.n8084 S.n8083 0.001
R14875 S.n7059 S.n7058 0.001
R14876 S.n7073 S.n7072 0.001
R14877 S.n6312 S.n6311 0.001
R14878 S.n6326 S.n6325 0.001
R14879 S.n5552 S.n5551 0.001
R14880 S.n5566 S.n5565 0.001
R14881 S.n4770 S.n4769 0.001
R14882 S.n4784 S.n4783 0.001
R14883 S.n3975 S.n3974 0.001
R14884 S.n3989 S.n3988 0.001
R14885 S.n3158 S.n3157 0.001
R14886 S.n3172 S.n3171 0.001
R14887 S.n2631 S.n2630 0.001
R14888 S.n2645 S.n2644 0.001
R14889 S.n1345 S.n1344 0.001
R14890 S.n1799 S.t320 0.001
R14891 S.n1808 S.n1801 0.001
R14892 S.t142 S.n1330 0.001
R14893 S.t142 S.n1333 0.001
R14894 S.t200 S.n2679 0.001
R14895 S.t200 S.n2682 0.001
R14896 S.n12935 S.n12928 0.001
R14897 S.t72 S.n12940 0.001
R14898 S.t72 S.n12943 0.001
R14899 S.t2 S.n12045 0.001
R14900 S.t2 S.n12048 0.001
R14901 S.t44 S.n11756 0.001
R14902 S.t44 S.n11759 0.001
R14903 S.n11188 S.n11181 0.001
R14904 S.t12 S.n11193 0.001
R14905 S.t12 S.n11196 0.001
R14906 S.n10565 S.n10558 0.001
R14907 S.t103 S.n10570 0.001
R14908 S.t103 S.n10573 0.001
R14909 S.n9907 S.n9900 0.001
R14910 S.t86 S.n9912 0.001
R14911 S.t86 S.n9915 0.001
R14912 S.n9230 S.n9223 0.001
R14913 S.t24 S.n9235 0.001
R14914 S.t24 S.n9238 0.001
R14915 S.n8826 S.n8819 0.001
R14916 S.t131 S.n8831 0.001
R14917 S.t131 S.n8834 0.001
R14918 S.n8114 S.n8107 0.001
R14919 S.t59 S.n8119 0.001
R14920 S.t59 S.n8122 0.001
R14921 S.n7103 S.n7096 0.001
R14922 S.t37 S.n7108 0.001
R14923 S.t37 S.n7111 0.001
R14924 S.n6356 S.n6349 0.001
R14925 S.t119 S.n6361 0.001
R14926 S.t119 S.n6364 0.001
R14927 S.n5596 S.n5589 0.001
R14928 S.t390 S.n5601 0.001
R14929 S.t390 S.n5604 0.001
R14930 S.n4814 S.n4807 0.001
R14931 S.t360 S.n4819 0.001
R14932 S.t360 S.n4822 0.001
R14933 S.n4022 S.n4015 0.001
R14934 S.t109 S.n3999 0.001
R14935 S.t109 S.n4027 0.001
R14936 S.n4027 S.n4024 0.001
R14937 S.n3493 S.t444 0.001
R14938 S.n3500 S.n3493 0.001
R14939 S.t240 S.n3505 0.001
R14940 S.t240 S.n3508 0.001
R14941 S.n2675 S.n2668 0.001
R14942 S.n2684 S.t200 0.001
R14943 S.n2692 S.n2684 0.001
R14944 S.t55 S.n2616 0.001
R14945 S.t55 S.n2619 0.001
R14946 S.t240 S.n3520 0.001
R14947 S.t240 S.n3523 0.001
R14948 S.t14 S.n12683 0.001
R14949 S.t14 S.n12686 0.001
R14950 S.t72 S.n12955 0.001
R14951 S.t72 S.n12958 0.001
R14952 S.t2 S.n12061 0.001
R14953 S.t2 S.n12064 0.001
R14954 S.t44 S.n11771 0.001
R14955 S.t44 S.n11774 0.001
R14956 S.t18 S.n11453 0.001
R14957 S.t18 S.n11456 0.001
R14958 S.t12 S.n11208 0.001
R14959 S.t12 S.n11211 0.001
R14960 S.t122 S.n10832 0.001
R14961 S.t122 S.n10835 0.001
R14962 S.t103 S.n10585 0.001
R14963 S.t103 S.n10588 0.001
R14964 S.t16 S.n10179 0.001
R14965 S.t16 S.n10182 0.001
R14966 S.t86 S.n9927 0.001
R14967 S.t86 S.n9930 0.001
R14968 S.t26 S.n9503 0.001
R14969 S.t26 S.n9506 0.001
R14970 S.t24 S.n9250 0.001
R14971 S.t24 S.n9253 0.001
R14972 S.t0 S.n8636 0.001
R14973 S.t0 S.n8639 0.001
R14974 S.t131 S.n8846 0.001
R14975 S.t131 S.n8849 0.001
R14976 S.t22 S.n7940 0.001
R14977 S.t22 S.n7943 0.001
R14978 S.t59 S.n8134 0.001
R14979 S.t59 S.n8137 0.001
R14980 S.t40 S.n7387 0.001
R14981 S.t40 S.n7390 0.001
R14982 S.t37 S.n7123 0.001
R14983 S.t37 S.n7126 0.001
R14984 S.t8 S.n6641 0.001
R14985 S.t8 S.n6644 0.001
R14986 S.t119 S.n6376 0.001
R14987 S.t119 S.n6379 0.001
R14988 S.t460 S.n5886 0.001
R14989 S.t460 S.n5889 0.001
R14990 S.t390 S.n5616 0.001
R14991 S.t390 S.n5619 0.001
R14992 S.t81 S.n5105 0.001
R14993 S.t81 S.n5108 0.001
R14994 S.t360 S.n4834 0.001
R14995 S.t360 S.n4837 0.001
R14996 S.t51 S.n4315 0.001
R14997 S.t51 S.n4318 0.001
R14998 S.t109 S.n4039 0.001
R14999 S.t109 S.n4042 0.001
R15000 S.t444 S.n3467 0.001
R15001 S.t444 S.n3470 0.001
R15002 S.n3525 S.t240 0.001
R15003 S.n3533 S.n3525 0.001
R15004 S.t444 S.n3487 0.001
R15005 S.t444 S.n3490 0.001
R15006 S.t109 S.n4352 0.001
R15007 S.t109 S.n4355 0.001
R15008 S.t14 S.n12699 0.001
R15009 S.t14 S.n12702 0.001
R15010 S.t72 S.n12970 0.001
R15011 S.t72 S.n12973 0.001
R15012 S.t2 S.n12077 0.001
R15013 S.t2 S.n12080 0.001
R15014 S.t44 S.n11786 0.001
R15015 S.t44 S.n11789 0.001
R15016 S.t18 S.n11469 0.001
R15017 S.t18 S.n11472 0.001
R15018 S.t12 S.n11223 0.001
R15019 S.t12 S.n11226 0.001
R15020 S.t122 S.n10848 0.001
R15021 S.t122 S.n10851 0.001
R15022 S.t103 S.n10600 0.001
R15023 S.t103 S.n10603 0.001
R15024 S.t16 S.n10195 0.001
R15025 S.t16 S.n10198 0.001
R15026 S.t86 S.n9942 0.001
R15027 S.t86 S.n9945 0.001
R15028 S.t26 S.n9519 0.001
R15029 S.t26 S.n9522 0.001
R15030 S.t24 S.n9265 0.001
R15031 S.t24 S.n9268 0.001
R15032 S.t0 S.n8652 0.001
R15033 S.t0 S.n8655 0.001
R15034 S.t131 S.n8861 0.001
R15035 S.t131 S.n8864 0.001
R15036 S.t22 S.n7956 0.001
R15037 S.t22 S.n7959 0.001
R15038 S.t59 S.n8149 0.001
R15039 S.t59 S.n8152 0.001
R15040 S.t40 S.n7403 0.001
R15041 S.t40 S.n7406 0.001
R15042 S.t37 S.n7138 0.001
R15043 S.t37 S.n7141 0.001
R15044 S.t8 S.n6657 0.001
R15045 S.t8 S.n6660 0.001
R15046 S.t119 S.n6391 0.001
R15047 S.t119 S.n6394 0.001
R15048 S.t460 S.n5902 0.001
R15049 S.t460 S.n5905 0.001
R15050 S.t390 S.n5631 0.001
R15051 S.t390 S.n5634 0.001
R15052 S.t81 S.n5121 0.001
R15053 S.t81 S.n5124 0.001
R15054 S.t360 S.n4849 0.001
R15055 S.t360 S.n4852 0.001
R15056 S.n4341 S.t51 0.001
R15057 S.n4348 S.n4341 0.001
R15058 S.n4357 S.t109 0.001
R15059 S.n4365 S.n4357 0.001
R15060 S.t51 S.n4335 0.001
R15061 S.t51 S.n4338 0.001
R15062 S.t360 S.n5158 0.001
R15063 S.t360 S.n5161 0.001
R15064 S.t14 S.n12715 0.001
R15065 S.t14 S.n12718 0.001
R15066 S.t72 S.n12985 0.001
R15067 S.t72 S.n12988 0.001
R15068 S.t2 S.n12093 0.001
R15069 S.t2 S.n12096 0.001
R15070 S.t44 S.n11801 0.001
R15071 S.t44 S.n11804 0.001
R15072 S.t18 S.n11485 0.001
R15073 S.t18 S.n11488 0.001
R15074 S.t12 S.n11238 0.001
R15075 S.t12 S.n11241 0.001
R15076 S.t122 S.n10864 0.001
R15077 S.t122 S.n10867 0.001
R15078 S.t103 S.n10615 0.001
R15079 S.t103 S.n10618 0.001
R15080 S.t16 S.n10211 0.001
R15081 S.t16 S.n10214 0.001
R15082 S.t86 S.n9957 0.001
R15083 S.t86 S.n9960 0.001
R15084 S.t26 S.n9535 0.001
R15085 S.t26 S.n9538 0.001
R15086 S.t24 S.n9280 0.001
R15087 S.t24 S.n9283 0.001
R15088 S.t0 S.n8668 0.001
R15089 S.t0 S.n8671 0.001
R15090 S.t131 S.n8876 0.001
R15091 S.t131 S.n8879 0.001
R15092 S.t22 S.n7972 0.001
R15093 S.t22 S.n7975 0.001
R15094 S.t59 S.n8164 0.001
R15095 S.t59 S.n8167 0.001
R15096 S.t40 S.n7419 0.001
R15097 S.t40 S.n7422 0.001
R15098 S.t37 S.n7153 0.001
R15099 S.t37 S.n7156 0.001
R15100 S.t8 S.n6673 0.001
R15101 S.t8 S.n6676 0.001
R15102 S.t119 S.n6406 0.001
R15103 S.t119 S.n6409 0.001
R15104 S.t460 S.n5918 0.001
R15105 S.t460 S.n5921 0.001
R15106 S.t390 S.n5646 0.001
R15107 S.t390 S.n5649 0.001
R15108 S.n5147 S.t81 0.001
R15109 S.n5154 S.n5147 0.001
R15110 S.n5163 S.t360 0.001
R15111 S.n5171 S.n5163 0.001
R15112 S.t81 S.n5141 0.001
R15113 S.t81 S.n5144 0.001
R15114 S.t390 S.n5955 0.001
R15115 S.t390 S.n5958 0.001
R15116 S.t14 S.n12731 0.001
R15117 S.t14 S.n12734 0.001
R15118 S.t72 S.n13000 0.001
R15119 S.t72 S.n13003 0.001
R15120 S.t2 S.n12109 0.001
R15121 S.t2 S.n12112 0.001
R15122 S.t44 S.n11816 0.001
R15123 S.t44 S.n11819 0.001
R15124 S.t18 S.n11501 0.001
R15125 S.t18 S.n11504 0.001
R15126 S.t12 S.n11253 0.001
R15127 S.t12 S.n11256 0.001
R15128 S.t122 S.n10880 0.001
R15129 S.t122 S.n10883 0.001
R15130 S.t103 S.n10630 0.001
R15131 S.t103 S.n10633 0.001
R15132 S.t16 S.n10227 0.001
R15133 S.t16 S.n10230 0.001
R15134 S.t86 S.n9972 0.001
R15135 S.t86 S.n9975 0.001
R15136 S.t26 S.n9551 0.001
R15137 S.t26 S.n9554 0.001
R15138 S.t24 S.n9295 0.001
R15139 S.t24 S.n9298 0.001
R15140 S.t0 S.n8684 0.001
R15141 S.t0 S.n8687 0.001
R15142 S.t131 S.n8891 0.001
R15143 S.t131 S.n8894 0.001
R15144 S.t22 S.n7988 0.001
R15145 S.t22 S.n7991 0.001
R15146 S.t59 S.n8179 0.001
R15147 S.t59 S.n8182 0.001
R15148 S.t40 S.n7435 0.001
R15149 S.t40 S.n7438 0.001
R15150 S.t37 S.n7168 0.001
R15151 S.t37 S.n7171 0.001
R15152 S.t8 S.n6689 0.001
R15153 S.t8 S.n6692 0.001
R15154 S.t119 S.n6421 0.001
R15155 S.t119 S.n6424 0.001
R15156 S.n5944 S.t460 0.001
R15157 S.n5951 S.n5944 0.001
R15158 S.n5960 S.t390 0.001
R15159 S.n5968 S.n5960 0.001
R15160 S.t460 S.n5938 0.001
R15161 S.t460 S.n5941 0.001
R15162 S.t119 S.n6726 0.001
R15163 S.t119 S.n6729 0.001
R15164 S.t14 S.n12747 0.001
R15165 S.t14 S.n12750 0.001
R15166 S.t72 S.n13015 0.001
R15167 S.t72 S.n13018 0.001
R15168 S.t2 S.n12125 0.001
R15169 S.t2 S.n12128 0.001
R15170 S.t44 S.n11831 0.001
R15171 S.t44 S.n11834 0.001
R15172 S.t18 S.n11517 0.001
R15173 S.t18 S.n11520 0.001
R15174 S.t12 S.n11268 0.001
R15175 S.t12 S.n11271 0.001
R15176 S.t122 S.n10896 0.001
R15177 S.t122 S.n10899 0.001
R15178 S.t103 S.n10645 0.001
R15179 S.t103 S.n10648 0.001
R15180 S.t16 S.n10243 0.001
R15181 S.t16 S.n10246 0.001
R15182 S.t86 S.n9987 0.001
R15183 S.t86 S.n9990 0.001
R15184 S.t26 S.n9567 0.001
R15185 S.t26 S.n9570 0.001
R15186 S.t24 S.n9310 0.001
R15187 S.t24 S.n9313 0.001
R15188 S.t0 S.n8700 0.001
R15189 S.t0 S.n8703 0.001
R15190 S.t131 S.n8906 0.001
R15191 S.t131 S.n8909 0.001
R15192 S.t22 S.n8004 0.001
R15193 S.t22 S.n8007 0.001
R15194 S.t59 S.n8194 0.001
R15195 S.t59 S.n8197 0.001
R15196 S.t40 S.n7451 0.001
R15197 S.t40 S.n7454 0.001
R15198 S.t37 S.n7183 0.001
R15199 S.t37 S.n7186 0.001
R15200 S.n6715 S.t8 0.001
R15201 S.n6722 S.n6715 0.001
R15202 S.n6731 S.t119 0.001
R15203 S.n6739 S.n6731 0.001
R15204 S.t8 S.n6709 0.001
R15205 S.t8 S.n6712 0.001
R15206 S.t37 S.n7488 0.001
R15207 S.t37 S.n7491 0.001
R15208 S.t14 S.n12763 0.001
R15209 S.t14 S.n12766 0.001
R15210 S.t72 S.n13030 0.001
R15211 S.t72 S.n13033 0.001
R15212 S.t2 S.n12141 0.001
R15213 S.t2 S.n12144 0.001
R15214 S.t44 S.n11846 0.001
R15215 S.t44 S.n11849 0.001
R15216 S.t18 S.n11533 0.001
R15217 S.t18 S.n11536 0.001
R15218 S.t12 S.n11283 0.001
R15219 S.t12 S.n11286 0.001
R15220 S.t122 S.n10912 0.001
R15221 S.t122 S.n10915 0.001
R15222 S.t103 S.n10660 0.001
R15223 S.t103 S.n10663 0.001
R15224 S.t16 S.n10259 0.001
R15225 S.t16 S.n10262 0.001
R15226 S.t86 S.n10002 0.001
R15227 S.t86 S.n10005 0.001
R15228 S.t26 S.n9583 0.001
R15229 S.t26 S.n9586 0.001
R15230 S.t24 S.n9325 0.001
R15231 S.t24 S.n9328 0.001
R15232 S.t0 S.n8716 0.001
R15233 S.t0 S.n8719 0.001
R15234 S.t131 S.n8921 0.001
R15235 S.t131 S.n8924 0.001
R15236 S.t22 S.n8020 0.001
R15237 S.t22 S.n8023 0.001
R15238 S.t59 S.n8209 0.001
R15239 S.t59 S.n8212 0.001
R15240 S.n7477 S.t40 0.001
R15241 S.n7484 S.n7477 0.001
R15242 S.n7493 S.t37 0.001
R15243 S.n7501 S.n7493 0.001
R15244 S.t40 S.n7471 0.001
R15245 S.t40 S.n7474 0.001
R15246 S.t59 S.n8224 0.001
R15247 S.t59 S.n8227 0.001
R15248 S.t14 S.n12779 0.001
R15249 S.t14 S.n12782 0.001
R15250 S.t72 S.n13045 0.001
R15251 S.t72 S.n13048 0.001
R15252 S.t2 S.n12157 0.001
R15253 S.t2 S.n12160 0.001
R15254 S.t44 S.n11861 0.001
R15255 S.t44 S.n11864 0.001
R15256 S.t18 S.n11549 0.001
R15257 S.t18 S.n11552 0.001
R15258 S.t12 S.n11298 0.001
R15259 S.t12 S.n11301 0.001
R15260 S.t122 S.n10928 0.001
R15261 S.t122 S.n10931 0.001
R15262 S.t103 S.n10675 0.001
R15263 S.t103 S.n10678 0.001
R15264 S.t16 S.n10275 0.001
R15265 S.t16 S.n10278 0.001
R15266 S.t86 S.n10017 0.001
R15267 S.t86 S.n10020 0.001
R15268 S.t26 S.n9599 0.001
R15269 S.t26 S.n9602 0.001
R15270 S.t24 S.n9340 0.001
R15271 S.t24 S.n9343 0.001
R15272 S.t0 S.n8732 0.001
R15273 S.t0 S.n8735 0.001
R15274 S.t131 S.n8936 0.001
R15275 S.t131 S.n8939 0.001
R15276 S.t22 S.n8035 0.001
R15277 S.t22 S.n8038 0.001
R15278 S.n8229 S.t59 0.001
R15279 S.n8237 S.n8229 0.001
R15280 S.t22 S.n8055 0.001
R15281 S.t22 S.n8058 0.001
R15282 S.t131 S.n8951 0.001
R15283 S.t131 S.n8954 0.001
R15284 S.t14 S.n12795 0.001
R15285 S.t14 S.n12798 0.001
R15286 S.t72 S.n13060 0.001
R15287 S.t72 S.n13063 0.001
R15288 S.t2 S.n12173 0.001
R15289 S.t2 S.n12176 0.001
R15290 S.t44 S.n11876 0.001
R15291 S.t44 S.n11879 0.001
R15292 S.t18 S.n11565 0.001
R15293 S.t18 S.n11568 0.001
R15294 S.t12 S.n11313 0.001
R15295 S.t12 S.n11316 0.001
R15296 S.t122 S.n10944 0.001
R15297 S.t122 S.n10947 0.001
R15298 S.t103 S.n10690 0.001
R15299 S.t103 S.n10693 0.001
R15300 S.t16 S.n10291 0.001
R15301 S.t16 S.n10294 0.001
R15302 S.t86 S.n10032 0.001
R15303 S.t86 S.n10035 0.001
R15304 S.t26 S.n9615 0.001
R15305 S.t26 S.n9618 0.001
R15306 S.t24 S.n9355 0.001
R15307 S.t24 S.n9358 0.001
R15308 S.t0 S.n8747 0.001
R15309 S.t0 S.n8750 0.001
R15310 S.n8956 S.t131 0.001
R15311 S.n8964 S.n8956 0.001
R15312 S.t0 S.n8767 0.001
R15313 S.t0 S.n8770 0.001
R15314 S.t24 S.n9652 0.001
R15315 S.t24 S.n9655 0.001
R15316 S.t14 S.n12811 0.001
R15317 S.t14 S.n12814 0.001
R15318 S.t72 S.n13075 0.001
R15319 S.t72 S.n13078 0.001
R15320 S.t2 S.n12189 0.001
R15321 S.t2 S.n12192 0.001
R15322 S.t44 S.n11891 0.001
R15323 S.t44 S.n11894 0.001
R15324 S.t18 S.n11581 0.001
R15325 S.t18 S.n11584 0.001
R15326 S.t12 S.n11328 0.001
R15327 S.t12 S.n11331 0.001
R15328 S.t122 S.n10960 0.001
R15329 S.t122 S.n10963 0.001
R15330 S.t103 S.n10705 0.001
R15331 S.t103 S.n10708 0.001
R15332 S.t16 S.n10307 0.001
R15333 S.t16 S.n10310 0.001
R15334 S.t86 S.n10047 0.001
R15335 S.t86 S.n10050 0.001
R15336 S.n9641 S.t26 0.001
R15337 S.n9648 S.n9641 0.001
R15338 S.n9657 S.t24 0.001
R15339 S.n9665 S.n9657 0.001
R15340 S.t26 S.n9635 0.001
R15341 S.t26 S.n9638 0.001
R15342 S.t86 S.n10344 0.001
R15343 S.t86 S.n10347 0.001
R15344 S.t14 S.n12827 0.001
R15345 S.t14 S.n12830 0.001
R15346 S.t72 S.n13090 0.001
R15347 S.t72 S.n13093 0.001
R15348 S.t2 S.n12205 0.001
R15349 S.t2 S.n12208 0.001
R15350 S.t44 S.n11906 0.001
R15351 S.t44 S.n11909 0.001
R15352 S.t18 S.n11597 0.001
R15353 S.t18 S.n11600 0.001
R15354 S.t12 S.n11343 0.001
R15355 S.t12 S.n11346 0.001
R15356 S.t122 S.n10976 0.001
R15357 S.t122 S.n10979 0.001
R15358 S.t103 S.n10720 0.001
R15359 S.t103 S.n10723 0.001
R15360 S.n10333 S.t16 0.001
R15361 S.n10340 S.n10333 0.001
R15362 S.n10349 S.t86 0.001
R15363 S.n10357 S.n10349 0.001
R15364 S.t16 S.n10327 0.001
R15365 S.t16 S.n10330 0.001
R15366 S.t103 S.n11013 0.001
R15367 S.t103 S.n11016 0.001
R15368 S.t14 S.n12843 0.001
R15369 S.t14 S.n12846 0.001
R15370 S.t72 S.n13105 0.001
R15371 S.t72 S.n13108 0.001
R15372 S.t2 S.n12221 0.001
R15373 S.t2 S.n12224 0.001
R15374 S.t44 S.n11921 0.001
R15375 S.t44 S.n11924 0.001
R15376 S.t18 S.n11613 0.001
R15377 S.t18 S.n11616 0.001
R15378 S.t12 S.n11358 0.001
R15379 S.t12 S.n11361 0.001
R15380 S.n11002 S.t122 0.001
R15381 S.n11009 S.n11002 0.001
R15382 S.n11018 S.t103 0.001
R15383 S.n11026 S.n11018 0.001
R15384 S.t122 S.n10996 0.001
R15385 S.t122 S.n10999 0.001
R15386 S.t12 S.n11653 0.001
R15387 S.t12 S.n11656 0.001
R15388 S.t14 S.n12859 0.001
R15389 S.t14 S.n12862 0.001
R15390 S.t72 S.n13120 0.001
R15391 S.t72 S.n13123 0.001
R15392 S.t2 S.n12237 0.001
R15393 S.t2 S.n12240 0.001
R15394 S.t44 S.n11936 0.001
R15395 S.t44 S.n11939 0.001
R15396 S.n11642 S.t18 0.001
R15397 S.n11649 S.n11642 0.001
R15398 S.n11658 S.t12 0.001
R15399 S.n11666 S.n11658 0.001
R15400 S.t18 S.n11636 0.001
R15401 S.t18 S.n11639 0.001
R15402 S.t44 S.n12268 0.001
R15403 S.t44 S.n12271 0.001
R15404 S.t14 S.n12875 0.001
R15405 S.t14 S.n12878 0.001
R15406 S.t72 S.n13138 0.001
R15407 S.t72 S.n13141 0.001
R15408 S.n12243 S.t2 0.001
R15409 S.n12251 S.n12246 0.001
R15410 S.t14 S.n12669 0.001
R15411 S.t14 S.n12666 0.001
R15412 S.n12666 S.n12663 0.001
R15413 S.n13144 S.t72 0.001
R15414 S.n13161 S.n13146 0.001
R15415 S.n104 S.n103 0.001
R15416 S.n108 S.n107 0.001
R15417 S.n13159 S.n13158 0.001
R15418 S.n12289 S.n12288 0.001
R15419 S.n872 S.n871 0.001
R15420 S.n995 S.n994 0.001
R15421 S.n1839 S.n1838 0.001
R15422 S.n2722 S.n2721 0.001
R15423 S.n3563 S.n3562 0.001
R15424 S.n4395 S.n4394 0.001
R15425 S.n5201 S.n5200 0.001
R15426 S.n5998 S.n5997 0.001
R15427 S.n6769 S.n6768 0.001
R15428 S.n7531 S.n7530 0.001
R15429 S.n8267 S.n8266 0.001
R15430 S.n8994 S.n8993 0.001
R15431 S.n9695 S.n9694 0.001
R15432 S.n10387 S.n10386 0.001
R15433 S.n11046 S.n11045 0.001
R15434 S.n12314 S.n12313 0.001
R15435 S.n12463 S.n12418 0.001
R15436 S.n12463 S.n12416 0.001
R15437 S.n12463 S.n12414 0.001
R15438 S.n12463 S.n12412 0.001
R15439 S.n12463 S.n12410 0.001
R15440 S.n12463 S.n12408 0.001
R15441 S.n12463 S.n12406 0.001
R15442 S.n12463 S.n12404 0.001
R15443 S.n12463 S.n12402 0.001
R15444 S.n12463 S.n12400 0.001
R15445 S.n12463 S.n12398 0.001
R15446 S.n12463 S.n12396 0.001
R15447 S.n12463 S.n12394 0.001
R15448 S.n12613 S.n12612 0.001
R15449 S.n12306 S.n12274 0.001
R15450 S.n12594 S.n12591 0.001
R15451 S.n11720 S.n11717 0.001
R15452 S.n11125 S.n11122 0.001
R15453 S.n901 S.n888 0.001
R15454 S.n765 S.n757 0.001
R15455 S.n10502 S.n10499 0.001
R15456 S.n9844 S.n9841 0.001
R15457 S.n9167 S.n9164 0.001
R15458 S.n8477 S.n8474 0.001
R15459 S.n7765 S.n7762 0.001
R15460 S.n7040 S.n7037 0.001
R15461 S.n6293 S.n6290 0.001
R15462 S.n5533 S.n5530 0.001
R15463 S.n59 S.n51 0.001
R15464 S.n4751 S.n4748 0.001
R15465 S.n3956 S.n3953 0.001
R15466 S.n1472 S.n1469 0.001
R15467 S.n3139 S.n3136 0.001
R15468 S.n2309 S.n2306 0.001
R15469 S.n854 S.n851 0.001
R15470 S.n13161 S.n13144 0.001
R15471 S.n883 S.n880 0.001
R15472 S.n12891 S.n12881 0.001
R15473 S.n12909 S.n12906 0.001
R15474 S.n12030 S.n12027 0.001
R15475 S.n11740 S.n11737 0.001
R15476 S.n11145 S.n11135 0.001
R15477 S.n11162 S.n11159 0.001
R15478 S.n10522 S.n10512 0.001
R15479 S.n10539 S.n10536 0.001
R15480 S.n9864 S.n9854 0.001
R15481 S.n9881 S.n9878 0.001
R15482 S.n9187 S.n9177 0.001
R15483 S.n9204 S.n9201 0.001
R15484 S.n8783 S.n8773 0.001
R15485 S.n8800 S.n8797 0.001
R15486 S.n8071 S.n8061 0.001
R15487 S.n8088 S.n8085 0.001
R15488 S.n7060 S.n7050 0.001
R15489 S.n7077 S.n7074 0.001
R15490 S.n6313 S.n6303 0.001
R15491 S.n6330 S.n6327 0.001
R15492 S.n5553 S.n5543 0.001
R15493 S.n5570 S.n5567 0.001
R15494 S.n4771 S.n4761 0.001
R15495 S.n4788 S.n4785 0.001
R15496 S.n3976 S.n3966 0.001
R15497 S.n3993 S.n3990 0.001
R15498 S.n3159 S.n3149 0.001
R15499 S.n3176 S.n3173 0.001
R15500 S.n2632 S.n2622 0.001
R15501 S.n2649 S.n2646 0.001
R15502 S.n1346 S.n1336 0.001
R15503 S.n751 S.n748 0.001
R15504 S.n1808 S.n1799 0.001
R15505 S.n12935 S.n12931 0.001
R15506 S.n12940 S.n12937 0.001
R15507 S.n12045 S.n12042 0.001
R15508 S.n11756 S.n11753 0.001
R15509 S.n11188 S.n11184 0.001
R15510 S.n11193 S.n11190 0.001
R15511 S.n10565 S.n10561 0.001
R15512 S.n10570 S.n10567 0.001
R15513 S.n9907 S.n9903 0.001
R15514 S.n9912 S.n9909 0.001
R15515 S.n9230 S.n9226 0.001
R15516 S.n9235 S.n9232 0.001
R15517 S.n8826 S.n8822 0.001
R15518 S.n8831 S.n8828 0.001
R15519 S.n8114 S.n8110 0.001
R15520 S.n8119 S.n8116 0.001
R15521 S.n7103 S.n7099 0.001
R15522 S.n7108 S.n7105 0.001
R15523 S.n6356 S.n6352 0.001
R15524 S.n6361 S.n6358 0.001
R15525 S.n5596 S.n5592 0.001
R15526 S.n5601 S.n5598 0.001
R15527 S.n4814 S.n4810 0.001
R15528 S.n4819 S.n4816 0.001
R15529 S.n4022 S.n4018 0.001
R15530 S.n3500 S.n3496 0.001
R15531 S.n3505 S.n3502 0.001
R15532 S.n2675 S.n2671 0.001
R15533 S.n2679 S.n2676 0.001
R15534 S.n1330 S.n1327 0.001
R15535 S.n2692 S.n2687 0.001
R15536 S.n2616 S.n2613 0.001
R15537 S.n3520 S.n3517 0.001
R15538 S.n3467 S.n3464 0.001
R15539 S.n4039 S.n4036 0.001
R15540 S.n4315 S.n4312 0.001
R15541 S.n4834 S.n4831 0.001
R15542 S.n5105 S.n5102 0.001
R15543 S.n5616 S.n5613 0.001
R15544 S.n5886 S.n5883 0.001
R15545 S.n6376 S.n6373 0.001
R15546 S.n6641 S.n6638 0.001
R15547 S.n7123 S.n7120 0.001
R15548 S.n7387 S.n7384 0.001
R15549 S.n8134 S.n8131 0.001
R15550 S.n7940 S.n7937 0.001
R15551 S.n8846 S.n8843 0.001
R15552 S.n8636 S.n8633 0.001
R15553 S.n9250 S.n9247 0.001
R15554 S.n9503 S.n9500 0.001
R15555 S.n9927 S.n9924 0.001
R15556 S.n10179 S.n10176 0.001
R15557 S.n10585 S.n10582 0.001
R15558 S.n10832 S.n10829 0.001
R15559 S.n11208 S.n11205 0.001
R15560 S.n11453 S.n11450 0.001
R15561 S.n11771 S.n11768 0.001
R15562 S.n12061 S.n12058 0.001
R15563 S.n12955 S.n12952 0.001
R15564 S.n12683 S.n12680 0.001
R15565 S.n3533 S.n3528 0.001
R15566 S.n3487 S.n3484 0.001
R15567 S.n4352 S.n4349 0.001
R15568 S.n4348 S.n4344 0.001
R15569 S.n4849 S.n4846 0.001
R15570 S.n5121 S.n5118 0.001
R15571 S.n5631 S.n5628 0.001
R15572 S.n5902 S.n5899 0.001
R15573 S.n6391 S.n6388 0.001
R15574 S.n6657 S.n6654 0.001
R15575 S.n7138 S.n7135 0.001
R15576 S.n7403 S.n7400 0.001
R15577 S.n8149 S.n8146 0.001
R15578 S.n7956 S.n7953 0.001
R15579 S.n8861 S.n8858 0.001
R15580 S.n8652 S.n8649 0.001
R15581 S.n9265 S.n9262 0.001
R15582 S.n9519 S.n9516 0.001
R15583 S.n9942 S.n9939 0.001
R15584 S.n10195 S.n10192 0.001
R15585 S.n10600 S.n10597 0.001
R15586 S.n10848 S.n10845 0.001
R15587 S.n11223 S.n11220 0.001
R15588 S.n11469 S.n11466 0.001
R15589 S.n11786 S.n11783 0.001
R15590 S.n12077 S.n12074 0.001
R15591 S.n12970 S.n12967 0.001
R15592 S.n12699 S.n12696 0.001
R15593 S.n4365 S.n4360 0.001
R15594 S.n4335 S.n4332 0.001
R15595 S.n5158 S.n5155 0.001
R15596 S.n5154 S.n5150 0.001
R15597 S.n5646 S.n5643 0.001
R15598 S.n5918 S.n5915 0.001
R15599 S.n6406 S.n6403 0.001
R15600 S.n6673 S.n6670 0.001
R15601 S.n7153 S.n7150 0.001
R15602 S.n7419 S.n7416 0.001
R15603 S.n8164 S.n8161 0.001
R15604 S.n7972 S.n7969 0.001
R15605 S.n8876 S.n8873 0.001
R15606 S.n8668 S.n8665 0.001
R15607 S.n9280 S.n9277 0.001
R15608 S.n9535 S.n9532 0.001
R15609 S.n9957 S.n9954 0.001
R15610 S.n10211 S.n10208 0.001
R15611 S.n10615 S.n10612 0.001
R15612 S.n10864 S.n10861 0.001
R15613 S.n11238 S.n11235 0.001
R15614 S.n11485 S.n11482 0.001
R15615 S.n11801 S.n11798 0.001
R15616 S.n12093 S.n12090 0.001
R15617 S.n12985 S.n12982 0.001
R15618 S.n12715 S.n12712 0.001
R15619 S.n5171 S.n5166 0.001
R15620 S.n5141 S.n5138 0.001
R15621 S.n5955 S.n5952 0.001
R15622 S.n5951 S.n5947 0.001
R15623 S.n6421 S.n6418 0.001
R15624 S.n6689 S.n6686 0.001
R15625 S.n7168 S.n7165 0.001
R15626 S.n7435 S.n7432 0.001
R15627 S.n8179 S.n8176 0.001
R15628 S.n7988 S.n7985 0.001
R15629 S.n8891 S.n8888 0.001
R15630 S.n8684 S.n8681 0.001
R15631 S.n9295 S.n9292 0.001
R15632 S.n9551 S.n9548 0.001
R15633 S.n9972 S.n9969 0.001
R15634 S.n10227 S.n10224 0.001
R15635 S.n10630 S.n10627 0.001
R15636 S.n10880 S.n10877 0.001
R15637 S.n11253 S.n11250 0.001
R15638 S.n11501 S.n11498 0.001
R15639 S.n11816 S.n11813 0.001
R15640 S.n12109 S.n12106 0.001
R15641 S.n13000 S.n12997 0.001
R15642 S.n12731 S.n12728 0.001
R15643 S.n5968 S.n5963 0.001
R15644 S.n5938 S.n5935 0.001
R15645 S.n6726 S.n6723 0.001
R15646 S.n6722 S.n6718 0.001
R15647 S.n7183 S.n7180 0.001
R15648 S.n7451 S.n7448 0.001
R15649 S.n8194 S.n8191 0.001
R15650 S.n8004 S.n8001 0.001
R15651 S.n8906 S.n8903 0.001
R15652 S.n8700 S.n8697 0.001
R15653 S.n9310 S.n9307 0.001
R15654 S.n9567 S.n9564 0.001
R15655 S.n9987 S.n9984 0.001
R15656 S.n10243 S.n10240 0.001
R15657 S.n10645 S.n10642 0.001
R15658 S.n10896 S.n10893 0.001
R15659 S.n11268 S.n11265 0.001
R15660 S.n11517 S.n11514 0.001
R15661 S.n11831 S.n11828 0.001
R15662 S.n12125 S.n12122 0.001
R15663 S.n13015 S.n13012 0.001
R15664 S.n12747 S.n12744 0.001
R15665 S.n6739 S.n6734 0.001
R15666 S.n6709 S.n6706 0.001
R15667 S.n7488 S.n7485 0.001
R15668 S.n7484 S.n7480 0.001
R15669 S.n8209 S.n8206 0.001
R15670 S.n8020 S.n8017 0.001
R15671 S.n8921 S.n8918 0.001
R15672 S.n8716 S.n8713 0.001
R15673 S.n9325 S.n9322 0.001
R15674 S.n9583 S.n9580 0.001
R15675 S.n10002 S.n9999 0.001
R15676 S.n10259 S.n10256 0.001
R15677 S.n10660 S.n10657 0.001
R15678 S.n10912 S.n10909 0.001
R15679 S.n11283 S.n11280 0.001
R15680 S.n11533 S.n11530 0.001
R15681 S.n11846 S.n11843 0.001
R15682 S.n12141 S.n12138 0.001
R15683 S.n13030 S.n13027 0.001
R15684 S.n12763 S.n12760 0.001
R15685 S.n7501 S.n7496 0.001
R15686 S.n7471 S.n7468 0.001
R15687 S.n8224 S.n8221 0.001
R15688 S.n8035 S.n8032 0.001
R15689 S.n8936 S.n8933 0.001
R15690 S.n8732 S.n8729 0.001
R15691 S.n9340 S.n9337 0.001
R15692 S.n9599 S.n9596 0.001
R15693 S.n10017 S.n10014 0.001
R15694 S.n10275 S.n10272 0.001
R15695 S.n10675 S.n10672 0.001
R15696 S.n10928 S.n10925 0.001
R15697 S.n11298 S.n11295 0.001
R15698 S.n11549 S.n11546 0.001
R15699 S.n11861 S.n11858 0.001
R15700 S.n12157 S.n12154 0.001
R15701 S.n13045 S.n13042 0.001
R15702 S.n12779 S.n12776 0.001
R15703 S.n8237 S.n8232 0.001
R15704 S.n8055 S.n8052 0.001
R15705 S.n8951 S.n8948 0.001
R15706 S.n8747 S.n8744 0.001
R15707 S.n9355 S.n9352 0.001
R15708 S.n9615 S.n9612 0.001
R15709 S.n10032 S.n10029 0.001
R15710 S.n10291 S.n10288 0.001
R15711 S.n10690 S.n10687 0.001
R15712 S.n10944 S.n10941 0.001
R15713 S.n11313 S.n11310 0.001
R15714 S.n11565 S.n11562 0.001
R15715 S.n11876 S.n11873 0.001
R15716 S.n12173 S.n12170 0.001
R15717 S.n13060 S.n13057 0.001
R15718 S.n12795 S.n12792 0.001
R15719 S.n8964 S.n8959 0.001
R15720 S.n8767 S.n8764 0.001
R15721 S.n9652 S.n9649 0.001
R15722 S.n9648 S.n9644 0.001
R15723 S.n10047 S.n10044 0.001
R15724 S.n10307 S.n10304 0.001
R15725 S.n10705 S.n10702 0.001
R15726 S.n10960 S.n10957 0.001
R15727 S.n11328 S.n11325 0.001
R15728 S.n11581 S.n11578 0.001
R15729 S.n11891 S.n11888 0.001
R15730 S.n12189 S.n12186 0.001
R15731 S.n13075 S.n13072 0.001
R15732 S.n12811 S.n12808 0.001
R15733 S.n9665 S.n9660 0.001
R15734 S.n9635 S.n9632 0.001
R15735 S.n10344 S.n10341 0.001
R15736 S.n10340 S.n10336 0.001
R15737 S.n10720 S.n10717 0.001
R15738 S.n10976 S.n10973 0.001
R15739 S.n11343 S.n11340 0.001
R15740 S.n11597 S.n11594 0.001
R15741 S.n11906 S.n11903 0.001
R15742 S.n12205 S.n12202 0.001
R15743 S.n13090 S.n13087 0.001
R15744 S.n12827 S.n12824 0.001
R15745 S.n10357 S.n10352 0.001
R15746 S.n10327 S.n10324 0.001
R15747 S.n11013 S.n11010 0.001
R15748 S.n11009 S.n11005 0.001
R15749 S.n11358 S.n11355 0.001
R15750 S.n11613 S.n11610 0.001
R15751 S.n11921 S.n11918 0.001
R15752 S.n12221 S.n12218 0.001
R15753 S.n13105 S.n13102 0.001
R15754 S.n12843 S.n12840 0.001
R15755 S.n11026 S.n11021 0.001
R15756 S.n10996 S.n10993 0.001
R15757 S.n11653 S.n11650 0.001
R15758 S.n11649 S.n11645 0.001
R15759 S.n11936 S.n11933 0.001
R15760 S.n12237 S.n12234 0.001
R15761 S.n13120 S.n13117 0.001
R15762 S.n12859 S.n12856 0.001
R15763 S.n11666 S.n11661 0.001
R15764 S.n11636 S.n11633 0.001
R15765 S.n12268 S.n12265 0.001
R15766 S.n12251 S.n12243 0.001
R15767 S.n13138 S.n13135 0.001
R15768 S.n12875 S.n12872 0.001
R15769 S.n12614 S.n12613 0.001
C0 DNW S 5943.07fF
C1 DNW G 9.27fF
C2 S G 3017.69fF
C3 DNW D 518.88fF
C4 S D 4783.55fF
C5 G D 2242.28fF
C6 D SUB -65.06fF
C7 G SUB -303.14fF
C8 S SUB 381.66fF $ **FLOATING
C9 DNW SUB 11261.70fF $ **FLOATING
C10 S.n0 SUB 0.96fF $ **FLOATING
C11 S.n1 SUB 0.94fF $ **FLOATING
C12 S.n2 SUB 0.34fF $ **FLOATING
C13 S.n3 SUB 0.46fF $ **FLOATING
C14 S.n4 SUB 0.33fF $ **FLOATING
C15 S.n5 SUB 1.49fF $ **FLOATING
C16 S.n6 SUB 2.63fF $ **FLOATING
C17 S.n7 SUB 8.97fF $ **FLOATING
C18 S.n8 SUB 8.97fF $ **FLOATING
C19 S.n9 SUB 5.38fF $ **FLOATING
C20 S.n10 SUB 2.17fF $ **FLOATING
C21 S.n11 SUB 0.96fF $ **FLOATING
C22 S.n12 SUB 0.94fF $ **FLOATING
C23 S.n13 SUB 0.34fF $ **FLOATING
C24 S.n14 SUB 0.46fF $ **FLOATING
C25 S.n15 SUB 0.33fF $ **FLOATING
C26 S.n16 SUB 1.49fF $ **FLOATING
C27 S.n17 SUB 2.63fF $ **FLOATING
C28 S.n18 SUB 8.97fF $ **FLOATING
C29 S.n19 SUB 8.97fF $ **FLOATING
C30 S.n20 SUB 5.38fF $ **FLOATING
C31 S.n21 SUB 2.17fF $ **FLOATING
C32 S.n22 SUB 0.96fF $ **FLOATING
C33 S.n23 SUB 0.94fF $ **FLOATING
C34 S.n24 SUB 0.34fF $ **FLOATING
C35 S.n25 SUB 0.46fF $ **FLOATING
C36 S.n26 SUB 0.33fF $ **FLOATING
C37 S.n27 SUB 9.44fF $ **FLOATING
C38 S.n28 SUB 1.49fF $ **FLOATING
C39 S.n29 SUB 2.63fF $ **FLOATING
C40 S.n30 SUB 8.97fF $ **FLOATING
C41 S.n31 SUB 8.97fF $ **FLOATING
C42 S.n32 SUB 5.38fF $ **FLOATING
C43 S.n33 SUB 2.17fF $ **FLOATING
C44 S.n34 SUB 0.96fF $ **FLOATING
C45 S.n35 SUB 0.94fF $ **FLOATING
C46 S.n36 SUB 0.34fF $ **FLOATING
C47 S.n37 SUB 0.46fF $ **FLOATING
C48 S.n38 SUB 0.33fF $ **FLOATING
C49 S.n39 SUB 9.44fF $ **FLOATING
C50 S.n40 SUB 0.18fF $ **FLOATING
C51 S.n41 SUB 0.10fF $ **FLOATING
C52 S.n42 SUB 0.77fF $ **FLOATING
C53 S.n43 SUB 0.21fF $ **FLOATING
C54 S.n44 SUB 0.36fF $ **FLOATING
C55 S.n45 SUB 0.53fF $ **FLOATING
C56 S.n46 SUB 0.12fF $ **FLOATING
C57 S.t2391 SUB 0.02fF
C58 S.n47 SUB 0.14fF $ **FLOATING
C59 S.t2461 SUB 0.02fF
C60 S.n49 SUB 0.12fF $ **FLOATING
C61 S.n50 SUB 0.14fF $ **FLOATING
C62 S.t1268 SUB 0.02fF
C63 S.n52 SUB 0.24fF $ **FLOATING
C64 S.n53 SUB 0.91fF $ **FLOATING
C65 S.n54 SUB 0.05fF $ **FLOATING
C66 S.t426 SUB 0.02fF
C67 S.n55 SUB 0.24fF $ **FLOATING
C68 S.n56 SUB 0.36fF $ **FLOATING
C69 S.n57 SUB 0.61fF $ **FLOATING
C70 S.n58 SUB 2.48fF $ **FLOATING
C71 S.n59 SUB 1.96fF $ **FLOATING
C72 S.n60 SUB 1.49fF $ **FLOATING
C73 S.n61 SUB 2.63fF $ **FLOATING
C74 S.n62 SUB 8.97fF $ **FLOATING
C75 S.n63 SUB 8.97fF $ **FLOATING
C76 S.n64 SUB 5.38fF $ **FLOATING
C77 S.n65 SUB 2.17fF $ **FLOATING
C78 S.n66 SUB 0.96fF $ **FLOATING
C79 S.n67 SUB 0.94fF $ **FLOATING
C80 S.n68 SUB 0.34fF $ **FLOATING
C81 S.n69 SUB 0.46fF $ **FLOATING
C82 S.n70 SUB 0.33fF $ **FLOATING
C83 S.n71 SUB 9.44fF $ **FLOATING
C84 S.n72 SUB 1.49fF $ **FLOATING
C85 S.n73 SUB 2.63fF $ **FLOATING
C86 S.n74 SUB 8.97fF $ **FLOATING
C87 S.n75 SUB 8.97fF $ **FLOATING
C88 S.n76 SUB 5.38fF $ **FLOATING
C89 S.n77 SUB 2.17fF $ **FLOATING
C90 S.n78 SUB 0.96fF $ **FLOATING
C91 S.n79 SUB 0.94fF $ **FLOATING
C92 S.n80 SUB 0.34fF $ **FLOATING
C93 S.n81 SUB 0.46fF $ **FLOATING
C94 S.n82 SUB 0.33fF $ **FLOATING
C95 S.n83 SUB 9.44fF $ **FLOATING
C96 S.n84 SUB 1.49fF $ **FLOATING
C97 S.n85 SUB 2.63fF $ **FLOATING
C98 S.n86 SUB 8.97fF $ **FLOATING
C99 S.n87 SUB 8.97fF $ **FLOATING
C100 S.n88 SUB 5.38fF $ **FLOATING
C101 S.n89 SUB 2.17fF $ **FLOATING
C102 S.n90 SUB 13.61fF $ **FLOATING
C103 S.n91 SUB 13.61fF $ **FLOATING
C104 S.n92 SUB 5.33fF $ **FLOATING
C105 S.n93 SUB 2.04fF $ **FLOATING
C106 S.n94 SUB 16.47fF $ **FLOATING
C107 S.n95 SUB 1.95fF $ **FLOATING
C108 S.n96 SUB 2.63fF $ **FLOATING
C109 S.n97 SUB 0.96fF $ **FLOATING
C110 S.n98 SUB 0.34fF $ **FLOATING
C111 S.n99 SUB 0.43fF $ **FLOATING
C112 S.n100 SUB 0.30fF $ **FLOATING
C113 S.n101 SUB 0.96fF $ **FLOATING
C114 S.t2099 SUB 0.02fF
C115 S.n102 SUB 1.31fF $ **FLOATING
C116 S.n103 SUB 54.08fF $ **FLOATING
C117 S.n104 SUB 2.23fF $ **FLOATING
C118 S.n105 SUB 0.35fF $ **FLOATING
C119 S.n106 SUB 0.62fF $ **FLOATING
C120 S.n107 SUB 0.53fF $ **FLOATING
C121 S.n108 SUB 3.66fF $ **FLOATING
C122 S.n109 SUB 4.25fF $ **FLOATING
C123 S.n110 SUB 4.22fF $ **FLOATING
C124 S.n111 SUB 4.22fF $ **FLOATING
C125 S.n112 SUB 4.22fF $ **FLOATING
C126 S.n113 SUB 4.22fF $ **FLOATING
C127 S.n114 SUB 4.22fF $ **FLOATING
C128 S.n115 SUB 4.22fF $ **FLOATING
C129 S.n116 SUB 4.70fF $ **FLOATING
C130 S.n117 SUB 4.30fF $ **FLOATING
C131 S.n118 SUB 4.28fF $ **FLOATING
C132 S.n119 SUB 130.19fF $ **FLOATING
C133 S.n120 SUB 2.19fF $ **FLOATING
C134 S.n121 SUB 12.90fF $ **FLOATING
C135 S.n122 SUB 1.90fF $ **FLOATING
C136 S.n123 SUB 9.41fF $ **FLOATING
C137 S.n124 SUB 0.25fF $ **FLOATING
C138 S.t1831 SUB 0.02fF
C139 S.n125 SUB 0.44fF $ **FLOATING
C140 S.n126 SUB 8.97fF $ **FLOATING
C141 S.n127 SUB 8.97fF $ **FLOATING
C142 S.n128 SUB 5.46fF $ **FLOATING
C143 S.n129 SUB 1.96fF $ **FLOATING
C144 S.t29 SUB 0.02fF
C145 S.n130 SUB 0.89fF $ **FLOATING
C146 S.t732 SUB 0.02fF
C147 S.n131 SUB 0.89fF $ **FLOATING
C148 S.n132 SUB 9.44fF $ **FLOATING
C149 S.n133 SUB 3.27fF $ **FLOATING
C150 S.n134 SUB 0.38fF $ **FLOATING
C151 S.n135 SUB 0.31fF $ **FLOATING
C152 S.n136 SUB 1.00fF $ **FLOATING
C153 S.n137 SUB 0.02fF $ **FLOATING
C154 S.t350 SUB 0.02fF
C155 S.n138 SUB 0.37fF $ **FLOATING
C156 S.n139 SUB 8.97fF $ **FLOATING
C157 S.n140 SUB 8.97fF $ **FLOATING
C158 S.n141 SUB 5.46fF $ **FLOATING
C159 S.n142 SUB 1.96fF $ **FLOATING
C160 S.t858 SUB 0.02fF
C161 S.n143 SUB 0.89fF $ **FLOATING
C162 S.t1642 SUB 0.02fF
C163 S.n144 SUB 0.89fF $ **FLOATING
C164 S.n145 SUB 9.44fF $ **FLOATING
C165 S.n146 SUB 3.27fF $ **FLOATING
C166 S.n147 SUB 0.38fF $ **FLOATING
C167 S.n148 SUB 0.31fF $ **FLOATING
C168 S.n149 SUB 1.00fF $ **FLOATING
C169 S.n150 SUB 0.02fF $ **FLOATING
C170 S.t1154 SUB 0.02fF
C171 S.n151 SUB 0.37fF $ **FLOATING
C172 S.n152 SUB 8.97fF $ **FLOATING
C173 S.n153 SUB 8.97fF $ **FLOATING
C174 S.n154 SUB 5.46fF $ **FLOATING
C175 S.n155 SUB 1.96fF $ **FLOATING
C176 S.t1626 SUB 0.02fF
C177 S.n156 SUB 0.89fF $ **FLOATING
C178 S.t2425 SUB 0.02fF
C179 S.n157 SUB 0.89fF $ **FLOATING
C180 S.n158 SUB 9.44fF $ **FLOATING
C181 S.n159 SUB 3.27fF $ **FLOATING
C182 S.n160 SUB 0.38fF $ **FLOATING
C183 S.n161 SUB 0.31fF $ **FLOATING
C184 S.n162 SUB 1.00fF $ **FLOATING
C185 S.n163 SUB 0.02fF $ **FLOATING
C186 S.t1942 SUB 0.02fF
C187 S.n164 SUB 0.37fF $ **FLOATING
C188 S.n165 SUB 8.97fF $ **FLOATING
C189 S.n166 SUB 8.97fF $ **FLOATING
C190 S.n167 SUB 5.46fF $ **FLOATING
C191 S.n168 SUB 1.96fF $ **FLOATING
C192 S.t729 SUB 0.02fF
C193 S.n169 SUB 0.89fF $ **FLOATING
C194 S.t696 SUB 0.02fF
C195 S.n170 SUB 0.89fF $ **FLOATING
C196 S.n171 SUB 9.44fF $ **FLOATING
C197 S.n172 SUB 3.27fF $ **FLOATING
C198 S.n173 SUB 0.38fF $ **FLOATING
C199 S.n174 SUB 0.31fF $ **FLOATING
C200 S.n175 SUB 1.00fF $ **FLOATING
C201 S.n176 SUB 0.02fF $ **FLOATING
C202 S.t2516 SUB 0.02fF
C203 S.n177 SUB 0.37fF $ **FLOATING
C204 S.n178 SUB 8.97fF $ **FLOATING
C205 S.n179 SUB 8.97fF $ **FLOATING
C206 S.n180 SUB 5.46fF $ **FLOATING
C207 S.n181 SUB 1.96fF $ **FLOATING
C208 S.t1528 SUB 0.02fF
C209 S.n182 SUB 0.89fF $ **FLOATING
C210 S.t2226 SUB 0.02fF
C211 S.n183 SUB 0.89fF $ **FLOATING
C212 S.n184 SUB 3.27fF $ **FLOATING
C213 S.n185 SUB 0.38fF $ **FLOATING
C214 S.n186 SUB 0.31fF $ **FLOATING
C215 S.n187 SUB 1.00fF $ **FLOATING
C216 S.n188 SUB 0.02fF $ **FLOATING
C217 S.t772 SUB 0.02fF
C218 S.n189 SUB 0.37fF $ **FLOATING
C219 S.n190 SUB 8.97fF $ **FLOATING
C220 S.n191 SUB 8.97fF $ **FLOATING
C221 S.n192 SUB 5.46fF $ **FLOATING
C222 S.n193 SUB 1.96fF $ **FLOATING
C223 S.t2322 SUB 0.02fF
C224 S.n194 SUB 0.89fF $ **FLOATING
C225 S.t491 SUB 0.02fF
C226 S.n195 SUB 0.89fF $ **FLOATING
C227 S.n196 SUB 3.27fF $ **FLOATING
C228 S.n197 SUB 0.38fF $ **FLOATING
C229 S.n198 SUB 0.31fF $ **FLOATING
C230 S.n199 SUB 1.00fF $ **FLOATING
C231 S.n200 SUB 0.02fF $ **FLOATING
C232 S.t1557 SUB 0.02fF
C233 S.n201 SUB 0.37fF $ **FLOATING
C234 S.n202 SUB 0.31fF $ **FLOATING
C235 S.n203 SUB 8.97fF $ **FLOATING
C236 S.n204 SUB 8.97fF $ **FLOATING
C237 S.n205 SUB 5.22fF $ **FLOATING
C238 S.n206 SUB 1.00fF $ **FLOATING
C239 S.n207 SUB 0.35fF $ **FLOATING
C240 S.t603 SUB 0.02fF
C241 S.n208 SUB 0.89fF $ **FLOATING
C242 S.t1409 SUB 0.02fF
C243 S.n209 SUB 0.89fF $ **FLOATING
C244 S.n210 SUB 3.26fF $ **FLOATING
C245 S.n211 SUB 0.27fF $ **FLOATING
C246 S.n212 SUB 1.05fF $ **FLOATING
C247 S.n213 SUB 1.14fF $ **FLOATING
C248 S.n214 SUB 0.42fF $ **FLOATING
C249 S.n215 SUB 0.02fF $ **FLOATING
C250 S.t2354 SUB 0.02fF
C251 S.n216 SUB 0.37fF $ **FLOATING
C252 S.n217 SUB 0.37fF $ **FLOATING
C253 S.n218 SUB 0.83fF $ **FLOATING
C254 S.t2256 SUB 0.02fF
C255 S.n219 SUB 0.89fF $ **FLOATING
C256 S.t543 SUB 0.02fF
C257 S.n220 SUB 0.89fF $ **FLOATING
C258 S.n221 SUB 0.04fF $ **FLOATING
C259 S.n222 SUB 0.49fF $ **FLOATING
C260 S.n223 SUB 0.38fF $ **FLOATING
C261 S.n224 SUB 0.12fF $ **FLOATING
C262 S.t1258 SUB 0.02fF
C263 S.n225 SUB 0.14fF $ **FLOATING
C264 S.n227 SUB 0.65fF $ **FLOATING
C265 S.n228 SUB 0.44fF $ **FLOATING
C266 S.n229 SUB 1.62fF $ **FLOATING
C267 S.n230 SUB 0.50fF $ **FLOATING
C268 S.n231 SUB 0.46fF $ **FLOATING
C269 S.n232 SUB 0.45fF $ **FLOATING
C270 S.n233 SUB 1.84fF $ **FLOATING
C271 S.n234 SUB 0.12fF $ **FLOATING
C272 S.t1563 SUB 0.02fF
C273 S.n235 SUB 0.14fF $ **FLOATING
C274 S.t2125 SUB 0.02fF
C275 S.n237 SUB 0.24fF $ **FLOATING
C276 S.n238 SUB 0.36fF $ **FLOATING
C277 S.n239 SUB 0.61fF $ **FLOATING
C278 S.n240 SUB 2.49fF $ **FLOATING
C279 S.n241 SUB 2.02fF $ **FLOATING
C280 S.t434 SUB 0.02fF
C281 S.n242 SUB 0.24fF $ **FLOATING
C282 S.n243 SUB 0.91fF $ **FLOATING
C283 S.n244 SUB 0.05fF $ **FLOATING
C284 S.t1789 SUB 0.02fF
C285 S.n245 SUB 0.12fF $ **FLOATING
C286 S.n246 SUB 0.14fF $ **FLOATING
C287 S.n248 SUB 0.18fF $ **FLOATING
C288 S.n249 SUB 0.10fF $ **FLOATING
C289 S.n250 SUB 0.77fF $ **FLOATING
C290 S.n251 SUB 0.21fF $ **FLOATING
C291 S.n252 SUB 0.36fF $ **FLOATING
C292 S.n253 SUB 0.53fF $ **FLOATING
C293 S.n254 SUB 0.12fF $ **FLOATING
C294 S.t831 SUB 0.02fF
C295 S.n255 SUB 0.14fF $ **FLOATING
C296 S.t1398 SUB 0.02fF
C297 S.n257 SUB 0.24fF $ **FLOATING
C298 S.n258 SUB 0.36fF $ **FLOATING
C299 S.n259 SUB 0.61fF $ **FLOATING
C300 S.n260 SUB 2.48fF $ **FLOATING
C301 S.n261 SUB 1.96fF $ **FLOATING
C302 S.t2225 SUB 0.02fF
C303 S.n262 SUB 0.24fF $ **FLOATING
C304 S.n263 SUB 0.91fF $ **FLOATING
C305 S.n264 SUB 0.05fF $ **FLOATING
C306 S.t919 SUB 0.02fF
C307 S.n265 SUB 0.12fF $ **FLOATING
C308 S.n266 SUB 0.14fF $ **FLOATING
C309 S.n268 SUB 0.65fF $ **FLOATING
C310 S.n269 SUB 0.44fF $ **FLOATING
C311 S.n270 SUB 1.62fF $ **FLOATING
C312 S.n271 SUB 0.50fF $ **FLOATING
C313 S.n272 SUB 0.46fF $ **FLOATING
C314 S.n273 SUB 0.45fF $ **FLOATING
C315 S.n274 SUB 1.84fF $ **FLOATING
C316 S.n275 SUB 0.12fF $ **FLOATING
C317 S.t2477 SUB 0.02fF
C318 S.n276 SUB 0.14fF $ **FLOATING
C319 S.t527 SUB 0.02fF
C320 S.n278 SUB 0.24fF $ **FLOATING
C321 S.n279 SUB 0.36fF $ **FLOATING
C322 S.n280 SUB 0.61fF $ **FLOATING
C323 S.n281 SUB 2.49fF $ **FLOATING
C324 S.n282 SUB 2.02fF $ **FLOATING
C325 S.t1364 SUB 0.02fF
C326 S.n283 SUB 0.24fF $ **FLOATING
C327 S.n284 SUB 0.91fF $ **FLOATING
C328 S.n285 SUB 0.05fF $ **FLOATING
C329 S.t2561 SUB 0.02fF
C330 S.n286 SUB 0.12fF $ **FLOATING
C331 S.n287 SUB 0.14fF $ **FLOATING
C332 S.n289 SUB 0.18fF $ **FLOATING
C333 S.n290 SUB 0.10fF $ **FLOATING
C334 S.n291 SUB 0.77fF $ **FLOATING
C335 S.n292 SUB 0.21fF $ **FLOATING
C336 S.n293 SUB 0.36fF $ **FLOATING
C337 S.n294 SUB 0.53fF $ **FLOATING
C338 S.n295 SUB 0.12fF $ **FLOATING
C339 S.t1606 SUB 0.02fF
C340 S.n296 SUB 0.14fF $ **FLOATING
C341 S.t2172 SUB 0.02fF
C342 S.n298 SUB 0.24fF $ **FLOATING
C343 S.n299 SUB 0.36fF $ **FLOATING
C344 S.n300 SUB 0.61fF $ **FLOATING
C345 S.n301 SUB 2.48fF $ **FLOATING
C346 S.n302 SUB 1.96fF $ **FLOATING
C347 S.t490 SUB 0.02fF
C348 S.n303 SUB 0.24fF $ **FLOATING
C349 S.n304 SUB 0.91fF $ **FLOATING
C350 S.n305 SUB 0.05fF $ **FLOATING
C351 S.t1687 SUB 0.02fF
C352 S.n306 SUB 0.12fF $ **FLOATING
C353 S.n307 SUB 0.14fF $ **FLOATING
C354 S.n309 SUB 0.65fF $ **FLOATING
C355 S.n310 SUB 0.44fF $ **FLOATING
C356 S.n311 SUB 1.62fF $ **FLOATING
C357 S.n312 SUB 0.50fF $ **FLOATING
C358 S.n313 SUB 0.46fF $ **FLOATING
C359 S.n314 SUB 0.45fF $ **FLOATING
C360 S.n315 SUB 1.84fF $ **FLOATING
C361 S.n316 SUB 0.12fF $ **FLOATING
C362 S.t742 SUB 0.02fF
C363 S.n317 SUB 0.14fF $ **FLOATING
C364 S.t1309 SUB 0.02fF
C365 S.n319 SUB 0.24fF $ **FLOATING
C366 S.n320 SUB 0.36fF $ **FLOATING
C367 S.n321 SUB 0.61fF $ **FLOATING
C368 S.n322 SUB 2.49fF $ **FLOATING
C369 S.n323 SUB 2.02fF $ **FLOATING
C370 S.t2133 SUB 0.02fF
C371 S.n324 SUB 0.24fF $ **FLOATING
C372 S.n325 SUB 0.91fF $ **FLOATING
C373 S.n326 SUB 0.05fF $ **FLOATING
C374 S.t814 SUB 0.02fF
C375 S.n327 SUB 0.12fF $ **FLOATING
C376 S.n328 SUB 0.14fF $ **FLOATING
C377 S.n330 SUB 0.65fF $ **FLOATING
C378 S.n331 SUB 0.44fF $ **FLOATING
C379 S.n332 SUB 1.62fF $ **FLOATING
C380 S.n333 SUB 0.50fF $ **FLOATING
C381 S.n334 SUB 0.46fF $ **FLOATING
C382 S.n335 SUB 0.45fF $ **FLOATING
C383 S.n336 SUB 1.84fF $ **FLOATING
C384 S.n337 SUB 0.12fF $ **FLOATING
C385 S.t1534 SUB 0.02fF
C386 S.n338 SUB 0.14fF $ **FLOATING
C387 S.t2074 SUB 0.02fF
C388 S.n340 SUB 0.24fF $ **FLOATING
C389 S.n341 SUB 0.36fF $ **FLOATING
C390 S.n342 SUB 0.61fF $ **FLOATING
C391 S.n343 SUB 2.49fF $ **FLOATING
C392 S.n344 SUB 2.02fF $ **FLOATING
C393 S.t386 SUB 0.02fF
C394 S.n345 SUB 0.24fF $ **FLOATING
C395 S.n346 SUB 0.91fF $ **FLOATING
C396 S.n347 SUB 0.05fF $ **FLOATING
C397 S.t1742 SUB 0.02fF
C398 S.n348 SUB 0.12fF $ **FLOATING
C399 S.n349 SUB 0.14fF $ **FLOATING
C400 S.n351 SUB 0.18fF $ **FLOATING
C401 S.n352 SUB 0.10fF $ **FLOATING
C402 S.n353 SUB 0.77fF $ **FLOATING
C403 S.n354 SUB 0.21fF $ **FLOATING
C404 S.n355 SUB 0.36fF $ **FLOATING
C405 S.n356 SUB 0.53fF $ **FLOATING
C406 S.n357 SUB 0.12fF $ **FLOATING
C407 S.t1299 SUB 0.02fF
C408 S.n358 SUB 0.14fF $ **FLOATING
C409 S.t1846 SUB 0.02fF
C410 S.n360 SUB 0.24fF $ **FLOATING
C411 S.n361 SUB 0.36fF $ **FLOATING
C412 S.n362 SUB 0.61fF $ **FLOATING
C413 S.n363 SUB 2.48fF $ **FLOATING
C414 S.n364 SUB 1.96fF $ **FLOATING
C415 S.t1728 SUB 0.02fF
C416 S.n365 SUB 0.24fF $ **FLOATING
C417 S.n366 SUB 0.91fF $ **FLOATING
C418 S.n367 SUB 0.05fF $ **FLOATING
C419 S.t1482 SUB 0.02fF
C420 S.n368 SUB 0.12fF $ **FLOATING
C421 S.n369 SUB 0.14fF $ **FLOATING
C422 S.n371 SUB 0.65fF $ **FLOATING
C423 S.n372 SUB 0.44fF $ **FLOATING
C424 S.n373 SUB 1.62fF $ **FLOATING
C425 S.n374 SUB 0.50fF $ **FLOATING
C426 S.n375 SUB 0.46fF $ **FLOATING
C427 S.n376 SUB 0.45fF $ **FLOATING
C428 S.n377 SUB 1.84fF $ **FLOATING
C429 S.n378 SUB 0.12fF $ **FLOATING
C430 S.t416 SUB 0.02fF
C431 S.n379 SUB 0.14fF $ **FLOATING
C432 S.t984 SUB 0.02fF
C433 S.n381 SUB 0.24fF $ **FLOATING
C434 S.n382 SUB 0.36fF $ **FLOATING
C435 S.n383 SUB 0.61fF $ **FLOATING
C436 S.n384 SUB 2.49fF $ **FLOATING
C437 S.n385 SUB 2.02fF $ **FLOATING
C438 S.t855 SUB 0.02fF
C439 S.n386 SUB 0.24fF $ **FLOATING
C440 S.n387 SUB 0.91fF $ **FLOATING
C441 S.n388 SUB 0.05fF $ **FLOATING
C442 S.t621 SUB 0.02fF
C443 S.n389 SUB 0.12fF $ **FLOATING
C444 S.n390 SUB 0.14fF $ **FLOATING
C445 S.n392 SUB 0.18fF $ **FLOATING
C446 S.n393 SUB 0.10fF $ **FLOATING
C447 S.n394 SUB 0.77fF $ **FLOATING
C448 S.n395 SUB 0.21fF $ **FLOATING
C449 S.n396 SUB 0.36fF $ **FLOATING
C450 S.n397 SUB 0.53fF $ **FLOATING
C451 S.n398 SUB 0.12fF $ **FLOATING
C452 S.t2066 SUB 0.02fF
C453 S.n399 SUB 0.14fF $ **FLOATING
C454 S.t62 SUB 0.02fF
C455 S.n401 SUB 0.24fF $ **FLOATING
C456 S.n402 SUB 0.36fF $ **FLOATING
C457 S.n403 SUB 0.61fF $ **FLOATING
C458 S.n404 SUB 2.48fF $ **FLOATING
C459 S.n405 SUB 1.96fF $ **FLOATING
C460 S.t2499 SUB 0.02fF
C461 S.n406 SUB 0.24fF $ **FLOATING
C462 S.n407 SUB 0.91fF $ **FLOATING
C463 S.n408 SUB 0.05fF $ **FLOATING
C464 S.t2279 SUB 0.02fF
C465 S.n409 SUB 0.12fF $ **FLOATING
C466 S.n410 SUB 0.14fF $ **FLOATING
C467 S.n412 SUB 0.65fF $ **FLOATING
C468 S.n413 SUB 0.44fF $ **FLOATING
C469 S.n414 SUB 1.62fF $ **FLOATING
C470 S.n415 SUB 0.50fF $ **FLOATING
C471 S.n416 SUB 0.46fF $ **FLOATING
C472 S.n417 SUB 0.45fF $ **FLOATING
C473 S.n418 SUB 1.84fF $ **FLOATING
C474 S.n419 SUB 0.12fF $ **FLOATING
C475 S.t1204 SUB 0.02fF
C476 S.n420 SUB 0.14fF $ **FLOATING
C477 S.t1749 SUB 0.02fF
C478 S.n422 SUB 0.24fF $ **FLOATING
C479 S.n423 SUB 0.36fF $ **FLOATING
C480 S.n424 SUB 0.61fF $ **FLOATING
C481 S.n425 SUB 2.49fF $ **FLOATING
C482 S.n426 SUB 2.02fF $ **FLOATING
C483 S.t1624 SUB 0.02fF
C484 S.n427 SUB 0.24fF $ **FLOATING
C485 S.n428 SUB 0.91fF $ **FLOATING
C486 S.n429 SUB 0.05fF $ **FLOATING
C487 S.t1424 SUB 0.02fF
C488 S.n430 SUB 0.12fF $ **FLOATING
C489 S.n431 SUB 0.14fF $ **FLOATING
C490 S.n433 SUB 0.18fF $ **FLOATING
C491 S.n434 SUB 0.10fF $ **FLOATING
C492 S.n435 SUB 0.77fF $ **FLOATING
C493 S.n436 SUB 0.21fF $ **FLOATING
C494 S.n437 SUB 0.36fF $ **FLOATING
C495 S.n438 SUB 0.53fF $ **FLOATING
C496 S.n439 SUB 0.12fF $ **FLOATING
C497 S.t473 SUB 0.02fF
C498 S.n440 SUB 0.14fF $ **FLOATING
C499 S.t1032 SUB 0.02fF
C500 S.n442 SUB 0.24fF $ **FLOATING
C501 S.n443 SUB 0.36fF $ **FLOATING
C502 S.n444 SUB 0.61fF $ **FLOATING
C503 S.n445 SUB 2.48fF $ **FLOATING
C504 S.n446 SUB 1.96fF $ **FLOATING
C505 S.t915 SUB 0.02fF
C506 S.n447 SUB 0.24fF $ **FLOATING
C507 S.n448 SUB 0.91fF $ **FLOATING
C508 S.n449 SUB 0.05fF $ **FLOATING
C509 S.t557 SUB 0.02fF
C510 S.n450 SUB 0.12fF $ **FLOATING
C511 S.n451 SUB 0.14fF $ **FLOATING
C512 S.n453 SUB 1.89fF $ **FLOATING
C513 S.n454 SUB 0.12fF $ **FLOATING
C514 S.t622 SUB 0.02fF
C515 S.n455 SUB 0.14fF $ **FLOATING
C516 S.t1828 SUB 0.02fF
C517 S.n457 SUB 1.22fF $ **FLOATING
C518 S.n458 SUB 2.29fF $ **FLOATING
C519 S.n459 SUB 0.61fF $ **FLOATING
C520 S.n460 SUB 0.35fF $ **FLOATING
C521 S.n461 SUB 0.63fF $ **FLOATING
C522 S.n462 SUB 1.15fF $ **FLOATING
C523 S.n463 SUB 3.03fF $ **FLOATING
C524 S.n464 SUB 0.59fF $ **FLOATING
C525 S.n465 SUB 0.02fF $ **FLOATING
C526 S.n466 SUB 0.97fF $ **FLOATING
C527 S.t20 SUB 21.38fF
C528 S.n467 SUB 20.25fF $ **FLOATING
C529 S.n469 SUB 0.38fF $ **FLOATING
C530 S.n470 SUB 0.23fF $ **FLOATING
C531 S.n471 SUB 2.89fF $ **FLOATING
C532 S.n472 SUB 2.46fF $ **FLOATING
C533 S.n473 SUB 4.30fF $ **FLOATING
C534 S.n474 SUB 0.25fF $ **FLOATING
C535 S.n475 SUB 0.01fF $ **FLOATING
C536 S.t1521 SUB 0.02fF
C537 S.n476 SUB 0.25fF $ **FLOATING
C538 S.t1276 SUB 0.02fF
C539 S.n477 SUB 0.95fF $ **FLOATING
C540 S.n478 SUB 0.70fF $ **FLOATING
C541 S.n479 SUB 1.89fF $ **FLOATING
C542 S.n480 SUB 1.78fF $ **FLOATING
C543 S.n481 SUB 0.12fF $ **FLOATING
C544 S.t659 SUB 0.02fF
C545 S.n482 SUB 0.14fF $ **FLOATING
C546 S.t962 SUB 0.02fF
C547 S.n484 SUB 0.24fF $ **FLOATING
C548 S.n485 SUB 0.36fF $ **FLOATING
C549 S.n486 SUB 0.61fF $ **FLOATING
C550 S.n487 SUB 2.74fF $ **FLOATING
C551 S.n488 SUB 2.05fF $ **FLOATING
C552 S.t389 SUB 0.02fF
C553 S.n489 SUB 0.24fF $ **FLOATING
C554 S.n490 SUB 0.91fF $ **FLOATING
C555 S.n491 SUB 0.05fF $ **FLOATING
C556 S.t1356 SUB 0.02fF
C557 S.n492 SUB 0.12fF $ **FLOATING
C558 S.n493 SUB 0.14fF $ **FLOATING
C559 S.n495 SUB 1.24fF $ **FLOATING
C560 S.n496 SUB 1.28fF $ **FLOATING
C561 S.n497 SUB 1.88fF $ **FLOATING
C562 S.n498 SUB 0.12fF $ **FLOATING
C563 S.t2313 SUB 0.02fF
C564 S.n499 SUB 0.14fF $ **FLOATING
C565 S.t21 SUB 0.02fF
C566 S.n501 SUB 0.24fF $ **FLOATING
C567 S.n502 SUB 0.36fF $ **FLOATING
C568 S.n503 SUB 0.61fF $ **FLOATING
C569 S.n504 SUB 2.75fF $ **FLOATING
C570 S.n505 SUB 2.17fF $ **FLOATING
C571 S.t2039 SUB 0.02fF
C572 S.n506 SUB 0.24fF $ **FLOATING
C573 S.n507 SUB 0.91fF $ **FLOATING
C574 S.n508 SUB 0.05fF $ **FLOATING
C575 S.t478 SUB 0.02fF
C576 S.n509 SUB 0.12fF $ **FLOATING
C577 S.n510 SUB 0.14fF $ **FLOATING
C578 S.n512 SUB 1.89fF $ **FLOATING
C579 S.n513 SUB 1.79fF $ **FLOATING
C580 S.n514 SUB 0.12fF $ **FLOATING
C581 S.t1455 SUB 0.02fF
C582 S.n515 SUB 0.14fF $ **FLOATING
C583 S.t1727 SUB 0.02fF
C584 S.n517 SUB 0.24fF $ **FLOATING
C585 S.n518 SUB 0.36fF $ **FLOATING
C586 S.n519 SUB 0.61fF $ **FLOATING
C587 S.n520 SUB 2.73fF $ **FLOATING
C588 S.n521 SUB 2.05fF $ **FLOATING
C589 S.t1185 SUB 0.02fF
C590 S.n522 SUB 0.24fF $ **FLOATING
C591 S.n523 SUB 0.91fF $ **FLOATING
C592 S.n524 SUB 0.05fF $ **FLOATING
C593 S.t2260 SUB 0.02fF
C594 S.n525 SUB 0.12fF $ **FLOATING
C595 S.n526 SUB 0.14fF $ **FLOATING
C596 S.n528 SUB 1.24fF $ **FLOATING
C597 S.n529 SUB 1.28fF $ **FLOATING
C598 S.n530 SUB 1.88fF $ **FLOATING
C599 S.n531 SUB 0.12fF $ **FLOATING
C600 S.t597 SUB 0.02fF
C601 S.n532 SUB 0.14fF $ **FLOATING
C602 S.t854 SUB 0.02fF
C603 S.n534 SUB 0.24fF $ **FLOATING
C604 S.n535 SUB 0.36fF $ **FLOATING
C605 S.n536 SUB 0.61fF $ **FLOATING
C606 S.n537 SUB 2.75fF $ **FLOATING
C607 S.n538 SUB 2.17fF $ **FLOATING
C608 S.t310 SUB 0.02fF
C609 S.n539 SUB 0.24fF $ **FLOATING
C610 S.n540 SUB 0.91fF $ **FLOATING
C611 S.n541 SUB 0.05fF $ **FLOATING
C612 S.t1403 SUB 0.02fF
C613 S.n542 SUB 0.12fF $ **FLOATING
C614 S.n543 SUB 0.14fF $ **FLOATING
C615 S.n545 SUB 1.89fF $ **FLOATING
C616 S.n546 SUB 1.79fF $ **FLOATING
C617 S.n547 SUB 0.12fF $ **FLOATING
C618 S.t2247 SUB 0.02fF
C619 S.n548 SUB 0.14fF $ **FLOATING
C620 S.t2497 SUB 0.02fF
C621 S.n550 SUB 0.24fF $ **FLOATING
C622 S.n551 SUB 0.36fF $ **FLOATING
C623 S.n552 SUB 0.61fF $ **FLOATING
C624 S.n553 SUB 2.73fF $ **FLOATING
C625 S.n554 SUB 2.05fF $ **FLOATING
C626 S.t1972 SUB 0.02fF
C627 S.n555 SUB 0.24fF $ **FLOATING
C628 S.n556 SUB 0.91fF $ **FLOATING
C629 S.n557 SUB 0.05fF $ **FLOATING
C630 S.t532 SUB 0.02fF
C631 S.n558 SUB 0.12fF $ **FLOATING
C632 S.n559 SUB 0.14fF $ **FLOATING
C633 S.n561 SUB 1.24fF $ **FLOATING
C634 S.n562 SUB 1.28fF $ **FLOATING
C635 S.n563 SUB 1.88fF $ **FLOATING
C636 S.n564 SUB 0.12fF $ **FLOATING
C637 S.t1388 SUB 0.02fF
C638 S.n565 SUB 0.14fF $ **FLOATING
C639 S.t1620 SUB 0.02fF
C640 S.n567 SUB 0.24fF $ **FLOATING
C641 S.n568 SUB 0.36fF $ **FLOATING
C642 S.n569 SUB 0.61fF $ **FLOATING
C643 S.n570 SUB 2.75fF $ **FLOATING
C644 S.n571 SUB 2.17fF $ **FLOATING
C645 S.t1117 SUB 0.02fF
C646 S.n572 SUB 0.24fF $ **FLOATING
C647 S.n573 SUB 0.91fF $ **FLOATING
C648 S.n574 SUB 0.05fF $ **FLOATING
C649 S.t2175 SUB 0.02fF
C650 S.n575 SUB 0.12fF $ **FLOATING
C651 S.n576 SUB 0.14fF $ **FLOATING
C652 S.n578 SUB 1.89fF $ **FLOATING
C653 S.n579 SUB 1.79fF $ **FLOATING
C654 S.n580 SUB 0.12fF $ **FLOATING
C655 S.t627 SUB 0.02fF
C656 S.n581 SUB 0.14fF $ **FLOATING
C657 S.t755 SUB 0.02fF
C658 S.n583 SUB 0.24fF $ **FLOATING
C659 S.n584 SUB 0.36fF $ **FLOATING
C660 S.n585 SUB 0.61fF $ **FLOATING
C661 S.n586 SUB 2.73fF $ **FLOATING
C662 S.n587 SUB 2.05fF $ **FLOATING
C663 S.t235 SUB 0.02fF
C664 S.n588 SUB 0.24fF $ **FLOATING
C665 S.n589 SUB 0.91fF $ **FLOATING
C666 S.n590 SUB 0.05fF $ **FLOATING
C667 S.t1311 SUB 0.02fF
C668 S.n591 SUB 0.12fF $ **FLOATING
C669 S.n592 SUB 0.14fF $ **FLOATING
C670 S.n594 SUB 1.24fF $ **FLOATING
C671 S.n595 SUB 1.28fF $ **FLOATING
C672 S.n596 SUB 1.88fF $ **FLOATING
C673 S.n597 SUB 0.12fF $ **FLOATING
C674 S.t2406 SUB 0.02fF
C675 S.n598 SUB 0.14fF $ **FLOATING
C676 S.t1678 SUB 0.02fF
C677 S.n600 SUB 0.24fF $ **FLOATING
C678 S.n601 SUB 0.36fF $ **FLOATING
C679 S.n602 SUB 0.61fF $ **FLOATING
C680 S.n603 SUB 2.75fF $ **FLOATING
C681 S.n604 SUB 2.17fF $ **FLOATING
C682 S.t90 SUB 0.02fF
C683 S.n605 SUB 0.24fF $ **FLOATING
C684 S.n606 SUB 0.91fF $ **FLOATING
C685 S.n607 SUB 0.05fF $ **FLOATING
C686 S.t431 SUB 0.02fF
C687 S.n608 SUB 0.12fF $ **FLOATING
C688 S.n609 SUB 0.14fF $ **FLOATING
C689 S.n611 SUB 1.89fF $ **FLOATING
C690 S.n612 SUB 1.79fF $ **FLOATING
C691 S.n613 SUB 0.12fF $ **FLOATING
C692 S.t1544 SUB 0.02fF
C693 S.n614 SUB 0.14fF $ **FLOATING
C694 S.t803 SUB 0.02fF
C695 S.n616 SUB 0.24fF $ **FLOATING
C696 S.n617 SUB 0.36fF $ **FLOATING
C697 S.n618 SUB 0.61fF $ **FLOATING
C698 S.n619 SUB 2.73fF $ **FLOATING
C699 S.n620 SUB 2.05fF $ **FLOATING
C700 S.t1765 SUB 0.02fF
C701 S.n621 SUB 0.24fF $ **FLOATING
C702 S.n622 SUB 0.91fF $ **FLOATING
C703 S.n623 SUB 0.05fF $ **FLOATING
C704 S.t2252 SUB 0.02fF
C705 S.n624 SUB 0.12fF $ **FLOATING
C706 S.n625 SUB 0.14fF $ **FLOATING
C707 S.n627 SUB 1.24fF $ **FLOATING
C708 S.n628 SUB 1.28fF $ **FLOATING
C709 S.n629 SUB 1.88fF $ **FLOATING
C710 S.n630 SUB 0.12fF $ **FLOATING
C711 S.t683 SUB 0.02fF
C712 S.n631 SUB 0.14fF $ **FLOATING
C713 S.t2453 SUB 0.02fF
C714 S.n633 SUB 0.24fF $ **FLOATING
C715 S.n634 SUB 0.36fF $ **FLOATING
C716 S.n635 SUB 0.61fF $ **FLOATING
C717 S.n636 SUB 2.75fF $ **FLOATING
C718 S.n637 SUB 2.17fF $ **FLOATING
C719 S.t891 SUB 0.02fF
C720 S.n638 SUB 0.24fF $ **FLOATING
C721 S.n639 SUB 0.91fF $ **FLOATING
C722 S.n640 SUB 0.05fF $ **FLOATING
C723 S.t1393 SUB 0.02fF
C724 S.n641 SUB 0.12fF $ **FLOATING
C725 S.n642 SUB 0.14fF $ **FLOATING
C726 S.n644 SUB 1.89fF $ **FLOATING
C727 S.n645 SUB 1.79fF $ **FLOATING
C728 S.n646 SUB 0.12fF $ **FLOATING
C729 S.t2342 SUB 0.02fF
C730 S.n647 SUB 0.14fF $ **FLOATING
C731 S.t1585 SUB 0.02fF
C732 S.n649 SUB 0.24fF $ **FLOATING
C733 S.n650 SUB 0.36fF $ **FLOATING
C734 S.n651 SUB 0.61fF $ **FLOATING
C735 S.n652 SUB 2.73fF $ **FLOATING
C736 S.n653 SUB 2.05fF $ **FLOATING
C737 S.t2534 SUB 0.02fF
C738 S.n654 SUB 0.24fF $ **FLOATING
C739 S.n655 SUB 0.91fF $ **FLOATING
C740 S.n656 SUB 0.05fF $ **FLOATING
C741 S.t521 SUB 0.02fF
C742 S.n657 SUB 0.12fF $ **FLOATING
C743 S.n658 SUB 0.14fF $ **FLOATING
C744 S.n660 SUB 1.24fF $ **FLOATING
C745 S.n661 SUB 1.28fF $ **FLOATING
C746 S.n662 SUB 1.88fF $ **FLOATING
C747 S.n663 SUB 0.12fF $ **FLOATING
C748 S.t1483 SUB 0.02fF
C749 S.n664 SUB 0.14fF $ **FLOATING
C750 S.t720 SUB 0.02fF
C751 S.n666 SUB 0.24fF $ **FLOATING
C752 S.n667 SUB 0.36fF $ **FLOATING
C753 S.n668 SUB 0.61fF $ **FLOATING
C754 S.n669 SUB 2.75fF $ **FLOATING
C755 S.n670 SUB 2.17fF $ **FLOATING
C756 S.t1662 SUB 0.02fF
C757 S.n671 SUB 0.24fF $ **FLOATING
C758 S.n672 SUB 0.91fF $ **FLOATING
C759 S.n673 SUB 0.05fF $ **FLOATING
C760 S.t2163 SUB 0.02fF
C761 S.n674 SUB 0.12fF $ **FLOATING
C762 S.n675 SUB 0.14fF $ **FLOATING
C763 S.n677 SUB 2.61fF $ **FLOATING
C764 S.n678 SUB 1.88fF $ **FLOATING
C765 S.n679 SUB 0.12fF $ **FLOATING
C766 S.t2280 SUB 0.02fF
C767 S.n680 SUB 0.14fF $ **FLOATING
C768 S.t1517 SUB 0.02fF
C769 S.n682 SUB 0.24fF $ **FLOATING
C770 S.n683 SUB 0.36fF $ **FLOATING
C771 S.n684 SUB 0.61fF $ **FLOATING
C772 S.n685 SUB 0.90fF $ **FLOATING
C773 S.n686 SUB 0.77fF $ **FLOATING
C774 S.n687 SUB 0.97fF $ **FLOATING
C775 S.n688 SUB 0.09fF $ **FLOATING
C776 S.n689 SUB 0.33fF $ **FLOATING
C777 S.n690 SUB 2.16fF $ **FLOATING
C778 S.t2440 SUB 0.02fF
C779 S.n691 SUB 0.24fF $ **FLOATING
C780 S.n692 SUB 0.91fF $ **FLOATING
C781 S.n693 SUB 0.05fF $ **FLOATING
C782 S.t570 SUB 0.02fF
C783 S.n694 SUB 0.12fF $ **FLOATING
C784 S.n695 SUB 0.14fF $ **FLOATING
C785 S.n697 SUB 2.30fF $ **FLOATING
C786 S.n698 SUB 1.88fF $ **FLOATING
C787 S.n699 SUB 0.12fF $ **FLOATING
C788 S.t1425 SUB 0.02fF
C789 S.n700 SUB 0.14fF $ **FLOATING
C790 S.t656 SUB 0.02fF
C791 S.n702 SUB 0.24fF $ **FLOATING
C792 S.n703 SUB 0.36fF $ **FLOATING
C793 S.n704 SUB 0.61fF $ **FLOATING
C794 S.n705 SUB 0.77fF $ **FLOATING
C795 S.n706 SUB 0.48fF $ **FLOATING
C796 S.n707 SUB 0.09fF $ **FLOATING
C797 S.n708 SUB 0.33fF $ **FLOATING
C798 S.n709 SUB 2.03fF $ **FLOATING
C799 S.t1575 SUB 0.02fF
C800 S.n710 SUB 0.24fF $ **FLOATING
C801 S.n711 SUB 0.91fF $ **FLOATING
C802 S.n712 SUB 0.05fF $ **FLOATING
C803 S.t2214 SUB 0.02fF
C804 S.n713 SUB 0.12fF $ **FLOATING
C805 S.n714 SUB 0.14fF $ **FLOATING
C806 S.n716 SUB 1.89fF $ **FLOATING
C807 S.n717 SUB 0.25fF $ **FLOATING
C808 S.n718 SUB 0.09fF $ **FLOATING
C809 S.n719 SUB 0.23fF $ **FLOATING
C810 S.n720 SUB 1.16fF $ **FLOATING
C811 S.n721 SUB 0.22fF $ **FLOATING
C812 S.n722 SUB 0.12fF $ **FLOATING
C813 S.t559 SUB 0.02fF
C814 S.n723 SUB 0.14fF $ **FLOATING
C815 S.t2310 SUB 0.02fF
C816 S.n725 SUB 0.24fF $ **FLOATING
C817 S.n726 SUB 0.36fF $ **FLOATING
C818 S.n727 SUB 0.61fF $ **FLOATING
C819 S.n728 SUB 2.73fF $ **FLOATING
C820 S.n729 SUB 1.88fF $ **FLOATING
C821 S.t706 SUB 0.02fF
C822 S.n730 SUB 0.24fF $ **FLOATING
C823 S.n731 SUB 0.91fF $ **FLOATING
C824 S.n732 SUB 0.05fF $ **FLOATING
C825 S.t1353 SUB 0.02fF
C826 S.n733 SUB 0.12fF $ **FLOATING
C827 S.n734 SUB 0.14fF $ **FLOATING
C828 S.n736 SUB 20.78fF $ **FLOATING
C829 S.n737 SUB 2.72fF $ **FLOATING
C830 S.n738 SUB 1.95fF $ **FLOATING
C831 S.n739 SUB 0.12fF $ **FLOATING
C832 S.t2289 SUB 0.02fF
C833 S.n740 SUB 0.14fF $ **FLOATING
C834 S.t2366 SUB 0.02fF
C835 S.n742 SUB 0.24fF $ **FLOATING
C836 S.n743 SUB 0.36fF $ **FLOATING
C837 S.n744 SUB 0.61fF $ **FLOATING
C838 S.n745 SUB 1.56fF $ **FLOATING
C839 S.n746 SUB 0.70fF $ **FLOATING
C840 S.n747 SUB 0.28fF $ **FLOATING
C841 S.n748 SUB 2.10fF $ **FLOATING
C842 S.t537 SUB 0.02fF
C843 S.n749 SUB 0.12fF $ **FLOATING
C844 S.n750 SUB 0.14fF $ **FLOATING
C845 S.t197 SUB 0.02fF
C846 S.n752 SUB 0.24fF $ **FLOATING
C847 S.n753 SUB 0.91fF $ **FLOATING
C848 S.n754 SUB 0.05fF $ **FLOATING
C849 S.t430 SUB 48.31fF
C850 S.t1434 SUB 0.02fF
C851 S.n755 SUB 0.12fF $ **FLOATING
C852 S.n756 SUB 0.14fF $ **FLOATING
C853 S.t791 SUB 0.02fF
C854 S.n758 SUB 0.24fF $ **FLOATING
C855 S.n759 SUB 0.91fF $ **FLOATING
C856 S.n760 SUB 0.05fF $ **FLOATING
C857 S.t2373 SUB 0.02fF
C858 S.n761 SUB 0.24fF $ **FLOATING
C859 S.n762 SUB 0.36fF $ **FLOATING
C860 S.n763 SUB 0.61fF $ **FLOATING
C861 S.n764 SUB 2.24fF $ **FLOATING
C862 S.n765 SUB 2.70fF $ **FLOATING
C863 S.n766 SUB 2.65fF $ **FLOATING
C864 S.n767 SUB 2.36fF $ **FLOATING
C865 S.n768 SUB 1.84fF $ **FLOATING
C866 S.n769 SUB 0.12fF $ **FLOATING
C867 S.t2123 SUB 0.02fF
C868 S.n770 SUB 0.14fF $ **FLOATING
C869 S.t135 SUB 0.02fF
C870 S.n772 SUB 0.24fF $ **FLOATING
C871 S.n773 SUB 0.36fF $ **FLOATING
C872 S.n774 SUB 0.61fF $ **FLOATING
C873 S.n775 SUB 0.67fF $ **FLOATING
C874 S.n776 SUB 0.40fF $ **FLOATING
C875 S.n777 SUB 0.55fF $ **FLOATING
C876 S.n778 SUB 0.33fF $ **FLOATING
C877 S.n779 SUB 1.07fF $ **FLOATING
C878 S.n780 SUB 2.13fF $ **FLOATING
C879 S.t2555 SUB 0.02fF
C880 S.n781 SUB 0.24fF $ **FLOATING
C881 S.n782 SUB 0.91fF $ **FLOATING
C882 S.n783 SUB 0.05fF $ **FLOATING
C883 S.t2194 SUB 0.02fF
C884 S.n784 SUB 0.12fF $ **FLOATING
C885 S.n785 SUB 0.14fF $ **FLOATING
C886 S.n787 SUB 0.25fF $ **FLOATING
C887 S.n788 SUB 0.09fF $ **FLOATING
C888 S.n789 SUB 0.12fF $ **FLOATING
C889 S.t373 SUB 0.02fF
C890 S.n790 SUB 0.14fF $ **FLOATING
C891 S.t937 SUB 0.02fF
C892 S.n792 SUB 0.24fF $ **FLOATING
C893 S.n793 SUB 0.36fF $ **FLOATING
C894 S.n794 SUB 0.61fF $ **FLOATING
C895 S.n795 SUB 0.83fF $ **FLOATING
C896 S.n796 SUB 0.32fF $ **FLOATING
C897 S.n797 SUB 0.29fF $ **FLOATING
C898 S.n798 SUB 0.25fF $ **FLOATING
C899 S.n799 SUB 0.22fF $ **FLOATING
C900 S.n800 SUB 0.60fF $ **FLOATING
C901 S.n801 SUB 0.28fF $ **FLOATING
C902 S.n802 SUB 1.94fF $ **FLOATING
C903 S.t809 SUB 0.02fF
C904 S.n803 SUB 0.24fF $ **FLOATING
C905 S.n804 SUB 0.91fF $ **FLOATING
C906 S.n805 SUB 0.05fF $ **FLOATING
C907 S.t459 SUB 0.02fF
C908 S.n806 SUB 0.12fF $ **FLOATING
C909 S.n807 SUB 0.14fF $ **FLOATING
C910 S.n809 SUB 0.19fF $ **FLOATING
C911 S.n810 SUB 0.10fF $ **FLOATING
C912 S.n811 SUB 0.68fF $ **FLOATING
C913 S.n812 SUB 0.28fF $ **FLOATING
C914 S.n813 SUB 1.74fF $ **FLOATING
C915 S.n814 SUB 0.21fF $ **FLOATING
C916 S.n815 SUB 1.84fF $ **FLOATING
C917 S.n816 SUB 0.12fF $ **FLOATING
C918 S.t2422 SUB 0.02fF
C919 S.n817 SUB 0.14fF $ **FLOATING
C920 S.t1202 SUB 0.02fF
C921 S.n819 SUB 0.24fF $ **FLOATING
C922 S.n820 SUB 0.36fF $ **FLOATING
C923 S.n821 SUB 0.61fF $ **FLOATING
C924 S.n822 SUB 2.49fF $ **FLOATING
C925 S.n823 SUB 1.86fF $ **FLOATING
C926 S.t2483 SUB 0.02fF
C927 S.n824 SUB 0.24fF $ **FLOATING
C928 S.n825 SUB 0.91fF $ **FLOATING
C929 S.n826 SUB 0.05fF $ **FLOATING
C930 S.t2105 SUB 0.02fF
C931 S.n827 SUB 0.12fF $ **FLOATING
C932 S.n828 SUB 0.14fF $ **FLOATING
C933 S.n830 SUB 20.78fF $ **FLOATING
C934 S.n831 SUB 0.06fF $ **FLOATING
C935 S.n832 SUB 0.20fF $ **FLOATING
C936 S.n833 SUB 0.09fF $ **FLOATING
C937 S.n834 SUB 0.21fF $ **FLOATING
C938 S.n835 SUB 0.10fF $ **FLOATING
C939 S.n836 SUB 0.30fF $ **FLOATING
C940 S.n837 SUB 1.01fF $ **FLOATING
C941 S.n838 SUB 0.45fF $ **FLOATING
C942 S.n839 SUB 0.12fF $ **FLOATING
C943 S.t2427 SUB 0.02fF
C944 S.n840 SUB 0.14fF $ **FLOATING
C945 S.t475 SUB 0.02fF
C946 S.n842 SUB 0.24fF $ **FLOATING
C947 S.n843 SUB 0.36fF $ **FLOATING
C948 S.n844 SUB 0.61fF $ **FLOATING
C949 S.n845 SUB 0.79fF $ **FLOATING
C950 S.n846 SUB 0.18fF $ **FLOATING
C951 S.n847 SUB 0.39fF $ **FLOATING
C952 S.n848 SUB 0.44fF $ **FLOATING
C953 S.n849 SUB 0.25fF $ **FLOATING
C954 S.n850 SUB 0.09fF $ **FLOATING
C955 S.n851 SUB 1.81fF $ **FLOATING
C956 S.t117 SUB 0.02fF
C957 S.n852 SUB 0.12fF $ **FLOATING
C958 S.n853 SUB 0.14fF $ **FLOATING
C959 S.t1313 SUB 0.02fF
C960 S.n855 SUB 0.24fF $ **FLOATING
C961 S.n856 SUB 0.91fF $ **FLOATING
C962 S.n857 SUB 0.05fF $ **FLOATING
C963 S.n858 SUB 1.14fF $ **FLOATING
C964 S.n859 SUB 8.97fF $ **FLOATING
C965 S.n860 SUB 20.36fF $ **FLOATING
C966 S.n861 SUB 8.97fF $ **FLOATING
C967 S.n862 SUB 20.36fF $ **FLOATING
C968 S.n863 SUB 0.60fF $ **FLOATING
C969 S.n864 SUB 0.22fF $ **FLOATING
C970 S.n865 SUB 0.88fF $ **FLOATING
C971 S.n866 SUB 0.88fF $ **FLOATING
C972 S.n867 SUB 3.43fF $ **FLOATING
C973 S.n868 SUB 0.29fF $ **FLOATING
C974 S.t61 SUB 21.38fF
C975 S.n869 SUB 21.67fF $ **FLOATING
C976 S.n870 SUB 0.21fF $ **FLOATING
C977 S.n871 SUB 1.41fF $ **FLOATING
C978 S.n872 SUB 4.25fF $ **FLOATING
C979 S.n873 SUB 1.80fF $ **FLOATING
C980 S.t1004 SUB 0.02fF
C981 S.n874 SUB 0.64fF $ **FLOATING
C982 S.n875 SUB 0.61fF $ **FLOATING
C983 S.n876 SUB 1.21fF $ **FLOATING
C984 S.n877 SUB 0.37fF $ **FLOATING
C985 S.n878 SUB 1.18fF $ **FLOATING
C986 S.n879 SUB 0.38fF $ **FLOATING
C987 S.n880 SUB 4.22fF $ **FLOATING
C988 S.t1688 SUB 0.02fF
C989 S.n881 SUB 0.01fF $ **FLOATING
C990 S.n882 SUB 0.26fF $ **FLOATING
C991 S.t886 SUB 0.02fF
C992 S.n884 SUB 1.19fF $ **FLOATING
C993 S.n885 SUB 0.05fF $ **FLOATING
C994 S.t116 SUB 47.92fF
C995 S.t1338 SUB 0.02fF
C996 S.n886 SUB 0.12fF $ **FLOATING
C997 S.n887 SUB 0.14fF $ **FLOATING
C998 S.t1683 SUB 0.02fF
C999 S.n889 SUB 0.24fF $ **FLOATING
C1000 S.n890 SUB 0.91fF $ **FLOATING
C1001 S.n891 SUB 0.05fF $ **FLOATING
C1002 S.t1804 SUB 0.02fF
C1003 S.n892 SUB 0.24fF $ **FLOATING
C1004 S.n893 SUB 0.36fF $ **FLOATING
C1005 S.n894 SUB 0.61fF $ **FLOATING
C1006 S.n895 SUB 0.35fF $ **FLOATING
C1007 S.n896 SUB 0.54fF $ **FLOATING
C1008 S.n897 SUB 0.38fF $ **FLOATING
C1009 S.n898 SUB 0.18fF $ **FLOATING
C1010 S.n899 SUB 0.25fF $ **FLOATING
C1011 S.n900 SUB 0.09fF $ **FLOATING
C1012 S.n901 SUB 1.96fF $ **FLOATING
C1013 S.n902 SUB 1.49fF $ **FLOATING
C1014 S.n903 SUB 2.63fF $ **FLOATING
C1015 S.n904 SUB 8.97fF $ **FLOATING
C1016 S.n905 SUB 8.97fF $ **FLOATING
C1017 S.n906 SUB 5.75fF $ **FLOATING
C1018 S.n907 SUB 0.03fF $ **FLOATING
C1019 S.n908 SUB 0.03fF $ **FLOATING
C1020 S.n909 SUB 0.10fF $ **FLOATING
C1021 S.n910 SUB 0.36fF $ **FLOATING
C1022 S.n911 SUB 0.38fF $ **FLOATING
C1023 S.n912 SUB 0.11fF $ **FLOATING
C1024 S.n913 SUB 0.12fF $ **FLOATING
C1025 S.n914 SUB 0.03fF $ **FLOATING
C1026 S.n915 SUB 0.07fF $ **FLOATING
C1027 S.n916 SUB 1.40fF $ **FLOATING
C1028 S.n917 SUB 1.77fF $ **FLOATING
C1029 S.n918 SUB 1.13fF $ **FLOATING
C1030 S.n919 SUB 0.00fF $ **FLOATING
C1031 S.n920 SUB 0.39fF $ **FLOATING
C1032 S.n921 SUB 0.02fF $ **FLOATING
C1033 S.t1496 SUB 0.02fF
C1034 S.n922 SUB 0.37fF $ **FLOATING
C1035 S.n923 SUB 0.14fF $ **FLOATING
C1036 S.n924 SUB 1.74fF $ **FLOATING
C1037 S.n925 SUB 1.61fF $ **FLOATING
C1038 S.t1396 SUB 0.02fF
C1039 S.n926 SUB 0.89fF $ **FLOATING
C1040 S.t2184 SUB 0.02fF
C1041 S.n927 SUB 0.89fF $ **FLOATING
C1042 S.n928 SUB 1.50fF $ **FLOATING
C1043 S.n929 SUB 2.63fF $ **FLOATING
C1044 S.n930 SUB 0.44fF $ **FLOATING
C1045 S.n931 SUB 0.78fF $ **FLOATING
C1046 S.n932 SUB 0.21fF $ **FLOATING
C1047 S.n933 SUB 1.73fF $ **FLOATING
C1048 S.n934 SUB 8.97fF $ **FLOATING
C1049 S.n935 SUB 8.97fF $ **FLOATING
C1050 S.n936 SUB 5.52fF $ **FLOATING
C1051 S.n937 SUB 1.51fF $ **FLOATING
C1052 S.n938 SUB 0.02fF $ **FLOATING
C1053 S.t633 SUB 0.02fF
C1054 S.n939 SUB 0.37fF $ **FLOATING
C1055 S.n940 SUB 20.80fF $ **FLOATING
C1056 S.n941 SUB 20.80fF $ **FLOATING
C1057 S.n942 SUB 5.78fF $ **FLOATING
C1058 S.n943 SUB 1.96fF $ **FLOATING
C1059 S.t1142 SUB 0.02fF
C1060 S.n944 SUB 0.89fF $ **FLOATING
C1061 S.t1901 SUB 0.02fF
C1062 S.n945 SUB 0.89fF $ **FLOATING
C1063 S.n946 SUB 1.62fF $ **FLOATING
C1064 S.n947 SUB 0.02fF $ **FLOATING
C1065 S.t1277 SUB 0.02fF
C1066 S.n948 SUB 0.37fF $ **FLOATING
C1067 S.t278 SUB 24.03fF
C1068 S.t1595 SUB 0.02fF
C1069 S.n949 SUB 0.89fF $ **FLOATING
C1070 S.n950 SUB 0.02fF $ **FLOATING
C1071 S.t1233 SUB 0.02fF
C1072 S.n951 SUB 0.37fF $ **FLOATING
C1073 S.t965 SUB 0.02fF
C1074 S.n952 SUB 0.89fF $ **FLOATING
C1075 S.t2519 SUB 0.02fF
C1076 S.n953 SUB 0.89fF $ **FLOATING
C1077 S.n954 SUB 0.02fF $ **FLOATING
C1078 S.t2007 SUB 0.02fF
C1079 S.n955 SUB 0.37fF $ **FLOATING
C1080 S.t1730 SUB 0.02fF
C1081 S.n956 SUB 0.89fF $ **FLOATING
C1082 S.t774 SUB 0.02fF
C1083 S.n957 SUB 0.89fF $ **FLOATING
C1084 S.n958 SUB 0.02fF $ **FLOATING
C1085 S.t279 SUB 0.02fF
C1086 S.n959 SUB 0.37fF $ **FLOATING
C1087 S.t2502 SUB 0.02fF
C1088 S.n960 SUB 0.89fF $ **FLOATING
C1089 S.t1560 SUB 0.02fF
C1090 S.n961 SUB 0.89fF $ **FLOATING
C1091 S.n962 SUB 0.02fF $ **FLOATING
C1092 S.t1081 SUB 0.02fF
C1093 S.n963 SUB 0.37fF $ **FLOATING
C1094 S.t914 SUB 0.02fF
C1095 S.n964 SUB 0.89fF $ **FLOATING
C1096 S.t580 SUB 0.02fF
C1097 S.n965 SUB 0.89fF $ **FLOATING
C1098 S.n966 SUB 0.02fF $ **FLOATING
C1099 S.t1639 SUB 0.02fF
C1100 S.n967 SUB 0.37fF $ **FLOATING
C1101 S.t2382 SUB 0.02fF
C1102 S.n968 SUB 0.89fF $ **FLOATING
C1103 S.t1365 SUB 0.02fF
C1104 S.n969 SUB 0.89fF $ **FLOATING
C1105 S.n970 SUB 0.02fF $ **FLOATING
C1106 S.t2423 SUB 0.02fF
C1107 S.n971 SUB 0.37fF $ **FLOATING
C1108 S.t668 SUB 0.02fF
C1109 S.n972 SUB 0.89fF $ **FLOATING
C1110 S.t2268 SUB 0.02fF
C1111 S.n973 SUB 0.89fF $ **FLOATING
C1112 S.n974 SUB 0.02fF $ **FLOATING
C1113 S.t695 SUB 0.02fF
C1114 S.n975 SUB 0.37fF $ **FLOATING
C1115 S.t1460 SUB 0.02fF
C1116 S.n976 SUB 0.89fF $ **FLOATING
C1117 S.t28 SUB 128.28fF
C1118 S.n977 SUB 3.27fF $ **FLOATING
C1119 S.n978 SUB 9.44fF $ **FLOATING
C1120 S.n979 SUB 9.44fF $ **FLOATING
C1121 S.n980 SUB 9.44fF $ **FLOATING
C1122 S.n981 SUB 9.44fF $ **FLOATING
C1123 S.n982 SUB 9.44fF $ **FLOATING
C1124 S.n983 SUB 9.44fF $ **FLOATING
C1125 S.n984 SUB 9.44fF $ **FLOATING
C1126 S.n985 SUB 7.74fF $ **FLOATING
C1127 S.n986 SUB 0.24fF $ **FLOATING
C1128 S.n987 SUB 0.60fF $ **FLOATING
C1129 S.n988 SUB 0.22fF $ **FLOATING
C1130 S.n989 SUB 0.59fF $ **FLOATING
C1131 S.n990 SUB 3.43fF $ **FLOATING
C1132 S.n991 SUB 0.29fF $ **FLOATING
C1133 S.t33 SUB 21.38fF
C1134 S.n992 SUB 21.67fF $ **FLOATING
C1135 S.n993 SUB 0.77fF $ **FLOATING
C1136 S.n994 SUB 0.28fF $ **FLOATING
C1137 S.n995 SUB 4.00fF $ **FLOATING
C1138 S.n996 SUB 1.50fF $ **FLOATING
C1139 S.n997 SUB 1.30fF $ **FLOATING
C1140 S.n998 SUB 0.28fF $ **FLOATING
C1141 S.n999 SUB 0.01fF $ **FLOATING
C1142 S.n1000 SUB 0.01fF $ **FLOATING
C1143 S.n1001 SUB 0.01fF $ **FLOATING
C1144 S.n1002 SUB 0.07fF $ **FLOATING
C1145 S.n1003 SUB 0.07fF $ **FLOATING
C1146 S.n1004 SUB 0.04fF $ **FLOATING
C1147 S.n1005 SUB 0.05fF $ **FLOATING
C1148 S.n1006 SUB 0.41fF $ **FLOATING
C1149 S.n1007 SUB 0.58fF $ **FLOATING
C1150 S.n1008 SUB 0.19fF $ **FLOATING
C1151 S.n1009 SUB 0.18fF $ **FLOATING
C1152 S.n1010 SUB 0.21fF $ **FLOATING
C1153 S.n1011 SUB 0.47fF $ **FLOATING
C1154 S.n1012 SUB 0.33fF $ **FLOATING
C1155 S.n1013 SUB 1.89fF $ **FLOATING
C1156 S.n1014 SUB 0.70fF $ **FLOATING
C1157 S.n1015 SUB 0.23fF $ **FLOATING
C1158 S.n1016 SUB 0.95fF $ **FLOATING
C1159 S.n1017 SUB 0.59fF $ **FLOATING
C1160 S.n1018 SUB 0.25fF $ **FLOATING
C1161 S.n1019 SUB 0.09fF $ **FLOATING
C1162 S.n1020 SUB 0.24fF $ **FLOATING
C1163 S.t169 SUB 0.02fF
C1164 S.n1021 SUB 0.92fF $ **FLOATING
C1165 S.t2590 SUB 0.02fF
C1166 S.n1022 SUB 0.24fF $ **FLOATING
C1167 S.n1023 SUB 0.92fF $ **FLOATING
C1168 S.n1024 SUB 1.88fF $ **FLOATING
C1169 S.n1025 SUB 0.12fF $ **FLOATING
C1170 S.t2227 SUB 0.02fF
C1171 S.n1026 SUB 0.14fF $ **FLOATING
C1172 S.t1518 SUB 0.02fF
C1173 S.n1028 SUB 1.22fF $ **FLOATING
C1174 S.n1029 SUB 0.61fF $ **FLOATING
C1175 S.n1030 SUB 0.35fF $ **FLOATING
C1176 S.n1031 SUB 0.63fF $ **FLOATING
C1177 S.n1032 SUB 1.15fF $ **FLOATING
C1178 S.n1033 SUB 3.03fF $ **FLOATING
C1179 S.n1034 SUB 0.59fF $ **FLOATING
C1180 S.n1035 SUB 0.02fF $ **FLOATING
C1181 S.n1036 SUB 0.97fF $ **FLOATING
C1182 S.t509 SUB 21.38fF
C1183 S.n1037 SUB 20.25fF $ **FLOATING
C1184 S.n1039 SUB 0.38fF $ **FLOATING
C1185 S.n1040 SUB 0.23fF $ **FLOATING
C1186 S.n1041 SUB 2.90fF $ **FLOATING
C1187 S.n1042 SUB 2.46fF $ **FLOATING
C1188 S.n1043 SUB 1.96fF $ **FLOATING
C1189 S.n1044 SUB 3.94fF $ **FLOATING
C1190 S.n1045 SUB 0.25fF $ **FLOATING
C1191 S.n1046 SUB 0.01fF $ **FLOATING
C1192 S.t1249 SUB 0.02fF
C1193 S.n1047 SUB 0.25fF $ **FLOATING
C1194 S.t1002 SUB 0.02fF
C1195 S.n1048 SUB 0.95fF $ **FLOATING
C1196 S.n1049 SUB 0.70fF $ **FLOATING
C1197 S.n1050 SUB 0.78fF $ **FLOATING
C1198 S.n1051 SUB 1.93fF $ **FLOATING
C1199 S.n1052 SUB 1.88fF $ **FLOATING
C1200 S.n1053 SUB 0.12fF $ **FLOATING
C1201 S.t367 SUB 0.02fF
C1202 S.n1054 SUB 0.14fF $ **FLOATING
C1203 S.t657 SUB 0.02fF
C1204 S.n1056 SUB 0.24fF $ **FLOATING
C1205 S.n1057 SUB 0.36fF $ **FLOATING
C1206 S.n1058 SUB 0.61fF $ **FLOATING
C1207 S.n1059 SUB 1.52fF $ **FLOATING
C1208 S.n1060 SUB 2.99fF $ **FLOATING
C1209 S.t97 SUB 0.02fF
C1210 S.n1061 SUB 0.24fF $ **FLOATING
C1211 S.n1062 SUB 0.91fF $ **FLOATING
C1212 S.n1063 SUB 0.05fF $ **FLOATING
C1213 S.t1069 SUB 0.02fF
C1214 S.n1064 SUB 0.12fF $ **FLOATING
C1215 S.n1065 SUB 0.14fF $ **FLOATING
C1216 S.n1067 SUB 1.89fF $ **FLOATING
C1217 S.n1068 SUB 1.88fF $ **FLOATING
C1218 S.t2311 SUB 0.02fF
C1219 S.n1069 SUB 0.24fF $ **FLOATING
C1220 S.n1070 SUB 0.36fF $ **FLOATING
C1221 S.n1071 SUB 0.61fF $ **FLOATING
C1222 S.n1072 SUB 0.12fF $ **FLOATING
C1223 S.t2019 SUB 0.02fF
C1224 S.n1073 SUB 0.14fF $ **FLOATING
C1225 S.n1075 SUB 1.16fF $ **FLOATING
C1226 S.n1076 SUB 0.22fF $ **FLOATING
C1227 S.n1077 SUB 1.88fF $ **FLOATING
C1228 S.t1773 SUB 0.02fF
C1229 S.n1078 SUB 0.24fF $ **FLOATING
C1230 S.n1079 SUB 0.91fF $ **FLOATING
C1231 S.n1080 SUB 0.05fF $ **FLOATING
C1232 S.t190 SUB 0.02fF
C1233 S.n1081 SUB 0.12fF $ **FLOATING
C1234 S.n1082 SUB 0.14fF $ **FLOATING
C1235 S.n1084 SUB 0.78fF $ **FLOATING
C1236 S.n1085 SUB 1.94fF $ **FLOATING
C1237 S.n1086 SUB 1.88fF $ **FLOATING
C1238 S.n1087 SUB 0.12fF $ **FLOATING
C1239 S.t1165 SUB 0.02fF
C1240 S.n1088 SUB 0.14fF $ **FLOATING
C1241 S.t1453 SUB 0.02fF
C1242 S.n1090 SUB 0.24fF $ **FLOATING
C1243 S.n1091 SUB 0.36fF $ **FLOATING
C1244 S.n1092 SUB 0.61fF $ **FLOATING
C1245 S.n1093 SUB 1.84fF $ **FLOATING
C1246 S.n1094 SUB 2.99fF $ **FLOATING
C1247 S.t899 SUB 0.02fF
C1248 S.n1095 SUB 0.24fF $ **FLOATING
C1249 S.n1096 SUB 0.91fF $ **FLOATING
C1250 S.n1097 SUB 0.05fF $ **FLOATING
C1251 S.t1965 SUB 0.02fF
C1252 S.n1098 SUB 0.12fF $ **FLOATING
C1253 S.n1099 SUB 0.14fF $ **FLOATING
C1254 S.n1101 SUB 1.89fF $ **FLOATING
C1255 S.n1102 SUB 1.88fF $ **FLOATING
C1256 S.t595 SUB 0.02fF
C1257 S.n1103 SUB 0.24fF $ **FLOATING
C1258 S.n1104 SUB 0.36fF $ **FLOATING
C1259 S.n1105 SUB 0.61fF $ **FLOATING
C1260 S.n1106 SUB 0.12fF $ **FLOATING
C1261 S.t292 SUB 0.02fF
C1262 S.n1107 SUB 0.14fF $ **FLOATING
C1263 S.n1109 SUB 1.16fF $ **FLOATING
C1264 S.n1110 SUB 0.22fF $ **FLOATING
C1265 S.n1111 SUB 1.88fF $ **FLOATING
C1266 S.t2542 SUB 0.02fF
C1267 S.n1112 SUB 0.24fF $ **FLOATING
C1268 S.n1113 SUB 0.91fF $ **FLOATING
C1269 S.n1114 SUB 0.05fF $ **FLOATING
C1270 S.t1111 SUB 0.02fF
C1271 S.n1115 SUB 0.12fF $ **FLOATING
C1272 S.n1116 SUB 0.14fF $ **FLOATING
C1273 S.n1118 SUB 0.78fF $ **FLOATING
C1274 S.n1119 SUB 1.94fF $ **FLOATING
C1275 S.n1120 SUB 1.88fF $ **FLOATING
C1276 S.n1121 SUB 0.12fF $ **FLOATING
C1277 S.t1955 SUB 0.02fF
C1278 S.n1122 SUB 0.14fF $ **FLOATING
C1279 S.t2244 SUB 0.02fF
C1280 S.n1124 SUB 0.24fF $ **FLOATING
C1281 S.n1125 SUB 0.36fF $ **FLOATING
C1282 S.n1126 SUB 0.61fF $ **FLOATING
C1283 S.n1127 SUB 1.84fF $ **FLOATING
C1284 S.n1128 SUB 2.99fF $ **FLOATING
C1285 S.t1670 SUB 0.02fF
C1286 S.n1129 SUB 0.24fF $ **FLOATING
C1287 S.n1130 SUB 0.91fF $ **FLOATING
C1288 S.n1131 SUB 0.05fF $ **FLOATING
C1289 S.t233 SUB 0.02fF
C1290 S.n1132 SUB 0.12fF $ **FLOATING
C1291 S.n1133 SUB 0.14fF $ **FLOATING
C1292 S.n1135 SUB 1.89fF $ **FLOATING
C1293 S.n1136 SUB 1.88fF $ **FLOATING
C1294 S.t1385 SUB 0.02fF
C1295 S.n1137 SUB 0.24fF $ **FLOATING
C1296 S.n1138 SUB 0.36fF $ **FLOATING
C1297 S.n1139 SUB 0.61fF $ **FLOATING
C1298 S.n1140 SUB 0.12fF $ **FLOATING
C1299 S.t1095 SUB 0.02fF
C1300 S.n1141 SUB 0.14fF $ **FLOATING
C1301 S.n1143 SUB 1.16fF $ **FLOATING
C1302 S.n1144 SUB 0.22fF $ **FLOATING
C1303 S.n1145 SUB 1.88fF $ **FLOATING
C1304 S.t795 SUB 0.02fF
C1305 S.n1146 SUB 0.24fF $ **FLOATING
C1306 S.n1147 SUB 0.91fF $ **FLOATING
C1307 S.n1148 SUB 0.05fF $ **FLOATING
C1308 S.t1899 SUB 0.02fF
C1309 S.n1149 SUB 0.12fF $ **FLOATING
C1310 S.n1150 SUB 0.14fF $ **FLOATING
C1311 S.n1152 SUB 0.78fF $ **FLOATING
C1312 S.n1153 SUB 1.94fF $ **FLOATING
C1313 S.n1154 SUB 1.88fF $ **FLOATING
C1314 S.n1155 SUB 0.12fF $ **FLOATING
C1315 S.t326 SUB 0.02fF
C1316 S.n1156 SUB 0.14fF $ **FLOATING
C1317 S.t510 SUB 0.02fF
C1318 S.n1158 SUB 0.24fF $ **FLOATING
C1319 S.n1159 SUB 0.36fF $ **FLOATING
C1320 S.n1160 SUB 0.61fF $ **FLOATING
C1321 S.n1161 SUB 1.84fF $ **FLOATING
C1322 S.n1162 SUB 2.99fF $ **FLOATING
C1323 S.t2443 SUB 0.02fF
C1324 S.n1163 SUB 0.24fF $ **FLOATING
C1325 S.n1164 SUB 0.91fF $ **FLOATING
C1326 S.n1165 SUB 0.05fF $ **FLOATING
C1327 S.t1039 SUB 0.02fF
C1328 S.n1166 SUB 0.12fF $ **FLOATING
C1329 S.n1167 SUB 0.14fF $ **FLOATING
C1330 S.n1169 SUB 1.89fF $ **FLOATING
C1331 S.n1170 SUB 1.88fF $ **FLOATING
C1332 S.t834 SUB 0.02fF
C1333 S.n1171 SUB 0.24fF $ **FLOATING
C1334 S.n1172 SUB 0.36fF $ **FLOATING
C1335 S.n1173 SUB 0.61fF $ **FLOATING
C1336 S.n1174 SUB 0.12fF $ **FLOATING
C1337 S.t1566 SUB 0.02fF
C1338 S.n1175 SUB 0.14fF $ **FLOATING
C1339 S.n1177 SUB 1.16fF $ **FLOATING
C1340 S.n1178 SUB 0.22fF $ **FLOATING
C1341 S.n1179 SUB 1.88fF $ **FLOATING
C1342 S.t1795 SUB 0.02fF
C1343 S.n1180 SUB 0.24fF $ **FLOATING
C1344 S.n1181 SUB 0.91fF $ **FLOATING
C1345 S.n1182 SUB 0.05fF $ **FLOATING
C1346 S.t143 SUB 0.02fF
C1347 S.n1183 SUB 0.12fF $ **FLOATING
C1348 S.n1184 SUB 0.14fF $ **FLOATING
C1349 S.n1186 SUB 0.78fF $ **FLOATING
C1350 S.n1187 SUB 1.94fF $ **FLOATING
C1351 S.n1188 SUB 1.88fF $ **FLOATING
C1352 S.n1189 SUB 0.12fF $ **FLOATING
C1353 S.t700 SUB 0.02fF
C1354 S.n1190 SUB 0.14fF $ **FLOATING
C1355 S.t2479 SUB 0.02fF
C1356 S.n1192 SUB 0.24fF $ **FLOATING
C1357 S.n1193 SUB 0.36fF $ **FLOATING
C1358 S.n1194 SUB 0.61fF $ **FLOATING
C1359 S.n1195 SUB 1.84fF $ **FLOATING
C1360 S.n1196 SUB 2.99fF $ **FLOATING
C1361 S.t925 SUB 0.02fF
C1362 S.n1197 SUB 0.24fF $ **FLOATING
C1363 S.n1198 SUB 0.91fF $ **FLOATING
C1364 S.n1199 SUB 0.05fF $ **FLOATING
C1365 S.t1420 SUB 0.02fF
C1366 S.n1200 SUB 0.12fF $ **FLOATING
C1367 S.n1201 SUB 0.14fF $ **FLOATING
C1368 S.n1203 SUB 1.89fF $ **FLOATING
C1369 S.n1204 SUB 1.88fF $ **FLOATING
C1370 S.t1608 SUB 0.02fF
C1371 S.n1205 SUB 0.24fF $ **FLOATING
C1372 S.n1206 SUB 0.36fF $ **FLOATING
C1373 S.n1207 SUB 0.61fF $ **FLOATING
C1374 S.n1208 SUB 0.12fF $ **FLOATING
C1375 S.t2359 SUB 0.02fF
C1376 S.n1209 SUB 0.14fF $ **FLOATING
C1377 S.n1211 SUB 1.16fF $ **FLOATING
C1378 S.n1212 SUB 0.22fF $ **FLOATING
C1379 S.n1213 SUB 1.88fF $ **FLOATING
C1380 S.t2565 SUB 0.02fF
C1381 S.n1214 SUB 0.24fF $ **FLOATING
C1382 S.n1215 SUB 0.91fF $ **FLOATING
C1383 S.n1216 SUB 0.05fF $ **FLOATING
C1384 S.t554 SUB 0.02fF
C1385 S.n1217 SUB 0.12fF $ **FLOATING
C1386 S.n1218 SUB 0.14fF $ **FLOATING
C1387 S.n1220 SUB 0.78fF $ **FLOATING
C1388 S.n1221 SUB 1.94fF $ **FLOATING
C1389 S.n1222 SUB 1.88fF $ **FLOATING
C1390 S.n1223 SUB 0.12fF $ **FLOATING
C1391 S.t1502 SUB 0.02fF
C1392 S.n1224 SUB 0.14fF $ **FLOATING
C1393 S.t744 SUB 0.02fF
C1394 S.n1226 SUB 0.24fF $ **FLOATING
C1395 S.n1227 SUB 0.36fF $ **FLOATING
C1396 S.n1228 SUB 0.61fF $ **FLOATING
C1397 S.n1229 SUB 0.06fF $ **FLOATING
C1398 S.n1230 SUB 0.90fF $ **FLOATING
C1399 S.n1231 SUB 1.11fF $ **FLOATING
C1400 S.n1232 SUB 2.98fF $ **FLOATING
C1401 S.t1692 SUB 0.02fF
C1402 S.n1233 SUB 0.24fF $ **FLOATING
C1403 S.n1234 SUB 0.91fF $ **FLOATING
C1404 S.n1235 SUB 0.05fF $ **FLOATING
C1405 S.t2192 SUB 0.02fF
C1406 S.n1236 SUB 0.12fF $ **FLOATING
C1407 S.n1237 SUB 0.14fF $ **FLOATING
C1408 S.n1239 SUB 1.16fF $ **FLOATING
C1409 S.n1240 SUB 0.22fF $ **FLOATING
C1410 S.n1241 SUB 1.89fF $ **FLOATING
C1411 S.n1242 SUB 0.12fF $ **FLOATING
C1412 S.t641 SUB 0.02fF
C1413 S.n1243 SUB 0.14fF $ **FLOATING
C1414 S.t2395 SUB 0.02fF
C1415 S.n1245 SUB 0.24fF $ **FLOATING
C1416 S.n1246 SUB 0.36fF $ **FLOATING
C1417 S.n1247 SUB 0.61fF $ **FLOATING
C1418 S.n1248 SUB 1.10fF $ **FLOATING
C1419 S.n1249 SUB 0.68fF $ **FLOATING
C1420 S.n1250 SUB 0.55fF $ **FLOATING
C1421 S.n1251 SUB 0.32fF $ **FLOATING
C1422 S.n1252 SUB 1.83fF $ **FLOATING
C1423 S.t820 SUB 0.02fF
C1424 S.n1253 SUB 0.24fF $ **FLOATING
C1425 S.n1254 SUB 0.91fF $ **FLOATING
C1426 S.n1255 SUB 0.05fF $ **FLOATING
C1427 S.t1332 SUB 0.02fF
C1428 S.n1256 SUB 0.12fF $ **FLOATING
C1429 S.n1257 SUB 0.14fF $ **FLOATING
C1430 S.n1259 SUB 1.88fF $ **FLOATING
C1431 S.n1260 SUB 0.48fF $ **FLOATING
C1432 S.n1261 SUB 0.09fF $ **FLOATING
C1433 S.n1262 SUB 0.33fF $ **FLOATING
C1434 S.n1263 SUB 0.30fF $ **FLOATING
C1435 S.n1264 SUB 0.77fF $ **FLOATING
C1436 S.n1265 SUB 0.59fF $ **FLOATING
C1437 S.t1535 SUB 0.02fF
C1438 S.n1266 SUB 0.24fF $ **FLOATING
C1439 S.n1267 SUB 0.36fF $ **FLOATING
C1440 S.n1268 SUB 0.61fF $ **FLOATING
C1441 S.n1269 SUB 0.12fF $ **FLOATING
C1442 S.t2299 SUB 0.02fF
C1443 S.n1270 SUB 0.14fF $ **FLOATING
C1444 S.n1272 SUB 2.61fF $ **FLOATING
C1445 S.n1273 SUB 2.16fF $ **FLOATING
C1446 S.t2465 SUB 0.02fF
C1447 S.n1274 SUB 0.24fF $ **FLOATING
C1448 S.n1275 SUB 0.91fF $ **FLOATING
C1449 S.n1276 SUB 0.05fF $ **FLOATING
C1450 S.t592 SUB 0.02fF
C1451 S.n1277 SUB 0.12fF $ **FLOATING
C1452 S.n1278 SUB 0.14fF $ **FLOATING
C1453 S.n1280 SUB 1.88fF $ **FLOATING
C1454 S.n1281 SUB 0.48fF $ **FLOATING
C1455 S.n1282 SUB 0.35fF $ **FLOATING
C1456 S.n1283 SUB 0.30fF $ **FLOATING
C1457 S.n1284 SUB 1.27fF $ **FLOATING
C1458 S.t675 SUB 0.02fF
C1459 S.n1285 SUB 0.24fF $ **FLOATING
C1460 S.n1286 SUB 0.36fF $ **FLOATING
C1461 S.n1287 SUB 0.61fF $ **FLOATING
C1462 S.n1288 SUB 0.12fF $ **FLOATING
C1463 S.t1443 SUB 0.02fF
C1464 S.n1289 SUB 0.14fF $ **FLOATING
C1465 S.n1291 SUB 0.78fF $ **FLOATING
C1466 S.n1292 SUB 2.30fF $ **FLOATING
C1467 S.n1293 SUB 2.03fF $ **FLOATING
C1468 S.t1596 SUB 0.02fF
C1469 S.n1294 SUB 0.24fF $ **FLOATING
C1470 S.n1295 SUB 0.91fF $ **FLOATING
C1471 S.n1296 SUB 0.05fF $ **FLOATING
C1472 S.t2239 SUB 0.02fF
C1473 S.n1297 SUB 0.12fF $ **FLOATING
C1474 S.n1298 SUB 0.14fF $ **FLOATING
C1475 S.n1300 SUB 1.89fF $ **FLOATING
C1476 S.n1301 SUB 2.68fF $ **FLOATING
C1477 S.t2333 SUB 0.02fF
C1478 S.n1302 SUB 0.24fF $ **FLOATING
C1479 S.n1303 SUB 0.36fF $ **FLOATING
C1480 S.n1304 SUB 0.61fF $ **FLOATING
C1481 S.n1305 SUB 0.12fF $ **FLOATING
C1482 S.t581 SUB 0.02fF
C1483 S.n1306 SUB 0.14fF $ **FLOATING
C1484 S.n1308 SUB 1.16fF $ **FLOATING
C1485 S.n1309 SUB 0.22fF $ **FLOATING
C1486 S.n1310 SUB 1.88fF $ **FLOATING
C1487 S.t734 SUB 0.02fF
C1488 S.n1311 SUB 0.24fF $ **FLOATING
C1489 S.n1312 SUB 0.91fF $ **FLOATING
C1490 S.n1313 SUB 0.05fF $ **FLOATING
C1491 S.t1381 SUB 0.02fF
C1492 S.n1314 SUB 0.12fF $ **FLOATING
C1493 S.n1315 SUB 0.14fF $ **FLOATING
C1494 S.n1317 SUB 20.78fF $ **FLOATING
C1495 S.n1318 SUB 2.72fF $ **FLOATING
C1496 S.n1319 SUB 1.81fF $ **FLOATING
C1497 S.n1320 SUB 0.12fF $ **FLOATING
C1498 S.t931 SUB 0.02fF
C1499 S.n1321 SUB 0.14fF $ **FLOATING
C1500 S.t1011 SUB 0.02fF
C1501 S.n1323 SUB 0.24fF $ **FLOATING
C1502 S.n1324 SUB 0.36fF $ **FLOATING
C1503 S.n1325 SUB 0.61fF $ **FLOATING
C1504 S.n1326 SUB 2.36fF $ **FLOATING
C1505 S.n1327 SUB 2.30fF $ **FLOATING
C1506 S.t1647 SUB 0.02fF
C1507 S.n1328 SUB 0.12fF $ **FLOATING
C1508 S.n1329 SUB 0.14fF $ **FLOATING
C1509 S.t1329 SUB 0.02fF
C1510 S.n1331 SUB 0.24fF $ **FLOATING
C1511 S.n1332 SUB 0.91fF $ **FLOATING
C1512 S.n1333 SUB 0.05fF $ **FLOATING
C1513 S.t142 SUB 48.31fF
C1514 S.t506 SUB 0.02fF
C1515 S.n1334 SUB 0.12fF $ **FLOATING
C1516 S.n1335 SUB 0.14fF $ **FLOATING
C1517 S.t2384 SUB 0.02fF
C1518 S.n1337 SUB 0.24fF $ **FLOATING
C1519 S.n1338 SUB 0.91fF $ **FLOATING
C1520 S.n1339 SUB 0.05fF $ **FLOATING
C1521 S.t1476 SUB 0.02fF
C1522 S.n1340 SUB 0.24fF $ **FLOATING
C1523 S.n1341 SUB 0.36fF $ **FLOATING
C1524 S.n1342 SUB 0.61fF $ **FLOATING
C1525 S.n1343 SUB 0.32fF $ **FLOATING
C1526 S.n1344 SUB 1.55fF $ **FLOATING
C1527 S.n1345 SUB 0.15fF $ **FLOATING
C1528 S.n1346 SUB 4.98fF $ **FLOATING
C1529 S.n1347 SUB 1.88fF $ **FLOATING
C1530 S.n1348 SUB 0.12fF $ **FLOATING
C1531 S.t1099 SUB 0.02fF
C1532 S.n1349 SUB 0.14fF $ **FLOATING
C1533 S.t2348 SUB 0.02fF
C1534 S.n1351 SUB 0.24fF $ **FLOATING
C1535 S.n1352 SUB 0.36fF $ **FLOATING
C1536 S.n1353 SUB 0.61fF $ **FLOATING
C1537 S.n1354 SUB 1.27fF $ **FLOATING
C1538 S.n1355 SUB 5.97fF $ **FLOATING
C1539 S.t1148 SUB 0.02fF
C1540 S.n1356 SUB 0.24fF $ **FLOATING
C1541 S.n1357 SUB 0.91fF $ **FLOATING
C1542 S.n1358 SUB 0.05fF $ **FLOATING
C1543 S.t1269 SUB 0.02fF
C1544 S.n1359 SUB 0.12fF $ **FLOATING
C1545 S.n1360 SUB 0.14fF $ **FLOATING
C1546 S.n1362 SUB 1.72fF $ **FLOATING
C1547 S.n1363 SUB 3.06fF $ **FLOATING
C1548 S.t187 SUB 0.02fF
C1549 S.n1364 SUB 0.24fF $ **FLOATING
C1550 S.n1365 SUB 0.36fF $ **FLOATING
C1551 S.n1366 SUB 0.61fF $ **FLOATING
C1552 S.n1367 SUB 0.12fF $ **FLOATING
C1553 S.t2178 SUB 0.02fF
C1554 S.n1368 SUB 0.14fF $ **FLOATING
C1555 S.n1370 SUB 0.28fF $ **FLOATING
C1556 S.n1371 SUB 0.74fF $ **FLOATING
C1557 S.n1372 SUB 0.60fF $ **FLOATING
C1558 S.n1373 SUB 0.21fF $ **FLOATING
C1559 S.n1374 SUB 0.20fF $ **FLOATING
C1560 S.n1375 SUB 0.06fF $ **FLOATING
C1561 S.n1376 SUB 0.09fF $ **FLOATING
C1562 S.n1377 SUB 0.10fF $ **FLOATING
C1563 S.n1378 SUB 1.99fF $ **FLOATING
C1564 S.t1042 SUB 0.02fF
C1565 S.n1379 SUB 0.24fF $ **FLOATING
C1566 S.n1380 SUB 0.91fF $ **FLOATING
C1567 S.n1381 SUB 0.05fF $ **FLOATING
C1568 S.t2351 SUB 0.02fF
C1569 S.n1382 SUB 0.12fF $ **FLOATING
C1570 S.n1383 SUB 0.14fF $ **FLOATING
C1571 S.n1385 SUB 1.88fF $ **FLOATING
C1572 S.n1386 SUB 0.25fF $ **FLOATING
C1573 S.n1387 SUB 0.09fF $ **FLOATING
C1574 S.n1388 SUB 0.21fF $ **FLOATING
C1575 S.n1389 SUB 0.79fF $ **FLOATING
C1576 S.n1390 SUB 0.44fF $ **FLOATING
C1577 S.n1391 SUB 0.12fF $ **FLOATING
C1578 S.t1316 SUB 0.02fF
C1579 S.n1392 SUB 0.14fF $ **FLOATING
C1580 S.t1854 SUB 0.02fF
C1581 S.n1394 SUB 0.24fF $ **FLOATING
C1582 S.n1395 SUB 0.36fF $ **FLOATING
C1583 S.n1396 SUB 0.61fF $ **FLOATING
C1584 S.n1397 SUB 0.02fF $ **FLOATING
C1585 S.n1398 SUB 0.01fF $ **FLOATING
C1586 S.n1399 SUB 0.02fF $ **FLOATING
C1587 S.n1400 SUB 0.08fF $ **FLOATING
C1588 S.n1401 SUB 0.06fF $ **FLOATING
C1589 S.n1402 SUB 0.03fF $ **FLOATING
C1590 S.n1403 SUB 0.04fF $ **FLOATING
C1591 S.n1404 SUB 1.00fF $ **FLOATING
C1592 S.n1405 SUB 0.36fF $ **FLOATING
C1593 S.n1406 SUB 1.85fF $ **FLOATING
C1594 S.n1407 SUB 1.99fF $ **FLOATING
C1595 S.t148 SUB 0.02fF
C1596 S.n1408 SUB 0.24fF $ **FLOATING
C1597 S.n1409 SUB 0.91fF $ **FLOATING
C1598 S.n1410 SUB 0.05fF $ **FLOATING
C1599 S.t1493 SUB 0.02fF
C1600 S.n1411 SUB 0.12fF $ **FLOATING
C1601 S.n1412 SUB 0.14fF $ **FLOATING
C1602 S.n1414 SUB 1.89fF $ **FLOATING
C1603 S.n1415 SUB 0.06fF $ **FLOATING
C1604 S.n1416 SUB 0.03fF $ **FLOATING
C1605 S.n1417 SUB 0.04fF $ **FLOATING
C1606 S.n1418 SUB 0.99fF $ **FLOATING
C1607 S.n1419 SUB 0.02fF $ **FLOATING
C1608 S.n1420 SUB 0.01fF $ **FLOATING
C1609 S.n1421 SUB 0.02fF $ **FLOATING
C1610 S.n1422 SUB 0.08fF $ **FLOATING
C1611 S.n1423 SUB 0.36fF $ **FLOATING
C1612 S.n1424 SUB 1.86fF $ **FLOATING
C1613 S.t1106 SUB 0.02fF
C1614 S.n1425 SUB 0.24fF $ **FLOATING
C1615 S.n1426 SUB 0.36fF $ **FLOATING
C1616 S.n1427 SUB 0.61fF $ **FLOATING
C1617 S.n1428 SUB 0.12fF $ **FLOATING
C1618 S.t582 SUB 0.02fF
C1619 S.n1429 SUB 0.14fF $ **FLOATING
C1620 S.n1431 SUB 0.95fF $ **FLOATING
C1621 S.n1432 SUB 0.59fF $ **FLOATING
C1622 S.n1433 SUB 0.25fF $ **FLOATING
C1623 S.n1434 SUB 0.70fF $ **FLOATING
C1624 S.n1435 SUB 0.23fF $ **FLOATING
C1625 S.n1436 SUB 0.09fF $ **FLOATING
C1626 S.n1437 SUB 1.89fF $ **FLOATING
C1627 S.t1934 SUB 0.02fF
C1628 S.n1438 SUB 0.24fF $ **FLOATING
C1629 S.n1439 SUB 0.91fF $ **FLOATING
C1630 S.n1440 SUB 0.05fF $ **FLOATING
C1631 S.t630 SUB 0.02fF
C1632 S.n1441 SUB 0.12fF $ **FLOATING
C1633 S.n1442 SUB 0.14fF $ **FLOATING
C1634 S.n1444 SUB 1.88fF $ **FLOATING
C1635 S.n1445 SUB 0.25fF $ **FLOATING
C1636 S.n1446 SUB 0.09fF $ **FLOATING
C1637 S.n1447 SUB 0.21fF $ **FLOATING
C1638 S.n1448 SUB 0.79fF $ **FLOATING
C1639 S.n1449 SUB 0.44fF $ **FLOATING
C1640 S.n1450 SUB 0.12fF $ **FLOATING
C1641 S.t2228 SUB 0.02fF
C1642 S.n1451 SUB 0.14fF $ **FLOATING
C1643 S.t1075 SUB 0.02fF
C1644 S.n1453 SUB 0.24fF $ **FLOATING
C1645 S.n1454 SUB 0.91fF $ **FLOATING
C1646 S.n1455 SUB 0.05fF $ **FLOATING
C1647 S.t230 SUB 0.02fF
C1648 S.n1456 SUB 0.24fF $ **FLOATING
C1649 S.n1457 SUB 0.36fF $ **FLOATING
C1650 S.n1458 SUB 0.61fF $ **FLOATING
C1651 S.n1459 SUB 0.02fF $ **FLOATING
C1652 S.n1460 SUB 0.01fF $ **FLOATING
C1653 S.n1461 SUB 0.02fF $ **FLOATING
C1654 S.n1462 SUB 0.08fF $ **FLOATING
C1655 S.n1463 SUB 0.06fF $ **FLOATING
C1656 S.n1464 SUB 0.03fF $ **FLOATING
C1657 S.n1465 SUB 0.04fF $ **FLOATING
C1658 S.n1466 SUB 1.00fF $ **FLOATING
C1659 S.n1467 SUB 0.36fF $ **FLOATING
C1660 S.n1468 SUB 1.85fF $ **FLOATING
C1661 S.n1469 SUB 1.99fF $ **FLOATING
C1662 S.t2286 SUB 0.02fF
C1663 S.n1470 SUB 0.12fF $ **FLOATING
C1664 S.n1471 SUB 0.14fF $ **FLOATING
C1665 S.n1473 SUB 1.89fF $ **FLOATING
C1666 S.n1474 SUB 0.06fF $ **FLOATING
C1667 S.n1475 SUB 0.03fF $ **FLOATING
C1668 S.n1476 SUB 0.04fF $ **FLOATING
C1669 S.n1477 SUB 0.99fF $ **FLOATING
C1670 S.n1478 SUB 0.02fF $ **FLOATING
C1671 S.n1479 SUB 0.01fF $ **FLOATING
C1672 S.n1480 SUB 0.02fF $ **FLOATING
C1673 S.n1481 SUB 0.08fF $ **FLOATING
C1674 S.n1482 SUB 0.36fF $ **FLOATING
C1675 S.n1483 SUB 1.86fF $ **FLOATING
C1676 S.t1895 SUB 0.02fF
C1677 S.n1484 SUB 0.24fF $ **FLOATING
C1678 S.n1485 SUB 0.36fF $ **FLOATING
C1679 S.n1486 SUB 0.61fF $ **FLOATING
C1680 S.n1487 SUB 0.12fF $ **FLOATING
C1681 S.t1366 SUB 0.02fF
C1682 S.n1488 SUB 0.14fF $ **FLOATING
C1683 S.n1490 SUB 0.70fF $ **FLOATING
C1684 S.n1491 SUB 0.23fF $ **FLOATING
C1685 S.n1492 SUB 0.95fF $ **FLOATING
C1686 S.n1493 SUB 0.59fF $ **FLOATING
C1687 S.n1494 SUB 0.25fF $ **FLOATING
C1688 S.n1495 SUB 0.09fF $ **FLOATING
C1689 S.n1496 SUB 1.89fF $ **FLOATING
C1690 S.t198 SUB 0.02fF
C1691 S.n1497 SUB 0.24fF $ **FLOATING
C1692 S.n1498 SUB 0.91fF $ **FLOATING
C1693 S.n1499 SUB 0.05fF $ **FLOATING
C1694 S.t1433 SUB 0.02fF
C1695 S.n1500 SUB 0.12fF $ **FLOATING
C1696 S.n1501 SUB 0.14fF $ **FLOATING
C1697 S.n1503 SUB 1.88fF $ **FLOATING
C1698 S.n1504 SUB 0.25fF $ **FLOATING
C1699 S.n1505 SUB 0.09fF $ **FLOATING
C1700 S.n1506 SUB 0.21fF $ **FLOATING
C1701 S.n1507 SUB 0.79fF $ **FLOATING
C1702 S.n1508 SUB 0.44fF $ **FLOATING
C1703 S.n1509 SUB 0.12fF $ **FLOATING
C1704 S.t492 SUB 0.02fF
C1705 S.n1510 SUB 0.14fF $ **FLOATING
C1706 S.t1035 SUB 0.02fF
C1707 S.n1512 SUB 0.24fF $ **FLOATING
C1708 S.n1513 SUB 0.36fF $ **FLOATING
C1709 S.n1514 SUB 0.61fF $ **FLOATING
C1710 S.n1515 SUB 0.02fF $ **FLOATING
C1711 S.n1516 SUB 0.01fF $ **FLOATING
C1712 S.n1517 SUB 0.02fF $ **FLOATING
C1713 S.n1518 SUB 0.08fF $ **FLOATING
C1714 S.n1519 SUB 0.06fF $ **FLOATING
C1715 S.n1520 SUB 0.03fF $ **FLOATING
C1716 S.n1521 SUB 0.04fF $ **FLOATING
C1717 S.n1522 SUB 1.00fF $ **FLOATING
C1718 S.n1523 SUB 0.36fF $ **FLOATING
C1719 S.n1524 SUB 1.85fF $ **FLOATING
C1720 S.n1525 SUB 1.99fF $ **FLOATING
C1721 S.t1865 SUB 0.02fF
C1722 S.n1526 SUB 0.24fF $ **FLOATING
C1723 S.n1527 SUB 0.91fF $ **FLOATING
C1724 S.n1528 SUB 0.05fF $ **FLOATING
C1725 S.t569 SUB 0.02fF
C1726 S.n1529 SUB 0.12fF $ **FLOATING
C1727 S.n1530 SUB 0.14fF $ **FLOATING
C1728 S.n1532 SUB 1.89fF $ **FLOATING
C1729 S.n1533 SUB 0.06fF $ **FLOATING
C1730 S.n1534 SUB 0.03fF $ **FLOATING
C1731 S.n1535 SUB 0.04fF $ **FLOATING
C1732 S.n1536 SUB 0.99fF $ **FLOATING
C1733 S.n1537 SUB 0.02fF $ **FLOATING
C1734 S.n1538 SUB 0.01fF $ **FLOATING
C1735 S.n1539 SUB 0.02fF $ **FLOATING
C1736 S.n1540 SUB 0.08fF $ **FLOATING
C1737 S.n1541 SUB 0.36fF $ **FLOATING
C1738 S.n1542 SUB 1.86fF $ **FLOATING
C1739 S.t138 SUB 0.02fF
C1740 S.n1543 SUB 0.24fF $ **FLOATING
C1741 S.n1544 SUB 0.36fF $ **FLOATING
C1742 S.n1545 SUB 0.61fF $ **FLOATING
C1743 S.n1546 SUB 0.12fF $ **FLOATING
C1744 S.t2137 SUB 0.02fF
C1745 S.n1547 SUB 0.14fF $ **FLOATING
C1746 S.n1549 SUB 0.70fF $ **FLOATING
C1747 S.n1550 SUB 0.23fF $ **FLOATING
C1748 S.n1551 SUB 0.95fF $ **FLOATING
C1749 S.n1552 SUB 0.59fF $ **FLOATING
C1750 S.n1553 SUB 0.25fF $ **FLOATING
C1751 S.n1554 SUB 0.09fF $ **FLOATING
C1752 S.n1555 SUB 1.89fF $ **FLOATING
C1753 S.t996 SUB 0.02fF
C1754 S.n1556 SUB 0.24fF $ **FLOATING
C1755 S.n1557 SUB 0.91fF $ **FLOATING
C1756 S.n1558 SUB 0.05fF $ **FLOATING
C1757 S.t2213 SUB 0.02fF
C1758 S.n1559 SUB 0.12fF $ **FLOATING
C1759 S.n1560 SUB 0.14fF $ **FLOATING
C1760 S.n1562 SUB 1.88fF $ **FLOATING
C1761 S.n1563 SUB 0.25fF $ **FLOATING
C1762 S.n1564 SUB 0.09fF $ **FLOATING
C1763 S.n1565 SUB 0.21fF $ **FLOATING
C1764 S.n1566 SUB 0.79fF $ **FLOATING
C1765 S.n1567 SUB 0.44fF $ **FLOATING
C1766 S.n1568 SUB 0.12fF $ **FLOATING
C1767 S.t1272 SUB 0.02fF
C1768 S.n1569 SUB 0.14fF $ **FLOATING
C1769 S.t1807 SUB 0.02fF
C1770 S.n1571 SUB 0.24fF $ **FLOATING
C1771 S.n1572 SUB 0.36fF $ **FLOATING
C1772 S.n1573 SUB 0.61fF $ **FLOATING
C1773 S.n1574 SUB 0.02fF $ **FLOATING
C1774 S.n1575 SUB 0.01fF $ **FLOATING
C1775 S.n1576 SUB 0.02fF $ **FLOATING
C1776 S.n1577 SUB 0.08fF $ **FLOATING
C1777 S.n1578 SUB 0.06fF $ **FLOATING
C1778 S.n1579 SUB 0.03fF $ **FLOATING
C1779 S.n1580 SUB 0.04fF $ **FLOATING
C1780 S.n1581 SUB 1.00fF $ **FLOATING
C1781 S.n1582 SUB 0.36fF $ **FLOATING
C1782 S.n1583 SUB 1.85fF $ **FLOATING
C1783 S.n1584 SUB 1.99fF $ **FLOATING
C1784 S.t89 SUB 0.02fF
C1785 S.n1585 SUB 0.24fF $ **FLOATING
C1786 S.n1586 SUB 0.91fF $ **FLOATING
C1787 S.n1587 SUB 0.05fF $ **FLOATING
C1788 S.t1464 SUB 0.02fF
C1789 S.n1588 SUB 0.12fF $ **FLOATING
C1790 S.n1589 SUB 0.14fF $ **FLOATING
C1791 S.n1591 SUB 1.89fF $ **FLOATING
C1792 S.n1592 SUB 0.06fF $ **FLOATING
C1793 S.n1593 SUB 0.03fF $ **FLOATING
C1794 S.n1594 SUB 0.04fF $ **FLOATING
C1795 S.n1595 SUB 0.99fF $ **FLOATING
C1796 S.n1596 SUB 0.02fF $ **FLOATING
C1797 S.n1597 SUB 0.01fF $ **FLOATING
C1798 S.n1598 SUB 0.02fF $ **FLOATING
C1799 S.n1599 SUB 0.08fF $ **FLOATING
C1800 S.n1600 SUB 0.36fF $ **FLOATING
C1801 S.n1601 SUB 1.86fF $ **FLOATING
C1802 S.t1007 SUB 0.02fF
C1803 S.n1602 SUB 0.24fF $ **FLOATING
C1804 S.n1603 SUB 0.36fF $ **FLOATING
C1805 S.n1604 SUB 0.61fF $ **FLOATING
C1806 S.n1605 SUB 0.12fF $ **FLOATING
C1807 S.t451 SUB 0.02fF
C1808 S.n1606 SUB 0.14fF $ **FLOATING
C1809 S.n1608 SUB 0.70fF $ **FLOATING
C1810 S.n1609 SUB 0.23fF $ **FLOATING
C1811 S.n1610 SUB 0.95fF $ **FLOATING
C1812 S.n1611 SUB 0.59fF $ **FLOATING
C1813 S.n1612 SUB 0.25fF $ **FLOATING
C1814 S.n1613 SUB 0.09fF $ **FLOATING
C1815 S.n1614 SUB 1.89fF $ **FLOATING
C1816 S.t888 SUB 0.02fF
C1817 S.n1615 SUB 0.24fF $ **FLOATING
C1818 S.n1616 SUB 0.91fF $ **FLOATING
C1819 S.n1617 SUB 0.05fF $ **FLOATING
C1820 S.t639 SUB 0.02fF
C1821 S.n1618 SUB 0.12fF $ **FLOATING
C1822 S.n1619 SUB 0.14fF $ **FLOATING
C1823 S.n1621 SUB 1.88fF $ **FLOATING
C1824 S.n1622 SUB 0.25fF $ **FLOATING
C1825 S.n1623 SUB 0.09fF $ **FLOATING
C1826 S.n1624 SUB 0.21fF $ **FLOATING
C1827 S.n1625 SUB 0.79fF $ **FLOATING
C1828 S.n1626 SUB 0.44fF $ **FLOATING
C1829 S.n1627 SUB 0.12fF $ **FLOATING
C1830 S.t2096 SUB 0.02fF
C1831 S.n1628 SUB 0.14fF $ **FLOATING
C1832 S.t107 SUB 0.02fF
C1833 S.n1630 SUB 0.24fF $ **FLOATING
C1834 S.n1631 SUB 0.36fF $ **FLOATING
C1835 S.n1632 SUB 0.61fF $ **FLOATING
C1836 S.n1633 SUB 0.02fF $ **FLOATING
C1837 S.n1634 SUB 0.01fF $ **FLOATING
C1838 S.n1635 SUB 0.02fF $ **FLOATING
C1839 S.n1636 SUB 0.08fF $ **FLOATING
C1840 S.n1637 SUB 0.06fF $ **FLOATING
C1841 S.n1638 SUB 0.03fF $ **FLOATING
C1842 S.n1639 SUB 0.04fF $ **FLOATING
C1843 S.n1640 SUB 1.00fF $ **FLOATING
C1844 S.n1641 SUB 0.36fF $ **FLOATING
C1845 S.n1642 SUB 1.85fF $ **FLOATING
C1846 S.n1643 SUB 1.99fF $ **FLOATING
C1847 S.t2530 SUB 0.02fF
C1848 S.n1644 SUB 0.24fF $ **FLOATING
C1849 S.n1645 SUB 0.91fF $ **FLOATING
C1850 S.n1646 SUB 0.05fF $ **FLOATING
C1851 S.t2298 SUB 0.02fF
C1852 S.n1647 SUB 0.12fF $ **FLOATING
C1853 S.n1648 SUB 0.14fF $ **FLOATING
C1854 S.n1650 SUB 1.89fF $ **FLOATING
C1855 S.n1651 SUB 0.06fF $ **FLOATING
C1856 S.n1652 SUB 0.03fF $ **FLOATING
C1857 S.n1653 SUB 0.04fF $ **FLOATING
C1858 S.n1654 SUB 0.99fF $ **FLOATING
C1859 S.n1655 SUB 0.02fF $ **FLOATING
C1860 S.n1656 SUB 0.01fF $ **FLOATING
C1861 S.n1657 SUB 0.02fF $ **FLOATING
C1862 S.n1658 SUB 0.08fF $ **FLOATING
C1863 S.n1659 SUB 0.36fF $ **FLOATING
C1864 S.n1660 SUB 1.86fF $ **FLOATING
C1865 S.t1780 SUB 0.02fF
C1866 S.n1661 SUB 0.24fF $ **FLOATING
C1867 S.n1662 SUB 0.36fF $ **FLOATING
C1868 S.n1663 SUB 0.61fF $ **FLOATING
C1869 S.n1664 SUB 0.12fF $ **FLOATING
C1870 S.t1231 SUB 0.02fF
C1871 S.n1665 SUB 0.14fF $ **FLOATING
C1872 S.n1667 SUB 0.70fF $ **FLOATING
C1873 S.n1668 SUB 0.23fF $ **FLOATING
C1874 S.n1669 SUB 0.95fF $ **FLOATING
C1875 S.n1670 SUB 0.59fF $ **FLOATING
C1876 S.n1671 SUB 0.25fF $ **FLOATING
C1877 S.n1672 SUB 0.09fF $ **FLOATING
C1878 S.n1673 SUB 1.89fF $ **FLOATING
C1879 S.t1657 SUB 0.02fF
C1880 S.n1674 SUB 0.24fF $ **FLOATING
C1881 S.n1675 SUB 0.91fF $ **FLOATING
C1882 S.n1676 SUB 0.05fF $ **FLOATING
C1883 S.t1442 SUB 0.02fF
C1884 S.n1677 SUB 0.12fF $ **FLOATING
C1885 S.n1678 SUB 0.14fF $ **FLOATING
C1886 S.n1680 SUB 1.88fF $ **FLOATING
C1887 S.n1681 SUB 0.25fF $ **FLOATING
C1888 S.n1682 SUB 0.09fF $ **FLOATING
C1889 S.n1683 SUB 0.21fF $ **FLOATING
C1890 S.n1684 SUB 0.79fF $ **FLOATING
C1891 S.n1685 SUB 0.44fF $ **FLOATING
C1892 S.n1686 SUB 0.12fF $ **FLOATING
C1893 S.t348 SUB 0.02fF
C1894 S.n1687 SUB 0.14fF $ **FLOATING
C1895 S.t908 SUB 0.02fF
C1896 S.n1689 SUB 0.24fF $ **FLOATING
C1897 S.n1690 SUB 0.36fF $ **FLOATING
C1898 S.n1691 SUB 0.61fF $ **FLOATING
C1899 S.n1692 SUB 0.02fF $ **FLOATING
C1900 S.n1693 SUB 0.01fF $ **FLOATING
C1901 S.n1694 SUB 0.02fF $ **FLOATING
C1902 S.n1695 SUB 0.08fF $ **FLOATING
C1903 S.n1696 SUB 0.03fF $ **FLOATING
C1904 S.n1697 SUB 0.04fF $ **FLOATING
C1905 S.n1698 SUB 1.02fF $ **FLOATING
C1906 S.n1699 SUB 0.36fF $ **FLOATING
C1907 S.n1700 SUB 1.85fF $ **FLOATING
C1908 S.n1701 SUB 1.99fF $ **FLOATING
C1909 S.t788 SUB 0.02fF
C1910 S.n1702 SUB 0.24fF $ **FLOATING
C1911 S.n1703 SUB 0.91fF $ **FLOATING
C1912 S.n1704 SUB 0.05fF $ **FLOATING
C1913 S.t579 SUB 0.02fF
C1914 S.n1705 SUB 0.12fF $ **FLOATING
C1915 S.n1706 SUB 0.14fF $ **FLOATING
C1916 S.n1708 SUB 0.04fF $ **FLOATING
C1917 S.n1709 SUB 0.03fF $ **FLOATING
C1918 S.n1710 SUB 0.03fF $ **FLOATING
C1919 S.n1711 SUB 0.10fF $ **FLOATING
C1920 S.n1712 SUB 0.36fF $ **FLOATING
C1921 S.n1713 SUB 0.38fF $ **FLOATING
C1922 S.n1714 SUB 0.11fF $ **FLOATING
C1923 S.n1715 SUB 0.12fF $ **FLOATING
C1924 S.n1716 SUB 0.07fF $ **FLOATING
C1925 S.n1717 SUB 0.12fF $ **FLOATING
C1926 S.n1718 SUB 0.18fF $ **FLOATING
C1927 S.n1719 SUB 1.88fF $ **FLOATING
C1928 S.n1720 SUB 0.12fF $ **FLOATING
C1929 S.t1291 SUB 0.02fF
C1930 S.n1721 SUB 0.14fF $ **FLOATING
C1931 S.t1832 SUB 0.02fF
C1932 S.n1723 SUB 0.24fF $ **FLOATING
C1933 S.n1724 SUB 0.36fF $ **FLOATING
C1934 S.n1725 SUB 0.61fF $ **FLOATING
C1935 S.n1726 SUB 0.42fF $ **FLOATING
C1936 S.n1727 SUB 0.21fF $ **FLOATING
C1937 S.n1728 SUB 0.16fF $ **FLOATING
C1938 S.n1729 SUB 0.28fF $ **FLOATING
C1939 S.n1730 SUB 0.21fF $ **FLOATING
C1940 S.n1731 SUB 0.79fF $ **FLOATING
C1941 S.n1732 SUB 0.31fF $ **FLOATING
C1942 S.n1733 SUB 0.22fF $ **FLOATING
C1943 S.n1734 SUB 0.38fF $ **FLOATING
C1944 S.n1735 SUB 3.61fF $ **FLOATING
C1945 S.t1714 SUB 0.02fF
C1946 S.n1736 SUB 0.24fF $ **FLOATING
C1947 S.n1737 SUB 0.91fF $ **FLOATING
C1948 S.n1738 SUB 0.05fF $ **FLOATING
C1949 S.t1361 SUB 0.02fF
C1950 S.n1739 SUB 0.12fF $ **FLOATING
C1951 S.n1740 SUB 0.14fF $ **FLOATING
C1952 S.n1742 SUB 0.25fF $ **FLOATING
C1953 S.n1743 SUB 0.09fF $ **FLOATING
C1954 S.n1744 SUB 0.21fF $ **FLOATING
C1955 S.n1745 SUB 1.28fF $ **FLOATING
C1956 S.n1746 SUB 0.53fF $ **FLOATING
C1957 S.n1747 SUB 1.88fF $ **FLOATING
C1958 S.n1748 SUB 0.12fF $ **FLOATING
C1959 S.t404 SUB 0.02fF
C1960 S.n1749 SUB 0.14fF $ **FLOATING
C1961 S.t966 SUB 0.02fF
C1962 S.n1751 SUB 0.24fF $ **FLOATING
C1963 S.n1752 SUB 0.36fF $ **FLOATING
C1964 S.n1753 SUB 0.61fF $ **FLOATING
C1965 S.n1754 SUB 0.42fF $ **FLOATING
C1966 S.n1755 SUB 0.21fF $ **FLOATING
C1967 S.n1756 SUB 0.16fF $ **FLOATING
C1968 S.n1757 SUB 0.28fF $ **FLOATING
C1969 S.n1758 SUB 0.21fF $ **FLOATING
C1970 S.n1759 SUB 0.30fF $ **FLOATING
C1971 S.n1760 SUB 0.36fF $ **FLOATING
C1972 S.n1761 SUB 0.22fF $ **FLOATING
C1973 S.n1762 SUB 0.38fF $ **FLOATING
C1974 S.n1763 SUB 2.42fF $ **FLOATING
C1975 S.t843 SUB 0.02fF
C1976 S.n1764 SUB 0.24fF $ **FLOATING
C1977 S.n1765 SUB 0.91fF $ **FLOATING
C1978 S.n1766 SUB 0.05fF $ **FLOATING
C1979 S.t488 SUB 0.02fF
C1980 S.n1767 SUB 0.12fF $ **FLOATING
C1981 S.n1768 SUB 0.14fF $ **FLOATING
C1982 S.n1770 SUB 1.89fF $ **FLOATING
C1983 S.n1771 SUB 2.67fF $ **FLOATING
C1984 S.t34 SUB 0.02fF
C1985 S.n1772 SUB 0.24fF $ **FLOATING
C1986 S.n1773 SUB 0.36fF $ **FLOATING
C1987 S.n1774 SUB 0.61fF $ **FLOATING
C1988 S.n1775 SUB 0.12fF $ **FLOATING
C1989 S.t2052 SUB 0.02fF
C1990 S.n1776 SUB 0.14fF $ **FLOATING
C1991 S.n1778 SUB 0.70fF $ **FLOATING
C1992 S.n1779 SUB 0.23fF $ **FLOATING
C1993 S.n1780 SUB 0.70fF $ **FLOATING
C1994 S.n1781 SUB 1.16fF $ **FLOATING
C1995 S.n1782 SUB 0.22fF $ **FLOATING
C1996 S.n1783 SUB 0.25fF $ **FLOATING
C1997 S.n1784 SUB 0.09fF $ **FLOATING
C1998 S.n1785 SUB 1.89fF $ **FLOATING
C1999 S.t2487 SUB 0.02fF
C2000 S.n1786 SUB 0.24fF $ **FLOATING
C2001 S.n1787 SUB 0.91fF $ **FLOATING
C2002 S.n1788 SUB 0.05fF $ **FLOATING
C2003 S.t2135 SUB 0.02fF
C2004 S.n1789 SUB 0.12fF $ **FLOATING
C2005 S.n1790 SUB 0.14fF $ **FLOATING
C2006 S.n1792 SUB 20.78fF $ **FLOATING
C2007 S.n1793 SUB 0.12fF $ **FLOATING
C2008 S.t2223 SUB 0.02fF
C2009 S.n1794 SUB 0.14fF $ **FLOATING
C2010 S.t2151 SUB 0.02fF
C2011 S.n1795 SUB 0.12fF $ **FLOATING
C2012 S.n1796 SUB 0.14fF $ **FLOATING
C2013 S.t320 SUB 49.98fF
C2014 S.t321 SUB 0.02fF
C2015 S.n1797 SUB 0.01fF $ **FLOATING
C2016 S.n1798 SUB 0.26fF $ **FLOATING
C2017 S.t2562 SUB 0.02fF
C2018 S.n1800 SUB 1.19fF $ **FLOATING
C2019 S.n1801 SUB 0.05fF $ **FLOATING
C2020 S.t139 SUB 0.02fF
C2021 S.n1802 SUB 0.64fF $ **FLOATING
C2022 S.n1803 SUB 0.61fF $ **FLOATING
C2023 S.n1804 SUB 1.50fF $ **FLOATING
C2024 S.n1805 SUB 0.35fF $ **FLOATING
C2025 S.n1806 SUB 1.30fF $ **FLOATING
C2026 S.n1807 SUB 0.16fF $ **FLOATING
C2027 S.n1808 SUB 1.75fF $ **FLOATING
C2028 S.n1809 SUB 2.29fF $ **FLOATING
C2029 S.n1810 SUB 0.01fF $ **FLOATING
C2030 S.n1811 SUB 0.02fF $ **FLOATING
C2031 S.n1812 SUB 0.03fF $ **FLOATING
C2032 S.n1813 SUB 0.04fF $ **FLOATING
C2033 S.n1814 SUB 0.17fF $ **FLOATING
C2034 S.n1815 SUB 0.01fF $ **FLOATING
C2035 S.n1816 SUB 0.02fF $ **FLOATING
C2036 S.n1817 SUB 0.01fF $ **FLOATING
C2037 S.n1818 SUB 0.01fF $ **FLOATING
C2038 S.n1819 SUB 0.01fF $ **FLOATING
C2039 S.n1820 SUB 0.01fF $ **FLOATING
C2040 S.n1821 SUB 0.02fF $ **FLOATING
C2041 S.n1822 SUB 0.01fF $ **FLOATING
C2042 S.n1823 SUB 0.02fF $ **FLOATING
C2043 S.n1824 SUB 0.05fF $ **FLOATING
C2044 S.n1825 SUB 0.04fF $ **FLOATING
C2045 S.n1826 SUB 0.11fF $ **FLOATING
C2046 S.n1827 SUB 0.38fF $ **FLOATING
C2047 S.n1828 SUB 0.20fF $ **FLOATING
C2048 S.n1829 SUB 8.97fF $ **FLOATING
C2049 S.n1830 SUB 8.97fF $ **FLOATING
C2050 S.n1831 SUB 0.60fF $ **FLOATING
C2051 S.n1832 SUB 0.22fF $ **FLOATING
C2052 S.n1833 SUB 0.59fF $ **FLOATING
C2053 S.n1834 SUB 3.43fF $ **FLOATING
C2054 S.n1835 SUB 0.29fF $ **FLOATING
C2055 S.t63 SUB 21.38fF
C2056 S.n1836 SUB 21.67fF $ **FLOATING
C2057 S.n1837 SUB 0.77fF $ **FLOATING
C2058 S.n1838 SUB 0.28fF $ **FLOATING
C2059 S.n1839 SUB 4.00fF $ **FLOATING
C2060 S.n1840 SUB 1.35fF $ **FLOATING
C2061 S.t158 SUB 0.02fF
C2062 S.n1841 SUB 0.64fF $ **FLOATING
C2063 S.n1842 SUB 0.61fF $ **FLOATING
C2064 S.n1843 SUB 1.89fF $ **FLOATING
C2065 S.n1844 SUB 0.06fF $ **FLOATING
C2066 S.n1845 SUB 0.03fF $ **FLOATING
C2067 S.n1846 SUB 0.04fF $ **FLOATING
C2068 S.n1847 SUB 0.99fF $ **FLOATING
C2069 S.n1848 SUB 0.02fF $ **FLOATING
C2070 S.n1849 SUB 0.01fF $ **FLOATING
C2071 S.n1850 SUB 0.02fF $ **FLOATING
C2072 S.n1851 SUB 0.08fF $ **FLOATING
C2073 S.n1852 SUB 0.36fF $ **FLOATING
C2074 S.n1853 SUB 1.85fF $ **FLOATING
C2075 S.t1271 SUB 0.02fF
C2076 S.n1854 SUB 0.24fF $ **FLOATING
C2077 S.n1855 SUB 0.36fF $ **FLOATING
C2078 S.n1856 SUB 0.61fF $ **FLOATING
C2079 S.n1857 SUB 0.12fF $ **FLOATING
C2080 S.t1043 SUB 0.02fF
C2081 S.n1858 SUB 0.14fF $ **FLOATING
C2082 S.n1860 SUB 0.70fF $ **FLOATING
C2083 S.n1861 SUB 0.23fF $ **FLOATING
C2084 S.n1862 SUB 0.25fF $ **FLOATING
C2085 S.n1863 SUB 0.09fF $ **FLOATING
C2086 S.n1864 SUB 0.23fF $ **FLOATING
C2087 S.n1865 SUB 0.70fF $ **FLOATING
C2088 S.n1866 SUB 1.16fF $ **FLOATING
C2089 S.n1867 SUB 0.22fF $ **FLOATING
C2090 S.n1868 SUB 0.25fF $ **FLOATING
C2091 S.n1869 SUB 0.09fF $ **FLOATING
C2092 S.n1870 SUB 1.88fF $ **FLOATING
C2093 S.t2363 SUB 0.02fF
C2094 S.n1871 SUB 0.24fF $ **FLOATING
C2095 S.n1872 SUB 0.91fF $ **FLOATING
C2096 S.n1873 SUB 0.05fF $ **FLOATING
C2097 S.t1211 SUB 0.02fF
C2098 S.n1874 SUB 0.12fF $ **FLOATING
C2099 S.n1875 SUB 0.14fF $ **FLOATING
C2100 S.n1877 SUB 0.25fF $ **FLOATING
C2101 S.n1878 SUB 0.09fF $ **FLOATING
C2102 S.n1879 SUB 0.21fF $ **FLOATING
C2103 S.n1880 SUB 0.92fF $ **FLOATING
C2104 S.n1881 SUB 0.44fF $ **FLOATING
C2105 S.n1882 SUB 1.88fF $ **FLOATING
C2106 S.n1883 SUB 0.12fF $ **FLOATING
C2107 S.t272 SUB 0.02fF
C2108 S.n1884 SUB 0.14fF $ **FLOATING
C2109 S.t544 SUB 0.02fF
C2110 S.n1886 SUB 0.24fF $ **FLOATING
C2111 S.n1887 SUB 0.36fF $ **FLOATING
C2112 S.n1888 SUB 0.61fF $ **FLOATING
C2113 S.n1889 SUB 0.02fF $ **FLOATING
C2114 S.n1890 SUB 0.01fF $ **FLOATING
C2115 S.n1891 SUB 0.02fF $ **FLOATING
C2116 S.n1892 SUB 0.08fF $ **FLOATING
C2117 S.n1893 SUB 0.06fF $ **FLOATING
C2118 S.n1894 SUB 0.03fF $ **FLOATING
C2119 S.n1895 SUB 0.04fF $ **FLOATING
C2120 S.n1896 SUB 1.00fF $ **FLOATING
C2121 S.n1897 SUB 0.36fF $ **FLOATING
C2122 S.n1898 SUB 1.87fF $ **FLOATING
C2123 S.n1899 SUB 1.99fF $ **FLOATING
C2124 S.t1613 SUB 0.02fF
C2125 S.n1900 SUB 0.24fF $ **FLOATING
C2126 S.n1901 SUB 0.91fF $ **FLOATING
C2127 S.n1902 SUB 0.05fF $ **FLOATING
C2128 S.t332 SUB 0.02fF
C2129 S.n1903 SUB 0.12fF $ **FLOATING
C2130 S.n1904 SUB 0.14fF $ **FLOATING
C2131 S.n1906 SUB 1.89fF $ **FLOATING
C2132 S.n1907 SUB 0.06fF $ **FLOATING
C2133 S.n1908 SUB 0.03fF $ **FLOATING
C2134 S.n1909 SUB 0.04fF $ **FLOATING
C2135 S.n1910 SUB 0.99fF $ **FLOATING
C2136 S.n1911 SUB 0.02fF $ **FLOATING
C2137 S.n1912 SUB 0.01fF $ **FLOATING
C2138 S.n1913 SUB 0.02fF $ **FLOATING
C2139 S.n1914 SUB 0.08fF $ **FLOATING
C2140 S.n1915 SUB 0.36fF $ **FLOATING
C2141 S.n1916 SUB 1.85fF $ **FLOATING
C2142 S.t2185 SUB 0.02fF
C2143 S.n1917 SUB 0.24fF $ **FLOATING
C2144 S.n1918 SUB 0.36fF $ **FLOATING
C2145 S.n1919 SUB 0.61fF $ **FLOATING
C2146 S.n1920 SUB 0.12fF $ **FLOATING
C2147 S.t1935 SUB 0.02fF
C2148 S.n1921 SUB 0.14fF $ **FLOATING
C2149 S.n1923 SUB 0.70fF $ **FLOATING
C2150 S.n1924 SUB 0.23fF $ **FLOATING
C2151 S.n1925 SUB 0.25fF $ **FLOATING
C2152 S.n1926 SUB 0.09fF $ **FLOATING
C2153 S.n1927 SUB 0.23fF $ **FLOATING
C2154 S.n1928 SUB 0.70fF $ **FLOATING
C2155 S.n1929 SUB 1.16fF $ **FLOATING
C2156 S.n1930 SUB 0.22fF $ **FLOATING
C2157 S.n1931 SUB 0.25fF $ **FLOATING
C2158 S.n1932 SUB 0.09fF $ **FLOATING
C2159 S.n1933 SUB 1.88fF $ **FLOATING
C2160 S.t750 SUB 0.02fF
C2161 S.n1934 SUB 0.24fF $ **FLOATING
C2162 S.n1935 SUB 0.91fF $ **FLOATING
C2163 S.n1936 SUB 0.05fF $ **FLOATING
C2164 S.t1989 SUB 0.02fF
C2165 S.n1937 SUB 0.12fF $ **FLOATING
C2166 S.n1938 SUB 0.14fF $ **FLOATING
C2167 S.n1940 SUB 0.25fF $ **FLOATING
C2168 S.n1941 SUB 0.09fF $ **FLOATING
C2169 S.n1942 SUB 0.21fF $ **FLOATING
C2170 S.n1943 SUB 0.92fF $ **FLOATING
C2171 S.n1944 SUB 0.44fF $ **FLOATING
C2172 S.n1945 SUB 1.88fF $ **FLOATING
C2173 S.n1946 SUB 0.12fF $ **FLOATING
C2174 S.t1077 SUB 0.02fF
C2175 S.n1947 SUB 0.14fF $ **FLOATING
C2176 S.t1321 SUB 0.02fF
C2177 S.n1949 SUB 0.24fF $ **FLOATING
C2178 S.n1950 SUB 0.36fF $ **FLOATING
C2179 S.n1951 SUB 0.61fF $ **FLOATING
C2180 S.n1952 SUB 0.02fF $ **FLOATING
C2181 S.n1953 SUB 0.01fF $ **FLOATING
C2182 S.n1954 SUB 0.02fF $ **FLOATING
C2183 S.n1955 SUB 0.08fF $ **FLOATING
C2184 S.n1956 SUB 0.06fF $ **FLOATING
C2185 S.n1957 SUB 0.03fF $ **FLOATING
C2186 S.n1958 SUB 0.04fF $ **FLOATING
C2187 S.n1959 SUB 1.00fF $ **FLOATING
C2188 S.n1960 SUB 0.36fF $ **FLOATING
C2189 S.n1961 SUB 1.87fF $ **FLOATING
C2190 S.n1962 SUB 1.99fF $ **FLOATING
C2191 S.t2402 SUB 0.02fF
C2192 S.n1963 SUB 0.24fF $ **FLOATING
C2193 S.n1964 SUB 0.91fF $ **FLOATING
C2194 S.n1965 SUB 0.05fF $ **FLOATING
C2195 S.t1139 SUB 0.02fF
C2196 S.n1966 SUB 0.12fF $ **FLOATING
C2197 S.n1967 SUB 0.14fF $ **FLOATING
C2198 S.n1969 SUB 1.89fF $ **FLOATING
C2199 S.n1970 SUB 0.06fF $ **FLOATING
C2200 S.n1971 SUB 0.03fF $ **FLOATING
C2201 S.n1972 SUB 0.04fF $ **FLOATING
C2202 S.n1973 SUB 0.99fF $ **FLOATING
C2203 S.n1974 SUB 0.02fF $ **FLOATING
C2204 S.n1975 SUB 0.01fF $ **FLOATING
C2205 S.n1976 SUB 0.02fF $ **FLOATING
C2206 S.n1977 SUB 0.08fF $ **FLOATING
C2207 S.n1978 SUB 0.36fF $ **FLOATING
C2208 S.n1979 SUB 1.85fF $ **FLOATING
C2209 S.t441 SUB 0.02fF
C2210 S.n1980 SUB 0.24fF $ **FLOATING
C2211 S.n1981 SUB 0.36fF $ **FLOATING
C2212 S.n1982 SUB 0.61fF $ **FLOATING
C2213 S.n1983 SUB 0.12fF $ **FLOATING
C2214 S.t201 SUB 0.02fF
C2215 S.n1984 SUB 0.14fF $ **FLOATING
C2216 S.n1986 SUB 0.70fF $ **FLOATING
C2217 S.n1987 SUB 0.23fF $ **FLOATING
C2218 S.n1988 SUB 0.25fF $ **FLOATING
C2219 S.n1989 SUB 0.09fF $ **FLOATING
C2220 S.n1990 SUB 0.23fF $ **FLOATING
C2221 S.n1991 SUB 0.70fF $ **FLOATING
C2222 S.n1992 SUB 1.16fF $ **FLOATING
C2223 S.n1993 SUB 0.22fF $ **FLOATING
C2224 S.n1994 SUB 0.25fF $ **FLOATING
C2225 S.n1995 SUB 0.09fF $ **FLOATING
C2226 S.n1996 SUB 1.88fF $ **FLOATING
C2227 S.t1539 SUB 0.02fF
C2228 S.n1997 SUB 0.24fF $ **FLOATING
C2229 S.n1998 SUB 0.91fF $ **FLOATING
C2230 S.n1999 SUB 0.05fF $ **FLOATING
C2231 S.t263 SUB 0.02fF
C2232 S.n2000 SUB 0.12fF $ **FLOATING
C2233 S.n2001 SUB 0.14fF $ **FLOATING
C2234 S.n2003 SUB 0.25fF $ **FLOATING
C2235 S.n2004 SUB 0.09fF $ **FLOATING
C2236 S.n2005 SUB 0.21fF $ **FLOATING
C2237 S.n2006 SUB 0.92fF $ **FLOATING
C2238 S.n2007 SUB 0.44fF $ **FLOATING
C2239 S.n2008 SUB 1.88fF $ **FLOATING
C2240 S.n2009 SUB 0.12fF $ **FLOATING
C2241 S.t1866 SUB 0.02fF
C2242 S.n2010 SUB 0.14fF $ **FLOATING
C2243 S.t2086 SUB 0.02fF
C2244 S.n2012 SUB 0.24fF $ **FLOATING
C2245 S.n2013 SUB 0.36fF $ **FLOATING
C2246 S.n2014 SUB 0.61fF $ **FLOATING
C2247 S.n2015 SUB 0.02fF $ **FLOATING
C2248 S.n2016 SUB 0.01fF $ **FLOATING
C2249 S.n2017 SUB 0.02fF $ **FLOATING
C2250 S.n2018 SUB 0.08fF $ **FLOATING
C2251 S.n2019 SUB 0.06fF $ **FLOATING
C2252 S.n2020 SUB 0.03fF $ **FLOATING
C2253 S.n2021 SUB 0.04fF $ **FLOATING
C2254 S.n2022 SUB 1.00fF $ **FLOATING
C2255 S.n2023 SUB 0.36fF $ **FLOATING
C2256 S.n2024 SUB 1.87fF $ **FLOATING
C2257 S.n2025 SUB 1.99fF $ **FLOATING
C2258 S.t678 SUB 0.02fF
C2259 S.n2026 SUB 0.24fF $ **FLOATING
C2260 S.n2027 SUB 0.91fF $ **FLOATING
C2261 S.n2028 SUB 0.05fF $ **FLOATING
C2262 S.t1927 SUB 0.02fF
C2263 S.n2029 SUB 0.12fF $ **FLOATING
C2264 S.n2030 SUB 0.14fF $ **FLOATING
C2265 S.n2032 SUB 1.89fF $ **FLOATING
C2266 S.n2033 SUB 0.06fF $ **FLOATING
C2267 S.n2034 SUB 0.03fF $ **FLOATING
C2268 S.n2035 SUB 0.04fF $ **FLOATING
C2269 S.n2036 SUB 0.99fF $ **FLOATING
C2270 S.n2037 SUB 0.02fF $ **FLOATING
C2271 S.n2038 SUB 0.01fF $ **FLOATING
C2272 S.n2039 SUB 0.02fF $ **FLOATING
C2273 S.n2040 SUB 0.08fF $ **FLOATING
C2274 S.n2041 SUB 0.36fF $ **FLOATING
C2275 S.n2042 SUB 1.85fF $ **FLOATING
C2276 S.t1224 SUB 0.02fF
C2277 S.n2043 SUB 0.24fF $ **FLOATING
C2278 S.n2044 SUB 0.36fF $ **FLOATING
C2279 S.n2045 SUB 0.61fF $ **FLOATING
C2280 S.n2046 SUB 0.12fF $ **FLOATING
C2281 S.t999 SUB 0.02fF
C2282 S.n2047 SUB 0.14fF $ **FLOATING
C2283 S.n2049 SUB 0.70fF $ **FLOATING
C2284 S.n2050 SUB 0.23fF $ **FLOATING
C2285 S.n2051 SUB 0.25fF $ **FLOATING
C2286 S.n2052 SUB 0.09fF $ **FLOATING
C2287 S.n2053 SUB 0.23fF $ **FLOATING
C2288 S.n2054 SUB 0.70fF $ **FLOATING
C2289 S.n2055 SUB 1.16fF $ **FLOATING
C2290 S.n2056 SUB 0.22fF $ **FLOATING
C2291 S.n2057 SUB 0.25fF $ **FLOATING
C2292 S.n2058 SUB 0.09fF $ **FLOATING
C2293 S.n2059 SUB 1.88fF $ **FLOATING
C2294 S.t2338 SUB 0.02fF
C2295 S.n2060 SUB 0.24fF $ **FLOATING
C2296 S.n2061 SUB 0.91fF $ **FLOATING
C2297 S.n2062 SUB 0.05fF $ **FLOATING
C2298 S.t1172 SUB 0.02fF
C2299 S.n2063 SUB 0.12fF $ **FLOATING
C2300 S.n2064 SUB 0.14fF $ **FLOATING
C2301 S.n2066 SUB 0.25fF $ **FLOATING
C2302 S.n2067 SUB 0.09fF $ **FLOATING
C2303 S.n2068 SUB 0.21fF $ **FLOATING
C2304 S.n2069 SUB 0.92fF $ **FLOATING
C2305 S.n2070 SUB 0.44fF $ **FLOATING
C2306 S.n2071 SUB 1.88fF $ **FLOATING
C2307 S.n2072 SUB 0.12fF $ **FLOATING
C2308 S.t2128 SUB 0.02fF
C2309 S.n2073 SUB 0.14fF $ **FLOATING
C2310 S.t1025 SUB 0.02fF
C2311 S.n2075 SUB 0.24fF $ **FLOATING
C2312 S.n2076 SUB 0.36fF $ **FLOATING
C2313 S.n2077 SUB 0.61fF $ **FLOATING
C2314 S.n2078 SUB 0.02fF $ **FLOATING
C2315 S.n2079 SUB 0.01fF $ **FLOATING
C2316 S.n2080 SUB 0.02fF $ **FLOATING
C2317 S.n2081 SUB 0.08fF $ **FLOATING
C2318 S.n2082 SUB 0.06fF $ **FLOATING
C2319 S.n2083 SUB 0.03fF $ **FLOATING
C2320 S.n2084 SUB 0.04fF $ **FLOATING
C2321 S.n2085 SUB 1.00fF $ **FLOATING
C2322 S.n2086 SUB 0.36fF $ **FLOATING
C2323 S.n2087 SUB 1.87fF $ **FLOATING
C2324 S.n2088 SUB 1.99fF $ **FLOATING
C2325 S.t2563 SUB 0.02fF
C2326 S.n2089 SUB 0.24fF $ **FLOATING
C2327 S.n2090 SUB 0.91fF $ **FLOATING
C2328 S.n2091 SUB 0.05fF $ **FLOATING
C2329 S.t2316 SUB 0.02fF
C2330 S.n2092 SUB 0.12fF $ **FLOATING
C2331 S.n2093 SUB 0.14fF $ **FLOATING
C2332 S.n2095 SUB 1.89fF $ **FLOATING
C2333 S.n2096 SUB 0.06fF $ **FLOATING
C2334 S.n2097 SUB 0.03fF $ **FLOATING
C2335 S.n2098 SUB 0.04fF $ **FLOATING
C2336 S.n2099 SUB 0.99fF $ **FLOATING
C2337 S.n2100 SUB 0.02fF $ **FLOATING
C2338 S.n2101 SUB 0.01fF $ **FLOATING
C2339 S.n2102 SUB 0.02fF $ **FLOATING
C2340 S.n2103 SUB 0.08fF $ **FLOATING
C2341 S.n2104 SUB 0.36fF $ **FLOATING
C2342 S.n2105 SUB 1.85fF $ **FLOATING
C2343 S.t121 SUB 0.02fF
C2344 S.n2106 SUB 0.24fF $ **FLOATING
C2345 S.n2107 SUB 0.36fF $ **FLOATING
C2346 S.n2108 SUB 0.61fF $ **FLOATING
C2347 S.n2109 SUB 0.12fF $ **FLOATING
C2348 S.t1264 SUB 0.02fF
C2349 S.n2110 SUB 0.14fF $ **FLOATING
C2350 S.n2112 SUB 0.70fF $ **FLOATING
C2351 S.n2113 SUB 0.23fF $ **FLOATING
C2352 S.n2114 SUB 0.25fF $ **FLOATING
C2353 S.n2115 SUB 0.09fF $ **FLOATING
C2354 S.n2116 SUB 0.23fF $ **FLOATING
C2355 S.n2117 SUB 0.70fF $ **FLOATING
C2356 S.n2118 SUB 1.16fF $ **FLOATING
C2357 S.n2119 SUB 0.22fF $ **FLOATING
C2358 S.n2120 SUB 0.25fF $ **FLOATING
C2359 S.n2121 SUB 0.09fF $ **FLOATING
C2360 S.n2122 SUB 1.88fF $ **FLOATING
C2361 S.t1689 SUB 0.02fF
C2362 S.n2123 SUB 0.24fF $ **FLOATING
C2363 S.n2124 SUB 0.91fF $ **FLOATING
C2364 S.n2125 SUB 0.05fF $ **FLOATING
C2365 S.t1456 SUB 0.02fF
C2366 S.n2126 SUB 0.12fF $ **FLOATING
C2367 S.n2127 SUB 0.14fF $ **FLOATING
C2368 S.n2129 SUB 0.25fF $ **FLOATING
C2369 S.n2130 SUB 0.09fF $ **FLOATING
C2370 S.n2131 SUB 0.21fF $ **FLOATING
C2371 S.n2132 SUB 0.92fF $ **FLOATING
C2372 S.n2133 SUB 0.44fF $ **FLOATING
C2373 S.n2134 SUB 1.88fF $ **FLOATING
C2374 S.n2135 SUB 0.12fF $ **FLOATING
C2375 S.t381 SUB 0.02fF
C2376 S.n2136 SUB 0.14fF $ **FLOATING
C2377 S.t1792 SUB 0.02fF
C2378 S.n2138 SUB 0.24fF $ **FLOATING
C2379 S.n2139 SUB 0.36fF $ **FLOATING
C2380 S.n2140 SUB 0.61fF $ **FLOATING
C2381 S.n2141 SUB 0.02fF $ **FLOATING
C2382 S.n2142 SUB 0.01fF $ **FLOATING
C2383 S.n2143 SUB 0.02fF $ **FLOATING
C2384 S.n2144 SUB 0.08fF $ **FLOATING
C2385 S.n2145 SUB 0.06fF $ **FLOATING
C2386 S.n2146 SUB 0.03fF $ **FLOATING
C2387 S.n2147 SUB 0.04fF $ **FLOATING
C2388 S.n2148 SUB 1.00fF $ **FLOATING
C2389 S.n2149 SUB 0.36fF $ **FLOATING
C2390 S.n2150 SUB 1.83fF $ **FLOATING
C2391 S.n2151 SUB 1.99fF $ **FLOATING
C2392 S.t815 SUB 0.02fF
C2393 S.n2152 SUB 0.24fF $ **FLOATING
C2394 S.n2153 SUB 0.91fF $ **FLOATING
C2395 S.n2154 SUB 0.05fF $ **FLOATING
C2396 S.t598 SUB 0.02fF
C2397 S.n2155 SUB 0.12fF $ **FLOATING
C2398 S.n2156 SUB 0.14fF $ **FLOATING
C2399 S.n2158 SUB 1.89fF $ **FLOATING
C2400 S.n2159 SUB 0.63fF $ **FLOATING
C2401 S.n2160 SUB 0.04fF $ **FLOATING
C2402 S.n2161 SUB 0.07fF $ **FLOATING
C2403 S.n2162 SUB 0.05fF $ **FLOATING
C2404 S.n2163 SUB 0.87fF $ **FLOATING
C2405 S.n2164 SUB 0.01fF $ **FLOATING
C2406 S.n2165 SUB 0.01fF $ **FLOATING
C2407 S.n2166 SUB 0.01fF $ **FLOATING
C2408 S.n2167 SUB 0.07fF $ **FLOATING
C2409 S.n2168 SUB 0.68fF $ **FLOATING
C2410 S.n2169 SUB 0.13fF $ **FLOATING
C2411 S.t923 SUB 0.02fF
C2412 S.n2170 SUB 0.24fF $ **FLOATING
C2413 S.n2171 SUB 0.36fF $ **FLOATING
C2414 S.n2172 SUB 0.61fF $ **FLOATING
C2415 S.n2173 SUB 0.12fF $ **FLOATING
C2416 S.t2032 SUB 0.02fF
C2417 S.n2174 SUB 0.14fF $ **FLOATING
C2418 S.n2176 SUB 0.70fF $ **FLOATING
C2419 S.n2177 SUB 0.23fF $ **FLOATING
C2420 S.n2178 SUB 0.25fF $ **FLOATING
C2421 S.n2179 SUB 0.09fF $ **FLOATING
C2422 S.n2180 SUB 0.23fF $ **FLOATING
C2423 S.n2181 SUB 0.70fF $ **FLOATING
C2424 S.n2182 SUB 1.16fF $ **FLOATING
C2425 S.n2183 SUB 0.22fF $ **FLOATING
C2426 S.n2184 SUB 0.25fF $ **FLOATING
C2427 S.n2185 SUB 0.09fF $ **FLOATING
C2428 S.n2186 SUB 2.31fF $ **FLOATING
C2429 S.t2463 SUB 0.02fF
C2430 S.n2187 SUB 0.24fF $ **FLOATING
C2431 S.n2188 SUB 0.91fF $ **FLOATING
C2432 S.n2189 SUB 0.05fF $ **FLOATING
C2433 S.t2249 SUB 0.02fF
C2434 S.n2190 SUB 0.12fF $ **FLOATING
C2435 S.n2191 SUB 0.14fF $ **FLOATING
C2436 S.n2193 SUB 1.88fF $ **FLOATING
C2437 S.n2194 SUB 0.46fF $ **FLOATING
C2438 S.n2195 SUB 0.22fF $ **FLOATING
C2439 S.n2196 SUB 0.38fF $ **FLOATING
C2440 S.n2197 SUB 0.16fF $ **FLOATING
C2441 S.n2198 SUB 0.28fF $ **FLOATING
C2442 S.n2199 SUB 0.21fF $ **FLOATING
C2443 S.n2200 SUB 0.30fF $ **FLOATING
C2444 S.n2201 SUB 0.42fF $ **FLOATING
C2445 S.n2202 SUB 0.21fF $ **FLOATING
C2446 S.t183 SUB 0.02fF
C2447 S.n2203 SUB 0.24fF $ **FLOATING
C2448 S.n2204 SUB 0.36fF $ **FLOATING
C2449 S.n2205 SUB 0.61fF $ **FLOATING
C2450 S.n2206 SUB 0.12fF $ **FLOATING
C2451 S.t1317 SUB 0.02fF
C2452 S.n2207 SUB 0.14fF $ **FLOATING
C2453 S.n2209 SUB 0.04fF $ **FLOATING
C2454 S.n2210 SUB 0.03fF $ **FLOATING
C2455 S.n2211 SUB 0.03fF $ **FLOATING
C2456 S.n2212 SUB 0.10fF $ **FLOATING
C2457 S.n2213 SUB 0.36fF $ **FLOATING
C2458 S.n2214 SUB 0.38fF $ **FLOATING
C2459 S.n2215 SUB 0.11fF $ **FLOATING
C2460 S.n2216 SUB 0.12fF $ **FLOATING
C2461 S.n2217 SUB 0.07fF $ **FLOATING
C2462 S.n2218 SUB 0.12fF $ **FLOATING
C2463 S.n2219 SUB 0.18fF $ **FLOATING
C2464 S.n2220 SUB 4.00fF $ **FLOATING
C2465 S.t1750 SUB 0.02fF
C2466 S.n2221 SUB 0.24fF $ **FLOATING
C2467 S.n2222 SUB 0.91fF $ **FLOATING
C2468 S.n2223 SUB 0.05fF $ **FLOATING
C2469 S.t1391 SUB 0.02fF
C2470 S.n2224 SUB 0.12fF $ **FLOATING
C2471 S.n2225 SUB 0.14fF $ **FLOATING
C2472 S.n2227 SUB 0.25fF $ **FLOATING
C2473 S.n2228 SUB 0.09fF $ **FLOATING
C2474 S.n2229 SUB 0.21fF $ **FLOATING
C2475 S.n2230 SUB 1.28fF $ **FLOATING
C2476 S.n2231 SUB 0.53fF $ **FLOATING
C2477 S.n2232 SUB 1.88fF $ **FLOATING
C2478 S.n2233 SUB 0.12fF $ **FLOATING
C2479 S.t438 SUB 0.02fF
C2480 S.n2234 SUB 0.14fF $ **FLOATING
C2481 S.t1847 SUB 0.02fF
C2482 S.n2236 SUB 0.24fF $ **FLOATING
C2483 S.n2237 SUB 0.36fF $ **FLOATING
C2484 S.n2238 SUB 0.61fF $ **FLOATING
C2485 S.n2239 SUB 0.71fF $ **FLOATING
C2486 S.n2240 SUB 1.58fF $ **FLOATING
C2487 S.n2241 SUB 2.45fF $ **FLOATING
C2488 S.t871 SUB 0.02fF
C2489 S.n2242 SUB 0.24fF $ **FLOATING
C2490 S.n2243 SUB 0.91fF $ **FLOATING
C2491 S.n2244 SUB 0.05fF $ **FLOATING
C2492 S.t519 SUB 0.02fF
C2493 S.n2245 SUB 0.12fF $ **FLOATING
C2494 S.n2246 SUB 0.14fF $ **FLOATING
C2495 S.n2248 SUB 1.89fF $ **FLOATING
C2496 S.n2249 SUB 0.06fF $ **FLOATING
C2497 S.n2250 SUB 0.03fF $ **FLOATING
C2498 S.n2251 SUB 0.04fF $ **FLOATING
C2499 S.n2252 SUB 0.99fF $ **FLOATING
C2500 S.n2253 SUB 0.02fF $ **FLOATING
C2501 S.n2254 SUB 0.01fF $ **FLOATING
C2502 S.n2255 SUB 0.02fF $ **FLOATING
C2503 S.n2256 SUB 0.08fF $ **FLOATING
C2504 S.n2257 SUB 0.36fF $ **FLOATING
C2505 S.n2258 SUB 1.85fF $ **FLOATING
C2506 S.t985 SUB 0.02fF
C2507 S.n2259 SUB 0.24fF $ **FLOATING
C2508 S.n2260 SUB 0.36fF $ **FLOATING
C2509 S.n2261 SUB 0.61fF $ **FLOATING
C2510 S.n2262 SUB 0.12fF $ **FLOATING
C2511 S.t2082 SUB 0.02fF
C2512 S.n2263 SUB 0.14fF $ **FLOATING
C2513 S.n2265 SUB 0.70fF $ **FLOATING
C2514 S.n2266 SUB 0.23fF $ **FLOATING
C2515 S.n2267 SUB 0.25fF $ **FLOATING
C2516 S.n2268 SUB 0.09fF $ **FLOATING
C2517 S.n2269 SUB 0.23fF $ **FLOATING
C2518 S.n2270 SUB 0.70fF $ **FLOATING
C2519 S.n2271 SUB 1.16fF $ **FLOATING
C2520 S.n2272 SUB 0.22fF $ **FLOATING
C2521 S.n2273 SUB 0.25fF $ **FLOATING
C2522 S.n2274 SUB 0.09fF $ **FLOATING
C2523 S.n2275 SUB 1.88fF $ **FLOATING
C2524 S.t2517 SUB 0.02fF
C2525 S.n2276 SUB 0.24fF $ **FLOATING
C2526 S.n2277 SUB 0.91fF $ **FLOATING
C2527 S.n2278 SUB 0.05fF $ **FLOATING
C2528 S.t2164 SUB 0.02fF
C2529 S.n2279 SUB 0.12fF $ **FLOATING
C2530 S.n2280 SUB 0.14fF $ **FLOATING
C2531 S.n2282 SUB 20.78fF $ **FLOATING
C2532 S.n2283 SUB 0.06fF $ **FLOATING
C2533 S.n2284 SUB 0.20fF $ **FLOATING
C2534 S.n2285 SUB 0.09fF $ **FLOATING
C2535 S.n2286 SUB 0.21fF $ **FLOATING
C2536 S.n2287 SUB 0.10fF $ **FLOATING
C2537 S.n2288 SUB 0.30fF $ **FLOATING
C2538 S.n2289 SUB 0.69fF $ **FLOATING
C2539 S.n2290 SUB 0.45fF $ **FLOATING
C2540 S.n2291 SUB 2.33fF $ **FLOATING
C2541 S.n2292 SUB 0.12fF $ **FLOATING
C2542 S.t1902 SUB 0.02fF
C2543 S.n2293 SUB 0.14fF $ **FLOATING
C2544 S.t2136 SUB 0.02fF
C2545 S.n2295 SUB 0.24fF $ **FLOATING
C2546 S.n2296 SUB 0.36fF $ **FLOATING
C2547 S.n2297 SUB 0.61fF $ **FLOATING
C2548 S.n2298 SUB 1.90fF $ **FLOATING
C2549 S.n2299 SUB 0.17fF $ **FLOATING
C2550 S.n2300 SUB 0.76fF $ **FLOATING
C2551 S.n2301 SUB 0.32fF $ **FLOATING
C2552 S.n2302 SUB 0.25fF $ **FLOATING
C2553 S.n2303 SUB 0.30fF $ **FLOATING
C2554 S.n2304 SUB 0.47fF $ **FLOATING
C2555 S.n2305 SUB 0.16fF $ **FLOATING
C2556 S.n2306 SUB 1.93fF $ **FLOATING
C2557 S.t2072 SUB 0.02fF
C2558 S.n2307 SUB 0.12fF $ **FLOATING
C2559 S.n2308 SUB 0.14fF $ **FLOATING
C2560 S.t705 SUB 0.02fF
C2561 S.n2310 SUB 0.24fF $ **FLOATING
C2562 S.n2311 SUB 0.91fF $ **FLOATING
C2563 S.n2312 SUB 0.05fF $ **FLOATING
C2564 S.n2313 SUB 1.88fF $ **FLOATING
C2565 S.n2314 SUB 0.12fF $ **FLOATING
C2566 S.t2253 SUB 0.02fF
C2567 S.n2315 SUB 0.14fF $ **FLOATING
C2568 S.t1245 SUB 0.02fF
C2569 S.n2317 SUB 1.22fF $ **FLOATING
C2570 S.n2318 SUB 0.36fF $ **FLOATING
C2571 S.n2319 SUB 1.22fF $ **FLOATING
C2572 S.n2320 SUB 0.61fF $ **FLOATING
C2573 S.n2321 SUB 0.35fF $ **FLOATING
C2574 S.n2322 SUB 0.63fF $ **FLOATING
C2575 S.n2323 SUB 1.15fF $ **FLOATING
C2576 S.n2324 SUB 3.03fF $ **FLOATING
C2577 S.n2325 SUB 0.59fF $ **FLOATING
C2578 S.n2326 SUB 0.02fF $ **FLOATING
C2579 S.n2327 SUB 0.97fF $ **FLOATING
C2580 S.t215 SUB 21.38fF
C2581 S.n2328 SUB 20.25fF $ **FLOATING
C2582 S.n2330 SUB 0.38fF $ **FLOATING
C2583 S.n2331 SUB 0.23fF $ **FLOATING
C2584 S.n2332 SUB 2.79fF $ **FLOATING
C2585 S.n2333 SUB 2.46fF $ **FLOATING
C2586 S.n2334 SUB 4.00fF $ **FLOATING
C2587 S.n2335 SUB 0.25fF $ **FLOATING
C2588 S.n2336 SUB 0.01fF $ **FLOATING
C2589 S.t982 SUB 0.02fF
C2590 S.n2337 SUB 0.25fF $ **FLOATING
C2591 S.t406 SUB 0.02fF
C2592 S.n2338 SUB 0.95fF $ **FLOATING
C2593 S.n2339 SUB 0.70fF $ **FLOATING
C2594 S.n2340 SUB 1.89fF $ **FLOATING
C2595 S.n2341 SUB 1.88fF $ **FLOATING
C2596 S.t363 SUB 0.02fF
C2597 S.n2342 SUB 0.24fF $ **FLOATING
C2598 S.n2343 SUB 0.36fF $ **FLOATING
C2599 S.n2344 SUB 0.61fF $ **FLOATING
C2600 S.n2345 SUB 0.12fF $ **FLOATING
C2601 S.t56 SUB 0.02fF
C2602 S.n2346 SUB 0.14fF $ **FLOATING
C2603 S.n2348 SUB 1.16fF $ **FLOATING
C2604 S.n2349 SUB 0.22fF $ **FLOATING
C2605 S.n2350 SUB 0.25fF $ **FLOATING
C2606 S.n2351 SUB 0.09fF $ **FLOATING
C2607 S.n2352 SUB 1.88fF $ **FLOATING
C2608 S.t2054 SUB 0.02fF
C2609 S.n2353 SUB 0.24fF $ **FLOATING
C2610 S.n2354 SUB 0.91fF $ **FLOATING
C2611 S.n2355 SUB 0.05fF $ **FLOATING
C2612 S.t743 SUB 0.02fF
C2613 S.n2356 SUB 0.12fF $ **FLOATING
C2614 S.n2357 SUB 0.14fF $ **FLOATING
C2615 S.n2359 SUB 0.78fF $ **FLOATING
C2616 S.n2360 SUB 1.94fF $ **FLOATING
C2617 S.n2361 SUB 1.88fF $ **FLOATING
C2618 S.n2362 SUB 0.12fF $ **FLOATING
C2619 S.t1746 SUB 0.02fF
C2620 S.n2363 SUB 0.14fF $ **FLOATING
C2621 S.t2015 SUB 0.02fF
C2622 S.n2365 SUB 0.24fF $ **FLOATING
C2623 S.n2366 SUB 0.36fF $ **FLOATING
C2624 S.n2367 SUB 0.61fF $ **FLOATING
C2625 S.n2368 SUB 1.84fF $ **FLOATING
C2626 S.n2369 SUB 2.99fF $ **FLOATING
C2627 S.t1194 SUB 0.02fF
C2628 S.n2370 SUB 0.24fF $ **FLOATING
C2629 S.n2371 SUB 0.91fF $ **FLOATING
C2630 S.n2372 SUB 0.05fF $ **FLOATING
C2631 S.t2394 SUB 0.02fF
C2632 S.n2373 SUB 0.12fF $ **FLOATING
C2633 S.n2374 SUB 0.14fF $ **FLOATING
C2634 S.n2376 SUB 1.89fF $ **FLOATING
C2635 S.n2377 SUB 1.88fF $ **FLOATING
C2636 S.t1162 SUB 0.02fF
C2637 S.n2378 SUB 0.24fF $ **FLOATING
C2638 S.n2379 SUB 0.36fF $ **FLOATING
C2639 S.n2380 SUB 0.61fF $ **FLOATING
C2640 S.n2381 SUB 0.12fF $ **FLOATING
C2641 S.t870 SUB 0.02fF
C2642 S.n2382 SUB 0.14fF $ **FLOATING
C2643 S.n2384 SUB 1.16fF $ **FLOATING
C2644 S.n2385 SUB 0.22fF $ **FLOATING
C2645 S.n2386 SUB 0.25fF $ **FLOATING
C2646 S.n2387 SUB 0.09fF $ **FLOATING
C2647 S.n2388 SUB 1.88fF $ **FLOATING
C2648 S.t315 SUB 0.02fF
C2649 S.n2389 SUB 0.24fF $ **FLOATING
C2650 S.n2390 SUB 0.91fF $ **FLOATING
C2651 S.n2391 SUB 0.05fF $ **FLOATING
C2652 S.t1656 SUB 0.02fF
C2653 S.n2392 SUB 0.12fF $ **FLOATING
C2654 S.n2393 SUB 0.14fF $ **FLOATING
C2655 S.n2395 SUB 0.78fF $ **FLOATING
C2656 S.n2396 SUB 1.94fF $ **FLOATING
C2657 S.n2397 SUB 1.88fF $ **FLOATING
C2658 S.n2398 SUB 0.12fF $ **FLOATING
C2659 S.t2514 SUB 0.02fF
C2660 S.n2399 SUB 0.14fF $ **FLOATING
C2661 S.t290 SUB 0.02fF
C2662 S.n2401 SUB 0.24fF $ **FLOATING
C2663 S.n2402 SUB 0.36fF $ **FLOATING
C2664 S.n2403 SUB 0.61fF $ **FLOATING
C2665 S.n2404 SUB 1.84fF $ **FLOATING
C2666 S.n2405 SUB 2.99fF $ **FLOATING
C2667 S.t1980 SUB 0.02fF
C2668 S.n2406 SUB 0.24fF $ **FLOATING
C2669 S.n2407 SUB 0.91fF $ **FLOATING
C2670 S.n2408 SUB 0.05fF $ **FLOATING
C2671 S.t786 SUB 0.02fF
C2672 S.n2409 SUB 0.12fF $ **FLOATING
C2673 S.n2410 SUB 0.14fF $ **FLOATING
C2674 S.n2412 SUB 1.89fF $ **FLOATING
C2675 S.n2413 SUB 1.88fF $ **FLOATING
C2676 S.t1953 SUB 0.02fF
C2677 S.n2414 SUB 0.24fF $ **FLOATING
C2678 S.n2415 SUB 0.36fF $ **FLOATING
C2679 S.n2416 SUB 0.61fF $ **FLOATING
C2680 S.n2417 SUB 0.12fF $ **FLOATING
C2681 S.t1638 SUB 0.02fF
C2682 S.n2418 SUB 0.14fF $ **FLOATING
C2683 S.n2420 SUB 1.16fF $ **FLOATING
C2684 S.n2421 SUB 0.22fF $ **FLOATING
C2685 S.n2422 SUB 0.25fF $ **FLOATING
C2686 S.n2423 SUB 0.09fF $ **FLOATING
C2687 S.n2424 SUB 1.88fF $ **FLOATING
C2688 S.t1127 SUB 0.02fF
C2689 S.n2425 SUB 0.24fF $ **FLOATING
C2690 S.n2426 SUB 0.91fF $ **FLOATING
C2691 S.n2427 SUB 0.05fF $ **FLOATING
C2692 S.t2437 SUB 0.02fF
C2693 S.n2428 SUB 0.12fF $ **FLOATING
C2694 S.n2429 SUB 0.14fF $ **FLOATING
C2695 S.n2431 SUB 0.78fF $ **FLOATING
C2696 S.n2432 SUB 1.94fF $ **FLOATING
C2697 S.n2433 SUB 1.88fF $ **FLOATING
C2698 S.n2434 SUB 0.12fF $ **FLOATING
C2699 S.t771 SUB 0.02fF
C2700 S.n2435 SUB 0.14fF $ **FLOATING
C2701 S.t1093 SUB 0.02fF
C2702 S.n2437 SUB 0.24fF $ **FLOATING
C2703 S.n2438 SUB 0.36fF $ **FLOATING
C2704 S.n2439 SUB 0.61fF $ **FLOATING
C2705 S.n2440 SUB 1.84fF $ **FLOATING
C2706 S.n2441 SUB 2.99fF $ **FLOATING
C2707 S.t249 SUB 0.02fF
C2708 S.n2442 SUB 0.24fF $ **FLOATING
C2709 S.n2443 SUB 0.91fF $ **FLOATING
C2710 S.n2444 SUB 0.05fF $ **FLOATING
C2711 S.t1573 SUB 0.02fF
C2712 S.n2445 SUB 0.12fF $ **FLOATING
C2713 S.n2446 SUB 0.14fF $ **FLOATING
C2714 S.n2448 SUB 1.89fF $ **FLOATING
C2715 S.n2449 SUB 1.88fF $ **FLOATING
C2716 S.t216 SUB 0.02fF
C2717 S.n2450 SUB 0.24fF $ **FLOATING
C2718 S.n2451 SUB 0.36fF $ **FLOATING
C2719 S.n2452 SUB 0.61fF $ **FLOATING
C2720 S.n2453 SUB 0.12fF $ **FLOATING
C2721 S.t2571 SUB 0.02fF
C2722 S.n2454 SUB 0.14fF $ **FLOATING
C2723 S.n2456 SUB 1.16fF $ **FLOATING
C2724 S.n2457 SUB 0.22fF $ **FLOATING
C2725 S.n2458 SUB 0.25fF $ **FLOATING
C2726 S.n2459 SUB 0.09fF $ **FLOATING
C2727 S.n2460 SUB 1.88fF $ **FLOATING
C2728 S.t1913 SUB 0.02fF
C2729 S.n2461 SUB 0.24fF $ **FLOATING
C2730 S.n2462 SUB 0.91fF $ **FLOATING
C2731 S.n2463 SUB 0.05fF $ **FLOATING
C2732 S.t703 SUB 0.02fF
C2733 S.n2464 SUB 0.12fF $ **FLOATING
C2734 S.n2465 SUB 0.14fF $ **FLOATING
C2735 S.n2467 SUB 0.78fF $ **FLOATING
C2736 S.n2468 SUB 1.94fF $ **FLOATING
C2737 S.n2469 SUB 1.88fF $ **FLOATING
C2738 S.n2470 SUB 0.12fF $ **FLOATING
C2739 S.t727 SUB 0.02fF
C2740 S.n2471 SUB 0.14fF $ **FLOATING
C2741 S.t2509 SUB 0.02fF
C2742 S.n2473 SUB 0.24fF $ **FLOATING
C2743 S.n2474 SUB 0.36fF $ **FLOATING
C2744 S.n2475 SUB 0.61fF $ **FLOATING
C2745 S.n2476 SUB 1.84fF $ **FLOATING
C2746 S.n2477 SUB 2.99fF $ **FLOATING
C2747 S.t1814 SUB 0.02fF
C2748 S.n2478 SUB 0.24fF $ **FLOATING
C2749 S.n2479 SUB 0.91fF $ **FLOATING
C2750 S.n2480 SUB 0.05fF $ **FLOATING
C2751 S.t2362 SUB 0.02fF
C2752 S.n2481 SUB 0.12fF $ **FLOATING
C2753 S.n2482 SUB 0.14fF $ **FLOATING
C2754 S.n2484 SUB 1.89fF $ **FLOATING
C2755 S.n2485 SUB 1.88fF $ **FLOATING
C2756 S.t1633 SUB 0.02fF
C2757 S.n2486 SUB 0.24fF $ **FLOATING
C2758 S.n2487 SUB 0.36fF $ **FLOATING
C2759 S.n2488 SUB 0.61fF $ **FLOATING
C2760 S.n2489 SUB 0.12fF $ **FLOATING
C2761 S.t2379 SUB 0.02fF
C2762 S.n2490 SUB 0.14fF $ **FLOATING
C2763 S.n2492 SUB 1.16fF $ **FLOATING
C2764 S.n2493 SUB 0.22fF $ **FLOATING
C2765 S.n2494 SUB 0.25fF $ **FLOATING
C2766 S.n2495 SUB 0.09fF $ **FLOATING
C2767 S.n2496 SUB 1.88fF $ **FLOATING
C2768 S.t947 SUB 0.02fF
C2769 S.n2497 SUB 0.24fF $ **FLOATING
C2770 S.n2498 SUB 0.91fF $ **FLOATING
C2771 S.n2499 SUB 0.05fF $ **FLOATING
C2772 S.t574 SUB 0.02fF
C2773 S.n2500 SUB 0.12fF $ **FLOATING
C2774 S.n2501 SUB 0.14fF $ **FLOATING
C2775 S.n2503 SUB 0.78fF $ **FLOATING
C2776 S.n2504 SUB 1.94fF $ **FLOATING
C2777 S.n2505 SUB 1.88fF $ **FLOATING
C2778 S.n2506 SUB 0.12fF $ **FLOATING
C2779 S.t1523 SUB 0.02fF
C2780 S.n2507 SUB 0.14fF $ **FLOATING
C2781 S.t769 SUB 0.02fF
C2782 S.n2509 SUB 0.24fF $ **FLOATING
C2783 S.n2510 SUB 0.36fF $ **FLOATING
C2784 S.n2511 SUB 0.61fF $ **FLOATING
C2785 S.n2512 SUB 1.84fF $ **FLOATING
C2786 S.n2513 SUB 2.99fF $ **FLOATING
C2787 S.t2586 SUB 0.02fF
C2788 S.n2514 SUB 0.24fF $ **FLOATING
C2789 S.n2515 SUB 0.91fF $ **FLOATING
C2790 S.n2516 SUB 0.05fF $ **FLOATING
C2791 S.t2219 SUB 0.02fF
C2792 S.n2517 SUB 0.12fF $ **FLOATING
C2793 S.n2518 SUB 0.14fF $ **FLOATING
C2794 S.n2520 SUB 1.89fF $ **FLOATING
C2795 S.n2521 SUB 1.75fF $ **FLOATING
C2796 S.t2420 SUB 0.02fF
C2797 S.n2522 SUB 0.24fF $ **FLOATING
C2798 S.n2523 SUB 0.36fF $ **FLOATING
C2799 S.n2524 SUB 0.61fF $ **FLOATING
C2800 S.n2525 SUB 0.12fF $ **FLOATING
C2801 S.t662 SUB 0.02fF
C2802 S.n2526 SUB 0.14fF $ **FLOATING
C2803 S.n2528 SUB 1.16fF $ **FLOATING
C2804 S.n2529 SUB 0.22fF $ **FLOATING
C2805 S.n2530 SUB 0.25fF $ **FLOATING
C2806 S.n2531 SUB 0.09fF $ **FLOATING
C2807 S.n2532 SUB 2.44fF $ **FLOATING
C2808 S.t1709 SUB 0.02fF
C2809 S.n2533 SUB 0.24fF $ **FLOATING
C2810 S.n2534 SUB 0.91fF $ **FLOATING
C2811 S.n2535 SUB 0.05fF $ **FLOATING
C2812 S.t1359 SUB 0.02fF
C2813 S.n2536 SUB 0.12fF $ **FLOATING
C2814 S.n2537 SUB 0.14fF $ **FLOATING
C2815 S.n2539 SUB 1.88fF $ **FLOATING
C2816 S.n2540 SUB 0.48fF $ **FLOATING
C2817 S.n2541 SUB 0.09fF $ **FLOATING
C2818 S.n2542 SUB 0.33fF $ **FLOATING
C2819 S.n2543 SUB 0.30fF $ **FLOATING
C2820 S.n2544 SUB 0.77fF $ **FLOATING
C2821 S.n2545 SUB 0.59fF $ **FLOATING
C2822 S.t1554 SUB 0.02fF
C2823 S.n2546 SUB 0.24fF $ **FLOATING
C2824 S.n2547 SUB 0.36fF $ **FLOATING
C2825 S.n2548 SUB 0.61fF $ **FLOATING
C2826 S.n2549 SUB 0.12fF $ **FLOATING
C2827 S.t2317 SUB 0.02fF
C2828 S.n2550 SUB 0.14fF $ **FLOATING
C2829 S.n2552 SUB 2.61fF $ **FLOATING
C2830 S.n2553 SUB 2.16fF $ **FLOATING
C2831 S.t839 SUB 0.02fF
C2832 S.n2554 SUB 0.24fF $ **FLOATING
C2833 S.n2555 SUB 0.91fF $ **FLOATING
C2834 S.n2556 SUB 0.05fF $ **FLOATING
C2835 S.t482 SUB 0.02fF
C2836 S.n2557 SUB 0.12fF $ **FLOATING
C2837 S.n2558 SUB 0.14fF $ **FLOATING
C2838 S.n2560 SUB 0.78fF $ **FLOATING
C2839 S.n2561 SUB 2.30fF $ **FLOATING
C2840 S.n2562 SUB 1.88fF $ **FLOATING
C2841 S.n2563 SUB 0.12fF $ **FLOATING
C2842 S.t1457 SUB 0.02fF
C2843 S.n2564 SUB 0.14fF $ **FLOATING
C2844 S.t691 SUB 0.02fF
C2845 S.n2566 SUB 0.24fF $ **FLOATING
C2846 S.n2567 SUB 0.36fF $ **FLOATING
C2847 S.n2568 SUB 0.61fF $ **FLOATING
C2848 S.n2569 SUB 1.39fF $ **FLOATING
C2849 S.n2570 SUB 0.71fF $ **FLOATING
C2850 S.n2571 SUB 1.14fF $ **FLOATING
C2851 S.n2572 SUB 0.35fF $ **FLOATING
C2852 S.n2573 SUB 2.03fF $ **FLOATING
C2853 S.t2482 SUB 0.02fF
C2854 S.n2574 SUB 0.24fF $ **FLOATING
C2855 S.n2575 SUB 0.91fF $ **FLOATING
C2856 S.n2576 SUB 0.05fF $ **FLOATING
C2857 S.t2263 SUB 0.02fF
C2858 S.n2577 SUB 0.12fF $ **FLOATING
C2859 S.n2578 SUB 0.14fF $ **FLOATING
C2860 S.n2580 SUB 1.89fF $ **FLOATING
C2861 S.n2581 SUB 1.88fF $ **FLOATING
C2862 S.t2352 SUB 0.02fF
C2863 S.n2582 SUB 0.24fF $ **FLOATING
C2864 S.n2583 SUB 0.36fF $ **FLOATING
C2865 S.n2584 SUB 0.61fF $ **FLOATING
C2866 S.n2585 SUB 0.12fF $ **FLOATING
C2867 S.t599 SUB 0.02fF
C2868 S.n2586 SUB 0.14fF $ **FLOATING
C2869 S.n2588 SUB 1.16fF $ **FLOATING
C2870 S.n2589 SUB 0.22fF $ **FLOATING
C2871 S.n2590 SUB 0.25fF $ **FLOATING
C2872 S.n2591 SUB 0.09fF $ **FLOATING
C2873 S.n2592 SUB 1.88fF $ **FLOATING
C2874 S.t1609 SUB 0.02fF
C2875 S.n2593 SUB 0.24fF $ **FLOATING
C2876 S.n2594 SUB 0.91fF $ **FLOATING
C2877 S.n2595 SUB 0.05fF $ **FLOATING
C2878 S.t1405 SUB 0.02fF
C2879 S.n2596 SUB 0.12fF $ **FLOATING
C2880 S.n2597 SUB 0.14fF $ **FLOATING
C2881 S.n2599 SUB 20.78fF $ **FLOATING
C2882 S.n2600 SUB 2.73fF $ **FLOATING
C2883 S.n2601 SUB 1.59fF $ **FLOATING
C2884 S.n2602 SUB 0.12fF $ **FLOATING
C2885 S.t2069 SUB 0.02fF
C2886 S.n2603 SUB 0.14fF $ **FLOATING
C2887 S.t2116 SUB 0.02fF
C2888 S.n2605 SUB 0.24fF $ **FLOATING
C2889 S.n2606 SUB 0.36fF $ **FLOATING
C2890 S.n2607 SUB 0.61fF $ **FLOATING
C2891 S.n2608 SUB 0.07fF $ **FLOATING
C2892 S.n2609 SUB 0.01fF $ **FLOATING
C2893 S.n2610 SUB 0.24fF $ **FLOATING
C2894 S.n2611 SUB 1.16fF $ **FLOATING
C2895 S.n2612 SUB 1.35fF $ **FLOATING
C2896 S.n2613 SUB 2.30fF $ **FLOATING
C2897 S.t296 SUB 0.02fF
C2898 S.n2614 SUB 0.12fF $ **FLOATING
C2899 S.n2615 SUB 0.14fF $ **FLOATING
C2900 S.t586 SUB 0.02fF
C2901 S.n2617 SUB 0.24fF $ **FLOATING
C2902 S.n2618 SUB 0.91fF $ **FLOATING
C2903 S.n2619 SUB 0.05fF $ **FLOATING
C2904 S.t55 SUB 48.31fF
C2905 S.t536 SUB 0.02fF
C2906 S.n2620 SUB 0.12fF $ **FLOATING
C2907 S.n2621 SUB 0.14fF $ **FLOATING
C2908 S.t745 SUB 0.02fF
C2909 S.n2623 SUB 0.24fF $ **FLOATING
C2910 S.n2624 SUB 0.91fF $ **FLOATING
C2911 S.n2625 SUB 0.05fF $ **FLOATING
C2912 S.t1494 SUB 0.02fF
C2913 S.n2626 SUB 0.24fF $ **FLOATING
C2914 S.n2627 SUB 0.36fF $ **FLOATING
C2915 S.n2628 SUB 0.61fF $ **FLOATING
C2916 S.n2629 SUB 0.32fF $ **FLOATING
C2917 S.n2630 SUB 1.09fF $ **FLOATING
C2918 S.n2631 SUB 0.15fF $ **FLOATING
C2919 S.n2632 SUB 2.10fF $ **FLOATING
C2920 S.n2633 SUB 2.94fF $ **FLOATING
C2921 S.n2634 SUB 1.88fF $ **FLOATING
C2922 S.n2635 SUB 0.12fF $ **FLOATING
C2923 S.t1220 SUB 0.02fF
C2924 S.n2636 SUB 0.14fF $ **FLOATING
C2925 S.t64 SUB 0.02fF
C2926 S.n2638 SUB 0.24fF $ **FLOATING
C2927 S.n2639 SUB 0.36fF $ **FLOATING
C2928 S.n2640 SUB 0.61fF $ **FLOATING
C2929 S.n2641 SUB 0.92fF $ **FLOATING
C2930 S.n2642 SUB 0.32fF $ **FLOATING
C2931 S.n2643 SUB 0.92fF $ **FLOATING
C2932 S.n2644 SUB 1.09fF $ **FLOATING
C2933 S.n2645 SUB 0.15fF $ **FLOATING
C2934 S.n2646 SUB 4.68fF $ **FLOATING
C2935 S.t1301 SUB 0.02fF
C2936 S.n2647 SUB 0.12fF $ **FLOATING
C2937 S.n2648 SUB 0.14fF $ **FLOATING
C2938 S.t1640 SUB 0.02fF
C2939 S.n2650 SUB 0.24fF $ **FLOATING
C2940 S.n2651 SUB 0.91fF $ **FLOATING
C2941 S.n2652 SUB 0.05fF $ **FLOATING
C2942 S.n2653 SUB 1.88fF $ **FLOATING
C2943 S.n2654 SUB 2.67fF $ **FLOATING
C2944 S.t345 SUB 0.02fF
C2945 S.n2655 SUB 0.24fF $ **FLOATING
C2946 S.n2656 SUB 0.36fF $ **FLOATING
C2947 S.n2657 SUB 0.61fF $ **FLOATING
C2948 S.n2658 SUB 0.12fF $ **FLOATING
C2949 S.t2250 SUB 0.02fF
C2950 S.n2659 SUB 0.14fF $ **FLOATING
C2951 S.n2661 SUB 1.88fF $ **FLOATING
C2952 S.n2662 SUB 2.68fF $ **FLOATING
C2953 S.t631 SUB 0.02fF
C2954 S.n2663 SUB 0.24fF $ **FLOATING
C2955 S.n2664 SUB 0.36fF $ **FLOATING
C2956 S.n2665 SUB 0.61fF $ **FLOATING
C2957 S.t2396 SUB 0.02fF
C2958 S.n2666 SUB 0.24fF $ **FLOATING
C2959 S.n2667 SUB 0.91fF $ **FLOATING
C2960 S.n2668 SUB 0.05fF $ **FLOATING
C2961 S.t2180 SUB 0.02fF
C2962 S.n2669 SUB 0.12fF $ **FLOATING
C2963 S.n2670 SUB 0.14fF $ **FLOATING
C2964 S.n2672 SUB 0.12fF $ **FLOATING
C2965 S.t1394 SUB 0.02fF
C2966 S.n2673 SUB 0.14fF $ **FLOATING
C2967 S.n2675 SUB 5.18fF $ **FLOATING
C2968 S.n2676 SUB 5.46fF $ **FLOATING
C2969 S.t417 SUB 0.02fF
C2970 S.n2677 SUB 0.12fF $ **FLOATING
C2971 S.n2678 SUB 0.14fF $ **FLOATING
C2972 S.t2296 SUB 0.02fF
C2973 S.n2680 SUB 0.24fF $ **FLOATING
C2974 S.n2681 SUB 0.91fF $ **FLOATING
C2975 S.n2682 SUB 0.05fF $ **FLOATING
C2976 S.t200 SUB 47.92fF
C2977 S.t1720 SUB 0.02fF
C2978 S.n2683 SUB 1.19fF $ **FLOATING
C2979 S.n2684 SUB 0.05fF $ **FLOATING
C2980 S.t1488 SUB 0.02fF
C2981 S.n2685 SUB 0.01fF $ **FLOATING
C2982 S.n2686 SUB 0.26fF $ **FLOATING
C2983 S.n2688 SUB 1.50fF $ **FLOATING
C2984 S.n2689 SUB 1.30fF $ **FLOATING
C2985 S.n2690 SUB 0.28fF $ **FLOATING
C2986 S.n2691 SUB 0.24fF $ **FLOATING
C2987 S.n2692 SUB 4.39fF $ **FLOATING
C2988 S.n2693 SUB 0.01fF $ **FLOATING
C2989 S.n2694 SUB 0.02fF $ **FLOATING
C2990 S.n2695 SUB 0.03fF $ **FLOATING
C2991 S.n2696 SUB 0.04fF $ **FLOATING
C2992 S.n2697 SUB 0.17fF $ **FLOATING
C2993 S.n2698 SUB 0.01fF $ **FLOATING
C2994 S.n2699 SUB 0.02fF $ **FLOATING
C2995 S.n2700 SUB 0.01fF $ **FLOATING
C2996 S.n2701 SUB 0.01fF $ **FLOATING
C2997 S.n2702 SUB 0.01fF $ **FLOATING
C2998 S.n2703 SUB 0.01fF $ **FLOATING
C2999 S.n2704 SUB 0.02fF $ **FLOATING
C3000 S.n2705 SUB 0.01fF $ **FLOATING
C3001 S.n2706 SUB 0.02fF $ **FLOATING
C3002 S.n2707 SUB 0.05fF $ **FLOATING
C3003 S.n2708 SUB 0.04fF $ **FLOATING
C3004 S.n2709 SUB 0.11fF $ **FLOATING
C3005 S.n2710 SUB 0.38fF $ **FLOATING
C3006 S.n2711 SUB 0.20fF $ **FLOATING
C3007 S.n2712 SUB 8.97fF $ **FLOATING
C3008 S.n2713 SUB 8.97fF $ **FLOATING
C3009 S.n2714 SUB 0.60fF $ **FLOATING
C3010 S.n2715 SUB 0.22fF $ **FLOATING
C3011 S.n2716 SUB 0.59fF $ **FLOATING
C3012 S.n2717 SUB 3.43fF $ **FLOATING
C3013 S.n2718 SUB 0.29fF $ **FLOATING
C3014 S.t10 SUB 21.38fF
C3015 S.n2719 SUB 21.67fF $ **FLOATING
C3016 S.n2720 SUB 0.77fF $ **FLOATING
C3017 S.n2721 SUB 0.28fF $ **FLOATING
C3018 S.n2722 SUB 4.00fF $ **FLOATING
C3019 S.n2723 SUB 1.35fF $ **FLOATING
C3020 S.t1855 SUB 0.02fF
C3021 S.n2724 SUB 0.64fF $ **FLOATING
C3022 S.n2725 SUB 0.61fF $ **FLOATING
C3023 S.n2726 SUB 0.25fF $ **FLOATING
C3024 S.n2727 SUB 0.09fF $ **FLOATING
C3025 S.n2728 SUB 0.21fF $ **FLOATING
C3026 S.n2729 SUB 0.92fF $ **FLOATING
C3027 S.n2730 SUB 0.44fF $ **FLOATING
C3028 S.n2731 SUB 1.88fF $ **FLOATING
C3029 S.n2732 SUB 0.12fF $ **FLOATING
C3030 S.t450 SUB 0.02fF
C3031 S.n2733 SUB 0.14fF $ **FLOATING
C3032 S.t998 SUB 0.02fF
C3033 S.n2735 SUB 0.24fF $ **FLOATING
C3034 S.n2736 SUB 0.36fF $ **FLOATING
C3035 S.n2737 SUB 0.61fF $ **FLOATING
C3036 S.n2738 SUB 0.02fF $ **FLOATING
C3037 S.n2739 SUB 0.01fF $ **FLOATING
C3038 S.n2740 SUB 0.02fF $ **FLOATING
C3039 S.n2741 SUB 0.08fF $ **FLOATING
C3040 S.n2742 SUB 0.06fF $ **FLOATING
C3041 S.n2743 SUB 0.03fF $ **FLOATING
C3042 S.n2744 SUB 0.04fF $ **FLOATING
C3043 S.n2745 SUB 1.00fF $ **FLOATING
C3044 S.n2746 SUB 0.36fF $ **FLOATING
C3045 S.n2747 SUB 1.87fF $ **FLOATING
C3046 S.n2748 SUB 1.99fF $ **FLOATING
C3047 S.t2093 SUB 0.02fF
C3048 S.n2749 SUB 0.24fF $ **FLOATING
C3049 S.n2750 SUB 0.91fF $ **FLOATING
C3050 S.n2751 SUB 0.05fF $ **FLOATING
C3051 S.t640 SUB 0.02fF
C3052 S.n2752 SUB 0.12fF $ **FLOATING
C3053 S.n2753 SUB 0.14fF $ **FLOATING
C3054 S.n2755 SUB 1.89fF $ **FLOATING
C3055 S.n2756 SUB 0.06fF $ **FLOATING
C3056 S.n2757 SUB 0.03fF $ **FLOATING
C3057 S.n2758 SUB 0.04fF $ **FLOATING
C3058 S.n2759 SUB 0.99fF $ **FLOATING
C3059 S.n2760 SUB 0.02fF $ **FLOATING
C3060 S.n2761 SUB 0.01fF $ **FLOATING
C3061 S.n2762 SUB 0.02fF $ **FLOATING
C3062 S.n2763 SUB 0.08fF $ **FLOATING
C3063 S.n2764 SUB 0.36fF $ **FLOATING
C3064 S.n2765 SUB 1.85fF $ **FLOATING
C3065 S.t238 SUB 0.02fF
C3066 S.n2766 SUB 0.24fF $ **FLOATING
C3067 S.n2767 SUB 0.36fF $ **FLOATING
C3068 S.n2768 SUB 0.61fF $ **FLOATING
C3069 S.n2769 SUB 0.12fF $ **FLOATING
C3070 S.t2237 SUB 0.02fF
C3071 S.n2770 SUB 0.14fF $ **FLOATING
C3072 S.n2772 SUB 0.70fF $ **FLOATING
C3073 S.n2773 SUB 0.23fF $ **FLOATING
C3074 S.n2774 SUB 0.23fF $ **FLOATING
C3075 S.n2775 SUB 0.70fF $ **FLOATING
C3076 S.n2776 SUB 1.16fF $ **FLOATING
C3077 S.n2777 SUB 0.22fF $ **FLOATING
C3078 S.n2778 SUB 0.25fF $ **FLOATING
C3079 S.n2779 SUB 0.09fF $ **FLOATING
C3080 S.n2780 SUB 1.88fF $ **FLOATING
C3081 S.t1374 SUB 0.02fF
C3082 S.n2781 SUB 0.24fF $ **FLOATING
C3083 S.n2782 SUB 0.91fF $ **FLOATING
C3084 S.n2783 SUB 0.05fF $ **FLOATING
C3085 S.t2297 SUB 0.02fF
C3086 S.n2784 SUB 0.12fF $ **FLOATING
C3087 S.n2785 SUB 0.14fF $ **FLOATING
C3088 S.n2787 SUB 0.25fF $ **FLOATING
C3089 S.n2788 SUB 0.09fF $ **FLOATING
C3090 S.n2789 SUB 0.21fF $ **FLOATING
C3091 S.n2790 SUB 0.92fF $ **FLOATING
C3092 S.n2791 SUB 0.44fF $ **FLOATING
C3093 S.n2792 SUB 1.88fF $ **FLOATING
C3094 S.n2793 SUB 0.12fF $ **FLOATING
C3095 S.t1378 SUB 0.02fF
C3096 S.n2794 SUB 0.14fF $ **FLOATING
C3097 S.t1905 SUB 0.02fF
C3098 S.n2796 SUB 0.24fF $ **FLOATING
C3099 S.n2797 SUB 0.36fF $ **FLOATING
C3100 S.n2798 SUB 0.61fF $ **FLOATING
C3101 S.n2799 SUB 0.02fF $ **FLOATING
C3102 S.n2800 SUB 0.01fF $ **FLOATING
C3103 S.n2801 SUB 0.02fF $ **FLOATING
C3104 S.n2802 SUB 0.08fF $ **FLOATING
C3105 S.n2803 SUB 0.06fF $ **FLOATING
C3106 S.n2804 SUB 0.03fF $ **FLOATING
C3107 S.n2805 SUB 0.04fF $ **FLOATING
C3108 S.n2806 SUB 1.00fF $ **FLOATING
C3109 S.n2807 SUB 0.36fF $ **FLOATING
C3110 S.n2808 SUB 1.87fF $ **FLOATING
C3111 S.n2809 SUB 1.99fF $ **FLOATING
C3112 S.t501 SUB 0.02fF
C3113 S.n2810 SUB 0.24fF $ **FLOATING
C3114 S.n2811 SUB 0.91fF $ **FLOATING
C3115 S.n2812 SUB 0.05fF $ **FLOATING
C3116 S.t1441 SUB 0.02fF
C3117 S.n2813 SUB 0.12fF $ **FLOATING
C3118 S.n2814 SUB 0.14fF $ **FLOATING
C3119 S.n2816 SUB 1.89fF $ **FLOATING
C3120 S.n2817 SUB 0.06fF $ **FLOATING
C3121 S.n2818 SUB 0.03fF $ **FLOATING
C3122 S.n2819 SUB 0.04fF $ **FLOATING
C3123 S.n2820 SUB 0.99fF $ **FLOATING
C3124 S.n2821 SUB 0.02fF $ **FLOATING
C3125 S.n2822 SUB 0.01fF $ **FLOATING
C3126 S.n2823 SUB 0.02fF $ **FLOATING
C3127 S.n2824 SUB 0.08fF $ **FLOATING
C3128 S.n2825 SUB 0.36fF $ **FLOATING
C3129 S.n2826 SUB 1.85fF $ **FLOATING
C3130 S.t1046 SUB 0.02fF
C3131 S.n2827 SUB 0.24fF $ **FLOATING
C3132 S.n2828 SUB 0.36fF $ **FLOATING
C3133 S.n2829 SUB 0.61fF $ **FLOATING
C3134 S.n2830 SUB 0.12fF $ **FLOATING
C3135 S.t504 SUB 0.02fF
C3136 S.n2831 SUB 0.14fF $ **FLOATING
C3137 S.n2833 SUB 0.70fF $ **FLOATING
C3138 S.n2834 SUB 0.23fF $ **FLOATING
C3139 S.n2835 SUB 0.23fF $ **FLOATING
C3140 S.n2836 SUB 0.70fF $ **FLOATING
C3141 S.n2837 SUB 1.16fF $ **FLOATING
C3142 S.n2838 SUB 0.22fF $ **FLOATING
C3143 S.n2839 SUB 0.25fF $ **FLOATING
C3144 S.n2840 SUB 0.09fF $ **FLOATING
C3145 S.n2841 SUB 1.88fF $ **FLOATING
C3146 S.t2146 SUB 0.02fF
C3147 S.n2842 SUB 0.24fF $ **FLOATING
C3148 S.n2843 SUB 0.91fF $ **FLOATING
C3149 S.n2844 SUB 0.05fF $ **FLOATING
C3150 S.t577 SUB 0.02fF
C3151 S.n2845 SUB 0.12fF $ **FLOATING
C3152 S.n2846 SUB 0.14fF $ **FLOATING
C3153 S.n2848 SUB 0.25fF $ **FLOATING
C3154 S.n2849 SUB 0.09fF $ **FLOATING
C3155 S.n2850 SUB 0.21fF $ **FLOATING
C3156 S.n2851 SUB 0.92fF $ **FLOATING
C3157 S.n2852 SUB 0.44fF $ **FLOATING
C3158 S.n2853 SUB 1.88fF $ **FLOATING
C3159 S.n2854 SUB 0.12fF $ **FLOATING
C3160 S.t2147 SUB 0.02fF
C3161 S.n2855 SUB 0.14fF $ **FLOATING
C3162 S.t155 SUB 0.02fF
C3163 S.n2857 SUB 0.24fF $ **FLOATING
C3164 S.n2858 SUB 0.36fF $ **FLOATING
C3165 S.n2859 SUB 0.61fF $ **FLOATING
C3166 S.n2860 SUB 0.02fF $ **FLOATING
C3167 S.n2861 SUB 0.01fF $ **FLOATING
C3168 S.n2862 SUB 0.02fF $ **FLOATING
C3169 S.n2863 SUB 0.08fF $ **FLOATING
C3170 S.n2864 SUB 0.06fF $ **FLOATING
C3171 S.n2865 SUB 0.03fF $ **FLOATING
C3172 S.n2866 SUB 0.04fF $ **FLOATING
C3173 S.n2867 SUB 1.00fF $ **FLOATING
C3174 S.n2868 SUB 0.36fF $ **FLOATING
C3175 S.n2869 SUB 1.87fF $ **FLOATING
C3176 S.n2870 SUB 1.99fF $ **FLOATING
C3177 S.t1283 SUB 0.02fF
C3178 S.n2871 SUB 0.24fF $ **FLOATING
C3179 S.n2872 SUB 0.91fF $ **FLOATING
C3180 S.n2873 SUB 0.05fF $ **FLOATING
C3181 S.t2222 SUB 0.02fF
C3182 S.n2874 SUB 0.12fF $ **FLOATING
C3183 S.n2875 SUB 0.14fF $ **FLOATING
C3184 S.n2877 SUB 1.89fF $ **FLOATING
C3185 S.n2878 SUB 0.06fF $ **FLOATING
C3186 S.n2879 SUB 0.03fF $ **FLOATING
C3187 S.n2880 SUB 0.04fF $ **FLOATING
C3188 S.n2881 SUB 0.99fF $ **FLOATING
C3189 S.n2882 SUB 0.02fF $ **FLOATING
C3190 S.n2883 SUB 0.01fF $ **FLOATING
C3191 S.n2884 SUB 0.02fF $ **FLOATING
C3192 S.n2885 SUB 0.08fF $ **FLOATING
C3193 S.n2886 SUB 0.36fF $ **FLOATING
C3194 S.n2887 SUB 1.85fF $ **FLOATING
C3195 S.t1819 SUB 0.02fF
C3196 S.n2888 SUB 0.24fF $ **FLOATING
C3197 S.n2889 SUB 0.36fF $ **FLOATING
C3198 S.n2890 SUB 0.61fF $ **FLOATING
C3199 S.n2891 SUB 0.12fF $ **FLOATING
C3200 S.t1287 SUB 0.02fF
C3201 S.n2892 SUB 0.14fF $ **FLOATING
C3202 S.n2894 SUB 0.70fF $ **FLOATING
C3203 S.n2895 SUB 0.23fF $ **FLOATING
C3204 S.n2896 SUB 0.23fF $ **FLOATING
C3205 S.n2897 SUB 0.70fF $ **FLOATING
C3206 S.n2898 SUB 1.16fF $ **FLOATING
C3207 S.n2899 SUB 0.22fF $ **FLOATING
C3208 S.n2900 SUB 0.25fF $ **FLOATING
C3209 S.n2901 SUB 0.09fF $ **FLOATING
C3210 S.n2902 SUB 1.88fF $ **FLOATING
C3211 S.t396 SUB 0.02fF
C3212 S.n2903 SUB 0.24fF $ **FLOATING
C3213 S.n2904 SUB 0.91fF $ **FLOATING
C3214 S.n2905 SUB 0.05fF $ **FLOATING
C3215 S.t1363 SUB 0.02fF
C3216 S.n2906 SUB 0.12fF $ **FLOATING
C3217 S.n2907 SUB 0.14fF $ **FLOATING
C3218 S.n2909 SUB 0.25fF $ **FLOATING
C3219 S.n2910 SUB 0.09fF $ **FLOATING
C3220 S.n2911 SUB 0.21fF $ **FLOATING
C3221 S.n2912 SUB 0.92fF $ **FLOATING
C3222 S.n2913 SUB 0.44fF $ **FLOATING
C3223 S.n2914 SUB 1.88fF $ **FLOATING
C3224 S.n2915 SUB 0.12fF $ **FLOATING
C3225 S.t400 SUB 0.02fF
C3226 S.n2916 SUB 0.14fF $ **FLOATING
C3227 S.t955 SUB 0.02fF
C3228 S.n2918 SUB 0.24fF $ **FLOATING
C3229 S.n2919 SUB 0.36fF $ **FLOATING
C3230 S.n2920 SUB 0.61fF $ **FLOATING
C3231 S.n2921 SUB 0.02fF $ **FLOATING
C3232 S.n2922 SUB 0.01fF $ **FLOATING
C3233 S.n2923 SUB 0.02fF $ **FLOATING
C3234 S.n2924 SUB 0.08fF $ **FLOATING
C3235 S.n2925 SUB 0.06fF $ **FLOATING
C3236 S.n2926 SUB 0.03fF $ **FLOATING
C3237 S.n2927 SUB 0.04fF $ **FLOATING
C3238 S.n2928 SUB 1.00fF $ **FLOATING
C3239 S.n2929 SUB 0.36fF $ **FLOATING
C3240 S.n2930 SUB 1.87fF $ **FLOATING
C3241 S.n2931 SUB 1.99fF $ **FLOATING
C3242 S.t2048 SUB 0.02fF
C3243 S.n2932 SUB 0.24fF $ **FLOATING
C3244 S.n2933 SUB 0.91fF $ **FLOATING
C3245 S.n2934 SUB 0.05fF $ **FLOATING
C3246 S.t612 SUB 0.02fF
C3247 S.n2935 SUB 0.12fF $ **FLOATING
C3248 S.n2936 SUB 0.14fF $ **FLOATING
C3249 S.n2938 SUB 1.89fF $ **FLOATING
C3250 S.n2939 SUB 0.06fF $ **FLOATING
C3251 S.n2940 SUB 0.03fF $ **FLOATING
C3252 S.n2941 SUB 0.04fF $ **FLOATING
C3253 S.n2942 SUB 0.99fF $ **FLOATING
C3254 S.n2943 SUB 0.02fF $ **FLOATING
C3255 S.n2944 SUB 0.01fF $ **FLOATING
C3256 S.n2945 SUB 0.02fF $ **FLOATING
C3257 S.n2946 SUB 0.08fF $ **FLOATING
C3258 S.n2947 SUB 0.36fF $ **FLOATING
C3259 S.n2948 SUB 1.85fF $ **FLOATING
C3260 S.t163 SUB 0.02fF
C3261 S.n2949 SUB 0.24fF $ **FLOATING
C3262 S.n2950 SUB 0.36fF $ **FLOATING
C3263 S.n2951 SUB 0.61fF $ **FLOATING
C3264 S.n2952 SUB 0.12fF $ **FLOATING
C3265 S.t2143 SUB 0.02fF
C3266 S.n2953 SUB 0.14fF $ **FLOATING
C3267 S.n2955 SUB 0.70fF $ **FLOATING
C3268 S.n2956 SUB 0.23fF $ **FLOATING
C3269 S.n2957 SUB 0.23fF $ **FLOATING
C3270 S.n2958 SUB 0.70fF $ **FLOATING
C3271 S.n2959 SUB 1.16fF $ **FLOATING
C3272 S.n2960 SUB 0.22fF $ **FLOATING
C3273 S.n2961 SUB 0.25fF $ **FLOATING
C3274 S.n2962 SUB 0.09fF $ **FLOATING
C3275 S.n2963 SUB 1.88fF $ **FLOATING
C3276 S.t1722 SUB 0.02fF
C3277 S.n2964 SUB 0.24fF $ **FLOATING
C3278 S.n2965 SUB 0.91fF $ **FLOATING
C3279 S.n2966 SUB 0.05fF $ **FLOATING
C3280 S.t2327 SUB 0.02fF
C3281 S.n2967 SUB 0.12fF $ **FLOATING
C3282 S.n2968 SUB 0.14fF $ **FLOATING
C3283 S.n2970 SUB 0.25fF $ **FLOATING
C3284 S.n2971 SUB 0.09fF $ **FLOATING
C3285 S.n2972 SUB 0.21fF $ **FLOATING
C3286 S.n2973 SUB 0.92fF $ **FLOATING
C3287 S.n2974 SUB 0.44fF $ **FLOATING
C3288 S.n2975 SUB 1.88fF $ **FLOATING
C3289 S.n2976 SUB 0.12fF $ **FLOATING
C3290 S.t1279 SUB 0.02fF
C3291 S.n2977 SUB 0.14fF $ **FLOATING
C3292 S.t1826 SUB 0.02fF
C3293 S.n2979 SUB 0.24fF $ **FLOATING
C3294 S.n2980 SUB 0.36fF $ **FLOATING
C3295 S.n2981 SUB 0.61fF $ **FLOATING
C3296 S.n2982 SUB 0.02fF $ **FLOATING
C3297 S.n2983 SUB 0.01fF $ **FLOATING
C3298 S.n2984 SUB 0.02fF $ **FLOATING
C3299 S.n2985 SUB 0.08fF $ **FLOATING
C3300 S.n2986 SUB 0.06fF $ **FLOATING
C3301 S.n2987 SUB 0.03fF $ **FLOATING
C3302 S.n2988 SUB 0.04fF $ **FLOATING
C3303 S.n2989 SUB 1.00fF $ **FLOATING
C3304 S.n2990 SUB 0.36fF $ **FLOATING
C3305 S.n2991 SUB 1.87fF $ **FLOATING
C3306 S.n2992 SUB 1.99fF $ **FLOATING
C3307 S.t850 SUB 0.02fF
C3308 S.n2993 SUB 0.24fF $ **FLOATING
C3309 S.n2994 SUB 0.91fF $ **FLOATING
C3310 S.n2995 SUB 0.05fF $ **FLOATING
C3311 S.t1468 SUB 0.02fF
C3312 S.n2996 SUB 0.12fF $ **FLOATING
C3313 S.n2997 SUB 0.14fF $ **FLOATING
C3314 S.n2999 SUB 1.89fF $ **FLOATING
C3315 S.n3000 SUB 0.04fF $ **FLOATING
C3316 S.n3001 SUB 0.07fF $ **FLOATING
C3317 S.n3002 SUB 0.05fF $ **FLOATING
C3318 S.n3003 SUB 0.87fF $ **FLOATING
C3319 S.n3004 SUB 0.01fF $ **FLOATING
C3320 S.n3005 SUB 0.01fF $ **FLOATING
C3321 S.n3006 SUB 0.01fF $ **FLOATING
C3322 S.n3007 SUB 0.07fF $ **FLOATING
C3323 S.n3008 SUB 0.68fF $ **FLOATING
C3324 S.n3009 SUB 0.72fF $ **FLOATING
C3325 S.t958 SUB 0.02fF
C3326 S.n3010 SUB 0.24fF $ **FLOATING
C3327 S.n3011 SUB 0.36fF $ **FLOATING
C3328 S.n3012 SUB 0.61fF $ **FLOATING
C3329 S.n3013 SUB 0.12fF $ **FLOATING
C3330 S.t393 SUB 0.02fF
C3331 S.n3014 SUB 0.14fF $ **FLOATING
C3332 S.n3016 SUB 0.70fF $ **FLOATING
C3333 S.n3017 SUB 0.23fF $ **FLOATING
C3334 S.n3018 SUB 0.23fF $ **FLOATING
C3335 S.n3019 SUB 0.70fF $ **FLOATING
C3336 S.n3020 SUB 1.16fF $ **FLOATING
C3337 S.n3021 SUB 0.22fF $ **FLOATING
C3338 S.n3022 SUB 0.25fF $ **FLOATING
C3339 S.n3023 SUB 0.09fF $ **FLOATING
C3340 S.n3024 SUB 2.31fF $ **FLOATING
C3341 S.t2494 SUB 0.02fF
C3342 S.n3025 SUB 0.24fF $ **FLOATING
C3343 S.n3026 SUB 0.91fF $ **FLOATING
C3344 S.n3027 SUB 0.05fF $ **FLOATING
C3345 S.t608 SUB 0.02fF
C3346 S.n3028 SUB 0.12fF $ **FLOATING
C3347 S.n3029 SUB 0.14fF $ **FLOATING
C3348 S.n3031 SUB 1.88fF $ **FLOATING
C3349 S.n3032 SUB 0.46fF $ **FLOATING
C3350 S.n3033 SUB 0.22fF $ **FLOATING
C3351 S.n3034 SUB 0.38fF $ **FLOATING
C3352 S.n3035 SUB 0.16fF $ **FLOATING
C3353 S.n3036 SUB 0.28fF $ **FLOATING
C3354 S.n3037 SUB 0.21fF $ **FLOATING
C3355 S.n3038 SUB 0.30fF $ **FLOATING
C3356 S.n3039 SUB 0.42fF $ **FLOATING
C3357 S.n3040 SUB 0.21fF $ **FLOATING
C3358 S.t11 SUB 0.02fF
C3359 S.n3041 SUB 0.24fF $ **FLOATING
C3360 S.n3042 SUB 0.36fF $ **FLOATING
C3361 S.n3043 SUB 0.61fF $ **FLOATING
C3362 S.n3044 SUB 0.12fF $ **FLOATING
C3363 S.t2045 SUB 0.02fF
C3364 S.n3045 SUB 0.14fF $ **FLOATING
C3365 S.n3047 SUB 0.04fF $ **FLOATING
C3366 S.n3048 SUB 0.03fF $ **FLOATING
C3367 S.n3049 SUB 0.03fF $ **FLOATING
C3368 S.n3050 SUB 0.10fF $ **FLOATING
C3369 S.n3051 SUB 0.36fF $ **FLOATING
C3370 S.n3052 SUB 0.38fF $ **FLOATING
C3371 S.n3053 SUB 0.11fF $ **FLOATING
C3372 S.n3054 SUB 0.12fF $ **FLOATING
C3373 S.n3055 SUB 0.07fF $ **FLOATING
C3374 S.n3056 SUB 0.12fF $ **FLOATING
C3375 S.n3057 SUB 0.18fF $ **FLOATING
C3376 S.n3058 SUB 4.00fF $ **FLOATING
C3377 S.t1618 SUB 0.02fF
C3378 S.n3059 SUB 0.24fF $ **FLOATING
C3379 S.n3060 SUB 0.91fF $ **FLOATING
C3380 S.n3061 SUB 0.05fF $ **FLOATING
C3381 S.t2261 SUB 0.02fF
C3382 S.n3062 SUB 0.12fF $ **FLOATING
C3383 S.n3063 SUB 0.14fF $ **FLOATING
C3384 S.n3065 SUB 0.25fF $ **FLOATING
C3385 S.n3066 SUB 0.09fF $ **FLOATING
C3386 S.n3067 SUB 0.21fF $ **FLOATING
C3387 S.n3068 SUB 1.28fF $ **FLOATING
C3388 S.n3069 SUB 0.53fF $ **FLOATING
C3389 S.n3070 SUB 1.88fF $ **FLOATING
C3390 S.n3071 SUB 0.12fF $ **FLOATING
C3391 S.t1333 SUB 0.02fF
C3392 S.n3072 SUB 0.14fF $ **FLOATING
C3393 S.t1876 SUB 0.02fF
C3394 S.n3074 SUB 0.24fF $ **FLOATING
C3395 S.n3075 SUB 0.36fF $ **FLOATING
C3396 S.n3076 SUB 0.61fF $ **FLOATING
C3397 S.n3077 SUB 1.58fF $ **FLOATING
C3398 S.n3078 SUB 2.45fF $ **FLOATING
C3399 S.t909 SUB 0.02fF
C3400 S.n3079 SUB 0.24fF $ **FLOATING
C3401 S.n3080 SUB 0.91fF $ **FLOATING
C3402 S.n3081 SUB 0.05fF $ **FLOATING
C3403 S.t1404 SUB 0.02fF
C3404 S.n3082 SUB 0.12fF $ **FLOATING
C3405 S.n3083 SUB 0.14fF $ **FLOATING
C3406 S.n3085 SUB 1.89fF $ **FLOATING
C3407 S.n3086 SUB 0.06fF $ **FLOATING
C3408 S.n3087 SUB 0.03fF $ **FLOATING
C3409 S.n3088 SUB 0.04fF $ **FLOATING
C3410 S.n3089 SUB 0.99fF $ **FLOATING
C3411 S.n3090 SUB 0.02fF $ **FLOATING
C3412 S.n3091 SUB 0.01fF $ **FLOATING
C3413 S.n3092 SUB 0.02fF $ **FLOATING
C3414 S.n3093 SUB 0.08fF $ **FLOATING
C3415 S.n3094 SUB 0.36fF $ **FLOATING
C3416 S.n3095 SUB 1.85fF $ **FLOATING
C3417 S.t1010 SUB 0.02fF
C3418 S.n3096 SUB 0.24fF $ **FLOATING
C3419 S.n3097 SUB 0.36fF $ **FLOATING
C3420 S.n3098 SUB 0.61fF $ **FLOATING
C3421 S.n3099 SUB 0.12fF $ **FLOATING
C3422 S.t453 SUB 0.02fF
C3423 S.n3100 SUB 0.14fF $ **FLOATING
C3424 S.n3102 SUB 0.70fF $ **FLOATING
C3425 S.n3103 SUB 0.23fF $ **FLOATING
C3426 S.n3104 SUB 0.23fF $ **FLOATING
C3427 S.n3105 SUB 0.70fF $ **FLOATING
C3428 S.n3106 SUB 1.16fF $ **FLOATING
C3429 S.n3107 SUB 0.22fF $ **FLOATING
C3430 S.n3108 SUB 0.25fF $ **FLOATING
C3431 S.n3109 SUB 0.09fF $ **FLOATING
C3432 S.n3110 SUB 1.88fF $ **FLOATING
C3433 S.t2550 SUB 0.02fF
C3434 S.n3111 SUB 0.24fF $ **FLOATING
C3435 S.n3112 SUB 0.91fF $ **FLOATING
C3436 S.n3113 SUB 0.05fF $ **FLOATING
C3437 S.t534 SUB 0.02fF
C3438 S.n3114 SUB 0.12fF $ **FLOATING
C3439 S.n3115 SUB 0.14fF $ **FLOATING
C3440 S.n3117 SUB 20.78fF $ **FLOATING
C3441 S.n3118 SUB 1.72fF $ **FLOATING
C3442 S.n3119 SUB 3.05fF $ **FLOATING
C3443 S.t1867 SUB 0.02fF
C3444 S.n3120 SUB 0.24fF $ **FLOATING
C3445 S.n3121 SUB 0.36fF $ **FLOATING
C3446 S.n3122 SUB 0.61fF $ **FLOATING
C3447 S.n3123 SUB 0.12fF $ **FLOATING
C3448 S.t1330 SUB 0.02fF
C3449 S.n3124 SUB 0.14fF $ **FLOATING
C3450 S.n3126 SUB 0.31fF $ **FLOATING
C3451 S.n3127 SUB 0.23fF $ **FLOATING
C3452 S.n3128 SUB 0.66fF $ **FLOATING
C3453 S.n3129 SUB 0.95fF $ **FLOATING
C3454 S.n3130 SUB 0.23fF $ **FLOATING
C3455 S.n3131 SUB 0.21fF $ **FLOATING
C3456 S.n3132 SUB 0.20fF $ **FLOATING
C3457 S.n3133 SUB 0.06fF $ **FLOATING
C3458 S.n3134 SUB 0.09fF $ **FLOATING
C3459 S.n3135 SUB 0.10fF $ **FLOATING
C3460 S.n3136 SUB 1.99fF $ **FLOATING
C3461 S.t1501 SUB 0.02fF
C3462 S.n3137 SUB 0.12fF $ **FLOATING
C3463 S.n3138 SUB 0.14fF $ **FLOATING
C3464 S.t448 SUB 0.02fF
C3465 S.n3140 SUB 0.24fF $ **FLOATING
C3466 S.n3141 SUB 0.91fF $ **FLOATING
C3467 S.n3142 SUB 0.05fF $ **FLOATING
C3468 S.n3143 SUB 1.88fF $ **FLOATING
C3469 S.n3144 SUB 0.12fF $ **FLOATING
C3470 S.t2277 SUB 0.02fF
C3471 S.n3145 SUB 0.14fF $ **FLOATING
C3472 S.t566 SUB 0.02fF
C3473 S.n3147 SUB 0.12fF $ **FLOATING
C3474 S.n3148 SUB 0.14fF $ **FLOATING
C3475 S.t770 SUB 0.02fF
C3476 S.n3150 SUB 0.24fF $ **FLOATING
C3477 S.n3151 SUB 0.91fF $ **FLOATING
C3478 S.n3152 SUB 0.05fF $ **FLOATING
C3479 S.t1511 SUB 0.02fF
C3480 S.n3153 SUB 0.24fF $ **FLOATING
C3481 S.n3154 SUB 0.36fF $ **FLOATING
C3482 S.n3155 SUB 0.61fF $ **FLOATING
C3483 S.n3156 SUB 0.32fF $ **FLOATING
C3484 S.n3157 SUB 1.09fF $ **FLOATING
C3485 S.n3158 SUB 0.15fF $ **FLOATING
C3486 S.n3159 SUB 2.10fF $ **FLOATING
C3487 S.n3160 SUB 2.94fF $ **FLOATING
C3488 S.n3161 SUB 1.88fF $ **FLOATING
C3489 S.n3162 SUB 0.12fF $ **FLOATING
C3490 S.t2098 SUB 0.02fF
C3491 S.n3163 SUB 0.14fF $ **FLOATING
C3492 S.t108 SUB 0.02fF
C3493 S.n3165 SUB 0.24fF $ **FLOATING
C3494 S.n3166 SUB 0.36fF $ **FLOATING
C3495 S.n3167 SUB 0.61fF $ **FLOATING
C3496 S.n3168 SUB 0.92fF $ **FLOATING
C3497 S.n3169 SUB 0.32fF $ **FLOATING
C3498 S.n3170 SUB 0.92fF $ **FLOATING
C3499 S.n3171 SUB 1.09fF $ **FLOATING
C3500 S.n3172 SUB 0.15fF $ **FLOATING
C3501 S.n3173 SUB 4.96fF $ **FLOATING
C3502 S.t2177 SUB 0.02fF
C3503 S.n3174 SUB 0.12fF $ **FLOATING
C3504 S.n3175 SUB 0.14fF $ **FLOATING
C3505 S.t1680 SUB 0.02fF
C3506 S.n3177 SUB 0.24fF $ **FLOATING
C3507 S.n3178 SUB 0.91fF $ **FLOATING
C3508 S.n3179 SUB 0.05fF $ **FLOATING
C3509 S.n3180 SUB 1.88fF $ **FLOATING
C3510 S.n3181 SUB 2.67fF $ **FLOATING
C3511 S.t1781 SUB 0.02fF
C3512 S.n3182 SUB 0.24fF $ **FLOATING
C3513 S.n3183 SUB 0.36fF $ **FLOATING
C3514 S.n3184 SUB 0.61fF $ **FLOATING
C3515 S.n3185 SUB 0.12fF $ **FLOATING
C3516 S.t1234 SUB 0.02fF
C3517 S.n3186 SUB 0.14fF $ **FLOATING
C3518 S.n3188 SUB 1.88fF $ **FLOATING
C3519 S.n3189 SUB 2.67fF $ **FLOATING
C3520 S.t654 SUB 0.02fF
C3521 S.n3190 SUB 0.24fF $ **FLOATING
C3522 S.n3191 SUB 0.36fF $ **FLOATING
C3523 S.n3192 SUB 0.61fF $ **FLOATING
C3524 S.t978 SUB 0.02fF
C3525 S.n3193 SUB 1.22fF $ **FLOATING
C3526 S.n3194 SUB 0.61fF $ **FLOATING
C3527 S.n3195 SUB 0.35fF $ **FLOATING
C3528 S.n3196 SUB 0.63fF $ **FLOATING
C3529 S.n3197 SUB 1.15fF $ **FLOATING
C3530 S.n3198 SUB 3.03fF $ **FLOATING
C3531 S.n3199 SUB 0.59fF $ **FLOATING
C3532 S.n3200 SUB 0.02fF $ **FLOATING
C3533 S.n3201 SUB 0.97fF $ **FLOATING
C3534 S.t46 SUB 21.38fF
C3535 S.n3202 SUB 20.25fF $ **FLOATING
C3536 S.n3204 SUB 0.38fF $ **FLOATING
C3537 S.n3205 SUB 0.23fF $ **FLOATING
C3538 S.n3206 SUB 2.90fF $ **FLOATING
C3539 S.n3207 SUB 2.46fF $ **FLOATING
C3540 S.n3208 SUB 1.96fF $ **FLOATING
C3541 S.n3209 SUB 3.94fF $ **FLOATING
C3542 S.n3210 SUB 0.25fF $ **FLOATING
C3543 S.n3211 SUB 0.01fF $ **FLOATING
C3544 S.t669 SUB 0.02fF
C3545 S.n3212 SUB 0.25fF $ **FLOATING
C3546 S.t112 SUB 0.02fF
C3547 S.n3213 SUB 0.95fF $ **FLOATING
C3548 S.n3214 SUB 0.70fF $ **FLOATING
C3549 S.n3215 SUB 0.78fF $ **FLOATING
C3550 S.n3216 SUB 1.93fF $ **FLOATING
C3551 S.n3217 SUB 1.88fF $ **FLOATING
C3552 S.n3218 SUB 0.12fF $ **FLOATING
C3553 S.t2323 SUB 0.02fF
C3554 S.n3219 SUB 0.14fF $ **FLOATING
C3555 S.t47 SUB 0.02fF
C3556 S.n3221 SUB 0.24fF $ **FLOATING
C3557 S.n3222 SUB 0.36fF $ **FLOATING
C3558 S.n3223 SUB 0.61fF $ **FLOATING
C3559 S.n3224 SUB 1.52fF $ **FLOATING
C3560 S.n3225 SUB 2.99fF $ **FLOATING
C3561 S.t1784 SUB 0.02fF
C3562 S.n3226 SUB 0.24fF $ **FLOATING
C3563 S.n3227 SUB 0.91fF $ **FLOATING
C3564 S.n3228 SUB 0.05fF $ **FLOATING
C3565 S.t493 SUB 0.02fF
C3566 S.n3229 SUB 0.12fF $ **FLOATING
C3567 S.n3230 SUB 0.14fF $ **FLOATING
C3568 S.n3232 SUB 1.89fF $ **FLOATING
C3569 S.n3233 SUB 1.88fF $ **FLOATING
C3570 S.t1739 SUB 0.02fF
C3571 S.n3234 SUB 0.24fF $ **FLOATING
C3572 S.n3235 SUB 0.36fF $ **FLOATING
C3573 S.n3236 SUB 0.61fF $ **FLOATING
C3574 S.n3237 SUB 0.12fF $ **FLOATING
C3575 S.t1465 SUB 0.02fF
C3576 S.n3238 SUB 0.14fF $ **FLOATING
C3577 S.n3240 SUB 1.16fF $ **FLOATING
C3578 S.n3241 SUB 0.22fF $ **FLOATING
C3579 S.n3242 SUB 0.25fF $ **FLOATING
C3580 S.n3243 SUB 0.09fF $ **FLOATING
C3581 S.n3244 SUB 1.88fF $ **FLOATING
C3582 S.t912 SUB 0.02fF
C3583 S.n3245 SUB 0.24fF $ **FLOATING
C3584 S.n3246 SUB 0.91fF $ **FLOATING
C3585 S.n3247 SUB 0.05fF $ **FLOATING
C3586 S.t2138 SUB 0.02fF
C3587 S.n3248 SUB 0.12fF $ **FLOATING
C3588 S.n3249 SUB 0.14fF $ **FLOATING
C3589 S.n3251 SUB 0.78fF $ **FLOATING
C3590 S.n3252 SUB 1.94fF $ **FLOATING
C3591 S.n3253 SUB 1.88fF $ **FLOATING
C3592 S.n3254 SUB 0.12fF $ **FLOATING
C3593 S.t606 SUB 0.02fF
C3594 S.n3255 SUB 0.14fF $ **FLOATING
C3595 S.t864 SUB 0.02fF
C3596 S.n3257 SUB 0.24fF $ **FLOATING
C3597 S.n3258 SUB 0.36fF $ **FLOATING
C3598 S.n3259 SUB 0.61fF $ **FLOATING
C3599 S.n3260 SUB 1.84fF $ **FLOATING
C3600 S.n3261 SUB 2.99fF $ **FLOATING
C3601 S.t2553 SUB 0.02fF
C3602 S.n3262 SUB 0.24fF $ **FLOATING
C3603 S.n3263 SUB 0.91fF $ **FLOATING
C3604 S.n3264 SUB 0.05fF $ **FLOATING
C3605 S.t1411 SUB 0.02fF
C3606 S.n3265 SUB 0.12fF $ **FLOATING
C3607 S.n3266 SUB 0.14fF $ **FLOATING
C3608 S.n3268 SUB 1.89fF $ **FLOATING
C3609 S.n3269 SUB 1.88fF $ **FLOATING
C3610 S.t2508 SUB 0.02fF
C3611 S.n3270 SUB 0.24fF $ **FLOATING
C3612 S.n3271 SUB 0.36fF $ **FLOATING
C3613 S.n3272 SUB 0.61fF $ **FLOATING
C3614 S.n3273 SUB 0.12fF $ **FLOATING
C3615 S.t2258 SUB 0.02fF
C3616 S.n3274 SUB 0.14fF $ **FLOATING
C3617 S.n3276 SUB 1.16fF $ **FLOATING
C3618 S.n3277 SUB 0.22fF $ **FLOATING
C3619 S.n3278 SUB 0.25fF $ **FLOATING
C3620 S.n3279 SUB 0.09fF $ **FLOATING
C3621 S.n3280 SUB 1.88fF $ **FLOATING
C3622 S.t1682 SUB 0.02fF
C3623 S.n3281 SUB 0.24fF $ **FLOATING
C3624 S.n3282 SUB 0.91fF $ **FLOATING
C3625 S.n3283 SUB 0.05fF $ **FLOATING
C3626 S.t546 SUB 0.02fF
C3627 S.n3284 SUB 0.12fF $ **FLOATING
C3628 S.n3285 SUB 0.14fF $ **FLOATING
C3629 S.n3287 SUB 0.78fF $ **FLOATING
C3630 S.n3288 SUB 1.94fF $ **FLOATING
C3631 S.n3289 SUB 1.88fF $ **FLOATING
C3632 S.n3290 SUB 0.12fF $ **FLOATING
C3633 S.t1397 SUB 0.02fF
C3634 S.n3291 SUB 0.14fF $ **FLOATING
C3635 S.t1636 SUB 0.02fF
C3636 S.n3293 SUB 0.24fF $ **FLOATING
C3637 S.n3294 SUB 0.36fF $ **FLOATING
C3638 S.n3295 SUB 0.61fF $ **FLOATING
C3639 S.n3296 SUB 1.84fF $ **FLOATING
C3640 S.n3297 SUB 2.99fF $ **FLOATING
C3641 S.t807 SUB 0.02fF
C3642 S.n3298 SUB 0.24fF $ **FLOATING
C3643 S.n3299 SUB 0.91fF $ **FLOATING
C3644 S.n3300 SUB 0.05fF $ **FLOATING
C3645 S.t2188 SUB 0.02fF
C3646 S.n3301 SUB 0.12fF $ **FLOATING
C3647 S.n3302 SUB 0.14fF $ **FLOATING
C3648 S.n3304 SUB 1.89fF $ **FLOATING
C3649 S.n3305 SUB 1.88fF $ **FLOATING
C3650 S.t768 SUB 0.02fF
C3651 S.n3306 SUB 0.24fF $ **FLOATING
C3652 S.n3307 SUB 0.36fF $ **FLOATING
C3653 S.n3308 SUB 0.61fF $ **FLOATING
C3654 S.n3309 SUB 0.12fF $ **FLOATING
C3655 S.t526 SUB 0.02fF
C3656 S.n3310 SUB 0.14fF $ **FLOATING
C3657 S.n3312 SUB 1.16fF $ **FLOATING
C3658 S.n3313 SUB 0.22fF $ **FLOATING
C3659 S.n3314 SUB 0.25fF $ **FLOATING
C3660 S.n3315 SUB 0.09fF $ **FLOATING
C3661 S.n3316 SUB 1.88fF $ **FLOATING
C3662 S.t2456 SUB 0.02fF
C3663 S.n3317 SUB 0.24fF $ **FLOATING
C3664 S.n3318 SUB 0.91fF $ **FLOATING
C3665 S.n3319 SUB 0.05fF $ **FLOATING
C3666 S.t1326 SUB 0.02fF
C3667 S.n3320 SUB 0.12fF $ **FLOATING
C3668 S.n3321 SUB 0.14fF $ **FLOATING
C3669 S.n3323 SUB 0.78fF $ **FLOATING
C3670 S.n3324 SUB 1.94fF $ **FLOATING
C3671 S.n3325 SUB 1.88fF $ **FLOATING
C3672 S.n3326 SUB 0.12fF $ **FLOATING
C3673 S.t2291 SUB 0.02fF
C3674 S.n3327 SUB 0.14fF $ **FLOATING
C3675 S.t2417 SUB 0.02fF
C3676 S.n3329 SUB 0.24fF $ **FLOATING
C3677 S.n3330 SUB 0.36fF $ **FLOATING
C3678 S.n3331 SUB 0.61fF $ **FLOATING
C3679 S.n3332 SUB 1.84fF $ **FLOATING
C3680 S.n3333 SUB 2.99fF $ **FLOATING
C3681 S.t1587 SUB 0.02fF
C3682 S.n3334 SUB 0.24fF $ **FLOATING
C3683 S.n3335 SUB 0.91fF $ **FLOATING
C3684 S.n3336 SUB 0.05fF $ **FLOATING
C3685 S.t445 SUB 0.02fF
C3686 S.n3337 SUB 0.12fF $ **FLOATING
C3687 S.n3338 SUB 0.14fF $ **FLOATING
C3688 S.n3340 SUB 1.89fF $ **FLOATING
C3689 S.n3341 SUB 1.88fF $ **FLOATING
C3690 S.t1672 SUB 0.02fF
C3691 S.n3342 SUB 0.24fF $ **FLOATING
C3692 S.n3343 SUB 0.36fF $ **FLOATING
C3693 S.n3344 SUB 0.61fF $ **FLOATING
C3694 S.n3345 SUB 0.12fF $ **FLOATING
C3695 S.t2403 SUB 0.02fF
C3696 S.n3346 SUB 0.14fF $ **FLOATING
C3697 S.n3348 SUB 1.16fF $ **FLOATING
C3698 S.n3349 SUB 0.22fF $ **FLOATING
C3699 S.n3350 SUB 0.25fF $ **FLOATING
C3700 S.n3351 SUB 0.09fF $ **FLOATING
C3701 S.n3352 SUB 1.88fF $ **FLOATING
C3702 S.t979 SUB 0.02fF
C3703 S.n3353 SUB 0.24fF $ **FLOATING
C3704 S.n3354 SUB 0.91fF $ **FLOATING
C3705 S.n3355 SUB 0.05fF $ **FLOATING
C3706 S.t2088 SUB 0.02fF
C3707 S.n3356 SUB 0.12fF $ **FLOATING
C3708 S.n3357 SUB 0.14fF $ **FLOATING
C3709 S.n3359 SUB 0.78fF $ **FLOATING
C3710 S.n3360 SUB 1.94fF $ **FLOATING
C3711 S.n3361 SUB 1.88fF $ **FLOATING
C3712 S.n3362 SUB 0.12fF $ **FLOATING
C3713 S.t1541 SUB 0.02fF
C3714 S.n3363 SUB 0.14fF $ **FLOATING
C3715 S.t797 SUB 0.02fF
C3716 S.n3365 SUB 0.24fF $ **FLOATING
C3717 S.n3366 SUB 0.36fF $ **FLOATING
C3718 S.n3367 SUB 0.61fF $ **FLOATING
C3719 S.n3368 SUB 1.84fF $ **FLOATING
C3720 S.n3369 SUB 2.99fF $ **FLOATING
C3721 S.t49 SUB 0.02fF
C3722 S.n3370 SUB 0.24fF $ **FLOATING
C3723 S.n3371 SUB 0.91fF $ **FLOATING
C3724 S.n3372 SUB 0.05fF $ **FLOATING
C3725 S.t2245 SUB 0.02fF
C3726 S.n3373 SUB 0.12fF $ **FLOATING
C3727 S.n3374 SUB 0.14fF $ **FLOATING
C3728 S.n3376 SUB 1.89fF $ **FLOATING
C3729 S.n3377 SUB 1.75fF $ **FLOATING
C3730 S.t2449 SUB 0.02fF
C3731 S.n3378 SUB 0.24fF $ **FLOATING
C3732 S.n3379 SUB 0.36fF $ **FLOATING
C3733 S.n3380 SUB 0.61fF $ **FLOATING
C3734 S.n3381 SUB 0.12fF $ **FLOATING
C3735 S.t681 SUB 0.02fF
C3736 S.n3382 SUB 0.14fF $ **FLOATING
C3737 S.n3384 SUB 1.16fF $ **FLOATING
C3738 S.n3385 SUB 0.22fF $ **FLOATING
C3739 S.n3386 SUB 0.25fF $ **FLOATING
C3740 S.n3387 SUB 0.09fF $ **FLOATING
C3741 S.n3388 SUB 2.44fF $ **FLOATING
C3742 S.t1743 SUB 0.02fF
C3743 S.n3389 SUB 0.24fF $ **FLOATING
C3744 S.n3390 SUB 0.91fF $ **FLOATING
C3745 S.n3391 SUB 0.05fF $ **FLOATING
C3746 S.t1386 SUB 0.02fF
C3747 S.n3392 SUB 0.12fF $ **FLOATING
C3748 S.n3393 SUB 0.14fF $ **FLOATING
C3749 S.n3395 SUB 1.88fF $ **FLOATING
C3750 S.n3396 SUB 0.48fF $ **FLOATING
C3751 S.n3397 SUB 0.09fF $ **FLOATING
C3752 S.n3398 SUB 0.33fF $ **FLOATING
C3753 S.n3399 SUB 0.30fF $ **FLOATING
C3754 S.n3400 SUB 0.77fF $ **FLOATING
C3755 S.n3401 SUB 0.59fF $ **FLOATING
C3756 S.t1581 SUB 0.02fF
C3757 S.n3402 SUB 0.24fF $ **FLOATING
C3758 S.n3403 SUB 0.36fF $ **FLOATING
C3759 S.n3404 SUB 0.61fF $ **FLOATING
C3760 S.n3405 SUB 0.12fF $ **FLOATING
C3761 S.t2340 SUB 0.02fF
C3762 S.n3406 SUB 0.14fF $ **FLOATING
C3763 S.n3408 SUB 2.61fF $ **FLOATING
C3764 S.n3409 SUB 2.16fF $ **FLOATING
C3765 S.t867 SUB 0.02fF
C3766 S.n3410 SUB 0.24fF $ **FLOATING
C3767 S.n3411 SUB 0.91fF $ **FLOATING
C3768 S.n3412 SUB 0.05fF $ **FLOATING
C3769 S.t515 SUB 0.02fF
C3770 S.n3413 SUB 0.12fF $ **FLOATING
C3771 S.n3414 SUB 0.14fF $ **FLOATING
C3772 S.n3416 SUB 0.78fF $ **FLOATING
C3773 S.n3417 SUB 2.30fF $ **FLOATING
C3774 S.n3418 SUB 1.88fF $ **FLOATING
C3775 S.n3419 SUB 0.12fF $ **FLOATING
C3776 S.t1481 SUB 0.02fF
C3777 S.n3420 SUB 0.14fF $ **FLOATING
C3778 S.t714 SUB 0.02fF
C3779 S.n3422 SUB 0.24fF $ **FLOATING
C3780 S.n3423 SUB 0.36fF $ **FLOATING
C3781 S.n3424 SUB 0.61fF $ **FLOATING
C3782 S.n3425 SUB 1.39fF $ **FLOATING
C3783 S.n3426 SUB 0.71fF $ **FLOATING
C3784 S.n3427 SUB 1.14fF $ **FLOATING
C3785 S.n3428 SUB 0.35fF $ **FLOATING
C3786 S.n3429 SUB 2.03fF $ **FLOATING
C3787 S.t2512 SUB 0.02fF
C3788 S.n3430 SUB 0.24fF $ **FLOATING
C3789 S.n3431 SUB 0.91fF $ **FLOATING
C3790 S.n3432 SUB 0.05fF $ **FLOATING
C3791 S.t2160 SUB 0.02fF
C3792 S.n3433 SUB 0.12fF $ **FLOATING
C3793 S.n3434 SUB 0.14fF $ **FLOATING
C3794 S.n3436 SUB 1.89fF $ **FLOATING
C3795 S.n3437 SUB 1.88fF $ **FLOATING
C3796 S.t2369 SUB 0.02fF
C3797 S.n3438 SUB 0.24fF $ **FLOATING
C3798 S.n3439 SUB 0.36fF $ **FLOATING
C3799 S.n3440 SUB 0.61fF $ **FLOATING
C3800 S.n3441 SUB 0.12fF $ **FLOATING
C3801 S.t619 SUB 0.02fF
C3802 S.n3442 SUB 0.14fF $ **FLOATING
C3803 S.n3444 SUB 1.16fF $ **FLOATING
C3804 S.n3445 SUB 0.22fF $ **FLOATING
C3805 S.n3446 SUB 0.25fF $ **FLOATING
C3806 S.n3447 SUB 0.09fF $ **FLOATING
C3807 S.n3448 SUB 1.88fF $ **FLOATING
C3808 S.t1637 SUB 0.02fF
C3809 S.n3449 SUB 0.24fF $ **FLOATING
C3810 S.n3450 SUB 0.91fF $ **FLOATING
C3811 S.n3451 SUB 0.05fF $ **FLOATING
C3812 S.t1431 SUB 0.02fF
C3813 S.n3452 SUB 0.12fF $ **FLOATING
C3814 S.n3453 SUB 0.14fF $ **FLOATING
C3815 S.n3455 SUB 20.78fF $ **FLOATING
C3816 S.n3456 SUB 1.88fF $ **FLOATING
C3817 S.n3457 SUB 2.68fF $ **FLOATING
C3818 S.t2308 SUB 0.02fF
C3819 S.n3458 SUB 0.24fF $ **FLOATING
C3820 S.n3459 SUB 0.36fF $ **FLOATING
C3821 S.n3460 SUB 0.61fF $ **FLOATING
C3822 S.n3461 SUB 0.12fF $ **FLOATING
C3823 S.t555 SUB 0.02fF
C3824 S.n3462 SUB 0.14fF $ **FLOATING
C3825 S.n3464 SUB 5.17fF $ **FLOATING
C3826 S.t1350 SUB 0.02fF
C3827 S.n3465 SUB 0.12fF $ **FLOATING
C3828 S.n3466 SUB 0.14fF $ **FLOATING
C3829 S.t1556 SUB 0.02fF
C3830 S.n3468 SUB 0.24fF $ **FLOATING
C3831 S.n3469 SUB 0.91fF $ **FLOATING
C3832 S.n3470 SUB 0.05fF $ **FLOATING
C3833 S.n3471 SUB 2.73fF $ **FLOATING
C3834 S.n3472 SUB 1.59fF $ **FLOATING
C3835 S.n3473 SUB 0.12fF $ **FLOATING
C3836 S.t690 SUB 0.02fF
C3837 S.n3474 SUB 0.14fF $ **FLOATING
C3838 S.t692 SUB 0.02fF
C3839 S.n3476 SUB 0.24fF $ **FLOATING
C3840 S.n3477 SUB 0.36fF $ **FLOATING
C3841 S.n3478 SUB 0.61fF $ **FLOATING
C3842 S.n3479 SUB 0.07fF $ **FLOATING
C3843 S.n3480 SUB 0.01fF $ **FLOATING
C3844 S.n3481 SUB 0.24fF $ **FLOATING
C3845 S.n3482 SUB 1.16fF $ **FLOATING
C3846 S.n3483 SUB 1.35fF $ **FLOATING
C3847 S.n3484 SUB 2.30fF $ **FLOATING
C3848 S.t1461 SUB 0.02fF
C3849 S.n3485 SUB 0.12fF $ **FLOATING
C3850 S.n3486 SUB 0.14fF $ **FLOATING
C3851 S.t1675 SUB 0.02fF
C3852 S.n3488 SUB 0.24fF $ **FLOATING
C3853 S.n3489 SUB 0.91fF $ **FLOATING
C3854 S.n3490 SUB 0.05fF $ **FLOATING
C3855 S.t444 SUB 48.31fF
C3856 S.t2421 SUB 0.02fF
C3857 S.n3491 SUB 0.24fF $ **FLOATING
C3858 S.n3492 SUB 0.91fF $ **FLOATING
C3859 S.n3493 SUB 0.05fF $ **FLOATING
C3860 S.t2209 SUB 0.02fF
C3861 S.n3494 SUB 0.12fF $ **FLOATING
C3862 S.n3495 SUB 0.14fF $ **FLOATING
C3863 S.n3497 SUB 0.12fF $ **FLOATING
C3864 S.t1421 SUB 0.02fF
C3865 S.n3498 SUB 0.14fF $ **FLOATING
C3866 S.n3500 SUB 2.30fF $ **FLOATING
C3867 S.n3501 SUB 2.94fF $ **FLOATING
C3868 S.n3502 SUB 4.88fF $ **FLOATING
C3869 S.t1315 SUB 0.02fF
C3870 S.n3503 SUB 0.12fF $ **FLOATING
C3871 S.n3504 SUB 0.14fF $ **FLOATING
C3872 S.t804 SUB 0.02fF
C3873 S.n3506 SUB 0.24fF $ **FLOATING
C3874 S.n3507 SUB 0.91fF $ **FLOATING
C3875 S.n3508 SUB 0.05fF $ **FLOATING
C3876 S.n3509 SUB 1.88fF $ **FLOATING
C3877 S.n3510 SUB 2.67fF $ **FLOATING
C3878 S.t1507 SUB 0.02fF
C3879 S.n3511 SUB 0.24fF $ **FLOATING
C3880 S.n3512 SUB 0.36fF $ **FLOATING
C3881 S.n3513 SUB 0.61fF $ **FLOATING
C3882 S.n3514 SUB 0.12fF $ **FLOATING
C3883 S.t241 SUB 0.02fF
C3884 S.n3515 SUB 0.14fF $ **FLOATING
C3885 S.n3517 SUB 5.44fF $ **FLOATING
C3886 S.t437 SUB 0.02fF
C3887 S.n3518 SUB 0.12fF $ **FLOATING
C3888 S.n3519 SUB 0.14fF $ **FLOATING
C3889 S.t938 SUB 0.02fF
C3890 S.n3521 SUB 0.24fF $ **FLOATING
C3891 S.n3522 SUB 0.91fF $ **FLOATING
C3892 S.n3523 SUB 0.05fF $ **FLOATING
C3893 S.t240 SUB 47.92fF
C3894 S.t877 SUB 0.02fF
C3895 S.n3524 SUB 1.19fF $ **FLOATING
C3896 S.n3525 SUB 0.05fF $ **FLOATING
C3897 S.t2000 SUB 0.02fF
C3898 S.n3526 SUB 0.01fF $ **FLOATING
C3899 S.n3527 SUB 0.26fF $ **FLOATING
C3900 S.n3529 SUB 1.50fF $ **FLOATING
C3901 S.n3530 SUB 1.30fF $ **FLOATING
C3902 S.n3531 SUB 0.28fF $ **FLOATING
C3903 S.n3532 SUB 0.24fF $ **FLOATING
C3904 S.n3533 SUB 4.39fF $ **FLOATING
C3905 S.n3534 SUB 0.01fF $ **FLOATING
C3906 S.n3535 SUB 0.02fF $ **FLOATING
C3907 S.n3536 SUB 0.03fF $ **FLOATING
C3908 S.n3537 SUB 0.04fF $ **FLOATING
C3909 S.n3538 SUB 0.17fF $ **FLOATING
C3910 S.n3539 SUB 0.01fF $ **FLOATING
C3911 S.n3540 SUB 0.02fF $ **FLOATING
C3912 S.n3541 SUB 0.01fF $ **FLOATING
C3913 S.n3542 SUB 0.01fF $ **FLOATING
C3914 S.n3543 SUB 0.01fF $ **FLOATING
C3915 S.n3544 SUB 0.01fF $ **FLOATING
C3916 S.n3545 SUB 0.02fF $ **FLOATING
C3917 S.n3546 SUB 0.01fF $ **FLOATING
C3918 S.n3547 SUB 0.02fF $ **FLOATING
C3919 S.n3548 SUB 0.05fF $ **FLOATING
C3920 S.n3549 SUB 0.04fF $ **FLOATING
C3921 S.n3550 SUB 0.11fF $ **FLOATING
C3922 S.n3551 SUB 0.38fF $ **FLOATING
C3923 S.n3552 SUB 0.20fF $ **FLOATING
C3924 S.n3553 SUB 8.97fF $ **FLOATING
C3925 S.n3554 SUB 8.97fF $ **FLOATING
C3926 S.n3555 SUB 0.60fF $ **FLOATING
C3927 S.n3556 SUB 0.22fF $ **FLOATING
C3928 S.n3557 SUB 0.59fF $ **FLOATING
C3929 S.n3558 SUB 3.43fF $ **FLOATING
C3930 S.n3559 SUB 0.29fF $ **FLOATING
C3931 S.t78 SUB 21.38fF
C3932 S.n3560 SUB 21.67fF $ **FLOATING
C3933 S.n3561 SUB 0.77fF $ **FLOATING
C3934 S.n3562 SUB 0.28fF $ **FLOATING
C3935 S.n3563 SUB 4.00fF $ **FLOATING
C3936 S.n3564 SUB 1.35fF $ **FLOATING
C3937 S.t1016 SUB 0.02fF
C3938 S.n3565 SUB 0.64fF $ **FLOATING
C3939 S.n3566 SUB 0.61fF $ **FLOATING
C3940 S.n3567 SUB 1.89fF $ **FLOATING
C3941 S.n3568 SUB 0.06fF $ **FLOATING
C3942 S.n3569 SUB 0.03fF $ **FLOATING
C3943 S.n3570 SUB 0.04fF $ **FLOATING
C3944 S.n3571 SUB 0.99fF $ **FLOATING
C3945 S.n3572 SUB 0.02fF $ **FLOATING
C3946 S.n3573 SUB 0.01fF $ **FLOATING
C3947 S.n3574 SUB 0.02fF $ **FLOATING
C3948 S.n3575 SUB 0.08fF $ **FLOATING
C3949 S.n3576 SUB 0.36fF $ **FLOATING
C3950 S.n3577 SUB 1.85fF $ **FLOATING
C3951 S.t680 SUB 0.02fF
C3952 S.n3578 SUB 0.24fF $ **FLOATING
C3953 S.n3579 SUB 0.36fF $ **FLOATING
C3954 S.n3580 SUB 0.61fF $ **FLOATING
C3955 S.n3581 SUB 0.12fF $ **FLOATING
C3956 S.t165 SUB 0.02fF
C3957 S.n3582 SUB 0.14fF $ **FLOATING
C3958 S.n3584 SUB 0.70fF $ **FLOATING
C3959 S.n3585 SUB 0.23fF $ **FLOATING
C3960 S.n3586 SUB 0.23fF $ **FLOATING
C3961 S.n3587 SUB 0.70fF $ **FLOATING
C3962 S.n3588 SUB 1.16fF $ **FLOATING
C3963 S.n3589 SUB 0.22fF $ **FLOATING
C3964 S.n3590 SUB 0.25fF $ **FLOATING
C3965 S.n3591 SUB 0.09fF $ **FLOATING
C3966 S.n3592 SUB 1.88fF $ **FLOATING
C3967 S.t1822 SUB 0.02fF
C3968 S.n3593 SUB 0.24fF $ **FLOATING
C3969 S.n3594 SUB 0.91fF $ **FLOATING
C3970 S.n3595 SUB 0.05fF $ **FLOATING
C3971 S.t341 SUB 0.02fF
C3972 S.n3596 SUB 0.12fF $ **FLOATING
C3973 S.n3597 SUB 0.14fF $ **FLOATING
C3974 S.n3599 SUB 0.25fF $ **FLOATING
C3975 S.n3600 SUB 0.09fF $ **FLOATING
C3976 S.n3601 SUB 0.21fF $ **FLOATING
C3977 S.n3602 SUB 0.92fF $ **FLOATING
C3978 S.n3603 SUB 0.44fF $ **FLOATING
C3979 S.n3604 SUB 1.88fF $ **FLOATING
C3980 S.n3605 SUB 0.12fF $ **FLOATING
C3981 S.t1945 SUB 0.02fF
C3982 S.n3606 SUB 0.14fF $ **FLOATING
C3983 S.t2446 SUB 0.02fF
C3984 S.n3608 SUB 0.24fF $ **FLOATING
C3985 S.n3609 SUB 0.36fF $ **FLOATING
C3986 S.n3610 SUB 0.61fF $ **FLOATING
C3987 S.n3611 SUB 0.02fF $ **FLOATING
C3988 S.n3612 SUB 0.01fF $ **FLOATING
C3989 S.n3613 SUB 0.02fF $ **FLOATING
C3990 S.n3614 SUB 0.08fF $ **FLOATING
C3991 S.n3615 SUB 0.06fF $ **FLOATING
C3992 S.n3616 SUB 0.03fF $ **FLOATING
C3993 S.n3617 SUB 0.04fF $ **FLOATING
C3994 S.n3618 SUB 1.00fF $ **FLOATING
C3995 S.n3619 SUB 0.36fF $ **FLOATING
C3996 S.n3620 SUB 1.87fF $ **FLOATING
C3997 S.n3621 SUB 1.99fF $ **FLOATING
C3998 S.t1083 SUB 0.02fF
C3999 S.n3622 SUB 0.24fF $ **FLOATING
C4000 S.n3623 SUB 0.91fF $ **FLOATING
C4001 S.n3624 SUB 0.05fF $ **FLOATING
C4002 S.t1999 SUB 0.02fF
C4003 S.n3625 SUB 0.12fF $ **FLOATING
C4004 S.n3626 SUB 0.14fF $ **FLOATING
C4005 S.n3628 SUB 1.89fF $ **FLOATING
C4006 S.n3629 SUB 0.06fF $ **FLOATING
C4007 S.n3630 SUB 0.03fF $ **FLOATING
C4008 S.n3631 SUB 0.04fF $ **FLOATING
C4009 S.n3632 SUB 0.99fF $ **FLOATING
C4010 S.n3633 SUB 0.02fF $ **FLOATING
C4011 S.n3634 SUB 0.01fF $ **FLOATING
C4012 S.n3635 SUB 0.02fF $ **FLOATING
C4013 S.n3636 SUB 0.08fF $ **FLOATING
C4014 S.n3637 SUB 0.36fF $ **FLOATING
C4015 S.n3638 SUB 1.85fF $ **FLOATING
C4016 S.t1579 SUB 0.02fF
C4017 S.n3639 SUB 0.24fF $ **FLOATING
C4018 S.n3640 SUB 0.36fF $ **FLOATING
C4019 S.n3641 SUB 0.61fF $ **FLOATING
C4020 S.n3642 SUB 0.12fF $ **FLOATING
C4021 S.t1088 SUB 0.02fF
C4022 S.n3643 SUB 0.14fF $ **FLOATING
C4023 S.n3645 SUB 0.70fF $ **FLOATING
C4024 S.n3646 SUB 0.23fF $ **FLOATING
C4025 S.n3647 SUB 0.23fF $ **FLOATING
C4026 S.n3648 SUB 0.70fF $ **FLOATING
C4027 S.n3649 SUB 1.16fF $ **FLOATING
C4028 S.n3650 SUB 0.22fF $ **FLOATING
C4029 S.n3651 SUB 0.25fF $ **FLOATING
C4030 S.n3652 SUB 0.09fF $ **FLOATING
C4031 S.n3653 SUB 1.88fF $ **FLOATING
C4032 S.t206 SUB 0.02fF
C4033 S.n3654 SUB 0.24fF $ **FLOATING
C4034 S.n3655 SUB 0.91fF $ **FLOATING
C4035 S.n3656 SUB 0.05fF $ **FLOATING
C4036 S.t1149 SUB 0.02fF
C4037 S.n3657 SUB 0.12fF $ **FLOATING
C4038 S.n3658 SUB 0.14fF $ **FLOATING
C4039 S.n3660 SUB 0.25fF $ **FLOATING
C4040 S.n3661 SUB 0.09fF $ **FLOATING
C4041 S.n3662 SUB 0.21fF $ **FLOATING
C4042 S.n3663 SUB 0.92fF $ **FLOATING
C4043 S.n3664 SUB 0.44fF $ **FLOATING
C4044 S.n3665 SUB 1.88fF $ **FLOATING
C4045 S.n3666 SUB 0.12fF $ **FLOATING
C4046 S.t210 SUB 0.02fF
C4047 S.n3667 SUB 0.14fF $ **FLOATING
C4048 S.t712 SUB 0.02fF
C4049 S.n3669 SUB 0.24fF $ **FLOATING
C4050 S.n3670 SUB 0.36fF $ **FLOATING
C4051 S.n3671 SUB 0.61fF $ **FLOATING
C4052 S.n3672 SUB 0.02fF $ **FLOATING
C4053 S.n3673 SUB 0.01fF $ **FLOATING
C4054 S.n3674 SUB 0.02fF $ **FLOATING
C4055 S.n3675 SUB 0.08fF $ **FLOATING
C4056 S.n3676 SUB 0.06fF $ **FLOATING
C4057 S.n3677 SUB 0.03fF $ **FLOATING
C4058 S.n3678 SUB 0.04fF $ **FLOATING
C4059 S.n3679 SUB 1.00fF $ **FLOATING
C4060 S.n3680 SUB 0.36fF $ **FLOATING
C4061 S.n3681 SUB 1.87fF $ **FLOATING
C4062 S.n3682 SUB 1.99fF $ **FLOATING
C4063 S.t1874 SUB 0.02fF
C4064 S.n3683 SUB 0.24fF $ **FLOATING
C4065 S.n3684 SUB 0.91fF $ **FLOATING
C4066 S.n3685 SUB 0.05fF $ **FLOATING
C4067 S.t271 SUB 0.02fF
C4068 S.n3686 SUB 0.12fF $ **FLOATING
C4069 S.n3687 SUB 0.14fF $ **FLOATING
C4070 S.n3689 SUB 1.89fF $ **FLOATING
C4071 S.n3690 SUB 0.06fF $ **FLOATING
C4072 S.n3691 SUB 0.03fF $ **FLOATING
C4073 S.n3692 SUB 0.04fF $ **FLOATING
C4074 S.n3693 SUB 0.99fF $ **FLOATING
C4075 S.n3694 SUB 0.02fF $ **FLOATING
C4076 S.n3695 SUB 0.01fF $ **FLOATING
C4077 S.n3696 SUB 0.02fF $ **FLOATING
C4078 S.n3697 SUB 0.08fF $ **FLOATING
C4079 S.n3698 SUB 0.36fF $ **FLOATING
C4080 S.n3699 SUB 1.85fF $ **FLOATING
C4081 S.t2367 SUB 0.02fF
C4082 S.n3700 SUB 0.24fF $ **FLOATING
C4083 S.n3701 SUB 0.36fF $ **FLOATING
C4084 S.n3702 SUB 0.61fF $ **FLOATING
C4085 S.n3703 SUB 0.12fF $ **FLOATING
C4086 S.t1878 SUB 0.02fF
C4087 S.n3704 SUB 0.14fF $ **FLOATING
C4088 S.n3706 SUB 0.70fF $ **FLOATING
C4089 S.n3707 SUB 0.23fF $ **FLOATING
C4090 S.n3708 SUB 0.23fF $ **FLOATING
C4091 S.n3709 SUB 0.70fF $ **FLOATING
C4092 S.n3710 SUB 1.16fF $ **FLOATING
C4093 S.n3711 SUB 0.22fF $ **FLOATING
C4094 S.n3712 SUB 0.25fF $ **FLOATING
C4095 S.n3713 SUB 0.09fF $ **FLOATING
C4096 S.n3714 SUB 1.88fF $ **FLOATING
C4097 S.t1005 SUB 0.02fF
C4098 S.n3715 SUB 0.24fF $ **FLOATING
C4099 S.n3716 SUB 0.91fF $ **FLOATING
C4100 S.n3717 SUB 0.05fF $ **FLOATING
C4101 S.t1933 SUB 0.02fF
C4102 S.n3718 SUB 0.12fF $ **FLOATING
C4103 S.n3719 SUB 0.14fF $ **FLOATING
C4104 S.n3721 SUB 0.25fF $ **FLOATING
C4105 S.n3722 SUB 0.09fF $ **FLOATING
C4106 S.n3723 SUB 0.21fF $ **FLOATING
C4107 S.n3724 SUB 0.92fF $ **FLOATING
C4108 S.n3725 SUB 0.44fF $ **FLOATING
C4109 S.n3726 SUB 1.88fF $ **FLOATING
C4110 S.n3727 SUB 0.12fF $ **FLOATING
C4111 S.t1013 SUB 0.02fF
C4112 S.n3728 SUB 0.14fF $ **FLOATING
C4113 S.t1510 SUB 0.02fF
C4114 S.n3730 SUB 0.24fF $ **FLOATING
C4115 S.n3731 SUB 0.36fF $ **FLOATING
C4116 S.n3732 SUB 0.61fF $ **FLOATING
C4117 S.n3733 SUB 0.02fF $ **FLOATING
C4118 S.n3734 SUB 0.01fF $ **FLOATING
C4119 S.n3735 SUB 0.02fF $ **FLOATING
C4120 S.n3736 SUB 0.08fF $ **FLOATING
C4121 S.n3737 SUB 0.06fF $ **FLOATING
C4122 S.n3738 SUB 0.03fF $ **FLOATING
C4123 S.n3739 SUB 0.04fF $ **FLOATING
C4124 S.n3740 SUB 1.00fF $ **FLOATING
C4125 S.n3741 SUB 0.36fF $ **FLOATING
C4126 S.n3742 SUB 1.87fF $ **FLOATING
C4127 S.n3743 SUB 1.99fF $ **FLOATING
C4128 S.t105 SUB 0.02fF
C4129 S.n3744 SUB 0.24fF $ **FLOATING
C4130 S.n3745 SUB 0.91fF $ **FLOATING
C4131 S.n3746 SUB 0.05fF $ **FLOATING
C4132 S.t1074 SUB 0.02fF
C4133 S.n3747 SUB 0.12fF $ **FLOATING
C4134 S.n3748 SUB 0.14fF $ **FLOATING
C4135 S.n3750 SUB 1.89fF $ **FLOATING
C4136 S.n3751 SUB 0.06fF $ **FLOATING
C4137 S.n3752 SUB 0.03fF $ **FLOATING
C4138 S.n3753 SUB 0.04fF $ **FLOATING
C4139 S.n3754 SUB 0.99fF $ **FLOATING
C4140 S.n3755 SUB 0.02fF $ **FLOATING
C4141 S.n3756 SUB 0.01fF $ **FLOATING
C4142 S.n3757 SUB 0.02fF $ **FLOATING
C4143 S.n3758 SUB 0.08fF $ **FLOATING
C4144 S.n3759 SUB 0.36fF $ **FLOATING
C4145 S.n3760 SUB 1.85fF $ **FLOATING
C4146 S.t650 SUB 0.02fF
C4147 S.n3761 SUB 0.24fF $ **FLOATING
C4148 S.n3762 SUB 0.36fF $ **FLOATING
C4149 S.n3763 SUB 0.61fF $ **FLOATING
C4150 S.n3764 SUB 0.12fF $ **FLOATING
C4151 S.t110 SUB 0.02fF
C4152 S.n3765 SUB 0.14fF $ **FLOATING
C4153 S.n3767 SUB 0.70fF $ **FLOATING
C4154 S.n3768 SUB 0.23fF $ **FLOATING
C4155 S.n3769 SUB 0.23fF $ **FLOATING
C4156 S.n3770 SUB 0.70fF $ **FLOATING
C4157 S.n3771 SUB 1.16fF $ **FLOATING
C4158 S.n3772 SUB 0.22fF $ **FLOATING
C4159 S.n3773 SUB 0.25fF $ **FLOATING
C4160 S.n3774 SUB 0.09fF $ **FLOATING
C4161 S.n3775 SUB 1.88fF $ **FLOATING
C4162 S.t1778 SUB 0.02fF
C4163 S.n3776 SUB 0.24fF $ **FLOATING
C4164 S.n3777 SUB 0.91fF $ **FLOATING
C4165 S.n3778 SUB 0.05fF $ **FLOATING
C4166 S.t308 SUB 0.02fF
C4167 S.n3779 SUB 0.12fF $ **FLOATING
C4168 S.n3780 SUB 0.14fF $ **FLOATING
C4169 S.n3782 SUB 0.25fF $ **FLOATING
C4170 S.n3783 SUB 0.09fF $ **FLOATING
C4171 S.n3784 SUB 0.21fF $ **FLOATING
C4172 S.n3785 SUB 0.92fF $ **FLOATING
C4173 S.n3786 SUB 0.44fF $ **FLOATING
C4174 S.n3787 SUB 1.88fF $ **FLOATING
C4175 S.n3788 SUB 0.12fF $ **FLOATING
C4176 S.t1305 SUB 0.02fF
C4177 S.n3789 SUB 0.14fF $ **FLOATING
C4178 S.t1858 SUB 0.02fF
C4179 S.n3791 SUB 0.24fF $ **FLOATING
C4180 S.n3792 SUB 0.36fF $ **FLOATING
C4181 S.n3793 SUB 0.61fF $ **FLOATING
C4182 S.n3794 SUB 0.02fF $ **FLOATING
C4183 S.n3795 SUB 0.01fF $ **FLOATING
C4184 S.n3796 SUB 0.02fF $ **FLOATING
C4185 S.n3797 SUB 0.08fF $ **FLOATING
C4186 S.n3798 SUB 0.06fF $ **FLOATING
C4187 S.n3799 SUB 0.03fF $ **FLOATING
C4188 S.n3800 SUB 0.04fF $ **FLOATING
C4189 S.n3801 SUB 1.00fF $ **FLOATING
C4190 S.n3802 SUB 0.36fF $ **FLOATING
C4191 S.n3803 SUB 1.87fF $ **FLOATING
C4192 S.n3804 SUB 1.99fF $ **FLOATING
C4193 S.t881 SUB 0.02fF
C4194 S.n3805 SUB 0.24fF $ **FLOATING
C4195 S.n3806 SUB 0.91fF $ **FLOATING
C4196 S.n3807 SUB 0.05fF $ **FLOATING
C4197 S.t1489 SUB 0.02fF
C4198 S.n3808 SUB 0.12fF $ **FLOATING
C4199 S.n3809 SUB 0.14fF $ **FLOATING
C4200 S.n3811 SUB 1.89fF $ **FLOATING
C4201 S.n3812 SUB 0.07fF $ **FLOATING
C4202 S.n3813 SUB 0.04fF $ **FLOATING
C4203 S.n3814 SUB 0.05fF $ **FLOATING
C4204 S.n3815 SUB 0.87fF $ **FLOATING
C4205 S.n3816 SUB 0.01fF $ **FLOATING
C4206 S.n3817 SUB 0.01fF $ **FLOATING
C4207 S.n3818 SUB 0.01fF $ **FLOATING
C4208 S.n3819 SUB 0.07fF $ **FLOATING
C4209 S.n3820 SUB 0.68fF $ **FLOATING
C4210 S.n3821 SUB 0.72fF $ **FLOATING
C4211 S.t991 SUB 0.02fF
C4212 S.n3822 SUB 0.24fF $ **FLOATING
C4213 S.n3823 SUB 0.36fF $ **FLOATING
C4214 S.n3824 SUB 0.61fF $ **FLOATING
C4215 S.n3825 SUB 0.12fF $ **FLOATING
C4216 S.t423 SUB 0.02fF
C4217 S.n3826 SUB 0.14fF $ **FLOATING
C4218 S.n3828 SUB 0.70fF $ **FLOATING
C4219 S.n3829 SUB 0.23fF $ **FLOATING
C4220 S.n3830 SUB 0.23fF $ **FLOATING
C4221 S.n3831 SUB 0.70fF $ **FLOATING
C4222 S.n3832 SUB 1.16fF $ **FLOATING
C4223 S.n3833 SUB 0.22fF $ **FLOATING
C4224 S.n3834 SUB 0.25fF $ **FLOATING
C4225 S.n3835 SUB 0.09fF $ **FLOATING
C4226 S.n3836 SUB 2.31fF $ **FLOATING
C4227 S.t2526 SUB 0.02fF
C4228 S.n3837 SUB 0.24fF $ **FLOATING
C4229 S.n3838 SUB 0.91fF $ **FLOATING
C4230 S.n3839 SUB 0.05fF $ **FLOATING
C4231 S.t624 SUB 0.02fF
C4232 S.n3840 SUB 0.12fF $ **FLOATING
C4233 S.n3841 SUB 0.14fF $ **FLOATING
C4234 S.n3843 SUB 1.88fF $ **FLOATING
C4235 S.n3844 SUB 0.46fF $ **FLOATING
C4236 S.n3845 SUB 0.22fF $ **FLOATING
C4237 S.n3846 SUB 0.38fF $ **FLOATING
C4238 S.n3847 SUB 0.16fF $ **FLOATING
C4239 S.n3848 SUB 0.28fF $ **FLOATING
C4240 S.n3849 SUB 0.21fF $ **FLOATING
C4241 S.n3850 SUB 0.30fF $ **FLOATING
C4242 S.n3851 SUB 0.42fF $ **FLOATING
C4243 S.n3852 SUB 0.21fF $ **FLOATING
C4244 S.t79 SUB 0.02fF
C4245 S.n3853 SUB 0.24fF $ **FLOATING
C4246 S.n3854 SUB 0.36fF $ **FLOATING
C4247 S.n3855 SUB 0.61fF $ **FLOATING
C4248 S.n3856 SUB 0.12fF $ **FLOATING
C4249 S.t2075 SUB 0.02fF
C4250 S.n3857 SUB 0.14fF $ **FLOATING
C4251 S.n3859 SUB 0.04fF $ **FLOATING
C4252 S.n3860 SUB 0.03fF $ **FLOATING
C4253 S.n3861 SUB 0.03fF $ **FLOATING
C4254 S.n3862 SUB 0.10fF $ **FLOATING
C4255 S.n3863 SUB 0.36fF $ **FLOATING
C4256 S.n3864 SUB 0.38fF $ **FLOATING
C4257 S.n3865 SUB 0.11fF $ **FLOATING
C4258 S.n3866 SUB 0.12fF $ **FLOATING
C4259 S.n3867 SUB 0.07fF $ **FLOATING
C4260 S.n3868 SUB 0.12fF $ **FLOATING
C4261 S.n3869 SUB 0.18fF $ **FLOATING
C4262 S.n3870 SUB 4.00fF $ **FLOATING
C4263 S.t1650 SUB 0.02fF
C4264 S.n3871 SUB 0.24fF $ **FLOATING
C4265 S.n3872 SUB 0.91fF $ **FLOATING
C4266 S.n3873 SUB 0.05fF $ **FLOATING
C4267 S.t2283 SUB 0.02fF
C4268 S.n3874 SUB 0.12fF $ **FLOATING
C4269 S.n3875 SUB 0.14fF $ **FLOATING
C4270 S.n3877 SUB 0.25fF $ **FLOATING
C4271 S.n3878 SUB 0.09fF $ **FLOATING
C4272 S.n3879 SUB 0.21fF $ **FLOATING
C4273 S.n3880 SUB 1.28fF $ **FLOATING
C4274 S.n3881 SUB 0.53fF $ **FLOATING
C4275 S.n3882 SUB 1.88fF $ **FLOATING
C4276 S.n3883 SUB 0.12fF $ **FLOATING
C4277 S.t1214 SUB 0.02fF
C4278 S.n3884 SUB 0.14fF $ **FLOATING
C4279 S.t1758 SUB 0.02fF
C4280 S.n3886 SUB 0.24fF $ **FLOATING
C4281 S.n3887 SUB 0.36fF $ **FLOATING
C4282 S.n3888 SUB 0.61fF $ **FLOATING
C4283 S.n3889 SUB 1.58fF $ **FLOATING
C4284 S.n3890 SUB 2.45fF $ **FLOATING
C4285 S.t779 SUB 0.02fF
C4286 S.n3891 SUB 0.24fF $ **FLOATING
C4287 S.n3892 SUB 0.91fF $ **FLOATING
C4288 S.n3893 SUB 0.05fF $ **FLOATING
C4289 S.t1429 SUB 0.02fF
C4290 S.n3894 SUB 0.12fF $ **FLOATING
C4291 S.n3895 SUB 0.14fF $ **FLOATING
C4292 S.n3897 SUB 1.89fF $ **FLOATING
C4293 S.n3898 SUB 0.06fF $ **FLOATING
C4294 S.n3899 SUB 0.03fF $ **FLOATING
C4295 S.n3900 SUB 0.04fF $ **FLOATING
C4296 S.n3901 SUB 0.99fF $ **FLOATING
C4297 S.n3902 SUB 0.02fF $ **FLOATING
C4298 S.n3903 SUB 0.01fF $ **FLOATING
C4299 S.n3904 SUB 0.02fF $ **FLOATING
C4300 S.n3905 SUB 0.08fF $ **FLOATING
C4301 S.n3906 SUB 0.36fF $ **FLOATING
C4302 S.n3907 SUB 1.85fF $ **FLOATING
C4303 S.t1040 SUB 0.02fF
C4304 S.n3908 SUB 0.24fF $ **FLOATING
C4305 S.n3909 SUB 0.36fF $ **FLOATING
C4306 S.n3910 SUB 0.61fF $ **FLOATING
C4307 S.n3911 SUB 0.12fF $ **FLOATING
C4308 S.t483 SUB 0.02fF
C4309 S.n3912 SUB 0.14fF $ **FLOATING
C4310 S.n3914 SUB 0.70fF $ **FLOATING
C4311 S.n3915 SUB 0.23fF $ **FLOATING
C4312 S.n3916 SUB 0.23fF $ **FLOATING
C4313 S.n3917 SUB 0.70fF $ **FLOATING
C4314 S.n3918 SUB 1.16fF $ **FLOATING
C4315 S.n3919 SUB 0.22fF $ **FLOATING
C4316 S.n3920 SUB 0.25fF $ **FLOATING
C4317 S.n3921 SUB 0.09fF $ **FLOATING
C4318 S.n3922 SUB 1.88fF $ **FLOATING
C4319 S.t2584 SUB 0.02fF
C4320 S.n3923 SUB 0.24fF $ **FLOATING
C4321 S.n3924 SUB 0.91fF $ **FLOATING
C4322 S.n3925 SUB 0.05fF $ **FLOATING
C4323 S.t564 SUB 0.02fF
C4324 S.n3926 SUB 0.12fF $ **FLOATING
C4325 S.n3927 SUB 0.14fF $ **FLOATING
C4326 S.n3929 SUB 20.78fF $ **FLOATING
C4327 S.n3930 SUB 0.06fF $ **FLOATING
C4328 S.n3931 SUB 0.20fF $ **FLOATING
C4329 S.n3932 SUB 0.09fF $ **FLOATING
C4330 S.n3933 SUB 0.21fF $ **FLOATING
C4331 S.n3934 SUB 0.10fF $ **FLOATING
C4332 S.n3935 SUB 0.30fF $ **FLOATING
C4333 S.n3936 SUB 0.69fF $ **FLOATING
C4334 S.n3937 SUB 0.45fF $ **FLOATING
C4335 S.n3938 SUB 2.33fF $ **FLOATING
C4336 S.n3939 SUB 0.12fF $ **FLOATING
C4337 S.t1053 SUB 0.02fF
C4338 S.n3940 SUB 0.14fF $ **FLOATING
C4339 S.t1540 SUB 0.02fF
C4340 S.n3942 SUB 0.24fF $ **FLOATING
C4341 S.n3943 SUB 0.36fF $ **FLOATING
C4342 S.n3944 SUB 0.61fF $ **FLOATING
C4343 S.n3945 SUB 1.90fF $ **FLOATING
C4344 S.n3946 SUB 0.17fF $ **FLOATING
C4345 S.n3947 SUB 0.76fF $ **FLOATING
C4346 S.n3948 SUB 0.32fF $ **FLOATING
C4347 S.n3949 SUB 0.25fF $ **FLOATING
C4348 S.n3950 SUB 0.30fF $ **FLOATING
C4349 S.n3951 SUB 0.47fF $ **FLOATING
C4350 S.n3952 SUB 0.16fF $ **FLOATING
C4351 S.n3953 SUB 1.93fF $ **FLOATING
C4352 S.t1222 SUB 0.02fF
C4353 S.n3954 SUB 0.12fF $ **FLOATING
C4354 S.n3955 SUB 0.14fF $ **FLOATING
C4355 S.t161 SUB 0.02fF
C4356 S.n3957 SUB 0.24fF $ **FLOATING
C4357 S.n3958 SUB 0.91fF $ **FLOATING
C4358 S.n3959 SUB 0.05fF $ **FLOATING
C4359 S.n3960 SUB 1.88fF $ **FLOATING
C4360 S.n3961 SUB 0.12fF $ **FLOATING
C4361 S.t2293 SUB 0.02fF
C4362 S.n3962 SUB 0.14fF $ **FLOATING
C4363 S.t588 SUB 0.02fF
C4364 S.n3964 SUB 0.12fF $ **FLOATING
C4365 S.n3965 SUB 0.14fF $ **FLOATING
C4366 S.t800 SUB 0.02fF
C4367 S.n3967 SUB 0.24fF $ **FLOATING
C4368 S.n3968 SUB 0.91fF $ **FLOATING
C4369 S.n3969 SUB 0.05fF $ **FLOATING
C4370 S.t1531 SUB 0.02fF
C4371 S.n3970 SUB 0.24fF $ **FLOATING
C4372 S.n3971 SUB 0.36fF $ **FLOATING
C4373 S.n3972 SUB 0.61fF $ **FLOATING
C4374 S.n3973 SUB 0.32fF $ **FLOATING
C4375 S.n3974 SUB 1.09fF $ **FLOATING
C4376 S.n3975 SUB 0.15fF $ **FLOATING
C4377 S.n3976 SUB 2.10fF $ **FLOATING
C4378 S.n3977 SUB 2.94fF $ **FLOATING
C4379 S.n3978 SUB 1.88fF $ **FLOATING
C4380 S.n3979 SUB 0.12fF $ **FLOATING
C4381 S.t2130 SUB 0.02fF
C4382 S.n3980 SUB 0.14fF $ **FLOATING
C4383 S.t145 SUB 0.02fF
C4384 S.n3982 SUB 0.24fF $ **FLOATING
C4385 S.n3983 SUB 0.36fF $ **FLOATING
C4386 S.n3984 SUB 0.61fF $ **FLOATING
C4387 S.n3985 SUB 0.92fF $ **FLOATING
C4388 S.n3986 SUB 0.32fF $ **FLOATING
C4389 S.n3987 SUB 0.92fF $ **FLOATING
C4390 S.n3988 SUB 1.09fF $ **FLOATING
C4391 S.n3989 SUB 0.15fF $ **FLOATING
C4392 S.n3990 SUB 4.96fF $ **FLOATING
C4393 S.t2206 SUB 0.02fF
C4394 S.n3991 SUB 0.12fF $ **FLOATING
C4395 S.n3992 SUB 0.14fF $ **FLOATING
C4396 S.t1707 SUB 0.02fF
C4397 S.n3994 SUB 0.24fF $ **FLOATING
C4398 S.n3995 SUB 0.91fF $ **FLOATING
C4399 S.n3996 SUB 0.05fF $ **FLOATING
C4400 S.t1348 SUB 0.02fF
C4401 S.n3997 SUB 0.12fF $ **FLOATING
C4402 S.n3998 SUB 0.14fF $ **FLOATING
C4403 S.n4000 SUB 1.88fF $ **FLOATING
C4404 S.n4001 SUB 2.67fF $ **FLOATING
C4405 S.t1815 SUB 0.02fF
C4406 S.n4002 SUB 0.24fF $ **FLOATING
C4407 S.n4003 SUB 0.36fF $ **FLOATING
C4408 S.n4004 SUB 0.61fF $ **FLOATING
C4409 S.n4005 SUB 0.12fF $ **FLOATING
C4410 S.t1266 SUB 0.02fF
C4411 S.n4006 SUB 0.14fF $ **FLOATING
C4412 S.n4008 SUB 1.88fF $ **FLOATING
C4413 S.n4009 SUB 2.67fF $ **FLOATING
C4414 S.t672 SUB 0.02fF
C4415 S.n4010 SUB 0.24fF $ **FLOATING
C4416 S.n4011 SUB 0.36fF $ **FLOATING
C4417 S.n4012 SUB 0.61fF $ **FLOATING
C4418 S.t2450 SUB 0.02fF
C4419 S.n4013 SUB 0.24fF $ **FLOATING
C4420 S.n4014 SUB 0.91fF $ **FLOATING
C4421 S.n4015 SUB 0.05fF $ **FLOATING
C4422 S.t2234 SUB 0.02fF
C4423 S.n4016 SUB 0.12fF $ **FLOATING
C4424 S.n4017 SUB 0.14fF $ **FLOATING
C4425 S.n4019 SUB 0.12fF $ **FLOATING
C4426 S.t1438 SUB 0.02fF
C4427 S.n4020 SUB 0.14fF $ **FLOATING
C4428 S.n4022 SUB 2.30fF $ **FLOATING
C4429 S.n4023 SUB 2.94fF $ **FLOATING
C4430 S.n4024 SUB 5.16fF $ **FLOATING
C4431 S.t836 SUB 0.02fF
C4432 S.n4025 SUB 0.24fF $ **FLOATING
C4433 S.n4026 SUB 0.91fF $ **FLOATING
C4434 S.n4027 SUB 0.05fF $ **FLOATING
C4435 S.n4028 SUB 1.88fF $ **FLOATING
C4436 S.n4029 SUB 2.67fF $ **FLOATING
C4437 S.t948 SUB 0.02fF
C4438 S.n4030 SUB 0.24fF $ **FLOATING
C4439 S.n4031 SUB 0.36fF $ **FLOATING
C4440 S.n4032 SUB 0.61fF $ **FLOATING
C4441 S.n4033 SUB 0.12fF $ **FLOATING
C4442 S.t383 SUB 0.02fF
C4443 S.n4034 SUB 0.14fF $ **FLOATING
C4444 S.n4036 SUB 4.90fF $ **FLOATING
C4445 S.t470 SUB 0.02fF
C4446 S.n4037 SUB 0.12fF $ **FLOATING
C4447 S.n4038 SUB 0.14fF $ **FLOATING
C4448 S.t2480 SUB 0.02fF
C4449 S.n4040 SUB 0.24fF $ **FLOATING
C4450 S.n4041 SUB 0.91fF $ **FLOATING
C4451 S.n4042 SUB 0.05fF $ **FLOATING
C4452 S.n4043 SUB 1.88fF $ **FLOATING
C4453 S.n4044 SUB 2.67fF $ **FLOATING
C4454 S.t146 SUB 0.02fF
C4455 S.n4045 SUB 0.24fF $ **FLOATING
C4456 S.n4046 SUB 0.36fF $ **FLOATING
C4457 S.n4047 SUB 0.61fF $ **FLOATING
C4458 S.n4048 SUB 0.12fF $ **FLOATING
C4459 S.t1413 SUB 0.02fF
C4460 S.n4049 SUB 0.14fF $ **FLOATING
C4461 S.n4051 SUB 1.88fF $ **FLOATING
C4462 S.n4052 SUB 2.68fF $ **FLOATING
C4463 S.t1470 SUB 0.02fF
C4464 S.n4053 SUB 0.24fF $ **FLOATING
C4465 S.n4054 SUB 0.36fF $ **FLOATING
C4466 S.n4055 SUB 0.61fF $ **FLOATING
C4467 S.t667 SUB 0.02fF
C4468 S.n4056 SUB 1.22fF $ **FLOATING
C4469 S.n4057 SUB 0.36fF $ **FLOATING
C4470 S.n4058 SUB 1.22fF $ **FLOATING
C4471 S.n4059 SUB 0.61fF $ **FLOATING
C4472 S.n4060 SUB 0.35fF $ **FLOATING
C4473 S.n4061 SUB 0.63fF $ **FLOATING
C4474 S.n4062 SUB 1.15fF $ **FLOATING
C4475 S.n4063 SUB 3.03fF $ **FLOATING
C4476 S.n4064 SUB 0.59fF $ **FLOATING
C4477 S.n4065 SUB 0.02fF $ **FLOATING
C4478 S.n4066 SUB 0.97fF $ **FLOATING
C4479 S.t522 SUB 21.38fF
C4480 S.n4067 SUB 20.25fF $ **FLOATING
C4481 S.n4069 SUB 0.38fF $ **FLOATING
C4482 S.n4070 SUB 0.23fF $ **FLOATING
C4483 S.n4071 SUB 2.79fF $ **FLOATING
C4484 S.n4072 SUB 2.46fF $ **FLOATING
C4485 S.n4073 SUB 4.00fF $ **FLOATING
C4486 S.n4074 SUB 0.25fF $ **FLOATING
C4487 S.n4075 SUB 0.01fF $ **FLOATING
C4488 S.t380 SUB 0.02fF
C4489 S.n4076 SUB 0.25fF $ **FLOATING
C4490 S.t2349 SUB 0.02fF
C4491 S.n4077 SUB 0.95fF $ **FLOATING
C4492 S.n4078 SUB 0.70fF $ **FLOATING
C4493 S.n4079 SUB 1.89fF $ **FLOATING
C4494 S.n4080 SUB 1.88fF $ **FLOATING
C4495 S.t2321 SUB 0.02fF
C4496 S.n4081 SUB 0.24fF $ **FLOATING
C4497 S.n4082 SUB 0.36fF $ **FLOATING
C4498 S.n4083 SUB 0.61fF $ **FLOATING
C4499 S.n4084 SUB 0.12fF $ **FLOATING
C4500 S.t2029 SUB 0.02fF
C4501 S.n4085 SUB 0.14fF $ **FLOATING
C4502 S.n4087 SUB 1.16fF $ **FLOATING
C4503 S.n4088 SUB 0.22fF $ **FLOATING
C4504 S.n4089 SUB 0.25fF $ **FLOATING
C4505 S.n4090 SUB 0.09fF $ **FLOATING
C4506 S.n4091 SUB 1.88fF $ **FLOATING
C4507 S.t1490 SUB 0.02fF
C4508 S.n4092 SUB 0.24fF $ **FLOATING
C4509 S.n4093 SUB 0.91fF $ **FLOATING
C4510 S.n4094 SUB 0.05fF $ **FLOATING
C4511 S.t202 SUB 0.02fF
C4512 S.n4095 SUB 0.12fF $ **FLOATING
C4513 S.n4096 SUB 0.14fF $ **FLOATING
C4514 S.n4098 SUB 0.78fF $ **FLOATING
C4515 S.n4099 SUB 1.94fF $ **FLOATING
C4516 S.n4100 SUB 1.88fF $ **FLOATING
C4517 S.n4101 SUB 0.12fF $ **FLOATING
C4518 S.t1174 SUB 0.02fF
C4519 S.n4102 SUB 0.14fF $ **FLOATING
C4520 S.t1459 SUB 0.02fF
C4521 S.n4104 SUB 0.24fF $ **FLOATING
C4522 S.n4105 SUB 0.36fF $ **FLOATING
C4523 S.n4106 SUB 0.61fF $ **FLOATING
C4524 S.n4107 SUB 1.84fF $ **FLOATING
C4525 S.n4108 SUB 2.99fF $ **FLOATING
C4526 S.t625 SUB 0.02fF
C4527 S.n4109 SUB 0.24fF $ **FLOATING
C4528 S.n4110 SUB 0.91fF $ **FLOATING
C4529 S.n4111 SUB 0.05fF $ **FLOATING
C4530 S.t1869 SUB 0.02fF
C4531 S.n4112 SUB 0.12fF $ **FLOATING
C4532 S.n4113 SUB 0.14fF $ **FLOATING
C4533 S.n4115 SUB 1.89fF $ **FLOATING
C4534 S.n4116 SUB 1.88fF $ **FLOATING
C4535 S.t601 SUB 0.02fF
C4536 S.n4117 SUB 0.24fF $ **FLOATING
C4537 S.n4118 SUB 0.36fF $ **FLOATING
C4538 S.n4119 SUB 0.61fF $ **FLOATING
C4539 S.n4120 SUB 0.12fF $ **FLOATING
C4540 S.t298 SUB 0.02fF
C4541 S.n4121 SUB 0.14fF $ **FLOATING
C4542 S.n4123 SUB 1.16fF $ **FLOATING
C4543 S.n4124 SUB 0.22fF $ **FLOATING
C4544 S.n4125 SUB 0.25fF $ **FLOATING
C4545 S.n4126 SUB 0.09fF $ **FLOATING
C4546 S.n4127 SUB 1.88fF $ **FLOATING
C4547 S.t2284 SUB 0.02fF
C4548 S.n4128 SUB 0.24fF $ **FLOATING
C4549 S.n4129 SUB 0.91fF $ **FLOATING
C4550 S.n4130 SUB 0.05fF $ **FLOATING
C4551 S.t1121 SUB 0.02fF
C4552 S.n4131 SUB 0.12fF $ **FLOATING
C4553 S.n4132 SUB 0.14fF $ **FLOATING
C4554 S.n4134 SUB 0.78fF $ **FLOATING
C4555 S.n4135 SUB 1.94fF $ **FLOATING
C4556 S.n4136 SUB 1.88fF $ **FLOATING
C4557 S.n4137 SUB 0.12fF $ **FLOATING
C4558 S.t1961 SUB 0.02fF
C4559 S.n4138 SUB 0.14fF $ **FLOATING
C4560 S.t2254 SUB 0.02fF
C4561 S.n4140 SUB 0.24fF $ **FLOATING
C4562 S.n4141 SUB 0.36fF $ **FLOATING
C4563 S.n4142 SUB 0.61fF $ **FLOATING
C4564 S.n4143 SUB 1.84fF $ **FLOATING
C4565 S.n4144 SUB 2.99fF $ **FLOATING
C4566 S.t1430 SUB 0.02fF
C4567 S.n4145 SUB 0.24fF $ **FLOATING
C4568 S.n4146 SUB 0.91fF $ **FLOATING
C4569 S.n4147 SUB 0.05fF $ **FLOATING
C4570 S.t242 SUB 0.02fF
C4571 S.n4148 SUB 0.12fF $ **FLOATING
C4572 S.n4149 SUB 0.14fF $ **FLOATING
C4573 S.n4151 SUB 1.89fF $ **FLOATING
C4574 S.n4152 SUB 1.88fF $ **FLOATING
C4575 S.t1395 SUB 0.02fF
C4576 S.n4153 SUB 0.24fF $ **FLOATING
C4577 S.n4154 SUB 0.36fF $ **FLOATING
C4578 S.n4155 SUB 0.61fF $ **FLOATING
C4579 S.n4156 SUB 0.12fF $ **FLOATING
C4580 S.t1105 SUB 0.02fF
C4581 S.n4157 SUB 0.14fF $ **FLOATING
C4582 S.n4159 SUB 1.16fF $ **FLOATING
C4583 S.n4160 SUB 0.22fF $ **FLOATING
C4584 S.n4161 SUB 0.25fF $ **FLOATING
C4585 S.n4162 SUB 0.09fF $ **FLOATING
C4586 S.n4163 SUB 1.88fF $ **FLOATING
C4587 S.t565 SUB 0.02fF
C4588 S.n4164 SUB 0.24fF $ **FLOATING
C4589 S.n4165 SUB 0.91fF $ **FLOATING
C4590 S.n4166 SUB 0.05fF $ **FLOATING
C4591 S.t1908 SUB 0.02fF
C4592 S.n4167 SUB 0.12fF $ **FLOATING
C4593 S.n4168 SUB 0.14fF $ **FLOATING
C4594 S.n4170 SUB 0.78fF $ **FLOATING
C4595 S.n4171 SUB 1.94fF $ **FLOATING
C4596 S.n4172 SUB 1.88fF $ **FLOATING
C4597 S.n4173 SUB 0.12fF $ **FLOATING
C4598 S.t229 SUB 0.02fF
C4599 S.n4174 SUB 0.14fF $ **FLOATING
C4600 S.t523 SUB 0.02fF
C4601 S.n4176 SUB 0.24fF $ **FLOATING
C4602 S.n4177 SUB 0.36fF $ **FLOATING
C4603 S.n4178 SUB 0.61fF $ **FLOATING
C4604 S.n4179 SUB 1.84fF $ **FLOATING
C4605 S.n4180 SUB 2.99fF $ **FLOATING
C4606 S.t2208 SUB 0.02fF
C4607 S.n4181 SUB 0.24fF $ **FLOATING
C4608 S.n4182 SUB 0.91fF $ **FLOATING
C4609 S.n4183 SUB 0.05fF $ **FLOATING
C4610 S.t1048 SUB 0.02fF
C4611 S.n4184 SUB 0.12fF $ **FLOATING
C4612 S.n4185 SUB 0.14fF $ **FLOATING
C4613 S.n4187 SUB 1.89fF $ **FLOATING
C4614 S.n4188 SUB 1.88fF $ **FLOATING
C4615 S.t2167 SUB 0.02fF
C4616 S.n4189 SUB 0.24fF $ **FLOATING
C4617 S.n4190 SUB 0.36fF $ **FLOATING
C4618 S.n4191 SUB 0.61fF $ **FLOATING
C4619 S.n4192 SUB 0.12fF $ **FLOATING
C4620 S.t1993 SUB 0.02fF
C4621 S.n4193 SUB 0.14fF $ **FLOATING
C4622 S.n4195 SUB 1.16fF $ **FLOATING
C4623 S.n4196 SUB 0.22fF $ **FLOATING
C4624 S.n4197 SUB 0.25fF $ **FLOATING
C4625 S.n4198 SUB 0.09fF $ **FLOATING
C4626 S.n4199 SUB 1.88fF $ **FLOATING
C4627 S.t1347 SUB 0.02fF
C4628 S.n4200 SUB 0.24fF $ **FLOATING
C4629 S.n4201 SUB 0.91fF $ **FLOATING
C4630 S.n4202 SUB 0.05fF $ **FLOATING
C4631 S.t160 SUB 0.02fF
C4632 S.n4203 SUB 0.12fF $ **FLOATING
C4633 S.n4204 SUB 0.14fF $ **FLOATING
C4634 S.n4206 SUB 0.78fF $ **FLOATING
C4635 S.n4207 SUB 1.94fF $ **FLOATING
C4636 S.n4208 SUB 1.88fF $ **FLOATING
C4637 S.n4209 SUB 0.12fF $ **FLOATING
C4638 S.t1561 SUB 0.02fF
C4639 S.n4210 SUB 0.14fF $ **FLOATING
C4640 S.t827 SUB 0.02fF
C4641 S.n4212 SUB 0.24fF $ **FLOATING
C4642 S.n4213 SUB 0.36fF $ **FLOATING
C4643 S.n4214 SUB 0.61fF $ **FLOATING
C4644 S.n4215 SUB 1.84fF $ **FLOATING
C4645 S.n4216 SUB 2.99fF $ **FLOATING
C4646 S.t98 SUB 0.02fF
C4647 S.n4217 SUB 0.24fF $ **FLOATING
C4648 S.n4218 SUB 0.91fF $ **FLOATING
C4649 S.n4219 SUB 0.05fF $ **FLOATING
C4650 S.t1821 SUB 0.02fF
C4651 S.n4220 SUB 0.12fF $ **FLOATING
C4652 S.n4221 SUB 0.14fF $ **FLOATING
C4653 S.n4223 SUB 1.89fF $ **FLOATING
C4654 S.n4224 SUB 1.75fF $ **FLOATING
C4655 S.t2474 SUB 0.02fF
C4656 S.n4225 SUB 0.24fF $ **FLOATING
C4657 S.n4226 SUB 0.36fF $ **FLOATING
C4658 S.n4227 SUB 0.61fF $ **FLOATING
C4659 S.n4228 SUB 0.12fF $ **FLOATING
C4660 S.t698 SUB 0.02fF
C4661 S.n4229 SUB 0.14fF $ **FLOATING
C4662 S.n4231 SUB 1.16fF $ **FLOATING
C4663 S.n4232 SUB 0.22fF $ **FLOATING
C4664 S.n4233 SUB 0.25fF $ **FLOATING
C4665 S.n4234 SUB 0.09fF $ **FLOATING
C4666 S.n4235 SUB 2.44fF $ **FLOATING
C4667 S.t1774 SUB 0.02fF
C4668 S.n4236 SUB 0.24fF $ **FLOATING
C4669 S.n4237 SUB 0.91fF $ **FLOATING
C4670 S.n4238 SUB 0.05fF $ **FLOATING
C4671 S.t1412 SUB 0.02fF
C4672 S.n4239 SUB 0.12fF $ **FLOATING
C4673 S.n4240 SUB 0.14fF $ **FLOATING
C4674 S.n4242 SUB 1.88fF $ **FLOATING
C4675 S.n4243 SUB 0.48fF $ **FLOATING
C4676 S.n4244 SUB 0.09fF $ **FLOATING
C4677 S.n4245 SUB 0.33fF $ **FLOATING
C4678 S.n4246 SUB 0.30fF $ **FLOATING
C4679 S.n4247 SUB 0.77fF $ **FLOATING
C4680 S.n4248 SUB 0.59fF $ **FLOATING
C4681 S.t1603 SUB 0.02fF
C4682 S.n4249 SUB 0.24fF $ **FLOATING
C4683 S.n4250 SUB 0.36fF $ **FLOATING
C4684 S.n4251 SUB 0.61fF $ **FLOATING
C4685 S.n4252 SUB 0.12fF $ **FLOATING
C4686 S.t2357 SUB 0.02fF
C4687 S.n4253 SUB 0.14fF $ **FLOATING
C4688 S.n4255 SUB 2.61fF $ **FLOATING
C4689 S.n4256 SUB 2.16fF $ **FLOATING
C4690 S.t904 SUB 0.02fF
C4691 S.n4257 SUB 0.24fF $ **FLOATING
C4692 S.n4258 SUB 0.91fF $ **FLOATING
C4693 S.n4259 SUB 0.05fF $ **FLOATING
C4694 S.t547 SUB 0.02fF
C4695 S.n4260 SUB 0.12fF $ **FLOATING
C4696 S.n4261 SUB 0.14fF $ **FLOATING
C4697 S.n4263 SUB 0.78fF $ **FLOATING
C4698 S.n4264 SUB 2.30fF $ **FLOATING
C4699 S.n4265 SUB 1.88fF $ **FLOATING
C4700 S.n4266 SUB 0.12fF $ **FLOATING
C4701 S.t1499 SUB 0.02fF
C4702 S.n4267 SUB 0.14fF $ **FLOATING
C4703 S.t739 SUB 0.02fF
C4704 S.n4269 SUB 0.24fF $ **FLOATING
C4705 S.n4270 SUB 0.36fF $ **FLOATING
C4706 S.n4271 SUB 0.61fF $ **FLOATING
C4707 S.n4272 SUB 1.39fF $ **FLOATING
C4708 S.n4273 SUB 0.71fF $ **FLOATING
C4709 S.n4274 SUB 1.14fF $ **FLOATING
C4710 S.n4275 SUB 0.35fF $ **FLOATING
C4711 S.n4276 SUB 2.03fF $ **FLOATING
C4712 S.t2547 SUB 0.02fF
C4713 S.n4277 SUB 0.24fF $ **FLOATING
C4714 S.n4278 SUB 0.91fF $ **FLOATING
C4715 S.n4279 SUB 0.05fF $ **FLOATING
C4716 S.t2189 SUB 0.02fF
C4717 S.n4280 SUB 0.12fF $ **FLOATING
C4718 S.n4281 SUB 0.14fF $ **FLOATING
C4719 S.n4283 SUB 1.89fF $ **FLOATING
C4720 S.n4284 SUB 1.88fF $ **FLOATING
C4721 S.t2389 SUB 0.02fF
C4722 S.n4285 SUB 0.24fF $ **FLOATING
C4723 S.n4286 SUB 0.36fF $ **FLOATING
C4724 S.n4287 SUB 0.61fF $ **FLOATING
C4725 S.n4288 SUB 0.12fF $ **FLOATING
C4726 S.t636 SUB 0.02fF
C4727 S.n4289 SUB 0.14fF $ **FLOATING
C4728 S.n4291 SUB 1.16fF $ **FLOATING
C4729 S.n4292 SUB 0.22fF $ **FLOATING
C4730 S.n4293 SUB 0.25fF $ **FLOATING
C4731 S.n4294 SUB 0.09fF $ **FLOATING
C4732 S.n4295 SUB 1.88fF $ **FLOATING
C4733 S.t1674 SUB 0.02fF
C4734 S.n4296 SUB 0.24fF $ **FLOATING
C4735 S.n4297 SUB 0.91fF $ **FLOATING
C4736 S.n4298 SUB 0.05fF $ **FLOATING
C4737 S.t1327 SUB 0.02fF
C4738 S.n4299 SUB 0.12fF $ **FLOATING
C4739 S.n4300 SUB 0.14fF $ **FLOATING
C4740 S.n4302 SUB 20.78fF $ **FLOATING
C4741 S.n4303 SUB 1.88fF $ **FLOATING
C4742 S.n4304 SUB 2.67fF $ **FLOATING
C4743 S.t2329 SUB 0.02fF
C4744 S.n4305 SUB 0.24fF $ **FLOATING
C4745 S.n4306 SUB 0.36fF $ **FLOATING
C4746 S.n4307 SUB 0.61fF $ **FLOATING
C4747 S.n4308 SUB 0.12fF $ **FLOATING
C4748 S.t575 SUB 0.02fF
C4749 S.n4309 SUB 0.14fF $ **FLOATING
C4750 S.n4311 SUB 2.80fF $ **FLOATING
C4751 S.n4312 SUB 2.30fF $ **FLOATING
C4752 S.t1372 SUB 0.02fF
C4753 S.n4313 SUB 0.12fF $ **FLOATING
C4754 S.n4314 SUB 0.14fF $ **FLOATING
C4755 S.t1583 SUB 0.02fF
C4756 S.n4316 SUB 0.24fF $ **FLOATING
C4757 S.n4317 SUB 0.91fF $ **FLOATING
C4758 S.n4318 SUB 0.05fF $ **FLOATING
C4759 S.n4319 SUB 2.73fF $ **FLOATING
C4760 S.n4320 SUB 1.59fF $ **FLOATING
C4761 S.n4321 SUB 0.12fF $ **FLOATING
C4762 S.t1881 SUB 0.02fF
C4763 S.n4322 SUB 0.14fF $ **FLOATING
C4764 S.t1852 SUB 0.02fF
C4765 S.n4324 SUB 0.24fF $ **FLOATING
C4766 S.n4325 SUB 0.36fF $ **FLOATING
C4767 S.n4326 SUB 0.61fF $ **FLOATING
C4768 S.n4327 SUB 0.07fF $ **FLOATING
C4769 S.n4328 SUB 0.01fF $ **FLOATING
C4770 S.n4329 SUB 0.24fF $ **FLOATING
C4771 S.n4330 SUB 1.16fF $ **FLOATING
C4772 S.n4331 SUB 1.35fF $ **FLOATING
C4773 S.n4332 SUB 2.30fF $ **FLOATING
C4774 S.t52 SUB 0.02fF
C4775 S.n4333 SUB 0.12fF $ **FLOATING
C4776 S.n4334 SUB 0.14fF $ **FLOATING
C4777 S.t287 SUB 0.02fF
C4778 S.n4336 SUB 0.24fF $ **FLOATING
C4779 S.n4337 SUB 0.91fF $ **FLOATING
C4780 S.n4338 SUB 0.05fF $ **FLOATING
C4781 S.t51 SUB 48.31fF
C4782 S.t716 SUB 0.02fF
C4783 S.n4339 SUB 0.24fF $ **FLOATING
C4784 S.n4340 SUB 0.91fF $ **FLOATING
C4785 S.n4341 SUB 0.05fF $ **FLOATING
C4786 S.t502 SUB 0.02fF
C4787 S.n4342 SUB 0.12fF $ **FLOATING
C4788 S.n4343 SUB 0.14fF $ **FLOATING
C4789 S.n4345 SUB 0.12fF $ **FLOATING
C4790 S.t2220 SUB 0.02fF
C4791 S.n4346 SUB 0.14fF $ **FLOATING
C4792 S.n4348 SUB 5.17fF $ **FLOATING
C4793 S.n4349 SUB 5.44fF $ **FLOATING
C4794 S.t2119 SUB 0.02fF
C4795 S.n4350 SUB 0.12fF $ **FLOATING
C4796 S.n4351 SUB 0.14fF $ **FLOATING
C4797 S.t2073 SUB 0.02fF
C4798 S.n4353 SUB 0.24fF $ **FLOATING
C4799 S.n4354 SUB 0.91fF $ **FLOATING
C4800 S.n4355 SUB 0.05fF $ **FLOATING
C4801 S.t109 SUB 47.92fF
C4802 S.t2556 SUB 0.02fF
C4803 S.n4356 SUB 1.19fF $ **FLOATING
C4804 S.n4357 SUB 0.05fF $ **FLOATING
C4805 S.t643 SUB 0.02fF
C4806 S.n4358 SUB 0.01fF $ **FLOATING
C4807 S.n4359 SUB 0.26fF $ **FLOATING
C4808 S.n4361 SUB 1.50fF $ **FLOATING
C4809 S.n4362 SUB 1.30fF $ **FLOATING
C4810 S.n4363 SUB 0.28fF $ **FLOATING
C4811 S.n4364 SUB 0.24fF $ **FLOATING
C4812 S.n4365 SUB 4.39fF $ **FLOATING
C4813 S.n4366 SUB 0.01fF $ **FLOATING
C4814 S.n4367 SUB 0.02fF $ **FLOATING
C4815 S.n4368 SUB 0.03fF $ **FLOATING
C4816 S.n4369 SUB 0.04fF $ **FLOATING
C4817 S.n4370 SUB 0.17fF $ **FLOATING
C4818 S.n4371 SUB 0.01fF $ **FLOATING
C4819 S.n4372 SUB 0.02fF $ **FLOATING
C4820 S.n4373 SUB 0.01fF $ **FLOATING
C4821 S.n4374 SUB 0.01fF $ **FLOATING
C4822 S.n4375 SUB 0.01fF $ **FLOATING
C4823 S.n4376 SUB 0.01fF $ **FLOATING
C4824 S.n4377 SUB 0.02fF $ **FLOATING
C4825 S.n4378 SUB 0.01fF $ **FLOATING
C4826 S.n4379 SUB 0.02fF $ **FLOATING
C4827 S.n4380 SUB 0.05fF $ **FLOATING
C4828 S.n4381 SUB 0.04fF $ **FLOATING
C4829 S.n4382 SUB 0.11fF $ **FLOATING
C4830 S.n4383 SUB 0.38fF $ **FLOATING
C4831 S.n4384 SUB 0.20fF $ **FLOATING
C4832 S.n4385 SUB 8.97fF $ **FLOATING
C4833 S.n4386 SUB 8.97fF $ **FLOATING
C4834 S.n4387 SUB 0.60fF $ **FLOATING
C4835 S.n4388 SUB 0.22fF $ **FLOATING
C4836 S.n4389 SUB 0.59fF $ **FLOATING
C4837 S.n4390 SUB 3.43fF $ **FLOATING
C4838 S.n4391 SUB 0.29fF $ **FLOATING
C4839 S.t53 SUB 21.38fF
C4840 S.n4392 SUB 21.67fF $ **FLOATING
C4841 S.n4393 SUB 0.77fF $ **FLOATING
C4842 S.n4394 SUB 0.28fF $ **FLOATING
C4843 S.n4395 SUB 4.00fF $ **FLOATING
C4844 S.n4396 SUB 1.35fF $ **FLOATING
C4845 S.t152 SUB 0.02fF
C4846 S.n4397 SUB 0.64fF $ **FLOATING
C4847 S.n4398 SUB 0.61fF $ **FLOATING
C4848 S.n4399 SUB 0.25fF $ **FLOATING
C4849 S.n4400 SUB 0.09fF $ **FLOATING
C4850 S.n4401 SUB 0.21fF $ **FLOATING
C4851 S.n4402 SUB 0.92fF $ **FLOATING
C4852 S.n4403 SUB 0.44fF $ **FLOATING
C4853 S.n4404 SUB 1.88fF $ **FLOATING
C4854 S.n4405 SUB 0.12fF $ **FLOATING
C4855 S.t2374 SUB 0.02fF
C4856 S.n4406 SUB 0.14fF $ **FLOATING
C4857 S.t399 SUB 0.02fF
C4858 S.n4408 SUB 0.24fF $ **FLOATING
C4859 S.n4409 SUB 0.36fF $ **FLOATING
C4860 S.n4410 SUB 0.61fF $ **FLOATING
C4861 S.n4411 SUB 0.02fF $ **FLOATING
C4862 S.n4412 SUB 0.01fF $ **FLOATING
C4863 S.n4413 SUB 0.02fF $ **FLOATING
C4864 S.n4414 SUB 0.08fF $ **FLOATING
C4865 S.n4415 SUB 0.06fF $ **FLOATING
C4866 S.n4416 SUB 0.03fF $ **FLOATING
C4867 S.n4417 SUB 0.04fF $ **FLOATING
C4868 S.n4418 SUB 1.00fF $ **FLOATING
C4869 S.n4419 SUB 0.36fF $ **FLOATING
C4870 S.n4420 SUB 1.87fF $ **FLOATING
C4871 S.n4421 SUB 1.99fF $ **FLOATING
C4872 S.t1514 SUB 0.02fF
C4873 S.n4422 SUB 0.24fF $ **FLOATING
C4874 S.n4423 SUB 0.91fF $ **FLOATING
C4875 S.n4424 SUB 0.05fF $ **FLOATING
C4876 S.t2589 SUB 0.02fF
C4877 S.n4425 SUB 0.12fF $ **FLOATING
C4878 S.n4426 SUB 0.14fF $ **FLOATING
C4879 S.n4428 SUB 1.89fF $ **FLOATING
C4880 S.n4429 SUB 0.06fF $ **FLOATING
C4881 S.n4430 SUB 0.03fF $ **FLOATING
C4882 S.n4431 SUB 0.04fF $ **FLOATING
C4883 S.n4432 SUB 0.99fF $ **FLOATING
C4884 S.n4433 SUB 0.02fF $ **FLOATING
C4885 S.n4434 SUB 0.01fF $ **FLOATING
C4886 S.n4435 SUB 0.02fF $ **FLOATING
C4887 S.n4436 SUB 0.08fF $ **FLOATING
C4888 S.n4437 SUB 0.36fF $ **FLOATING
C4889 S.n4438 SUB 1.85fF $ **FLOATING
C4890 S.t2193 SUB 0.02fF
C4891 S.n4439 SUB 0.24fF $ **FLOATING
C4892 S.n4440 SUB 0.36fF $ **FLOATING
C4893 S.n4441 SUB 0.61fF $ **FLOATING
C4894 S.n4442 SUB 0.12fF $ **FLOATING
C4895 S.t1627 SUB 0.02fF
C4896 S.n4443 SUB 0.14fF $ **FLOATING
C4897 S.n4445 SUB 0.70fF $ **FLOATING
C4898 S.n4446 SUB 0.23fF $ **FLOATING
C4899 S.n4447 SUB 0.23fF $ **FLOATING
C4900 S.n4448 SUB 0.70fF $ **FLOATING
C4901 S.n4449 SUB 1.16fF $ **FLOATING
C4902 S.n4450 SUB 0.22fF $ **FLOATING
C4903 S.n4451 SUB 0.25fF $ **FLOATING
C4904 S.n4452 SUB 0.09fF $ **FLOATING
C4905 S.n4453 SUB 1.88fF $ **FLOATING
C4906 S.t757 SUB 0.02fF
C4907 S.n4454 SUB 0.24fF $ **FLOATING
C4908 S.n4455 SUB 0.91fF $ **FLOATING
C4909 S.n4456 SUB 0.05fF $ **FLOATING
C4910 S.t1713 SUB 0.02fF
C4911 S.n4457 SUB 0.12fF $ **FLOATING
C4912 S.n4458 SUB 0.14fF $ **FLOATING
C4913 S.n4460 SUB 0.25fF $ **FLOATING
C4914 S.n4461 SUB 0.09fF $ **FLOATING
C4915 S.n4462 SUB 0.21fF $ **FLOATING
C4916 S.n4463 SUB 0.92fF $ **FLOATING
C4917 S.n4464 SUB 0.44fF $ **FLOATING
C4918 S.n4465 SUB 1.88fF $ **FLOATING
C4919 S.n4466 SUB 0.12fF $ **FLOATING
C4920 S.t760 SUB 0.02fF
C4921 S.n4467 SUB 0.14fF $ **FLOATING
C4922 S.t1337 SUB 0.02fF
C4923 S.n4469 SUB 0.24fF $ **FLOATING
C4924 S.n4470 SUB 0.36fF $ **FLOATING
C4925 S.n4471 SUB 0.61fF $ **FLOATING
C4926 S.n4472 SUB 0.02fF $ **FLOATING
C4927 S.n4473 SUB 0.01fF $ **FLOATING
C4928 S.n4474 SUB 0.02fF $ **FLOATING
C4929 S.n4475 SUB 0.08fF $ **FLOATING
C4930 S.n4476 SUB 0.06fF $ **FLOATING
C4931 S.n4477 SUB 0.03fF $ **FLOATING
C4932 S.n4478 SUB 0.04fF $ **FLOATING
C4933 S.n4479 SUB 1.00fF $ **FLOATING
C4934 S.n4480 SUB 0.36fF $ **FLOATING
C4935 S.n4481 SUB 1.87fF $ **FLOATING
C4936 S.n4482 SUB 1.99fF $ **FLOATING
C4937 S.t2411 SUB 0.02fF
C4938 S.n4483 SUB 0.24fF $ **FLOATING
C4939 S.n4484 SUB 0.91fF $ **FLOATING
C4940 S.n4485 SUB 0.05fF $ **FLOATING
C4941 S.t844 SUB 0.02fF
C4942 S.n4486 SUB 0.12fF $ **FLOATING
C4943 S.n4487 SUB 0.14fF $ **FLOATING
C4944 S.n4489 SUB 1.89fF $ **FLOATING
C4945 S.n4490 SUB 0.06fF $ **FLOATING
C4946 S.n4491 SUB 0.03fF $ **FLOATING
C4947 S.n4492 SUB 0.04fF $ **FLOATING
C4948 S.n4493 SUB 0.99fF $ **FLOATING
C4949 S.n4494 SUB 0.02fF $ **FLOATING
C4950 S.n4495 SUB 0.01fF $ **FLOATING
C4951 S.n4496 SUB 0.02fF $ **FLOATING
C4952 S.n4497 SUB 0.08fF $ **FLOATING
C4953 S.n4498 SUB 0.36fF $ **FLOATING
C4954 S.n4499 SUB 1.85fF $ **FLOATING
C4955 S.t457 SUB 0.02fF
C4956 S.n4500 SUB 0.24fF $ **FLOATING
C4957 S.n4501 SUB 0.36fF $ **FLOATING
C4958 S.n4502 SUB 0.61fF $ **FLOATING
C4959 S.n4503 SUB 0.12fF $ **FLOATING
C4960 S.t2413 SUB 0.02fF
C4961 S.n4504 SUB 0.14fF $ **FLOATING
C4962 S.n4506 SUB 0.70fF $ **FLOATING
C4963 S.n4507 SUB 0.23fF $ **FLOATING
C4964 S.n4508 SUB 0.23fF $ **FLOATING
C4965 S.n4509 SUB 0.70fF $ **FLOATING
C4966 S.n4510 SUB 1.16fF $ **FLOATING
C4967 S.n4511 SUB 0.22fF $ **FLOATING
C4968 S.n4512 SUB 0.25fF $ **FLOATING
C4969 S.n4513 SUB 0.09fF $ **FLOATING
C4970 S.n4514 SUB 1.88fF $ **FLOATING
C4971 S.t1547 SUB 0.02fF
C4972 S.n4515 SUB 0.24fF $ **FLOATING
C4973 S.n4516 SUB 0.91fF $ **FLOATING
C4974 S.n4517 SUB 0.05fF $ **FLOATING
C4975 S.t2488 SUB 0.02fF
C4976 S.n4518 SUB 0.12fF $ **FLOATING
C4977 S.n4519 SUB 0.14fF $ **FLOATING
C4978 S.n4521 SUB 0.25fF $ **FLOATING
C4979 S.n4522 SUB 0.09fF $ **FLOATING
C4980 S.n4523 SUB 0.21fF $ **FLOATING
C4981 S.n4524 SUB 0.92fF $ **FLOATING
C4982 S.n4525 SUB 0.44fF $ **FLOATING
C4983 S.n4526 SUB 1.88fF $ **FLOATING
C4984 S.n4527 SUB 0.12fF $ **FLOATING
C4985 S.t1549 SUB 0.02fF
C4986 S.n4528 SUB 0.14fF $ **FLOATING
C4987 S.t2103 SUB 0.02fF
C4988 S.n4530 SUB 0.24fF $ **FLOATING
C4989 S.n4531 SUB 0.36fF $ **FLOATING
C4990 S.n4532 SUB 0.61fF $ **FLOATING
C4991 S.n4533 SUB 0.02fF $ **FLOATING
C4992 S.n4534 SUB 0.01fF $ **FLOATING
C4993 S.n4535 SUB 0.02fF $ **FLOATING
C4994 S.n4536 SUB 0.08fF $ **FLOATING
C4995 S.n4537 SUB 0.06fF $ **FLOATING
C4996 S.n4538 SUB 0.03fF $ **FLOATING
C4997 S.n4539 SUB 0.04fF $ **FLOATING
C4998 S.n4540 SUB 1.00fF $ **FLOATING
C4999 S.n4541 SUB 0.36fF $ **FLOATING
C5000 S.n4542 SUB 1.87fF $ **FLOATING
C5001 S.n4543 SUB 1.99fF $ **FLOATING
C5002 S.t685 SUB 0.02fF
C5003 S.n4544 SUB 0.24fF $ **FLOATING
C5004 S.n4545 SUB 0.91fF $ **FLOATING
C5005 S.n4546 SUB 0.05fF $ **FLOATING
C5006 S.t1612 SUB 0.02fF
C5007 S.n4547 SUB 0.12fF $ **FLOATING
C5008 S.n4548 SUB 0.14fF $ **FLOATING
C5009 S.n4550 SUB 1.89fF $ **FLOATING
C5010 S.n4551 SUB 0.06fF $ **FLOATING
C5011 S.n4552 SUB 0.03fF $ **FLOATING
C5012 S.n4553 SUB 0.04fF $ **FLOATING
C5013 S.n4554 SUB 0.99fF $ **FLOATING
C5014 S.n4555 SUB 0.02fF $ **FLOATING
C5015 S.n4556 SUB 0.01fF $ **FLOATING
C5016 S.n4557 SUB 0.02fF $ **FLOATING
C5017 S.n4558 SUB 0.08fF $ **FLOATING
C5018 S.n4559 SUB 0.36fF $ **FLOATING
C5019 S.n4560 SUB 1.85fF $ **FLOATING
C5020 S.t1237 SUB 0.02fF
C5021 S.n4561 SUB 0.24fF $ **FLOATING
C5022 S.n4562 SUB 0.36fF $ **FLOATING
C5023 S.n4563 SUB 0.61fF $ **FLOATING
C5024 S.n4564 SUB 0.12fF $ **FLOATING
C5025 S.t687 SUB 0.02fF
C5026 S.n4565 SUB 0.14fF $ **FLOATING
C5027 S.n4567 SUB 0.70fF $ **FLOATING
C5028 S.n4568 SUB 0.23fF $ **FLOATING
C5029 S.n4569 SUB 0.23fF $ **FLOATING
C5030 S.n4570 SUB 0.70fF $ **FLOATING
C5031 S.n4571 SUB 1.16fF $ **FLOATING
C5032 S.n4572 SUB 0.22fF $ **FLOATING
C5033 S.n4573 SUB 0.25fF $ **FLOATING
C5034 S.n4574 SUB 0.09fF $ **FLOATING
C5035 S.n4575 SUB 1.88fF $ **FLOATING
C5036 S.t2343 SUB 0.02fF
C5037 S.n4576 SUB 0.24fF $ **FLOATING
C5038 S.n4577 SUB 0.91fF $ **FLOATING
C5039 S.n4578 SUB 0.05fF $ **FLOATING
C5040 S.t748 SUB 0.02fF
C5041 S.n4579 SUB 0.12fF $ **FLOATING
C5042 S.n4580 SUB 0.14fF $ **FLOATING
C5043 S.n4582 SUB 0.25fF $ **FLOATING
C5044 S.n4583 SUB 0.09fF $ **FLOATING
C5045 S.n4584 SUB 0.21fF $ **FLOATING
C5046 S.n4585 SUB 0.92fF $ **FLOATING
C5047 S.n4586 SUB 0.44fF $ **FLOATING
C5048 S.n4587 SUB 1.88fF $ **FLOATING
C5049 S.n4588 SUB 0.12fF $ **FLOATING
C5050 S.t2346 SUB 0.02fF
C5051 S.n4589 SUB 0.14fF $ **FLOATING
C5052 S.t354 SUB 0.02fF
C5053 S.n4591 SUB 0.24fF $ **FLOATING
C5054 S.n4592 SUB 0.36fF $ **FLOATING
C5055 S.n4593 SUB 0.61fF $ **FLOATING
C5056 S.n4594 SUB 0.02fF $ **FLOATING
C5057 S.n4595 SUB 0.01fF $ **FLOATING
C5058 S.n4596 SUB 0.02fF $ **FLOATING
C5059 S.n4597 SUB 0.08fF $ **FLOATING
C5060 S.n4598 SUB 0.06fF $ **FLOATING
C5061 S.n4599 SUB 0.03fF $ **FLOATING
C5062 S.n4600 SUB 0.04fF $ **FLOATING
C5063 S.n4601 SUB 1.00fF $ **FLOATING
C5064 S.n4602 SUB 0.36fF $ **FLOATING
C5065 S.n4603 SUB 1.87fF $ **FLOATING
C5066 S.n4604 SUB 1.99fF $ **FLOATING
C5067 S.t1487 SUB 0.02fF
C5068 S.n4605 SUB 0.24fF $ **FLOATING
C5069 S.n4606 SUB 0.91fF $ **FLOATING
C5070 S.n4607 SUB 0.05fF $ **FLOATING
C5071 S.t2540 SUB 0.02fF
C5072 S.n4608 SUB 0.12fF $ **FLOATING
C5073 S.n4609 SUB 0.14fF $ **FLOATING
C5074 S.n4611 SUB 1.89fF $ **FLOATING
C5075 S.n4612 SUB 0.07fF $ **FLOATING
C5076 S.n4613 SUB 0.04fF $ **FLOATING
C5077 S.n4614 SUB 0.05fF $ **FLOATING
C5078 S.n4615 SUB 0.87fF $ **FLOATING
C5079 S.n4616 SUB 0.01fF $ **FLOATING
C5080 S.n4617 SUB 0.01fF $ **FLOATING
C5081 S.n4618 SUB 0.01fF $ **FLOATING
C5082 S.n4619 SUB 0.07fF $ **FLOATING
C5083 S.n4620 SUB 0.68fF $ **FLOATING
C5084 S.n4621 SUB 0.72fF $ **FLOATING
C5085 S.t1019 SUB 0.02fF
C5086 S.n4622 SUB 0.24fF $ **FLOATING
C5087 S.n4623 SUB 0.36fF $ **FLOATING
C5088 S.n4624 SUB 0.61fF $ **FLOATING
C5089 S.n4625 SUB 0.12fF $ **FLOATING
C5090 S.t463 SUB 0.02fF
C5091 S.n4626 SUB 0.14fF $ **FLOATING
C5092 S.n4628 SUB 0.70fF $ **FLOATING
C5093 S.n4629 SUB 0.23fF $ **FLOATING
C5094 S.n4630 SUB 0.23fF $ **FLOATING
C5095 S.n4631 SUB 0.70fF $ **FLOATING
C5096 S.n4632 SUB 1.16fF $ **FLOATING
C5097 S.n4633 SUB 0.22fF $ **FLOATING
C5098 S.n4634 SUB 0.25fF $ **FLOATING
C5099 S.n4635 SUB 0.09fF $ **FLOATING
C5100 S.n4636 SUB 2.31fF $ **FLOATING
C5101 S.t2558 SUB 0.02fF
C5102 S.n4637 SUB 0.24fF $ **FLOATING
C5103 S.n4638 SUB 0.91fF $ **FLOATING
C5104 S.n4639 SUB 0.05fF $ **FLOATING
C5105 S.t646 SUB 0.02fF
C5106 S.n4640 SUB 0.12fF $ **FLOATING
C5107 S.n4641 SUB 0.14fF $ **FLOATING
C5108 S.n4643 SUB 1.88fF $ **FLOATING
C5109 S.n4644 SUB 0.46fF $ **FLOATING
C5110 S.n4645 SUB 0.22fF $ **FLOATING
C5111 S.n4646 SUB 0.38fF $ **FLOATING
C5112 S.n4647 SUB 0.16fF $ **FLOATING
C5113 S.n4648 SUB 0.28fF $ **FLOATING
C5114 S.n4649 SUB 0.21fF $ **FLOATING
C5115 S.n4650 SUB 0.30fF $ **FLOATING
C5116 S.n4651 SUB 0.42fF $ **FLOATING
C5117 S.n4652 SUB 0.21fF $ **FLOATING
C5118 S.t113 SUB 0.02fF
C5119 S.n4653 SUB 0.24fF $ **FLOATING
C5120 S.n4654 SUB 0.36fF $ **FLOATING
C5121 S.n4655 SUB 0.61fF $ **FLOATING
C5122 S.n4656 SUB 0.12fF $ **FLOATING
C5123 S.t2108 SUB 0.02fF
C5124 S.n4657 SUB 0.14fF $ **FLOATING
C5125 S.n4659 SUB 0.04fF $ **FLOATING
C5126 S.n4660 SUB 0.03fF $ **FLOATING
C5127 S.n4661 SUB 0.03fF $ **FLOATING
C5128 S.n4662 SUB 0.10fF $ **FLOATING
C5129 S.n4663 SUB 0.36fF $ **FLOATING
C5130 S.n4664 SUB 0.38fF $ **FLOATING
C5131 S.n4665 SUB 0.11fF $ **FLOATING
C5132 S.n4666 SUB 0.12fF $ **FLOATING
C5133 S.n4667 SUB 0.07fF $ **FLOATING
C5134 S.n4668 SUB 0.12fF $ **FLOATING
C5135 S.n4669 SUB 0.18fF $ **FLOATING
C5136 S.n4670 SUB 4.00fF $ **FLOATING
C5137 S.t1685 SUB 0.02fF
C5138 S.n4671 SUB 0.24fF $ **FLOATING
C5139 S.n4672 SUB 0.91fF $ **FLOATING
C5140 S.n4673 SUB 0.05fF $ **FLOATING
C5141 S.t2303 SUB 0.02fF
C5142 S.n4674 SUB 0.12fF $ **FLOATING
C5143 S.n4675 SUB 0.14fF $ **FLOATING
C5144 S.n4677 SUB 0.25fF $ **FLOATING
C5145 S.n4678 SUB 0.09fF $ **FLOATING
C5146 S.n4679 SUB 0.21fF $ **FLOATING
C5147 S.n4680 SUB 1.28fF $ **FLOATING
C5148 S.n4681 SUB 0.53fF $ **FLOATING
C5149 S.n4682 SUB 1.88fF $ **FLOATING
C5150 S.n4683 SUB 0.12fF $ **FLOATING
C5151 S.t1243 SUB 0.02fF
C5152 S.n4684 SUB 0.14fF $ **FLOATING
C5153 S.t1787 SUB 0.02fF
C5154 S.n4686 SUB 0.24fF $ **FLOATING
C5155 S.n4687 SUB 0.36fF $ **FLOATING
C5156 S.n4688 SUB 0.61fF $ **FLOATING
C5157 S.n4689 SUB 1.58fF $ **FLOATING
C5158 S.n4690 SUB 2.45fF $ **FLOATING
C5159 S.t811 SUB 0.02fF
C5160 S.n4691 SUB 0.24fF $ **FLOATING
C5161 S.n4692 SUB 0.91fF $ **FLOATING
C5162 S.n4693 SUB 0.05fF $ **FLOATING
C5163 S.t1448 SUB 0.02fF
C5164 S.n4694 SUB 0.12fF $ **FLOATING
C5165 S.n4695 SUB 0.14fF $ **FLOATING
C5166 S.n4697 SUB 1.89fF $ **FLOATING
C5167 S.n4698 SUB 0.06fF $ **FLOATING
C5168 S.n4699 SUB 0.03fF $ **FLOATING
C5169 S.n4700 SUB 0.04fF $ **FLOATING
C5170 S.n4701 SUB 0.99fF $ **FLOATING
C5171 S.n4702 SUB 0.02fF $ **FLOATING
C5172 S.n4703 SUB 0.01fF $ **FLOATING
C5173 S.n4704 SUB 0.02fF $ **FLOATING
C5174 S.n4705 SUB 0.08fF $ **FLOATING
C5175 S.n4706 SUB 0.36fF $ **FLOATING
C5176 S.n4707 SUB 1.85fF $ **FLOATING
C5177 S.t918 SUB 0.02fF
C5178 S.n4708 SUB 0.24fF $ **FLOATING
C5179 S.n4709 SUB 0.36fF $ **FLOATING
C5180 S.n4710 SUB 0.61fF $ **FLOATING
C5181 S.n4711 SUB 0.12fF $ **FLOATING
C5182 S.t361 SUB 0.02fF
C5183 S.n4712 SUB 0.14fF $ **FLOATING
C5184 S.n4714 SUB 0.70fF $ **FLOATING
C5185 S.n4715 SUB 0.23fF $ **FLOATING
C5186 S.n4716 SUB 0.23fF $ **FLOATING
C5187 S.n4717 SUB 0.70fF $ **FLOATING
C5188 S.n4718 SUB 1.16fF $ **FLOATING
C5189 S.n4719 SUB 0.22fF $ **FLOATING
C5190 S.n4720 SUB 0.25fF $ **FLOATING
C5191 S.n4721 SUB 0.09fF $ **FLOATING
C5192 S.n4722 SUB 1.88fF $ **FLOATING
C5193 S.t2459 SUB 0.02fF
C5194 S.n4723 SUB 0.24fF $ **FLOATING
C5195 S.n4724 SUB 0.91fF $ **FLOATING
C5196 S.n4725 SUB 0.05fF $ **FLOATING
C5197 S.t585 SUB 0.02fF
C5198 S.n4726 SUB 0.12fF $ **FLOATING
C5199 S.n4727 SUB 0.14fF $ **FLOATING
C5200 S.n4729 SUB 20.78fF $ **FLOATING
C5201 S.n4730 SUB 1.72fF $ **FLOATING
C5202 S.n4731 SUB 3.05fF $ **FLOATING
C5203 S.t1284 SUB 0.02fF
C5204 S.n4732 SUB 0.24fF $ **FLOATING
C5205 S.n4733 SUB 0.36fF $ **FLOATING
C5206 S.n4734 SUB 0.61fF $ **FLOATING
C5207 S.n4735 SUB 0.12fF $ **FLOATING
C5208 S.t719 SUB 0.02fF
C5209 S.n4736 SUB 0.14fF $ **FLOATING
C5210 S.n4738 SUB 0.31fF $ **FLOATING
C5211 S.n4739 SUB 0.23fF $ **FLOATING
C5212 S.n4740 SUB 0.66fF $ **FLOATING
C5213 S.n4741 SUB 0.95fF $ **FLOATING
C5214 S.n4742 SUB 0.23fF $ **FLOATING
C5215 S.n4743 SUB 0.21fF $ **FLOATING
C5216 S.n4744 SUB 0.20fF $ **FLOATING
C5217 S.n4745 SUB 0.06fF $ **FLOATING
C5218 S.n4746 SUB 0.09fF $ **FLOATING
C5219 S.n4747 SUB 0.10fF $ **FLOATING
C5220 S.n4748 SUB 1.99fF $ **FLOATING
C5221 S.t951 SUB 0.02fF
C5222 S.n4749 SUB 0.12fF $ **FLOATING
C5223 S.n4750 SUB 0.14fF $ **FLOATING
C5224 S.t2371 SUB 0.02fF
C5225 S.n4752 SUB 0.24fF $ **FLOATING
C5226 S.n4753 SUB 0.91fF $ **FLOATING
C5227 S.n4754 SUB 0.05fF $ **FLOATING
C5228 S.n4755 SUB 1.88fF $ **FLOATING
C5229 S.n4756 SUB 0.12fF $ **FLOATING
C5230 S.t2312 SUB 0.02fF
C5231 S.n4757 SUB 0.14fF $ **FLOATING
C5232 S.t477 SUB 0.02fF
C5233 S.n4759 SUB 0.12fF $ **FLOATING
C5234 S.n4760 SUB 0.14fF $ **FLOATING
C5235 S.t830 SUB 0.02fF
C5236 S.n4762 SUB 0.24fF $ **FLOATING
C5237 S.n4763 SUB 0.91fF $ **FLOATING
C5238 S.n4764 SUB 0.05fF $ **FLOATING
C5239 S.t1551 SUB 0.02fF
C5240 S.n4765 SUB 0.24fF $ **FLOATING
C5241 S.n4766 SUB 0.36fF $ **FLOATING
C5242 S.n4767 SUB 0.61fF $ **FLOATING
C5243 S.n4768 SUB 0.32fF $ **FLOATING
C5244 S.n4769 SUB 1.09fF $ **FLOATING
C5245 S.n4770 SUB 0.15fF $ **FLOATING
C5246 S.n4771 SUB 2.10fF $ **FLOATING
C5247 S.n4772 SUB 2.94fF $ **FLOATING
C5248 S.n4773 SUB 1.88fF $ **FLOATING
C5249 S.n4774 SUB 0.12fF $ **FLOATING
C5250 S.t2159 SUB 0.02fF
C5251 S.n4775 SUB 0.14fF $ **FLOATING
C5252 S.t179 SUB 0.02fF
C5253 S.n4777 SUB 0.24fF $ **FLOATING
C5254 S.n4778 SUB 0.36fF $ **FLOATING
C5255 S.n4779 SUB 0.61fF $ **FLOATING
C5256 S.n4780 SUB 0.92fF $ **FLOATING
C5257 S.n4781 SUB 0.32fF $ **FLOATING
C5258 S.n4782 SUB 0.92fF $ **FLOATING
C5259 S.n4783 SUB 1.09fF $ **FLOATING
C5260 S.n4784 SUB 0.15fF $ **FLOATING
C5261 S.n4785 SUB 4.96fF $ **FLOATING
C5262 S.t2232 SUB 0.02fF
C5263 S.n4786 SUB 0.12fF $ **FLOATING
C5264 S.n4787 SUB 0.14fF $ **FLOATING
C5265 S.t1740 SUB 0.02fF
C5266 S.n4789 SUB 0.24fF $ **FLOATING
C5267 S.n4790 SUB 0.91fF $ **FLOATING
C5268 S.n4791 SUB 0.05fF $ **FLOATING
C5269 S.n4792 SUB 1.88fF $ **FLOATING
C5270 S.n4793 SUB 2.67fF $ **FLOATING
C5271 S.t1844 SUB 0.02fF
C5272 S.n4794 SUB 0.24fF $ **FLOATING
C5273 S.n4795 SUB 0.36fF $ **FLOATING
C5274 S.n4796 SUB 0.61fF $ **FLOATING
C5275 S.n4797 SUB 0.12fF $ **FLOATING
C5276 S.t1296 SUB 0.02fF
C5277 S.n4798 SUB 0.14fF $ **FLOATING
C5278 S.n4800 SUB 1.88fF $ **FLOATING
C5279 S.n4801 SUB 2.67fF $ **FLOATING
C5280 S.t689 SUB 0.02fF
C5281 S.n4802 SUB 0.24fF $ **FLOATING
C5282 S.n4803 SUB 0.36fF $ **FLOATING
C5283 S.n4804 SUB 0.61fF $ **FLOATING
C5284 S.t2475 SUB 0.02fF
C5285 S.n4805 SUB 0.24fF $ **FLOATING
C5286 S.n4806 SUB 0.91fF $ **FLOATING
C5287 S.n4807 SUB 0.05fF $ **FLOATING
C5288 S.t2259 SUB 0.02fF
C5289 S.n4808 SUB 0.12fF $ **FLOATING
C5290 S.n4809 SUB 0.14fF $ **FLOATING
C5291 S.n4811 SUB 0.12fF $ **FLOATING
C5292 S.t1454 SUB 0.02fF
C5293 S.n4812 SUB 0.14fF $ **FLOATING
C5294 S.n4814 SUB 2.30fF $ **FLOATING
C5295 S.n4815 SUB 2.94fF $ **FLOATING
C5296 S.n4816 SUB 5.16fF $ **FLOATING
C5297 S.t1370 SUB 0.02fF
C5298 S.n4817 SUB 0.12fF $ **FLOATING
C5299 S.n4818 SUB 0.14fF $ **FLOATING
C5300 S.t866 SUB 0.02fF
C5301 S.n4820 SUB 0.24fF $ **FLOATING
C5302 S.n4821 SUB 0.91fF $ **FLOATING
C5303 S.n4822 SUB 0.05fF $ **FLOATING
C5304 S.n4823 SUB 1.88fF $ **FLOATING
C5305 S.n4824 SUB 2.67fF $ **FLOATING
C5306 S.t980 SUB 0.02fF
C5307 S.n4825 SUB 0.24fF $ **FLOATING
C5308 S.n4826 SUB 0.36fF $ **FLOATING
C5309 S.n4827 SUB 0.61fF $ **FLOATING
C5310 S.n4828 SUB 0.12fF $ **FLOATING
C5311 S.t412 SUB 0.02fF
C5312 S.n4829 SUB 0.14fF $ **FLOATING
C5313 S.n4831 SUB 5.17fF $ **FLOATING
C5314 S.t497 SUB 0.02fF
C5315 S.n4832 SUB 0.12fF $ **FLOATING
C5316 S.n4833 SUB 0.14fF $ **FLOATING
C5317 S.t2511 SUB 0.02fF
C5318 S.n4835 SUB 0.24fF $ **FLOATING
C5319 S.n4836 SUB 0.91fF $ **FLOATING
C5320 S.n4837 SUB 0.05fF $ **FLOATING
C5321 S.n4838 SUB 1.88fF $ **FLOATING
C5322 S.n4839 SUB 2.67fF $ **FLOATING
C5323 S.t54 SUB 0.02fF
C5324 S.n4840 SUB 0.24fF $ **FLOATING
C5325 S.n4841 SUB 0.36fF $ **FLOATING
C5326 S.n4842 SUB 0.61fF $ **FLOATING
C5327 S.n4843 SUB 0.12fF $ **FLOATING
C5328 S.t2060 SUB 0.02fF
C5329 S.n4844 SUB 0.14fF $ **FLOATING
C5330 S.n4846 SUB 4.90fF $ **FLOATING
C5331 S.t2145 SUB 0.02fF
C5332 S.n4847 SUB 0.12fF $ **FLOATING
C5333 S.n4848 SUB 0.14fF $ **FLOATING
C5334 S.t1634 SUB 0.02fF
C5335 S.n4850 SUB 0.24fF $ **FLOATING
C5336 S.n4851 SUB 0.91fF $ **FLOATING
C5337 S.n4852 SUB 0.05fF $ **FLOATING
C5338 S.n4853 SUB 1.88fF $ **FLOATING
C5339 S.n4854 SUB 2.67fF $ **FLOATING
C5340 S.t1314 SUB 0.02fF
C5341 S.n4855 SUB 0.24fF $ **FLOATING
C5342 S.n4856 SUB 0.36fF $ **FLOATING
C5343 S.n4857 SUB 0.61fF $ **FLOATING
C5344 S.n4858 SUB 0.12fF $ **FLOATING
C5345 S.t2532 SUB 0.02fF
C5346 S.n4859 SUB 0.14fF $ **FLOATING
C5347 S.n4861 SUB 1.88fF $ **FLOATING
C5348 S.n4862 SUB 2.68fF $ **FLOATING
C5349 S.t628 SUB 0.02fF
C5350 S.n4863 SUB 0.24fF $ **FLOATING
C5351 S.n4864 SUB 0.36fF $ **FLOATING
C5352 S.n4865 SUB 0.61fF $ **FLOATING
C5353 S.t376 SUB 0.02fF
C5354 S.n4866 SUB 1.22fF $ **FLOATING
C5355 S.n4867 SUB 0.61fF $ **FLOATING
C5356 S.n4868 SUB 0.35fF $ **FLOATING
C5357 S.n4869 SUB 0.63fF $ **FLOATING
C5358 S.n4870 SUB 1.15fF $ **FLOATING
C5359 S.n4871 SUB 3.03fF $ **FLOATING
C5360 S.n4872 SUB 0.59fF $ **FLOATING
C5361 S.n4873 SUB 0.02fF $ **FLOATING
C5362 S.n4874 SUB 0.97fF $ **FLOATING
C5363 S.t226 SUB 21.38fF
C5364 S.n4875 SUB 20.25fF $ **FLOATING
C5365 S.n4877 SUB 0.38fF $ **FLOATING
C5366 S.n4878 SUB 0.23fF $ **FLOATING
C5367 S.n4879 SUB 2.90fF $ **FLOATING
C5368 S.n4880 SUB 2.46fF $ **FLOATING
C5369 S.n4881 SUB 1.96fF $ **FLOATING
C5370 S.n4882 SUB 3.94fF $ **FLOATING
C5371 S.n4883 SUB 0.25fF $ **FLOATING
C5372 S.n4884 SUB 0.01fF $ **FLOATING
C5373 S.t82 SUB 0.02fF
C5374 S.n4885 SUB 0.25fF $ **FLOATING
C5375 S.t2065 SUB 0.02fF
C5376 S.n4886 SUB 0.95fF $ **FLOATING
C5377 S.n4887 SUB 0.70fF $ **FLOATING
C5378 S.n4888 SUB 0.78fF $ **FLOATING
C5379 S.n4889 SUB 1.93fF $ **FLOATING
C5380 S.n4890 SUB 1.88fF $ **FLOATING
C5381 S.n4891 SUB 0.12fF $ **FLOATING
C5382 S.t1759 SUB 0.02fF
C5383 S.n4892 SUB 0.14fF $ **FLOATING
C5384 S.t2027 SUB 0.02fF
C5385 S.n4894 SUB 0.24fF $ **FLOATING
C5386 S.n4895 SUB 0.36fF $ **FLOATING
C5387 S.n4896 SUB 0.61fF $ **FLOATING
C5388 S.n4897 SUB 1.52fF $ **FLOATING
C5389 S.n4898 SUB 2.99fF $ **FLOATING
C5390 S.t1203 SUB 0.02fF
C5391 S.n4899 SUB 0.24fF $ **FLOATING
C5392 S.n4900 SUB 0.91fF $ **FLOATING
C5393 S.n4901 SUB 0.05fF $ **FLOATING
C5394 S.t2404 SUB 0.02fF
C5395 S.n4902 SUB 0.12fF $ **FLOATING
C5396 S.n4903 SUB 0.14fF $ **FLOATING
C5397 S.n4905 SUB 1.89fF $ **FLOATING
C5398 S.n4906 SUB 1.88fF $ **FLOATING
C5399 S.t1171 SUB 0.02fF
C5400 S.n4907 SUB 0.24fF $ **FLOATING
C5401 S.n4908 SUB 0.36fF $ **FLOATING
C5402 S.n4909 SUB 0.61fF $ **FLOATING
C5403 S.n4910 SUB 0.12fF $ **FLOATING
C5404 S.t882 SUB 0.02fF
C5405 S.n4911 SUB 0.14fF $ **FLOATING
C5406 S.n4913 SUB 1.16fF $ **FLOATING
C5407 S.n4914 SUB 0.22fF $ **FLOATING
C5408 S.n4915 SUB 0.25fF $ **FLOATING
C5409 S.n4916 SUB 0.09fF $ **FLOATING
C5410 S.n4917 SUB 1.88fF $ **FLOATING
C5411 S.t323 SUB 0.02fF
C5412 S.n4918 SUB 0.24fF $ **FLOATING
C5413 S.n4919 SUB 0.91fF $ **FLOATING
C5414 S.n4920 SUB 0.05fF $ **FLOATING
C5415 S.t1542 SUB 0.02fF
C5416 S.n4921 SUB 0.12fF $ **FLOATING
C5417 S.n4922 SUB 0.14fF $ **FLOATING
C5418 S.n4924 SUB 0.78fF $ **FLOATING
C5419 S.n4925 SUB 1.94fF $ **FLOATING
C5420 S.n4926 SUB 1.88fF $ **FLOATING
C5421 S.n4927 SUB 0.12fF $ **FLOATING
C5422 S.t2527 SUB 0.02fF
C5423 S.n4928 SUB 0.14fF $ **FLOATING
C5424 S.t294 SUB 0.02fF
C5425 S.n4930 SUB 0.24fF $ **FLOATING
C5426 S.n4931 SUB 0.36fF $ **FLOATING
C5427 S.n4932 SUB 0.61fF $ **FLOATING
C5428 S.n4933 SUB 1.84fF $ **FLOATING
C5429 S.n4934 SUB 2.99fF $ **FLOATING
C5430 S.t1984 SUB 0.02fF
C5431 S.n4935 SUB 0.24fF $ **FLOATING
C5432 S.n4936 SUB 0.91fF $ **FLOATING
C5433 S.n4937 SUB 0.05fF $ **FLOATING
C5434 S.t801 SUB 0.02fF
C5435 S.n4938 SUB 0.12fF $ **FLOATING
C5436 S.n4939 SUB 0.14fF $ **FLOATING
C5437 S.n4941 SUB 1.89fF $ **FLOATING
C5438 S.n4942 SUB 1.88fF $ **FLOATING
C5439 S.t1960 SUB 0.02fF
C5440 S.n4943 SUB 0.24fF $ **FLOATING
C5441 S.n4944 SUB 0.36fF $ **FLOATING
C5442 S.n4945 SUB 0.61fF $ **FLOATING
C5443 S.n4946 SUB 0.12fF $ **FLOATING
C5444 S.t1651 SUB 0.02fF
C5445 S.n4947 SUB 0.14fF $ **FLOATING
C5446 S.n4949 SUB 1.16fF $ **FLOATING
C5447 S.n4950 SUB 0.22fF $ **FLOATING
C5448 S.n4951 SUB 0.25fF $ **FLOATING
C5449 S.n4952 SUB 0.09fF $ **FLOATING
C5450 S.n4953 SUB 1.88fF $ **FLOATING
C5451 S.t1136 SUB 0.02fF
C5452 S.n4954 SUB 0.24fF $ **FLOATING
C5453 S.n4955 SUB 0.91fF $ **FLOATING
C5454 S.n4956 SUB 0.05fF $ **FLOATING
C5455 S.t2451 SUB 0.02fF
C5456 S.n4957 SUB 0.12fF $ **FLOATING
C5457 S.n4958 SUB 0.14fF $ **FLOATING
C5458 S.n4960 SUB 0.78fF $ **FLOATING
C5459 S.n4961 SUB 1.94fF $ **FLOATING
C5460 S.n4962 SUB 1.88fF $ **FLOATING
C5461 S.n4963 SUB 0.12fF $ **FLOATING
C5462 S.t780 SUB 0.02fF
C5463 S.n4964 SUB 0.14fF $ **FLOATING
C5464 S.t1102 SUB 0.02fF
C5465 S.n4966 SUB 0.24fF $ **FLOATING
C5466 S.n4967 SUB 0.36fF $ **FLOATING
C5467 S.n4968 SUB 0.61fF $ **FLOATING
C5468 S.n4969 SUB 1.84fF $ **FLOATING
C5469 S.n4970 SUB 2.99fF $ **FLOATING
C5470 S.t257 SUB 0.02fF
C5471 S.n4971 SUB 0.24fF $ **FLOATING
C5472 S.n4972 SUB 0.91fF $ **FLOATING
C5473 S.n4973 SUB 0.05fF $ **FLOATING
C5474 S.t1582 SUB 0.02fF
C5475 S.n4974 SUB 0.12fF $ **FLOATING
C5476 S.n4975 SUB 0.14fF $ **FLOATING
C5477 S.n4977 SUB 1.89fF $ **FLOATING
C5478 S.n4978 SUB 1.88fF $ **FLOATING
C5479 S.t227 SUB 0.02fF
C5480 S.n4979 SUB 0.24fF $ **FLOATING
C5481 S.n4980 SUB 0.36fF $ **FLOATING
C5482 S.n4981 SUB 0.61fF $ **FLOATING
C5483 S.n4982 SUB 0.12fF $ **FLOATING
C5484 S.t2433 SUB 0.02fF
C5485 S.n4983 SUB 0.14fF $ **FLOATING
C5486 S.n4985 SUB 1.16fF $ **FLOATING
C5487 S.n4986 SUB 0.22fF $ **FLOATING
C5488 S.n4987 SUB 0.25fF $ **FLOATING
C5489 S.n4988 SUB 0.09fF $ **FLOATING
C5490 S.n4989 SUB 1.88fF $ **FLOATING
C5491 S.t1923 SUB 0.02fF
C5492 S.n4990 SUB 0.24fF $ **FLOATING
C5493 S.n4991 SUB 0.91fF $ **FLOATING
C5494 S.n4992 SUB 0.05fF $ **FLOATING
C5495 S.t715 SUB 0.02fF
C5496 S.n4993 SUB 0.12fF $ **FLOATING
C5497 S.n4994 SUB 0.14fF $ **FLOATING
C5498 S.n4996 SUB 0.78fF $ **FLOATING
C5499 S.n4997 SUB 1.94fF $ **FLOATING
C5500 S.n4998 SUB 1.88fF $ **FLOATING
C5501 S.n4999 SUB 0.12fF $ **FLOATING
C5502 S.t1706 SUB 0.02fF
C5503 S.n5000 SUB 0.14fF $ **FLOATING
C5504 S.t1893 SUB 0.02fF
C5505 S.n5002 SUB 0.24fF $ **FLOATING
C5506 S.n5003 SUB 0.36fF $ **FLOATING
C5507 S.n5004 SUB 0.61fF $ **FLOATING
C5508 S.n5005 SUB 1.84fF $ **FLOATING
C5509 S.n5006 SUB 2.99fF $ **FLOATING
C5510 S.t1061 SUB 0.02fF
C5511 S.n5007 SUB 0.24fF $ **FLOATING
C5512 S.n5008 SUB 0.91fF $ **FLOATING
C5513 S.n5009 SUB 0.05fF $ **FLOATING
C5514 S.t2370 SUB 0.02fF
C5515 S.n5010 SUB 0.12fF $ **FLOATING
C5516 S.n5011 SUB 0.14fF $ **FLOATING
C5517 S.n5013 SUB 1.89fF $ **FLOATING
C5518 S.n5014 SUB 1.75fF $ **FLOATING
C5519 S.t2504 SUB 0.02fF
C5520 S.n5015 SUB 0.24fF $ **FLOATING
C5521 S.n5016 SUB 0.36fF $ **FLOATING
C5522 S.n5017 SUB 0.61fF $ **FLOATING
C5523 S.n5018 SUB 0.12fF $ **FLOATING
C5524 S.t722 SUB 0.02fF
C5525 S.n5019 SUB 0.14fF $ **FLOATING
C5526 S.n5021 SUB 1.16fF $ **FLOATING
C5527 S.n5022 SUB 0.22fF $ **FLOATING
C5528 S.n5023 SUB 0.25fF $ **FLOATING
C5529 S.n5024 SUB 0.09fF $ **FLOATING
C5530 S.n5025 SUB 2.44fF $ **FLOATING
C5531 S.t1805 SUB 0.02fF
C5532 S.n5026 SUB 0.24fF $ **FLOATING
C5533 S.n5027 SUB 0.91fF $ **FLOATING
C5534 S.n5028 SUB 0.05fF $ **FLOATING
C5535 S.t1513 SUB 0.02fF
C5536 S.n5029 SUB 0.12fF $ **FLOATING
C5537 S.n5030 SUB 0.14fF $ **FLOATING
C5538 S.n5032 SUB 1.88fF $ **FLOATING
C5539 S.n5033 SUB 0.48fF $ **FLOATING
C5540 S.n5034 SUB 0.09fF $ **FLOATING
C5541 S.n5035 SUB 0.33fF $ **FLOATING
C5542 S.n5036 SUB 0.30fF $ **FLOATING
C5543 S.n5037 SUB 0.77fF $ **FLOATING
C5544 S.n5038 SUB 0.59fF $ **FLOATING
C5545 S.t1629 SUB 0.02fF
C5546 S.n5039 SUB 0.24fF $ **FLOATING
C5547 S.n5040 SUB 0.36fF $ **FLOATING
C5548 S.n5041 SUB 0.61fF $ **FLOATING
C5549 S.n5042 SUB 0.12fF $ **FLOATING
C5550 S.t2375 SUB 0.02fF
C5551 S.n5043 SUB 0.14fF $ **FLOATING
C5552 S.n5045 SUB 2.61fF $ **FLOATING
C5553 S.n5046 SUB 2.16fF $ **FLOATING
C5554 S.t940 SUB 0.02fF
C5555 S.n5047 SUB 0.24fF $ **FLOATING
C5556 S.n5048 SUB 0.91fF $ **FLOATING
C5557 S.n5049 SUB 0.05fF $ **FLOATING
C5558 S.t571 SUB 0.02fF
C5559 S.n5050 SUB 0.12fF $ **FLOATING
C5560 S.n5051 SUB 0.14fF $ **FLOATING
C5561 S.n5053 SUB 0.78fF $ **FLOATING
C5562 S.n5054 SUB 2.30fF $ **FLOATING
C5563 S.n5055 SUB 1.88fF $ **FLOATING
C5564 S.n5056 SUB 0.12fF $ **FLOATING
C5565 S.t1519 SUB 0.02fF
C5566 S.n5057 SUB 0.14fF $ **FLOATING
C5567 S.t762 SUB 0.02fF
C5568 S.n5059 SUB 0.24fF $ **FLOATING
C5569 S.n5060 SUB 0.36fF $ **FLOATING
C5570 S.n5061 SUB 0.61fF $ **FLOATING
C5571 S.n5062 SUB 1.39fF $ **FLOATING
C5572 S.n5063 SUB 0.71fF $ **FLOATING
C5573 S.n5064 SUB 1.14fF $ **FLOATING
C5574 S.n5065 SUB 0.35fF $ **FLOATING
C5575 S.n5066 SUB 2.03fF $ **FLOATING
C5576 S.t2580 SUB 0.02fF
C5577 S.n5067 SUB 0.24fF $ **FLOATING
C5578 S.n5068 SUB 0.91fF $ **FLOATING
C5579 S.n5069 SUB 0.05fF $ **FLOATING
C5580 S.t2216 SUB 0.02fF
C5581 S.n5070 SUB 0.12fF $ **FLOATING
C5582 S.n5071 SUB 0.14fF $ **FLOATING
C5583 S.n5073 SUB 1.89fF $ **FLOATING
C5584 S.n5074 SUB 1.88fF $ **FLOATING
C5585 S.t2415 SUB 0.02fF
C5586 S.n5075 SUB 0.24fF $ **FLOATING
C5587 S.n5076 SUB 0.36fF $ **FLOATING
C5588 S.n5077 SUB 0.61fF $ **FLOATING
C5589 S.n5078 SUB 0.12fF $ **FLOATING
C5590 S.t658 SUB 0.02fF
C5591 S.n5079 SUB 0.14fF $ **FLOATING
C5592 S.n5081 SUB 1.16fF $ **FLOATING
C5593 S.n5082 SUB 0.22fF $ **FLOATING
C5594 S.n5083 SUB 0.25fF $ **FLOATING
C5595 S.n5084 SUB 0.09fF $ **FLOATING
C5596 S.n5085 SUB 1.88fF $ **FLOATING
C5597 S.t1703 SUB 0.02fF
C5598 S.n5086 SUB 0.24fF $ **FLOATING
C5599 S.n5087 SUB 0.91fF $ **FLOATING
C5600 S.n5088 SUB 0.05fF $ **FLOATING
C5601 S.t1355 SUB 0.02fF
C5602 S.n5089 SUB 0.12fF $ **FLOATING
C5603 S.n5090 SUB 0.14fF $ **FLOATING
C5604 S.n5092 SUB 20.78fF $ **FLOATING
C5605 S.n5093 SUB 1.88fF $ **FLOATING
C5606 S.n5094 SUB 2.67fF $ **FLOATING
C5607 S.t2350 SUB 0.02fF
C5608 S.n5095 SUB 0.24fF $ **FLOATING
C5609 S.n5096 SUB 0.36fF $ **FLOATING
C5610 S.n5097 SUB 0.61fF $ **FLOATING
C5611 S.n5098 SUB 0.12fF $ **FLOATING
C5612 S.t596 SUB 0.02fF
C5613 S.n5099 SUB 0.14fF $ **FLOATING
C5614 S.n5101 SUB 2.80fF $ **FLOATING
C5615 S.n5102 SUB 2.30fF $ **FLOATING
C5616 S.t1401 SUB 0.02fF
C5617 S.n5103 SUB 0.12fF $ **FLOATING
C5618 S.n5104 SUB 0.14fF $ **FLOATING
C5619 S.t1605 SUB 0.02fF
C5620 S.n5106 SUB 0.24fF $ **FLOATING
C5621 S.n5107 SUB 0.91fF $ **FLOATING
C5622 S.n5108 SUB 0.05fF $ **FLOATING
C5623 S.n5109 SUB 1.88fF $ **FLOATING
C5624 S.n5110 SUB 2.67fF $ **FLOATING
C5625 S.t1491 SUB 0.02fF
C5626 S.n5111 SUB 0.24fF $ **FLOATING
C5627 S.n5112 SUB 0.36fF $ **FLOATING
C5628 S.n5113 SUB 0.61fF $ **FLOATING
C5629 S.n5114 SUB 0.12fF $ **FLOATING
C5630 S.t2246 SUB 0.02fF
C5631 S.n5115 SUB 0.14fF $ **FLOATING
C5632 S.n5117 SUB 2.80fF $ **FLOATING
C5633 S.n5118 SUB 2.30fF $ **FLOATING
C5634 S.t531 SUB 0.02fF
C5635 S.n5119 SUB 0.12fF $ **FLOATING
C5636 S.n5120 SUB 0.14fF $ **FLOATING
C5637 S.t741 SUB 0.02fF
C5638 S.n5122 SUB 0.24fF $ **FLOATING
C5639 S.n5123 SUB 0.91fF $ **FLOATING
C5640 S.n5124 SUB 0.05fF $ **FLOATING
C5641 S.n5125 SUB 2.73fF $ **FLOATING
C5642 S.n5126 SUB 1.59fF $ **FLOATING
C5643 S.n5127 SUB 0.12fF $ **FLOATING
C5644 S.t511 SUB 0.02fF
C5645 S.n5128 SUB 0.14fF $ **FLOATING
C5646 S.t436 SUB 0.02fF
C5647 S.n5130 SUB 0.24fF $ **FLOATING
C5648 S.n5131 SUB 0.36fF $ **FLOATING
C5649 S.n5132 SUB 0.61fF $ **FLOATING
C5650 S.n5133 SUB 0.07fF $ **FLOATING
C5651 S.n5134 SUB 0.01fF $ **FLOATING
C5652 S.n5135 SUB 0.24fF $ **FLOATING
C5653 S.n5136 SUB 1.16fF $ **FLOATING
C5654 S.n5137 SUB 1.35fF $ **FLOATING
C5655 S.n5138 SUB 2.30fF $ **FLOATING
C5656 S.t1250 SUB 0.02fF
C5657 S.n5139 SUB 0.12fF $ **FLOATING
C5658 S.n5140 SUB 0.14fF $ **FLOATING
C5659 S.t1432 SUB 0.02fF
C5660 S.n5142 SUB 0.24fF $ **FLOATING
C5661 S.n5143 SUB 0.91fF $ **FLOATING
C5662 S.n5144 SUB 0.05fF $ **FLOATING
C5663 S.t81 SUB 48.31fF
C5664 S.t2393 SUB 0.02fF
C5665 S.n5145 SUB 0.24fF $ **FLOATING
C5666 S.n5146 SUB 0.91fF $ **FLOATING
C5667 S.n5147 SUB 0.05fF $ **FLOATING
C5668 S.t2174 SUB 0.02fF
C5669 S.n5148 SUB 0.12fF $ **FLOATING
C5670 S.n5149 SUB 0.14fF $ **FLOATING
C5671 S.n5151 SUB 0.12fF $ **FLOATING
C5672 S.t1387 SUB 0.02fF
C5673 S.n5152 SUB 0.14fF $ **FLOATING
C5674 S.n5154 SUB 5.17fF $ **FLOATING
C5675 S.n5155 SUB 5.44fF $ **FLOATING
C5676 S.t1281 SUB 0.02fF
C5677 S.n5156 SUB 0.12fF $ **FLOATING
C5678 S.n5157 SUB 0.14fF $ **FLOATING
C5679 S.t694 SUB 0.02fF
C5680 S.n5159 SUB 0.24fF $ **FLOATING
C5681 S.n5160 SUB 0.91fF $ **FLOATING
C5682 S.n5161 SUB 0.05fF $ **FLOATING
C5683 S.t360 SUB 47.92fF
C5684 S.t1715 SUB 0.02fF
C5685 S.n5162 SUB 1.19fF $ **FLOATING
C5686 S.n5163 SUB 0.05fF $ **FLOATING
C5687 S.t1809 SUB 0.02fF
C5688 S.n5164 SUB 0.01fF $ **FLOATING
C5689 S.n5165 SUB 0.26fF $ **FLOATING
C5690 S.n5167 SUB 1.50fF $ **FLOATING
C5691 S.n5168 SUB 1.30fF $ **FLOATING
C5692 S.n5169 SUB 0.28fF $ **FLOATING
C5693 S.n5170 SUB 0.24fF $ **FLOATING
C5694 S.n5171 SUB 4.39fF $ **FLOATING
C5695 S.n5172 SUB 0.01fF $ **FLOATING
C5696 S.n5173 SUB 0.02fF $ **FLOATING
C5697 S.n5174 SUB 0.03fF $ **FLOATING
C5698 S.n5175 SUB 0.04fF $ **FLOATING
C5699 S.n5176 SUB 0.17fF $ **FLOATING
C5700 S.n5177 SUB 0.01fF $ **FLOATING
C5701 S.n5178 SUB 0.02fF $ **FLOATING
C5702 S.n5179 SUB 0.01fF $ **FLOATING
C5703 S.n5180 SUB 0.01fF $ **FLOATING
C5704 S.n5181 SUB 0.01fF $ **FLOATING
C5705 S.n5182 SUB 0.01fF $ **FLOATING
C5706 S.n5183 SUB 0.02fF $ **FLOATING
C5707 S.n5184 SUB 0.01fF $ **FLOATING
C5708 S.n5185 SUB 0.02fF $ **FLOATING
C5709 S.n5186 SUB 0.05fF $ **FLOATING
C5710 S.n5187 SUB 0.04fF $ **FLOATING
C5711 S.n5188 SUB 0.11fF $ **FLOATING
C5712 S.n5189 SUB 0.38fF $ **FLOATING
C5713 S.n5190 SUB 0.20fF $ **FLOATING
C5714 S.n5191 SUB 8.97fF $ **FLOATING
C5715 S.n5192 SUB 8.97fF $ **FLOATING
C5716 S.n5193 SUB 0.60fF $ **FLOATING
C5717 S.n5194 SUB 0.22fF $ **FLOATING
C5718 S.n5195 SUB 0.59fF $ **FLOATING
C5719 S.n5196 SUB 3.43fF $ **FLOATING
C5720 S.n5197 SUB 0.29fF $ **FLOATING
C5721 S.t4 SUB 21.38fF
C5722 S.n5198 SUB 21.67fF $ **FLOATING
C5723 S.n5199 SUB 0.77fF $ **FLOATING
C5724 S.n5200 SUB 0.28fF $ **FLOATING
C5725 S.n5201 SUB 4.00fF $ **FLOATING
C5726 S.n5202 SUB 1.35fF $ **FLOATING
C5727 S.t1849 SUB 0.02fF
C5728 S.n5203 SUB 0.64fF $ **FLOATING
C5729 S.n5204 SUB 0.61fF $ **FLOATING
C5730 S.n5205 SUB 1.89fF $ **FLOATING
C5731 S.n5206 SUB 0.06fF $ **FLOATING
C5732 S.n5207 SUB 0.03fF $ **FLOATING
C5733 S.n5208 SUB 0.04fF $ **FLOATING
C5734 S.n5209 SUB 0.99fF $ **FLOATING
C5735 S.n5210 SUB 0.02fF $ **FLOATING
C5736 S.n5211 SUB 0.01fF $ **FLOATING
C5737 S.n5212 SUB 0.02fF $ **FLOATING
C5738 S.n5213 SUB 0.08fF $ **FLOATING
C5739 S.n5214 SUB 0.36fF $ **FLOATING
C5740 S.n5215 SUB 1.85fF $ **FLOATING
C5741 S.t106 SUB 0.02fF
C5742 S.n5216 SUB 0.24fF $ **FLOATING
C5743 S.n5217 SUB 0.36fF $ **FLOATING
C5744 S.n5218 SUB 0.61fF $ **FLOATING
C5745 S.n5219 SUB 0.12fF $ **FLOATING
C5746 S.t2114 SUB 0.02fF
C5747 S.n5220 SUB 0.14fF $ **FLOATING
C5748 S.n5222 SUB 0.70fF $ **FLOATING
C5749 S.n5223 SUB 0.23fF $ **FLOATING
C5750 S.n5224 SUB 0.23fF $ **FLOATING
C5751 S.n5225 SUB 0.70fF $ **FLOATING
C5752 S.n5226 SUB 1.16fF $ **FLOATING
C5753 S.n5227 SUB 0.22fF $ **FLOATING
C5754 S.n5228 SUB 0.25fF $ **FLOATING
C5755 S.n5229 SUB 0.09fF $ **FLOATING
C5756 S.n5230 SUB 1.88fF $ **FLOATING
C5757 S.t1240 SUB 0.02fF
C5758 S.n5231 SUB 0.24fF $ **FLOATING
C5759 S.n5232 SUB 0.91fF $ **FLOATING
C5760 S.n5233 SUB 0.05fF $ **FLOATING
C5761 S.t2304 SUB 0.02fF
C5762 S.n5234 SUB 0.12fF $ **FLOATING
C5763 S.n5235 SUB 0.14fF $ **FLOATING
C5764 S.n5237 SUB 0.25fF $ **FLOATING
C5765 S.n5238 SUB 0.09fF $ **FLOATING
C5766 S.n5239 SUB 0.21fF $ **FLOATING
C5767 S.n5240 SUB 0.92fF $ **FLOATING
C5768 S.n5241 SUB 0.44fF $ **FLOATING
C5769 S.n5242 SUB 1.88fF $ **FLOATING
C5770 S.n5243 SUB 0.12fF $ **FLOATING
C5771 S.t1389 SUB 0.02fF
C5772 S.n5244 SUB 0.14fF $ **FLOATING
C5773 S.t1915 SUB 0.02fF
C5774 S.n5246 SUB 0.24fF $ **FLOATING
C5775 S.n5247 SUB 0.36fF $ **FLOATING
C5776 S.n5248 SUB 0.61fF $ **FLOATING
C5777 S.n5249 SUB 0.02fF $ **FLOATING
C5778 S.n5250 SUB 0.01fF $ **FLOATING
C5779 S.n5251 SUB 0.02fF $ **FLOATING
C5780 S.n5252 SUB 0.08fF $ **FLOATING
C5781 S.n5253 SUB 0.06fF $ **FLOATING
C5782 S.n5254 SUB 0.03fF $ **FLOATING
C5783 S.n5255 SUB 0.04fF $ **FLOATING
C5784 S.n5256 SUB 1.00fF $ **FLOATING
C5785 S.n5257 SUB 0.36fF $ **FLOATING
C5786 S.n5258 SUB 1.87fF $ **FLOATING
C5787 S.n5259 SUB 1.99fF $ **FLOATING
C5788 S.t514 SUB 0.02fF
C5789 S.n5260 SUB 0.24fF $ **FLOATING
C5790 S.n5261 SUB 0.91fF $ **FLOATING
C5791 S.n5262 SUB 0.05fF $ **FLOATING
C5792 S.t1449 SUB 0.02fF
C5793 S.n5263 SUB 0.12fF $ **FLOATING
C5794 S.n5264 SUB 0.14fF $ **FLOATING
C5795 S.n5266 SUB 1.89fF $ **FLOATING
C5796 S.n5267 SUB 0.06fF $ **FLOATING
C5797 S.n5268 SUB 0.03fF $ **FLOATING
C5798 S.n5269 SUB 0.04fF $ **FLOATING
C5799 S.n5270 SUB 0.99fF $ **FLOATING
C5800 S.n5271 SUB 0.02fF $ **FLOATING
C5801 S.n5272 SUB 0.01fF $ **FLOATING
C5802 S.n5273 SUB 0.02fF $ **FLOATING
C5803 S.n5274 SUB 0.08fF $ **FLOATING
C5804 S.n5275 SUB 0.36fF $ **FLOATING
C5805 S.n5276 SUB 1.85fF $ **FLOATING
C5806 S.t1055 SUB 0.02fF
C5807 S.n5277 SUB 0.24fF $ **FLOATING
C5808 S.n5278 SUB 0.36fF $ **FLOATING
C5809 S.n5279 SUB 0.61fF $ **FLOATING
C5810 S.n5280 SUB 0.12fF $ **FLOATING
C5811 S.t516 SUB 0.02fF
C5812 S.n5281 SUB 0.14fF $ **FLOATING
C5813 S.n5283 SUB 0.70fF $ **FLOATING
C5814 S.n5284 SUB 0.23fF $ **FLOATING
C5815 S.n5285 SUB 0.23fF $ **FLOATING
C5816 S.n5286 SUB 0.70fF $ **FLOATING
C5817 S.n5287 SUB 1.16fF $ **FLOATING
C5818 S.n5288 SUB 0.22fF $ **FLOATING
C5819 S.n5289 SUB 0.25fF $ **FLOATING
C5820 S.n5290 SUB 0.09fF $ **FLOATING
C5821 S.n5291 SUB 1.88fF $ **FLOATING
C5822 S.t2157 SUB 0.02fF
C5823 S.n5292 SUB 0.24fF $ **FLOATING
C5824 S.n5293 SUB 0.91fF $ **FLOATING
C5825 S.n5294 SUB 0.05fF $ **FLOATING
C5826 S.t587 SUB 0.02fF
C5827 S.n5295 SUB 0.12fF $ **FLOATING
C5828 S.n5296 SUB 0.14fF $ **FLOATING
C5829 S.n5298 SUB 0.25fF $ **FLOATING
C5830 S.n5299 SUB 0.09fF $ **FLOATING
C5831 S.n5300 SUB 0.21fF $ **FLOATING
C5832 S.n5301 SUB 0.92fF $ **FLOATING
C5833 S.n5302 SUB 0.44fF $ **FLOATING
C5834 S.n5303 SUB 1.88fF $ **FLOATING
C5835 S.n5304 SUB 0.12fF $ **FLOATING
C5836 S.t2161 SUB 0.02fF
C5837 S.n5305 SUB 0.14fF $ **FLOATING
C5838 S.t168 SUB 0.02fF
C5839 S.n5307 SUB 0.24fF $ **FLOATING
C5840 S.n5308 SUB 0.36fF $ **FLOATING
C5841 S.n5309 SUB 0.61fF $ **FLOATING
C5842 S.n5310 SUB 0.02fF $ **FLOATING
C5843 S.n5311 SUB 0.01fF $ **FLOATING
C5844 S.n5312 SUB 0.02fF $ **FLOATING
C5845 S.n5313 SUB 0.08fF $ **FLOATING
C5846 S.n5314 SUB 0.06fF $ **FLOATING
C5847 S.n5315 SUB 0.03fF $ **FLOATING
C5848 S.n5316 SUB 0.04fF $ **FLOATING
C5849 S.n5317 SUB 1.00fF $ **FLOATING
C5850 S.n5318 SUB 0.36fF $ **FLOATING
C5851 S.n5319 SUB 1.87fF $ **FLOATING
C5852 S.n5320 SUB 1.99fF $ **FLOATING
C5853 S.t1294 SUB 0.02fF
C5854 S.n5321 SUB 0.24fF $ **FLOATING
C5855 S.n5322 SUB 0.91fF $ **FLOATING
C5856 S.n5323 SUB 0.05fF $ **FLOATING
C5857 S.t2235 SUB 0.02fF
C5858 S.n5324 SUB 0.12fF $ **FLOATING
C5859 S.n5325 SUB 0.14fF $ **FLOATING
C5860 S.n5327 SUB 1.89fF $ **FLOATING
C5861 S.n5328 SUB 0.06fF $ **FLOATING
C5862 S.n5329 SUB 0.03fF $ **FLOATING
C5863 S.n5330 SUB 0.04fF $ **FLOATING
C5864 S.n5331 SUB 0.99fF $ **FLOATING
C5865 S.n5332 SUB 0.02fF $ **FLOATING
C5866 S.n5333 SUB 0.01fF $ **FLOATING
C5867 S.n5334 SUB 0.02fF $ **FLOATING
C5868 S.n5335 SUB 0.08fF $ **FLOATING
C5869 S.n5336 SUB 0.36fF $ **FLOATING
C5870 S.n5337 SUB 1.85fF $ **FLOATING
C5871 S.t1833 SUB 0.02fF
C5872 S.n5338 SUB 0.24fF $ **FLOATING
C5873 S.n5339 SUB 0.36fF $ **FLOATING
C5874 S.n5340 SUB 0.61fF $ **FLOATING
C5875 S.n5341 SUB 0.12fF $ **FLOATING
C5876 S.t1297 SUB 0.02fF
C5877 S.n5342 SUB 0.14fF $ **FLOATING
C5878 S.n5344 SUB 0.70fF $ **FLOATING
C5879 S.n5345 SUB 0.23fF $ **FLOATING
C5880 S.n5346 SUB 0.23fF $ **FLOATING
C5881 S.n5347 SUB 0.70fF $ **FLOATING
C5882 S.n5348 SUB 1.16fF $ **FLOATING
C5883 S.n5349 SUB 0.22fF $ **FLOATING
C5884 S.n5350 SUB 0.25fF $ **FLOATING
C5885 S.n5351 SUB 0.09fF $ **FLOATING
C5886 S.n5352 SUB 1.88fF $ **FLOATING
C5887 S.t410 SUB 0.02fF
C5888 S.n5353 SUB 0.24fF $ **FLOATING
C5889 S.n5354 SUB 0.91fF $ **FLOATING
C5890 S.n5355 SUB 0.05fF $ **FLOATING
C5891 S.t1373 SUB 0.02fF
C5892 S.n5356 SUB 0.12fF $ **FLOATING
C5893 S.n5357 SUB 0.14fF $ **FLOATING
C5894 S.n5359 SUB 0.25fF $ **FLOATING
C5895 S.n5360 SUB 0.09fF $ **FLOATING
C5896 S.n5361 SUB 0.21fF $ **FLOATING
C5897 S.n5362 SUB 0.92fF $ **FLOATING
C5898 S.n5363 SUB 0.44fF $ **FLOATING
C5899 S.n5364 SUB 1.88fF $ **FLOATING
C5900 S.n5365 SUB 0.12fF $ **FLOATING
C5901 S.t414 SUB 0.02fF
C5902 S.n5366 SUB 0.14fF $ **FLOATING
C5903 S.t967 SUB 0.02fF
C5904 S.n5368 SUB 0.24fF $ **FLOATING
C5905 S.n5369 SUB 0.36fF $ **FLOATING
C5906 S.n5370 SUB 0.61fF $ **FLOATING
C5907 S.n5371 SUB 0.02fF $ **FLOATING
C5908 S.n5372 SUB 0.01fF $ **FLOATING
C5909 S.n5373 SUB 0.02fF $ **FLOATING
C5910 S.n5374 SUB 0.08fF $ **FLOATING
C5911 S.n5375 SUB 0.06fF $ **FLOATING
C5912 S.n5376 SUB 0.03fF $ **FLOATING
C5913 S.n5377 SUB 0.04fF $ **FLOATING
C5914 S.n5378 SUB 1.00fF $ **FLOATING
C5915 S.n5379 SUB 0.36fF $ **FLOATING
C5916 S.n5380 SUB 1.87fF $ **FLOATING
C5917 S.n5381 SUB 1.99fF $ **FLOATING
C5918 S.t2058 SUB 0.02fF
C5919 S.n5382 SUB 0.24fF $ **FLOATING
C5920 S.n5383 SUB 0.91fF $ **FLOATING
C5921 S.n5384 SUB 0.05fF $ **FLOATING
C5922 S.t500 SUB 0.02fF
C5923 S.n5385 SUB 0.12fF $ **FLOATING
C5924 S.n5386 SUB 0.14fF $ **FLOATING
C5925 S.n5388 SUB 1.89fF $ **FLOATING
C5926 S.n5389 SUB 0.07fF $ **FLOATING
C5927 S.n5390 SUB 0.04fF $ **FLOATING
C5928 S.n5391 SUB 0.05fF $ **FLOATING
C5929 S.n5392 SUB 0.87fF $ **FLOATING
C5930 S.n5393 SUB 0.01fF $ **FLOATING
C5931 S.n5394 SUB 0.01fF $ **FLOATING
C5932 S.n5395 SUB 0.01fF $ **FLOATING
C5933 S.n5396 SUB 0.07fF $ **FLOATING
C5934 S.n5397 SUB 0.68fF $ **FLOATING
C5935 S.n5398 SUB 0.72fF $ **FLOATING
C5936 S.t32 SUB 0.02fF
C5937 S.n5399 SUB 0.24fF $ **FLOATING
C5938 S.n5400 SUB 0.36fF $ **FLOATING
C5939 S.n5401 SUB 0.61fF $ **FLOATING
C5940 S.n5402 SUB 0.12fF $ **FLOATING
C5941 S.t2061 SUB 0.02fF
C5942 S.n5403 SUB 0.14fF $ **FLOATING
C5943 S.n5405 SUB 0.70fF $ **FLOATING
C5944 S.n5406 SUB 0.23fF $ **FLOATING
C5945 S.n5407 SUB 0.23fF $ **FLOATING
C5946 S.n5408 SUB 0.70fF $ **FLOATING
C5947 S.n5409 SUB 1.16fF $ **FLOATING
C5948 S.n5410 SUB 0.22fF $ **FLOATING
C5949 S.n5411 SUB 0.25fF $ **FLOATING
C5950 S.n5412 SUB 0.09fF $ **FLOATING
C5951 S.n5413 SUB 2.31fF $ **FLOATING
C5952 S.t1197 SUB 0.02fF
C5953 S.n5414 SUB 0.24fF $ **FLOATING
C5954 S.n5415 SUB 0.91fF $ **FLOATING
C5955 S.n5416 SUB 0.05fF $ **FLOATING
C5956 S.t2276 SUB 0.02fF
C5957 S.n5417 SUB 0.12fF $ **FLOATING
C5958 S.n5418 SUB 0.14fF $ **FLOATING
C5959 S.n5420 SUB 1.88fF $ **FLOATING
C5960 S.n5421 SUB 0.46fF $ **FLOATING
C5961 S.n5422 SUB 0.22fF $ **FLOATING
C5962 S.n5423 SUB 0.38fF $ **FLOATING
C5963 S.n5424 SUB 0.16fF $ **FLOATING
C5964 S.n5425 SUB 0.28fF $ **FLOATING
C5965 S.n5426 SUB 0.21fF $ **FLOATING
C5966 S.n5427 SUB 0.30fF $ **FLOATING
C5967 S.n5428 SUB 0.42fF $ **FLOATING
C5968 S.n5429 SUB 0.21fF $ **FLOATING
C5969 S.t154 SUB 0.02fF
C5970 S.n5430 SUB 0.24fF $ **FLOATING
C5971 S.n5431 SUB 0.36fF $ **FLOATING
C5972 S.n5432 SUB 0.61fF $ **FLOATING
C5973 S.n5433 SUB 0.12fF $ **FLOATING
C5974 S.t2139 SUB 0.02fF
C5975 S.n5434 SUB 0.14fF $ **FLOATING
C5976 S.n5436 SUB 0.04fF $ **FLOATING
C5977 S.n5437 SUB 0.03fF $ **FLOATING
C5978 S.n5438 SUB 0.03fF $ **FLOATING
C5979 S.n5439 SUB 0.10fF $ **FLOATING
C5980 S.n5440 SUB 0.36fF $ **FLOATING
C5981 S.n5441 SUB 0.38fF $ **FLOATING
C5982 S.n5442 SUB 0.11fF $ **FLOATING
C5983 S.n5443 SUB 0.12fF $ **FLOATING
C5984 S.n5444 SUB 0.07fF $ **FLOATING
C5985 S.n5445 SUB 0.12fF $ **FLOATING
C5986 S.n5446 SUB 0.18fF $ **FLOATING
C5987 S.n5447 SUB 4.00fF $ **FLOATING
C5988 S.t1717 SUB 0.02fF
C5989 S.n5448 SUB 0.24fF $ **FLOATING
C5990 S.n5449 SUB 0.91fF $ **FLOATING
C5991 S.n5450 SUB 0.05fF $ **FLOATING
C5992 S.t2324 SUB 0.02fF
C5993 S.n5451 SUB 0.12fF $ **FLOATING
C5994 S.n5452 SUB 0.14fF $ **FLOATING
C5995 S.n5454 SUB 0.25fF $ **FLOATING
C5996 S.n5455 SUB 0.09fF $ **FLOATING
C5997 S.n5456 SUB 0.21fF $ **FLOATING
C5998 S.n5457 SUB 1.28fF $ **FLOATING
C5999 S.n5458 SUB 0.53fF $ **FLOATING
C6000 S.n5459 SUB 1.88fF $ **FLOATING
C6001 S.n5460 SUB 0.12fF $ **FLOATING
C6002 S.t1273 SUB 0.02fF
C6003 S.n5461 SUB 0.14fF $ **FLOATING
C6004 S.t1818 SUB 0.02fF
C6005 S.n5463 SUB 0.24fF $ **FLOATING
C6006 S.n5464 SUB 0.36fF $ **FLOATING
C6007 S.n5465 SUB 0.61fF $ **FLOATING
C6008 S.n5466 SUB 1.58fF $ **FLOATING
C6009 S.n5467 SUB 2.45fF $ **FLOATING
C6010 S.t846 SUB 0.02fF
C6011 S.n5468 SUB 0.24fF $ **FLOATING
C6012 S.n5469 SUB 0.91fF $ **FLOATING
C6013 S.n5470 SUB 0.05fF $ **FLOATING
C6014 S.t1466 SUB 0.02fF
C6015 S.n5471 SUB 0.12fF $ **FLOATING
C6016 S.n5472 SUB 0.14fF $ **FLOATING
C6017 S.n5474 SUB 1.89fF $ **FLOATING
C6018 S.n5475 SUB 0.06fF $ **FLOATING
C6019 S.n5476 SUB 0.03fF $ **FLOATING
C6020 S.n5477 SUB 0.04fF $ **FLOATING
C6021 S.n5478 SUB 0.99fF $ **FLOATING
C6022 S.n5479 SUB 0.02fF $ **FLOATING
C6023 S.n5480 SUB 0.01fF $ **FLOATING
C6024 S.n5481 SUB 0.02fF $ **FLOATING
C6025 S.n5482 SUB 0.08fF $ **FLOATING
C6026 S.n5483 SUB 0.36fF $ **FLOATING
C6027 S.n5484 SUB 1.85fF $ **FLOATING
C6028 S.t953 SUB 0.02fF
C6029 S.n5485 SUB 0.24fF $ **FLOATING
C6030 S.n5486 SUB 0.36fF $ **FLOATING
C6031 S.n5487 SUB 0.61fF $ **FLOATING
C6032 S.n5488 SUB 0.12fF $ **FLOATING
C6033 S.t391 SUB 0.02fF
C6034 S.n5489 SUB 0.14fF $ **FLOATING
C6035 S.n5491 SUB 0.70fF $ **FLOATING
C6036 S.n5492 SUB 0.23fF $ **FLOATING
C6037 S.n5493 SUB 0.23fF $ **FLOATING
C6038 S.n5494 SUB 0.70fF $ **FLOATING
C6039 S.n5495 SUB 1.16fF $ **FLOATING
C6040 S.n5496 SUB 0.22fF $ **FLOATING
C6041 S.n5497 SUB 0.25fF $ **FLOATING
C6042 S.n5498 SUB 0.09fF $ **FLOATING
C6043 S.n5499 SUB 1.88fF $ **FLOATING
C6044 S.t2489 SUB 0.02fF
C6045 S.n5500 SUB 0.24fF $ **FLOATING
C6046 S.n5501 SUB 0.91fF $ **FLOATING
C6047 S.n5502 SUB 0.05fF $ **FLOATING
C6048 S.t605 SUB 0.02fF
C6049 S.n5503 SUB 0.12fF $ **FLOATING
C6050 S.n5504 SUB 0.14fF $ **FLOATING
C6051 S.n5506 SUB 20.78fF $ **FLOATING
C6052 S.n5507 SUB 0.06fF $ **FLOATING
C6053 S.n5508 SUB 0.20fF $ **FLOATING
C6054 S.n5509 SUB 0.09fF $ **FLOATING
C6055 S.n5510 SUB 0.21fF $ **FLOATING
C6056 S.n5511 SUB 0.10fF $ **FLOATING
C6057 S.n5512 SUB 0.30fF $ **FLOATING
C6058 S.n5513 SUB 0.69fF $ **FLOATING
C6059 S.n5514 SUB 0.45fF $ **FLOATING
C6060 S.n5515 SUB 2.33fF $ **FLOATING
C6061 S.n5516 SUB 0.12fF $ **FLOATING
C6062 S.t467 SUB 0.02fF
C6063 S.n5517 SUB 0.14fF $ **FLOATING
C6064 S.t1009 SUB 0.02fF
C6065 S.n5519 SUB 0.24fF $ **FLOATING
C6066 S.n5520 SUB 0.36fF $ **FLOATING
C6067 S.n5521 SUB 0.61fF $ **FLOATING
C6068 S.n5522 SUB 1.90fF $ **FLOATING
C6069 S.n5523 SUB 0.17fF $ **FLOATING
C6070 S.n5524 SUB 0.76fF $ **FLOATING
C6071 S.n5525 SUB 0.25fF $ **FLOATING
C6072 S.n5526 SUB 0.30fF $ **FLOATING
C6073 S.n5527 SUB 0.32fF $ **FLOATING
C6074 S.n5528 SUB 0.47fF $ **FLOATING
C6075 S.n5529 SUB 0.16fF $ **FLOATING
C6076 S.n5530 SUB 1.93fF $ **FLOATING
C6077 S.t647 SUB 0.02fF
C6078 S.n5531 SUB 0.12fF $ **FLOATING
C6079 S.n5532 SUB 0.14fF $ **FLOATING
C6080 S.t2107 SUB 0.02fF
C6081 S.n5534 SUB 0.24fF $ **FLOATING
C6082 S.n5535 SUB 0.91fF $ **FLOATING
C6083 S.n5536 SUB 0.05fF $ **FLOATING
C6084 S.n5537 SUB 1.88fF $ **FLOATING
C6085 S.n5538 SUB 0.12fF $ **FLOATING
C6086 S.t2335 SUB 0.02fF
C6087 S.n5539 SUB 0.14fF $ **FLOATING
C6088 S.t508 SUB 0.02fF
C6089 S.n5541 SUB 0.12fF $ **FLOATING
C6090 S.n5542 SUB 0.14fF $ **FLOATING
C6091 S.t860 SUB 0.02fF
C6092 S.n5544 SUB 0.24fF $ **FLOATING
C6093 S.n5545 SUB 0.91fF $ **FLOATING
C6094 S.n5546 SUB 0.05fF $ **FLOATING
C6095 S.t1576 SUB 0.02fF
C6096 S.n5547 SUB 0.24fF $ **FLOATING
C6097 S.n5548 SUB 0.36fF $ **FLOATING
C6098 S.n5549 SUB 0.61fF $ **FLOATING
C6099 S.n5550 SUB 0.32fF $ **FLOATING
C6100 S.n5551 SUB 1.09fF $ **FLOATING
C6101 S.n5552 SUB 0.15fF $ **FLOATING
C6102 S.n5553 SUB 2.10fF $ **FLOATING
C6103 S.n5554 SUB 2.94fF $ **FLOATING
C6104 S.n5555 SUB 1.88fF $ **FLOATING
C6105 S.n5556 SUB 0.12fF $ **FLOATING
C6106 S.t2040 SUB 0.02fF
C6107 S.n5557 SUB 0.14fF $ **FLOATING
C6108 S.t5 SUB 0.02fF
C6109 S.n5559 SUB 0.24fF $ **FLOATING
C6110 S.n5560 SUB 0.36fF $ **FLOATING
C6111 S.n5561 SUB 0.61fF $ **FLOATING
C6112 S.n5562 SUB 0.92fF $ **FLOATING
C6113 S.n5563 SUB 0.32fF $ **FLOATING
C6114 S.n5564 SUB 0.92fF $ **FLOATING
C6115 S.n5565 SUB 1.09fF $ **FLOATING
C6116 S.n5566 SUB 0.15fF $ **FLOATING
C6117 S.n5567 SUB 4.96fF $ **FLOATING
C6118 S.t2257 SUB 0.02fF
C6119 S.n5568 SUB 0.12fF $ **FLOATING
C6120 S.n5569 SUB 0.14fF $ **FLOATING
C6121 S.t1615 SUB 0.02fF
C6122 S.n5571 SUB 0.24fF $ **FLOATING
C6123 S.n5572 SUB 0.91fF $ **FLOATING
C6124 S.n5573 SUB 0.05fF $ **FLOATING
C6125 S.n5574 SUB 1.88fF $ **FLOATING
C6126 S.n5575 SUB 2.67fF $ **FLOATING
C6127 S.t1871 SUB 0.02fF
C6128 S.n5576 SUB 0.24fF $ **FLOATING
C6129 S.n5577 SUB 0.36fF $ **FLOATING
C6130 S.n5578 SUB 0.61fF $ **FLOATING
C6131 S.n5579 SUB 0.12fF $ **FLOATING
C6132 S.t1325 SUB 0.02fF
C6133 S.n5580 SUB 0.14fF $ **FLOATING
C6134 S.n5582 SUB 1.88fF $ **FLOATING
C6135 S.n5583 SUB 2.67fF $ **FLOATING
C6136 S.t708 SUB 0.02fF
C6137 S.n5584 SUB 0.24fF $ **FLOATING
C6138 S.n5585 SUB 0.36fF $ **FLOATING
C6139 S.n5586 SUB 0.61fF $ **FLOATING
C6140 S.t2505 SUB 0.02fF
C6141 S.n5587 SUB 0.24fF $ **FLOATING
C6142 S.n5588 SUB 0.91fF $ **FLOATING
C6143 S.n5589 SUB 0.05fF $ **FLOATING
C6144 S.t2154 SUB 0.02fF
C6145 S.n5590 SUB 0.12fF $ **FLOATING
C6146 S.n5591 SUB 0.14fF $ **FLOATING
C6147 S.n5593 SUB 0.12fF $ **FLOATING
C6148 S.t1477 SUB 0.02fF
C6149 S.n5594 SUB 0.14fF $ **FLOATING
C6150 S.n5596 SUB 2.30fF $ **FLOATING
C6151 S.n5597 SUB 2.94fF $ **FLOATING
C6152 S.n5598 SUB 5.16fF $ **FLOATING
C6153 S.t1399 SUB 0.02fF
C6154 S.n5599 SUB 0.12fF $ **FLOATING
C6155 S.n5600 SUB 0.14fF $ **FLOATING
C6156 S.t903 SUB 0.02fF
C6157 S.n5602 SUB 0.24fF $ **FLOATING
C6158 S.n5603 SUB 0.91fF $ **FLOATING
C6159 S.n5604 SUB 0.05fF $ **FLOATING
C6160 S.n5605 SUB 1.88fF $ **FLOATING
C6161 S.n5606 SUB 2.67fF $ **FLOATING
C6162 S.t1003 SUB 0.02fF
C6163 S.n5607 SUB 0.24fF $ **FLOATING
C6164 S.n5608 SUB 0.36fF $ **FLOATING
C6165 S.n5609 SUB 0.61fF $ **FLOATING
C6166 S.n5610 SUB 0.12fF $ **FLOATING
C6167 S.t447 SUB 0.02fF
C6168 S.n5611 SUB 0.14fF $ **FLOATING
C6169 S.n5613 SUB 5.17fF $ **FLOATING
C6170 S.t528 SUB 0.02fF
C6171 S.n5614 SUB 0.12fF $ **FLOATING
C6172 S.n5615 SUB 0.14fF $ **FLOATING
C6173 S.t2546 SUB 0.02fF
C6174 S.n5617 SUB 0.24fF $ **FLOATING
C6175 S.n5618 SUB 0.91fF $ **FLOATING
C6176 S.n5619 SUB 0.05fF $ **FLOATING
C6177 S.n5620 SUB 1.88fF $ **FLOATING
C6178 S.n5621 SUB 2.67fF $ **FLOATING
C6179 S.t99 SUB 0.02fF
C6180 S.n5622 SUB 0.24fF $ **FLOATING
C6181 S.n5623 SUB 0.36fF $ **FLOATING
C6182 S.n5624 SUB 0.61fF $ **FLOATING
C6183 S.n5625 SUB 0.12fF $ **FLOATING
C6184 S.t2090 SUB 0.02fF
C6185 S.n5626 SUB 0.14fF $ **FLOATING
C6186 S.n5628 SUB 5.17fF $ **FLOATING
C6187 S.t2170 SUB 0.02fF
C6188 S.n5629 SUB 0.12fF $ **FLOATING
C6189 S.n5630 SUB 0.14fF $ **FLOATING
C6190 S.t1673 SUB 0.02fF
C6191 S.n5632 SUB 0.24fF $ **FLOATING
C6192 S.n5633 SUB 0.91fF $ **FLOATING
C6193 S.n5634 SUB 0.05fF $ **FLOATING
C6194 S.n5635 SUB 1.88fF $ **FLOATING
C6195 S.n5636 SUB 2.67fF $ **FLOATING
C6196 S.t1776 SUB 0.02fF
C6197 S.n5637 SUB 0.24fF $ **FLOATING
C6198 S.n5638 SUB 0.36fF $ **FLOATING
C6199 S.n5639 SUB 0.61fF $ **FLOATING
C6200 S.n5640 SUB 0.12fF $ **FLOATING
C6201 S.t1228 SUB 0.02fF
C6202 S.n5641 SUB 0.14fF $ **FLOATING
C6203 S.n5643 SUB 4.90fF $ **FLOATING
C6204 S.t1308 SUB 0.02fF
C6205 S.n5644 SUB 0.12fF $ **FLOATING
C6206 S.n5645 SUB 0.14fF $ **FLOATING
C6207 S.t798 SUB 0.02fF
C6208 S.n5647 SUB 0.24fF $ **FLOATING
C6209 S.n5648 SUB 0.91fF $ **FLOATING
C6210 S.n5649 SUB 0.05fF $ **FLOATING
C6211 S.n5650 SUB 1.88fF $ **FLOATING
C6212 S.n5651 SUB 2.67fF $ **FLOATING
C6213 S.t2426 SUB 0.02fF
C6214 S.n5652 SUB 0.24fF $ **FLOATING
C6215 S.n5653 SUB 0.36fF $ **FLOATING
C6216 S.n5654 SUB 0.61fF $ **FLOATING
C6217 S.n5655 SUB 0.12fF $ **FLOATING
C6218 S.t1179 SUB 0.02fF
C6219 S.n5656 SUB 0.14fF $ **FLOATING
C6220 S.n5658 SUB 1.88fF $ **FLOATING
C6221 S.n5659 SUB 2.68fF $ **FLOATING
C6222 S.t2305 SUB 0.02fF
C6223 S.n5660 SUB 0.24fF $ **FLOATING
C6224 S.n5661 SUB 0.36fF $ **FLOATING
C6225 S.n5662 SUB 0.61fF $ **FLOATING
C6226 S.t75 SUB 0.02fF
C6227 S.n5663 SUB 1.22fF $ **FLOATING
C6228 S.n5664 SUB 0.36fF $ **FLOATING
C6229 S.n5665 SUB 1.22fF $ **FLOATING
C6230 S.n5666 SUB 0.61fF $ **FLOATING
C6231 S.n5667 SUB 0.35fF $ **FLOATING
C6232 S.n5668 SUB 0.63fF $ **FLOATING
C6233 S.n5669 SUB 1.15fF $ **FLOATING
C6234 S.n5670 SUB 3.03fF $ **FLOATING
C6235 S.n5671 SUB 0.59fF $ **FLOATING
C6236 S.n5672 SUB 0.02fF $ **FLOATING
C6237 S.n5673 SUB 0.97fF $ **FLOATING
C6238 S.t74 SUB 21.38fF
C6239 S.n5674 SUB 20.25fF $ **FLOATING
C6240 S.n5676 SUB 0.38fF $ **FLOATING
C6241 S.n5677 SUB 0.23fF $ **FLOATING
C6242 S.n5678 SUB 2.79fF $ **FLOATING
C6243 S.n5679 SUB 2.46fF $ **FLOATING
C6244 S.n5680 SUB 4.00fF $ **FLOATING
C6245 S.n5681 SUB 0.25fF $ **FLOATING
C6246 S.n5682 SUB 0.01fF $ **FLOATING
C6247 S.t2332 SUB 0.02fF
C6248 S.n5683 SUB 0.25fF $ **FLOATING
C6249 S.t1797 SUB 0.02fF
C6250 S.n5684 SUB 0.95fF $ **FLOATING
C6251 S.n5685 SUB 0.70fF $ **FLOATING
C6252 S.n5686 SUB 1.89fF $ **FLOATING
C6253 S.n5687 SUB 1.88fF $ **FLOATING
C6254 S.t1755 SUB 0.02fF
C6255 S.n5688 SUB 0.24fF $ **FLOATING
C6256 S.n5689 SUB 0.36fF $ **FLOATING
C6257 S.n5690 SUB 0.61fF $ **FLOATING
C6258 S.n5691 SUB 0.12fF $ **FLOATING
C6259 S.t1475 SUB 0.02fF
C6260 S.n5692 SUB 0.14fF $ **FLOATING
C6261 S.n5694 SUB 1.16fF $ **FLOATING
C6262 S.n5695 SUB 0.22fF $ **FLOATING
C6263 S.n5696 SUB 0.25fF $ **FLOATING
C6264 S.n5697 SUB 0.09fF $ **FLOATING
C6265 S.n5698 SUB 1.88fF $ **FLOATING
C6266 S.t927 SUB 0.02fF
C6267 S.n5699 SUB 0.24fF $ **FLOATING
C6268 S.n5700 SUB 0.91fF $ **FLOATING
C6269 S.n5701 SUB 0.05fF $ **FLOATING
C6270 S.t2150 SUB 0.02fF
C6271 S.n5702 SUB 0.12fF $ **FLOATING
C6272 S.n5703 SUB 0.14fF $ **FLOATING
C6273 S.n5705 SUB 0.78fF $ **FLOATING
C6274 S.n5706 SUB 1.94fF $ **FLOATING
C6275 S.n5707 SUB 1.88fF $ **FLOATING
C6276 S.n5708 SUB 0.12fF $ **FLOATING
C6277 S.t614 SUB 0.02fF
C6278 S.n5709 SUB 0.14fF $ **FLOATING
C6279 S.t876 SUB 0.02fF
C6280 S.n5711 SUB 0.24fF $ **FLOATING
C6281 S.n5712 SUB 0.36fF $ **FLOATING
C6282 S.n5713 SUB 0.61fF $ **FLOATING
C6283 S.n5714 SUB 1.84fF $ **FLOATING
C6284 S.n5715 SUB 2.99fF $ **FLOATING
C6285 S.t2567 SUB 0.02fF
C6286 S.n5716 SUB 0.24fF $ **FLOATING
C6287 S.n5717 SUB 0.91fF $ **FLOATING
C6288 S.n5718 SUB 0.05fF $ **FLOATING
C6289 S.t1290 SUB 0.02fF
C6290 S.n5719 SUB 0.12fF $ **FLOATING
C6291 S.n5720 SUB 0.14fF $ **FLOATING
C6292 S.n5722 SUB 1.89fF $ **FLOATING
C6293 S.n5723 SUB 1.88fF $ **FLOATING
C6294 S.t2523 SUB 0.02fF
C6295 S.n5724 SUB 0.24fF $ **FLOATING
C6296 S.n5725 SUB 0.36fF $ **FLOATING
C6297 S.n5726 SUB 0.61fF $ **FLOATING
C6298 S.n5727 SUB 0.12fF $ **FLOATING
C6299 S.t2267 SUB 0.02fF
C6300 S.n5728 SUB 0.14fF $ **FLOATING
C6301 S.n5730 SUB 1.16fF $ **FLOATING
C6302 S.n5731 SUB 0.22fF $ **FLOATING
C6303 S.n5732 SUB 0.25fF $ **FLOATING
C6304 S.n5733 SUB 0.09fF $ **FLOATING
C6305 S.n5734 SUB 1.88fF $ **FLOATING
C6306 S.t1691 SUB 0.02fF
C6307 S.n5735 SUB 0.24fF $ **FLOATING
C6308 S.n5736 SUB 0.91fF $ **FLOATING
C6309 S.n5737 SUB 0.05fF $ **FLOATING
C6310 S.t558 SUB 0.02fF
C6311 S.n5738 SUB 0.12fF $ **FLOATING
C6312 S.n5739 SUB 0.14fF $ **FLOATING
C6313 S.n5741 SUB 0.78fF $ **FLOATING
C6314 S.n5742 SUB 1.94fF $ **FLOATING
C6315 S.n5743 SUB 1.88fF $ **FLOATING
C6316 S.n5744 SUB 0.12fF $ **FLOATING
C6317 S.t1408 SUB 0.02fF
C6318 S.n5745 SUB 0.14fF $ **FLOATING
C6319 S.t1648 SUB 0.02fF
C6320 S.n5747 SUB 0.24fF $ **FLOATING
C6321 S.n5748 SUB 0.36fF $ **FLOATING
C6322 S.n5749 SUB 0.61fF $ **FLOATING
C6323 S.n5750 SUB 1.84fF $ **FLOATING
C6324 S.n5751 SUB 2.99fF $ **FLOATING
C6325 S.t821 SUB 0.02fF
C6326 S.n5752 SUB 0.24fF $ **FLOATING
C6327 S.n5753 SUB 0.91fF $ **FLOATING
C6328 S.n5754 SUB 0.05fF $ **FLOATING
C6329 S.t2198 SUB 0.02fF
C6330 S.n5755 SUB 0.12fF $ **FLOATING
C6331 S.n5756 SUB 0.14fF $ **FLOATING
C6332 S.n5758 SUB 1.89fF $ **FLOATING
C6333 S.n5759 SUB 1.88fF $ **FLOATING
C6334 S.t776 SUB 0.02fF
C6335 S.n5760 SUB 0.24fF $ **FLOATING
C6336 S.n5761 SUB 0.36fF $ **FLOATING
C6337 S.n5762 SUB 0.61fF $ **FLOATING
C6338 S.n5763 SUB 0.12fF $ **FLOATING
C6339 S.t541 SUB 0.02fF
C6340 S.n5764 SUB 0.14fF $ **FLOATING
C6341 S.n5766 SUB 1.16fF $ **FLOATING
C6342 S.n5767 SUB 0.22fF $ **FLOATING
C6343 S.n5768 SUB 0.25fF $ **FLOATING
C6344 S.n5769 SUB 0.09fF $ **FLOATING
C6345 S.n5770 SUB 1.88fF $ **FLOATING
C6346 S.t2466 SUB 0.02fF
C6347 S.n5771 SUB 0.24fF $ **FLOATING
C6348 S.n5772 SUB 0.91fF $ **FLOATING
C6349 S.n5773 SUB 0.05fF $ **FLOATING
C6350 S.t1340 SUB 0.02fF
C6351 S.n5774 SUB 0.12fF $ **FLOATING
C6352 S.n5775 SUB 0.14fF $ **FLOATING
C6353 S.n5777 SUB 0.78fF $ **FLOATING
C6354 S.n5778 SUB 1.94fF $ **FLOATING
C6355 S.n5779 SUB 1.88fF $ **FLOATING
C6356 S.n5780 SUB 0.12fF $ **FLOATING
C6357 S.t2182 SUB 0.02fF
C6358 S.n5781 SUB 0.14fF $ **FLOATING
C6359 S.t2428 SUB 0.02fF
C6360 S.n5783 SUB 0.24fF $ **FLOATING
C6361 S.n5784 SUB 0.36fF $ **FLOATING
C6362 S.n5785 SUB 0.61fF $ **FLOATING
C6363 S.n5786 SUB 1.84fF $ **FLOATING
C6364 S.n5787 SUB 2.99fF $ **FLOATING
C6365 S.t1597 SUB 0.02fF
C6366 S.n5788 SUB 0.24fF $ **FLOATING
C6367 S.n5789 SUB 0.91fF $ **FLOATING
C6368 S.n5790 SUB 0.05fF $ **FLOATING
C6369 S.t461 SUB 0.02fF
C6370 S.n5791 SUB 0.12fF $ **FLOATING
C6371 S.n5792 SUB 0.14fF $ **FLOATING
C6372 S.n5794 SUB 1.89fF $ **FLOATING
C6373 S.n5795 SUB 1.75fF $ **FLOATING
C6374 S.t1562 SUB 0.02fF
C6375 S.n5796 SUB 0.24fF $ **FLOATING
C6376 S.n5797 SUB 0.36fF $ **FLOATING
C6377 S.n5798 SUB 0.61fF $ **FLOATING
C6378 S.n5799 SUB 0.12fF $ **FLOATING
C6379 S.t1445 SUB 0.02fF
C6380 S.n5800 SUB 0.14fF $ **FLOATING
C6381 S.n5802 SUB 1.16fF $ **FLOATING
C6382 S.n5803 SUB 0.22fF $ **FLOATING
C6383 S.n5804 SUB 0.25fF $ **FLOATING
C6384 S.n5805 SUB 0.09fF $ **FLOATING
C6385 S.n5806 SUB 2.44fF $ **FLOATING
C6386 S.t733 SUB 0.02fF
C6387 S.n5807 SUB 0.24fF $ **FLOATING
C6388 S.n5808 SUB 0.91fF $ **FLOATING
C6389 S.n5809 SUB 0.05fF $ **FLOATING
C6390 S.t2106 SUB 0.02fF
C6391 S.n5810 SUB 0.12fF $ **FLOATING
C6392 S.n5811 SUB 0.14fF $ **FLOATING
C6393 S.n5813 SUB 1.88fF $ **FLOATING
C6394 S.n5814 SUB 0.48fF $ **FLOATING
C6395 S.n5815 SUB 0.09fF $ **FLOATING
C6396 S.n5816 SUB 0.33fF $ **FLOATING
C6397 S.n5817 SUB 0.30fF $ **FLOATING
C6398 S.n5818 SUB 0.77fF $ **FLOATING
C6399 S.n5819 SUB 0.59fF $ **FLOATING
C6400 S.t1664 SUB 0.02fF
C6401 S.n5820 SUB 0.24fF $ **FLOATING
C6402 S.n5821 SUB 0.36fF $ **FLOATING
C6403 S.n5822 SUB 0.61fF $ **FLOATING
C6404 S.n5823 SUB 0.12fF $ **FLOATING
C6405 S.t2398 SUB 0.02fF
C6406 S.n5824 SUB 0.14fF $ **FLOATING
C6407 S.n5826 SUB 2.61fF $ **FLOATING
C6408 S.n5827 SUB 2.16fF $ **FLOATING
C6409 S.t973 SUB 0.02fF
C6410 S.n5828 SUB 0.24fF $ **FLOATING
C6411 S.n5829 SUB 0.91fF $ **FLOATING
C6412 S.n5830 SUB 0.05fF $ **FLOATING
C6413 S.t1239 SUB 0.02fF
C6414 S.n5831 SUB 0.12fF $ **FLOATING
C6415 S.n5832 SUB 0.14fF $ **FLOATING
C6416 S.n5834 SUB 0.78fF $ **FLOATING
C6417 S.n5835 SUB 2.30fF $ **FLOATING
C6418 S.n5836 SUB 1.88fF $ **FLOATING
C6419 S.n5837 SUB 0.12fF $ **FLOATING
C6420 S.t1536 SUB 0.02fF
C6421 S.n5838 SUB 0.14fF $ **FLOATING
C6422 S.t792 SUB 0.02fF
C6423 S.n5840 SUB 0.24fF $ **FLOATING
C6424 S.n5841 SUB 0.36fF $ **FLOATING
C6425 S.n5842 SUB 0.61fF $ **FLOATING
C6426 S.n5843 SUB 1.39fF $ **FLOATING
C6427 S.n5844 SUB 0.71fF $ **FLOATING
C6428 S.n5845 SUB 1.14fF $ **FLOATING
C6429 S.n5846 SUB 0.35fF $ **FLOATING
C6430 S.n5847 SUB 2.03fF $ **FLOATING
C6431 S.t39 SUB 0.02fF
C6432 S.n5848 SUB 0.24fF $ **FLOATING
C6433 S.n5849 SUB 0.91fF $ **FLOATING
C6434 S.n5850 SUB 0.05fF $ **FLOATING
C6435 S.t2242 SUB 0.02fF
C6436 S.n5851 SUB 0.12fF $ **FLOATING
C6437 S.n5852 SUB 0.14fF $ **FLOATING
C6438 S.n5854 SUB 1.89fF $ **FLOATING
C6439 S.n5855 SUB 1.88fF $ **FLOATING
C6440 S.t2441 SUB 0.02fF
C6441 S.n5856 SUB 0.24fF $ **FLOATING
C6442 S.n5857 SUB 0.36fF $ **FLOATING
C6443 S.n5858 SUB 0.61fF $ **FLOATING
C6444 S.n5859 SUB 0.12fF $ **FLOATING
C6445 S.t676 SUB 0.02fF
C6446 S.n5860 SUB 0.14fF $ **FLOATING
C6447 S.n5862 SUB 1.16fF $ **FLOATING
C6448 S.n5863 SUB 0.22fF $ **FLOATING
C6449 S.n5864 SUB 0.25fF $ **FLOATING
C6450 S.n5865 SUB 0.09fF $ **FLOATING
C6451 S.n5866 SUB 1.88fF $ **FLOATING
C6452 S.t1734 SUB 0.02fF
C6453 S.n5867 SUB 0.24fF $ **FLOATING
C6454 S.n5868 SUB 0.91fF $ **FLOATING
C6455 S.n5869 SUB 0.05fF $ **FLOATING
C6456 S.t1383 SUB 0.02fF
C6457 S.n5870 SUB 0.12fF $ **FLOATING
C6458 S.n5871 SUB 0.14fF $ **FLOATING
C6459 S.n5873 SUB 20.78fF $ **FLOATING
C6460 S.n5874 SUB 1.88fF $ **FLOATING
C6461 S.n5875 SUB 2.67fF $ **FLOATING
C6462 S.t2365 SUB 0.02fF
C6463 S.n5876 SUB 0.24fF $ **FLOATING
C6464 S.n5877 SUB 0.36fF $ **FLOATING
C6465 S.n5878 SUB 0.61fF $ **FLOATING
C6466 S.n5879 SUB 0.12fF $ **FLOATING
C6467 S.t615 SUB 0.02fF
C6468 S.n5880 SUB 0.14fF $ **FLOATING
C6469 S.n5882 SUB 2.80fF $ **FLOATING
C6470 S.n5883 SUB 2.30fF $ **FLOATING
C6471 S.t1428 SUB 0.02fF
C6472 S.n5884 SUB 0.12fF $ **FLOATING
C6473 S.n5885 SUB 0.14fF $ **FLOATING
C6474 S.t1630 SUB 0.02fF
C6475 S.n5887 SUB 0.24fF $ **FLOATING
C6476 S.n5888 SUB 0.91fF $ **FLOATING
C6477 S.n5889 SUB 0.05fF $ **FLOATING
C6478 S.n5890 SUB 1.88fF $ **FLOATING
C6479 S.n5891 SUB 2.67fF $ **FLOATING
C6480 S.t1509 SUB 0.02fF
C6481 S.n5892 SUB 0.24fF $ **FLOATING
C6482 S.n5893 SUB 0.36fF $ **FLOATING
C6483 S.n5894 SUB 0.61fF $ **FLOATING
C6484 S.n5895 SUB 0.12fF $ **FLOATING
C6485 S.t2270 SUB 0.02fF
C6486 S.n5896 SUB 0.14fF $ **FLOATING
C6487 S.n5898 SUB 2.80fF $ **FLOATING
C6488 S.n5899 SUB 2.30fF $ **FLOATING
C6489 S.t563 SUB 0.02fF
C6490 S.n5900 SUB 0.12fF $ **FLOATING
C6491 S.n5901 SUB 0.14fF $ **FLOATING
C6492 S.t764 SUB 0.02fF
C6493 S.n5903 SUB 0.24fF $ **FLOATING
C6494 S.n5904 SUB 0.91fF $ **FLOATING
C6495 S.n5905 SUB 0.05fF $ **FLOATING
C6496 S.n5906 SUB 1.88fF $ **FLOATING
C6497 S.n5907 SUB 2.67fF $ **FLOATING
C6498 S.t649 SUB 0.02fF
C6499 S.n5908 SUB 0.24fF $ **FLOATING
C6500 S.n5909 SUB 0.36fF $ **FLOATING
C6501 S.n5910 SUB 0.61fF $ **FLOATING
C6502 S.n5911 SUB 0.12fF $ **FLOATING
C6503 S.t1414 SUB 0.02fF
C6504 S.n5912 SUB 0.14fF $ **FLOATING
C6505 S.n5914 SUB 2.80fF $ **FLOATING
C6506 S.n5915 SUB 2.30fF $ **FLOATING
C6507 S.t2202 SUB 0.02fF
C6508 S.n5916 SUB 0.12fF $ **FLOATING
C6509 S.n5917 SUB 0.14fF $ **FLOATING
C6510 S.t2416 SUB 0.02fF
C6511 S.n5919 SUB 0.24fF $ **FLOATING
C6512 S.n5920 SUB 0.91fF $ **FLOATING
C6513 S.n5921 SUB 0.05fF $ **FLOATING
C6514 S.n5922 SUB 2.73fF $ **FLOATING
C6515 S.n5923 SUB 1.59fF $ **FLOATING
C6516 S.n5924 SUB 0.12fF $ **FLOATING
C6517 S.t1622 SUB 0.02fF
C6518 S.n5925 SUB 0.14fF $ **FLOATING
C6519 S.t1537 SUB 0.02fF
C6520 S.n5927 SUB 0.24fF $ **FLOATING
C6521 S.n5928 SUB 0.36fF $ **FLOATING
C6522 S.n5929 SUB 0.61fF $ **FLOATING
C6523 S.n5930 SUB 0.07fF $ **FLOATING
C6524 S.n5931 SUB 0.01fF $ **FLOATING
C6525 S.n5932 SUB 0.24fF $ **FLOATING
C6526 S.n5933 SUB 1.16fF $ **FLOATING
C6527 S.n5934 SUB 1.35fF $ **FLOATING
C6528 S.n5935 SUB 2.30fF $ **FLOATING
C6529 S.t2376 SUB 0.02fF
C6530 S.n5936 SUB 0.12fF $ **FLOATING
C6531 S.n5937 SUB 0.14fF $ **FLOATING
C6532 S.t2515 SUB 0.02fF
C6533 S.n5939 SUB 0.24fF $ **FLOATING
C6534 S.n5940 SUB 0.91fF $ **FLOATING
C6535 S.n5941 SUB 0.05fF $ **FLOATING
C6536 S.t460 SUB 48.31fF
C6537 S.t1552 SUB 0.02fF
C6538 S.n5942 SUB 0.24fF $ **FLOATING
C6539 S.n5943 SUB 0.91fF $ **FLOATING
C6540 S.n5944 SUB 0.05fF $ **FLOATING
C6541 S.t1345 SUB 0.02fF
C6542 S.n5945 SUB 0.12fF $ **FLOATING
C6543 S.n5946 SUB 0.14fF $ **FLOATING
C6544 S.n5948 SUB 0.12fF $ **FLOATING
C6545 S.t549 SUB 0.02fF
C6546 S.n5949 SUB 0.14fF $ **FLOATING
C6547 S.n5951 SUB 5.17fF $ **FLOATING
C6548 S.n5952 SUB 5.44fF $ **FLOATING
C6549 S.t425 SUB 0.02fF
C6550 S.n5953 SUB 0.12fF $ **FLOATING
C6551 S.n5954 SUB 0.14fF $ **FLOATING
C6552 S.t1885 SUB 0.02fF
C6553 S.n5956 SUB 0.24fF $ **FLOATING
C6554 S.n5957 SUB 0.91fF $ **FLOATING
C6555 S.n5958 SUB 0.05fF $ **FLOATING
C6556 S.t390 SUB 47.92fF
C6557 S.t872 SUB 0.02fF
C6558 S.n5959 SUB 1.19fF $ **FLOATING
C6559 S.n5960 SUB 0.05fF $ **FLOATING
C6560 S.t429 SUB 0.02fF
C6561 S.n5961 SUB 0.01fF $ **FLOATING
C6562 S.n5962 SUB 0.26fF $ **FLOATING
C6563 S.n5964 SUB 1.50fF $ **FLOATING
C6564 S.n5965 SUB 1.30fF $ **FLOATING
C6565 S.n5966 SUB 0.28fF $ **FLOATING
C6566 S.n5967 SUB 0.24fF $ **FLOATING
C6567 S.n5968 SUB 4.39fF $ **FLOATING
C6568 S.n5969 SUB 0.01fF $ **FLOATING
C6569 S.n5970 SUB 0.02fF $ **FLOATING
C6570 S.n5971 SUB 0.03fF $ **FLOATING
C6571 S.n5972 SUB 0.04fF $ **FLOATING
C6572 S.n5973 SUB 0.17fF $ **FLOATING
C6573 S.n5974 SUB 0.01fF $ **FLOATING
C6574 S.n5975 SUB 0.02fF $ **FLOATING
C6575 S.n5976 SUB 0.01fF $ **FLOATING
C6576 S.n5977 SUB 0.01fF $ **FLOATING
C6577 S.n5978 SUB 0.01fF $ **FLOATING
C6578 S.n5979 SUB 0.01fF $ **FLOATING
C6579 S.n5980 SUB 0.02fF $ **FLOATING
C6580 S.n5981 SUB 0.01fF $ **FLOATING
C6581 S.n5982 SUB 0.02fF $ **FLOATING
C6582 S.n5983 SUB 0.05fF $ **FLOATING
C6583 S.n5984 SUB 0.04fF $ **FLOATING
C6584 S.n5985 SUB 0.11fF $ **FLOATING
C6585 S.n5986 SUB 0.38fF $ **FLOATING
C6586 S.n5987 SUB 0.20fF $ **FLOATING
C6587 S.n5988 SUB 8.97fF $ **FLOATING
C6588 S.n5989 SUB 8.97fF $ **FLOATING
C6589 S.n5990 SUB 0.60fF $ **FLOATING
C6590 S.n5991 SUB 0.22fF $ **FLOATING
C6591 S.n5992 SUB 0.59fF $ **FLOATING
C6592 S.n5993 SUB 3.43fF $ **FLOATING
C6593 S.n5994 SUB 0.29fF $ **FLOATING
C6594 S.t69 SUB 21.38fF
C6595 S.n5995 SUB 21.67fF $ **FLOATING
C6596 S.n5996 SUB 0.77fF $ **FLOATING
C6597 S.n5997 SUB 0.28fF $ **FLOATING
C6598 S.n5998 SUB 4.00fF $ **FLOATING
C6599 S.n5999 SUB 1.35fF $ **FLOATING
C6600 S.t1014 SUB 0.02fF
C6601 S.n6000 SUB 0.64fF $ **FLOATING
C6602 S.n6001 SUB 0.61fF $ **FLOATING
C6603 S.n6002 SUB 0.25fF $ **FLOATING
C6604 S.n6003 SUB 0.09fF $ **FLOATING
C6605 S.n6004 SUB 0.21fF $ **FLOATING
C6606 S.n6005 SUB 0.92fF $ **FLOATING
C6607 S.n6006 SUB 0.44fF $ **FLOATING
C6608 S.n6007 SUB 1.88fF $ **FLOATING
C6609 S.n6008 SUB 0.12fF $ **FLOATING
C6610 S.t1841 SUB 0.02fF
C6611 S.n6009 SUB 0.14fF $ **FLOATING
C6612 S.t2345 SUB 0.02fF
C6613 S.n6011 SUB 0.24fF $ **FLOATING
C6614 S.n6012 SUB 0.36fF $ **FLOATING
C6615 S.n6013 SUB 0.61fF $ **FLOATING
C6616 S.n6014 SUB 0.02fF $ **FLOATING
C6617 S.n6015 SUB 0.01fF $ **FLOATING
C6618 S.n6016 SUB 0.02fF $ **FLOATING
C6619 S.n6017 SUB 0.08fF $ **FLOATING
C6620 S.n6018 SUB 0.06fF $ **FLOATING
C6621 S.n6019 SUB 0.03fF $ **FLOATING
C6622 S.n6020 SUB 0.04fF $ **FLOATING
C6623 S.n6021 SUB 1.00fF $ **FLOATING
C6624 S.n6022 SUB 0.36fF $ **FLOATING
C6625 S.n6023 SUB 1.87fF $ **FLOATING
C6626 S.n6024 SUB 1.99fF $ **FLOATING
C6627 S.t972 SUB 0.02fF
C6628 S.n6025 SUB 0.24fF $ **FLOATING
C6629 S.n6026 SUB 0.91fF $ **FLOATING
C6630 S.n6027 SUB 0.05fF $ **FLOATING
C6631 S.t2008 SUB 0.02fF
C6632 S.n6028 SUB 0.12fF $ **FLOATING
C6633 S.n6029 SUB 0.14fF $ **FLOATING
C6634 S.n6031 SUB 1.89fF $ **FLOATING
C6635 S.n6032 SUB 0.06fF $ **FLOATING
C6636 S.n6033 SUB 0.03fF $ **FLOATING
C6637 S.n6034 SUB 0.04fF $ **FLOATING
C6638 S.n6035 SUB 0.99fF $ **FLOATING
C6639 S.n6036 SUB 0.02fF $ **FLOATING
C6640 S.n6037 SUB 0.01fF $ **FLOATING
C6641 S.n6038 SUB 0.02fF $ **FLOATING
C6642 S.n6039 SUB 0.08fF $ **FLOATING
C6643 S.n6040 SUB 0.36fF $ **FLOATING
C6644 S.n6041 SUB 1.85fF $ **FLOATING
C6645 S.t1588 SUB 0.02fF
C6646 S.n6042 SUB 0.24fF $ **FLOATING
C6647 S.n6043 SUB 0.36fF $ **FLOATING
C6648 S.n6044 SUB 0.61fF $ **FLOATING
C6649 S.n6045 SUB 0.12fF $ **FLOATING
C6650 S.t1096 SUB 0.02fF
C6651 S.n6046 SUB 0.14fF $ **FLOATING
C6652 S.n6048 SUB 0.70fF $ **FLOATING
C6653 S.n6049 SUB 0.23fF $ **FLOATING
C6654 S.n6050 SUB 0.23fF $ **FLOATING
C6655 S.n6051 SUB 0.70fF $ **FLOATING
C6656 S.n6052 SUB 1.16fF $ **FLOATING
C6657 S.n6053 SUB 0.22fF $ **FLOATING
C6658 S.n6054 SUB 0.25fF $ **FLOATING
C6659 S.n6055 SUB 0.09fF $ **FLOATING
C6660 S.n6056 SUB 1.88fF $ **FLOATING
C6661 S.t217 SUB 0.02fF
C6662 S.n6057 SUB 0.24fF $ **FLOATING
C6663 S.n6058 SUB 0.91fF $ **FLOATING
C6664 S.n6059 SUB 0.05fF $ **FLOATING
C6665 S.t1155 SUB 0.02fF
C6666 S.n6060 SUB 0.12fF $ **FLOATING
C6667 S.n6061 SUB 0.14fF $ **FLOATING
C6668 S.n6063 SUB 0.25fF $ **FLOATING
C6669 S.n6064 SUB 0.09fF $ **FLOATING
C6670 S.n6065 SUB 0.21fF $ **FLOATING
C6671 S.n6066 SUB 0.92fF $ **FLOATING
C6672 S.n6067 SUB 0.44fF $ **FLOATING
C6673 S.n6068 SUB 1.88fF $ **FLOATING
C6674 S.n6069 SUB 0.12fF $ **FLOATING
C6675 S.t221 SUB 0.02fF
C6676 S.n6070 SUB 0.14fF $ **FLOATING
C6677 S.t723 SUB 0.02fF
C6678 S.n6072 SUB 0.24fF $ **FLOATING
C6679 S.n6073 SUB 0.36fF $ **FLOATING
C6680 S.n6074 SUB 0.61fF $ **FLOATING
C6681 S.n6075 SUB 0.02fF $ **FLOATING
C6682 S.n6076 SUB 0.01fF $ **FLOATING
C6683 S.n6077 SUB 0.02fF $ **FLOATING
C6684 S.n6078 SUB 0.08fF $ **FLOATING
C6685 S.n6079 SUB 0.06fF $ **FLOATING
C6686 S.n6080 SUB 0.03fF $ **FLOATING
C6687 S.n6081 SUB 0.04fF $ **FLOATING
C6688 S.n6082 SUB 1.00fF $ **FLOATING
C6689 S.n6083 SUB 0.36fF $ **FLOATING
C6690 S.n6084 SUB 1.87fF $ **FLOATING
C6691 S.n6085 SUB 1.99fF $ **FLOATING
C6692 S.t1882 SUB 0.02fF
C6693 S.n6086 SUB 0.24fF $ **FLOATING
C6694 S.n6087 SUB 0.91fF $ **FLOATING
C6695 S.n6088 SUB 0.05fF $ **FLOATING
C6696 S.t280 SUB 0.02fF
C6697 S.n6089 SUB 0.12fF $ **FLOATING
C6698 S.n6090 SUB 0.14fF $ **FLOATING
C6699 S.n6092 SUB 1.89fF $ **FLOATING
C6700 S.n6093 SUB 0.06fF $ **FLOATING
C6701 S.n6094 SUB 0.03fF $ **FLOATING
C6702 S.n6095 SUB 0.04fF $ **FLOATING
C6703 S.n6096 SUB 0.99fF $ **FLOATING
C6704 S.n6097 SUB 0.02fF $ **FLOATING
C6705 S.n6098 SUB 0.01fF $ **FLOATING
C6706 S.n6099 SUB 0.02fF $ **FLOATING
C6707 S.n6100 SUB 0.08fF $ **FLOATING
C6708 S.n6101 SUB 0.36fF $ **FLOATING
C6709 S.n6102 SUB 1.85fF $ **FLOATING
C6710 S.t2377 SUB 0.02fF
C6711 S.n6103 SUB 0.24fF $ **FLOATING
C6712 S.n6104 SUB 0.36fF $ **FLOATING
C6713 S.n6105 SUB 0.61fF $ **FLOATING
C6714 S.n6106 SUB 0.12fF $ **FLOATING
C6715 S.t1886 SUB 0.02fF
C6716 S.n6107 SUB 0.14fF $ **FLOATING
C6717 S.n6109 SUB 0.70fF $ **FLOATING
C6718 S.n6110 SUB 0.23fF $ **FLOATING
C6719 S.n6111 SUB 0.23fF $ **FLOATING
C6720 S.n6112 SUB 0.70fF $ **FLOATING
C6721 S.n6113 SUB 1.16fF $ **FLOATING
C6722 S.n6114 SUB 0.22fF $ **FLOATING
C6723 S.n6115 SUB 0.25fF $ **FLOATING
C6724 S.n6116 SUB 0.09fF $ **FLOATING
C6725 S.n6117 SUB 1.88fF $ **FLOATING
C6726 S.t1021 SUB 0.02fF
C6727 S.n6118 SUB 0.24fF $ **FLOATING
C6728 S.n6119 SUB 0.91fF $ **FLOATING
C6729 S.n6120 SUB 0.05fF $ **FLOATING
C6730 S.t1939 SUB 0.02fF
C6731 S.n6121 SUB 0.12fF $ **FLOATING
C6732 S.n6122 SUB 0.14fF $ **FLOATING
C6733 S.n6124 SUB 0.25fF $ **FLOATING
C6734 S.n6125 SUB 0.09fF $ **FLOATING
C6735 S.n6126 SUB 0.21fF $ **FLOATING
C6736 S.n6127 SUB 0.92fF $ **FLOATING
C6737 S.n6128 SUB 0.44fF $ **FLOATING
C6738 S.n6129 SUB 1.88fF $ **FLOATING
C6739 S.n6130 SUB 0.12fF $ **FLOATING
C6740 S.t1023 SUB 0.02fF
C6741 S.n6131 SUB 0.14fF $ **FLOATING
C6742 S.t1520 SUB 0.02fF
C6743 S.n6133 SUB 0.24fF $ **FLOATING
C6744 S.n6134 SUB 0.36fF $ **FLOATING
C6745 S.n6135 SUB 0.61fF $ **FLOATING
C6746 S.n6136 SUB 0.02fF $ **FLOATING
C6747 S.n6137 SUB 0.01fF $ **FLOATING
C6748 S.n6138 SUB 0.02fF $ **FLOATING
C6749 S.n6139 SUB 0.08fF $ **FLOATING
C6750 S.n6140 SUB 0.06fF $ **FLOATING
C6751 S.n6141 SUB 0.03fF $ **FLOATING
C6752 S.n6142 SUB 0.04fF $ **FLOATING
C6753 S.n6143 SUB 1.00fF $ **FLOATING
C6754 S.n6144 SUB 0.36fF $ **FLOATING
C6755 S.n6145 SUB 1.87fF $ **FLOATING
C6756 S.n6146 SUB 1.99fF $ **FLOATING
C6757 S.t118 SUB 0.02fF
C6758 S.n6147 SUB 0.24fF $ **FLOATING
C6759 S.n6148 SUB 0.91fF $ **FLOATING
C6760 S.n6149 SUB 0.05fF $ **FLOATING
C6761 S.t1082 SUB 0.02fF
C6762 S.n6150 SUB 0.12fF $ **FLOATING
C6763 S.n6151 SUB 0.14fF $ **FLOATING
C6764 S.n6153 SUB 1.89fF $ **FLOATING
C6765 S.n6154 SUB 0.04fF $ **FLOATING
C6766 S.n6155 SUB 0.07fF $ **FLOATING
C6767 S.n6156 SUB 0.05fF $ **FLOATING
C6768 S.n6157 SUB 0.87fF $ **FLOATING
C6769 S.n6158 SUB 0.01fF $ **FLOATING
C6770 S.n6159 SUB 0.01fF $ **FLOATING
C6771 S.n6160 SUB 0.01fF $ **FLOATING
C6772 S.n6161 SUB 0.07fF $ **FLOATING
C6773 S.n6162 SUB 0.68fF $ **FLOATING
C6774 S.n6163 SUB 0.72fF $ **FLOATING
C6775 S.t660 SUB 0.02fF
C6776 S.n6164 SUB 0.24fF $ **FLOATING
C6777 S.n6165 SUB 0.36fF $ **FLOATING
C6778 S.n6166 SUB 0.61fF $ **FLOATING
C6779 S.n6167 SUB 0.12fF $ **FLOATING
C6780 S.t120 SUB 0.02fF
C6781 S.n6168 SUB 0.14fF $ **FLOATING
C6782 S.n6170 SUB 0.70fF $ **FLOATING
C6783 S.n6171 SUB 0.23fF $ **FLOATING
C6784 S.n6172 SUB 0.23fF $ **FLOATING
C6785 S.n6173 SUB 0.70fF $ **FLOATING
C6786 S.n6174 SUB 1.16fF $ **FLOATING
C6787 S.n6175 SUB 0.22fF $ **FLOATING
C6788 S.n6176 SUB 0.25fF $ **FLOATING
C6789 S.n6177 SUB 0.09fF $ **FLOATING
C6790 S.n6178 SUB 2.31fF $ **FLOATING
C6791 S.t1790 SUB 0.02fF
C6792 S.n6179 SUB 0.24fF $ **FLOATING
C6793 S.n6180 SUB 0.91fF $ **FLOATING
C6794 S.n6181 SUB 0.05fF $ **FLOATING
C6795 S.t205 SUB 0.02fF
C6796 S.n6182 SUB 0.12fF $ **FLOATING
C6797 S.n6183 SUB 0.14fF $ **FLOATING
C6798 S.n6185 SUB 1.88fF $ **FLOATING
C6799 S.n6186 SUB 0.46fF $ **FLOATING
C6800 S.n6187 SUB 0.22fF $ **FLOATING
C6801 S.n6188 SUB 0.38fF $ **FLOATING
C6802 S.n6189 SUB 0.16fF $ **FLOATING
C6803 S.n6190 SUB 0.28fF $ **FLOATING
C6804 S.n6191 SUB 0.21fF $ **FLOATING
C6805 S.n6192 SUB 0.30fF $ **FLOATING
C6806 S.n6193 SUB 0.42fF $ **FLOATING
C6807 S.n6194 SUB 0.21fF $ **FLOATING
C6808 S.t2315 SUB 0.02fF
C6809 S.n6195 SUB 0.24fF $ **FLOATING
C6810 S.n6196 SUB 0.36fF $ **FLOATING
C6811 S.n6197 SUB 0.61fF $ **FLOATING
C6812 S.n6198 SUB 0.12fF $ **FLOATING
C6813 S.t1791 SUB 0.02fF
C6814 S.n6199 SUB 0.14fF $ **FLOATING
C6815 S.n6201 SUB 0.04fF $ **FLOATING
C6816 S.n6202 SUB 0.03fF $ **FLOATING
C6817 S.n6203 SUB 0.03fF $ **FLOATING
C6818 S.n6204 SUB 0.10fF $ **FLOATING
C6819 S.n6205 SUB 0.36fF $ **FLOATING
C6820 S.n6206 SUB 0.38fF $ **FLOATING
C6821 S.n6207 SUB 0.11fF $ **FLOATING
C6822 S.n6208 SUB 0.12fF $ **FLOATING
C6823 S.n6209 SUB 0.07fF $ **FLOATING
C6824 S.n6210 SUB 0.12fF $ **FLOATING
C6825 S.n6211 SUB 0.18fF $ **FLOATING
C6826 S.n6212 SUB 4.00fF $ **FLOATING
C6827 S.t921 SUB 0.02fF
C6828 S.n6213 SUB 0.24fF $ **FLOATING
C6829 S.n6214 SUB 0.91fF $ **FLOATING
C6830 S.n6215 SUB 0.05fF $ **FLOATING
C6831 S.t1979 SUB 0.02fF
C6832 S.n6216 SUB 0.12fF $ **FLOATING
C6833 S.n6217 SUB 0.14fF $ **FLOATING
C6834 S.n6219 SUB 0.25fF $ **FLOATING
C6835 S.n6220 SUB 0.09fF $ **FLOATING
C6836 S.n6221 SUB 0.21fF $ **FLOATING
C6837 S.n6222 SUB 1.28fF $ **FLOATING
C6838 S.n6223 SUB 0.53fF $ **FLOATING
C6839 S.n6224 SUB 1.88fF $ **FLOATING
C6840 S.n6225 SUB 0.12fF $ **FLOATING
C6841 S.t1303 SUB 0.02fF
C6842 S.n6226 SUB 0.14fF $ **FLOATING
C6843 S.t1851 SUB 0.02fF
C6844 S.n6228 SUB 0.24fF $ **FLOATING
C6845 S.n6229 SUB 0.36fF $ **FLOATING
C6846 S.n6230 SUB 0.61fF $ **FLOATING
C6847 S.n6231 SUB 1.58fF $ **FLOATING
C6848 S.n6232 SUB 2.45fF $ **FLOATING
C6849 S.t874 SUB 0.02fF
C6850 S.n6233 SUB 0.24fF $ **FLOATING
C6851 S.n6234 SUB 0.91fF $ **FLOATING
C6852 S.n6235 SUB 0.05fF $ **FLOATING
C6853 S.t1485 SUB 0.02fF
C6854 S.n6236 SUB 0.12fF $ **FLOATING
C6855 S.n6237 SUB 0.14fF $ **FLOATING
C6856 S.n6239 SUB 1.89fF $ **FLOATING
C6857 S.n6240 SUB 0.06fF $ **FLOATING
C6858 S.n6241 SUB 0.03fF $ **FLOATING
C6859 S.n6242 SUB 0.04fF $ **FLOATING
C6860 S.n6243 SUB 0.99fF $ **FLOATING
C6861 S.n6244 SUB 0.02fF $ **FLOATING
C6862 S.n6245 SUB 0.01fF $ **FLOATING
C6863 S.n6246 SUB 0.02fF $ **FLOATING
C6864 S.n6247 SUB 0.08fF $ **FLOATING
C6865 S.n6248 SUB 0.36fF $ **FLOATING
C6866 S.n6249 SUB 1.85fF $ **FLOATING
C6867 S.t988 SUB 0.02fF
C6868 S.n6250 SUB 0.24fF $ **FLOATING
C6869 S.n6251 SUB 0.36fF $ **FLOATING
C6870 S.n6252 SUB 0.61fF $ **FLOATING
C6871 S.n6253 SUB 0.12fF $ **FLOATING
C6872 S.t419 SUB 0.02fF
C6873 S.n6254 SUB 0.14fF $ **FLOATING
C6874 S.n6256 SUB 0.70fF $ **FLOATING
C6875 S.n6257 SUB 0.23fF $ **FLOATING
C6876 S.n6258 SUB 0.23fF $ **FLOATING
C6877 S.n6259 SUB 0.70fF $ **FLOATING
C6878 S.n6260 SUB 1.16fF $ **FLOATING
C6879 S.n6261 SUB 0.22fF $ **FLOATING
C6880 S.n6262 SUB 0.25fF $ **FLOATING
C6881 S.n6263 SUB 0.09fF $ **FLOATING
C6882 S.n6264 SUB 1.88fF $ **FLOATING
C6883 S.t2520 SUB 0.02fF
C6884 S.n6265 SUB 0.24fF $ **FLOATING
C6885 S.n6266 SUB 0.91fF $ **FLOATING
C6886 S.n6267 SUB 0.05fF $ **FLOATING
C6887 S.t623 SUB 0.02fF
C6888 S.n6268 SUB 0.12fF $ **FLOATING
C6889 S.n6269 SUB 0.14fF $ **FLOATING
C6890 S.n6271 SUB 20.78fF $ **FLOATING
C6891 S.n6272 SUB 1.72fF $ **FLOATING
C6892 S.n6273 SUB 3.05fF $ **FLOATING
C6893 S.t686 SUB 0.02fF
C6894 S.n6274 SUB 0.24fF $ **FLOATING
C6895 S.n6275 SUB 0.36fF $ **FLOATING
C6896 S.n6276 SUB 0.61fF $ **FLOATING
C6897 S.n6277 SUB 0.12fF $ **FLOATING
C6898 S.t176 SUB 0.02fF
C6899 S.n6278 SUB 0.14fF $ **FLOATING
C6900 S.n6280 SUB 0.31fF $ **FLOATING
C6901 S.n6281 SUB 0.23fF $ **FLOATING
C6902 S.n6282 SUB 0.66fF $ **FLOATING
C6903 S.n6283 SUB 0.95fF $ **FLOATING
C6904 S.n6284 SUB 0.23fF $ **FLOATING
C6905 S.n6285 SUB 0.21fF $ **FLOATING
C6906 S.n6286 SUB 0.20fF $ **FLOATING
C6907 S.n6287 SUB 0.06fF $ **FLOATING
C6908 S.n6288 SUB 0.09fF $ **FLOATING
C6909 S.n6289 SUB 0.10fF $ **FLOATING
C6910 S.n6290 SUB 1.99fF $ **FLOATING
C6911 S.t351 SUB 0.02fF
C6912 S.n6291 SUB 0.12fF $ **FLOATING
C6913 S.n6292 SUB 0.14fF $ **FLOATING
C6914 S.t1838 SUB 0.02fF
C6915 S.n6294 SUB 0.24fF $ **FLOATING
C6916 S.n6295 SUB 0.91fF $ **FLOATING
C6917 S.n6296 SUB 0.05fF $ **FLOATING
C6918 S.n6297 SUB 1.88fF $ **FLOATING
C6919 S.n6298 SUB 0.12fF $ **FLOATING
C6920 S.t228 SUB 0.02fF
C6921 S.n6299 SUB 0.14fF $ **FLOATING
C6922 S.t895 SUB 0.02fF
C6923 S.n6301 SUB 0.12fF $ **FLOATING
C6924 S.n6302 SUB 0.14fF $ **FLOATING
C6925 S.t896 SUB 0.02fF
C6926 S.n6304 SUB 0.24fF $ **FLOATING
C6927 S.n6305 SUB 0.91fF $ **FLOATING
C6928 S.n6306 SUB 0.05fF $ **FLOATING
C6929 S.t1995 SUB 0.02fF
C6930 S.n6307 SUB 0.24fF $ **FLOATING
C6931 S.n6308 SUB 0.36fF $ **FLOATING
C6932 S.n6309 SUB 0.61fF $ **FLOATING
C6933 S.n6310 SUB 0.32fF $ **FLOATING
C6934 S.n6311 SUB 1.09fF $ **FLOATING
C6935 S.n6312 SUB 0.15fF $ **FLOATING
C6936 S.n6313 SUB 2.10fF $ **FLOATING
C6937 S.n6314 SUB 2.94fF $ **FLOATING
C6938 S.n6315 SUB 1.88fF $ **FLOATING
C6939 S.n6316 SUB 0.12fF $ **FLOATING
C6940 S.t2070 SUB 0.02fF
C6941 S.n6317 SUB 0.14fF $ **FLOATING
C6942 S.t70 SUB 0.02fF
C6943 S.n6319 SUB 0.24fF $ **FLOATING
C6944 S.n6320 SUB 0.36fF $ **FLOATING
C6945 S.n6321 SUB 0.61fF $ **FLOATING
C6946 S.n6322 SUB 0.92fF $ **FLOATING
C6947 S.n6323 SUB 0.32fF $ **FLOATING
C6948 S.n6324 SUB 0.92fF $ **FLOATING
C6949 S.n6325 SUB 1.09fF $ **FLOATING
C6950 S.n6326 SUB 0.15fF $ **FLOATING
C6951 S.n6327 SUB 4.96fF $ **FLOATING
C6952 S.t2282 SUB 0.02fF
C6953 S.n6328 SUB 0.12fF $ **FLOATING
C6954 S.n6329 SUB 0.14fF $ **FLOATING
C6955 S.t1644 SUB 0.02fF
C6956 S.n6331 SUB 0.24fF $ **FLOATING
C6957 S.n6332 SUB 0.91fF $ **FLOATING
C6958 S.n6333 SUB 0.05fF $ **FLOATING
C6959 S.n6334 SUB 1.88fF $ **FLOATING
C6960 S.n6335 SUB 2.67fF $ **FLOATING
C6961 S.t1754 SUB 0.02fF
C6962 S.n6336 SUB 0.24fF $ **FLOATING
C6963 S.n6337 SUB 0.36fF $ **FLOATING
C6964 S.n6338 SUB 0.61fF $ **FLOATING
C6965 S.n6339 SUB 0.12fF $ **FLOATING
C6966 S.t1209 SUB 0.02fF
C6967 S.n6340 SUB 0.14fF $ **FLOATING
C6968 S.n6342 SUB 1.88fF $ **FLOATING
C6969 S.n6343 SUB 2.67fF $ **FLOATING
C6970 S.t1146 SUB 0.02fF
C6971 S.n6344 SUB 0.24fF $ **FLOATING
C6972 S.n6345 SUB 0.36fF $ **FLOATING
C6973 S.n6346 SUB 0.61fF $ **FLOATING
C6974 S.t2538 SUB 0.02fF
C6975 S.n6347 SUB 0.24fF $ **FLOATING
C6976 S.n6348 SUB 0.91fF $ **FLOATING
C6977 S.n6349 SUB 0.05fF $ **FLOATING
C6978 S.t2541 SUB 0.02fF
C6979 S.n6350 SUB 0.12fF $ **FLOATING
C6980 S.n6351 SUB 0.14fF $ **FLOATING
C6981 S.n6353 SUB 0.12fF $ **FLOATING
C6982 S.t1896 SUB 0.02fF
C6983 S.n6354 SUB 0.14fF $ **FLOATING
C6984 S.n6356 SUB 2.30fF $ **FLOATING
C6985 S.n6357 SUB 2.94fF $ **FLOATING
C6986 S.n6358 SUB 5.16fF $ **FLOATING
C6987 S.t1426 SUB 0.02fF
C6988 S.n6359 SUB 0.12fF $ **FLOATING
C6989 S.n6360 SUB 0.14fF $ **FLOATING
C6990 S.t775 SUB 0.02fF
C6991 S.n6362 SUB 0.24fF $ **FLOATING
C6992 S.n6363 SUB 0.91fF $ **FLOATING
C6993 S.n6364 SUB 0.05fF $ **FLOATING
C6994 S.n6365 SUB 1.88fF $ **FLOATING
C6995 S.n6366 SUB 2.67fF $ **FLOATING
C6996 S.t1033 SUB 0.02fF
C6997 S.n6367 SUB 0.24fF $ **FLOATING
C6998 S.n6368 SUB 0.36fF $ **FLOATING
C6999 S.n6369 SUB 0.61fF $ **FLOATING
C7000 S.n6370 SUB 0.12fF $ **FLOATING
C7001 S.t476 SUB 0.02fF
C7002 S.n6371 SUB 0.14fF $ **FLOATING
C7003 S.n6373 SUB 5.17fF $ **FLOATING
C7004 S.t561 SUB 0.02fF
C7005 S.n6374 SUB 0.12fF $ **FLOATING
C7006 S.n6375 SUB 0.14fF $ **FLOATING
C7007 S.t2579 SUB 0.02fF
C7008 S.n6377 SUB 0.24fF $ **FLOATING
C7009 S.n6378 SUB 0.91fF $ **FLOATING
C7010 S.n6379 SUB 0.05fF $ **FLOATING
C7011 S.n6380 SUB 1.88fF $ **FLOATING
C7012 S.n6381 SUB 2.67fF $ **FLOATING
C7013 S.t136 SUB 0.02fF
C7014 S.n6382 SUB 0.24fF $ **FLOATING
C7015 S.n6383 SUB 0.36fF $ **FLOATING
C7016 S.n6384 SUB 0.61fF $ **FLOATING
C7017 S.n6385 SUB 0.12fF $ **FLOATING
C7018 S.t2127 SUB 0.02fF
C7019 S.n6386 SUB 0.14fF $ **FLOATING
C7020 S.n6388 SUB 5.17fF $ **FLOATING
C7021 S.t2200 SUB 0.02fF
C7022 S.n6389 SUB 0.12fF $ **FLOATING
C7023 S.n6390 SUB 0.14fF $ **FLOATING
C7024 S.t1702 SUB 0.02fF
C7025 S.n6392 SUB 0.24fF $ **FLOATING
C7026 S.n6393 SUB 0.91fF $ **FLOATING
C7027 S.n6394 SUB 0.05fF $ **FLOATING
C7028 S.n6395 SUB 1.88fF $ **FLOATING
C7029 S.n6396 SUB 2.67fF $ **FLOATING
C7030 S.t1806 SUB 0.02fF
C7031 S.n6397 SUB 0.24fF $ **FLOATING
C7032 S.n6398 SUB 0.36fF $ **FLOATING
C7033 S.n6399 SUB 0.61fF $ **FLOATING
C7034 S.n6400 SUB 0.12fF $ **FLOATING
C7035 S.t1261 SUB 0.02fF
C7036 S.n6401 SUB 0.14fF $ **FLOATING
C7037 S.n6403 SUB 5.17fF $ **FLOATING
C7038 S.t1343 SUB 0.02fF
C7039 S.n6404 SUB 0.12fF $ **FLOATING
C7040 S.n6405 SUB 0.14fF $ **FLOATING
C7041 S.t829 SUB 0.02fF
C7042 S.n6407 SUB 0.24fF $ **FLOATING
C7043 S.n6408 SUB 0.91fF $ **FLOATING
C7044 S.n6409 SUB 0.05fF $ **FLOATING
C7045 S.n6410 SUB 1.88fF $ **FLOATING
C7046 S.n6411 SUB 2.67fF $ **FLOATING
C7047 S.t941 SUB 0.02fF
C7048 S.n6412 SUB 0.24fF $ **FLOATING
C7049 S.n6413 SUB 0.36fF $ **FLOATING
C7050 S.n6414 SUB 0.61fF $ **FLOATING
C7051 S.n6415 SUB 0.12fF $ **FLOATING
C7052 S.t378 SUB 0.02fF
C7053 S.n6416 SUB 0.14fF $ **FLOATING
C7054 S.n6418 SUB 4.90fF $ **FLOATING
C7055 S.t466 SUB 0.02fF
C7056 S.n6419 SUB 0.12fF $ **FLOATING
C7057 S.n6420 SUB 0.14fF $ **FLOATING
C7058 S.t2476 SUB 0.02fF
C7059 S.n6422 SUB 0.24fF $ **FLOATING
C7060 S.n6423 SUB 0.91fF $ **FLOATING
C7061 S.n6424 SUB 0.05fF $ **FLOATING
C7062 S.n6425 SUB 1.88fF $ **FLOATING
C7063 S.n6426 SUB 2.67fF $ **FLOATING
C7064 S.t1101 SUB 0.02fF
C7065 S.n6427 SUB 0.24fF $ **FLOATING
C7066 S.n6428 SUB 0.36fF $ **FLOATING
C7067 S.n6429 SUB 0.61fF $ **FLOATING
C7068 S.n6430 SUB 0.12fF $ **FLOATING
C7069 S.t2328 SUB 0.02fF
C7070 S.n6431 SUB 0.14fF $ **FLOATING
C7071 S.n6433 SUB 1.88fF $ **FLOATING
C7072 S.n6434 SUB 2.68fF $ **FLOATING
C7073 S.t1861 SUB 0.02fF
C7074 S.n6435 SUB 0.24fF $ **FLOATING
C7075 S.n6436 SUB 0.36fF $ **FLOATING
C7076 S.n6437 SUB 0.61fF $ **FLOATING
C7077 S.t2529 SUB 0.02fF
C7078 S.n6438 SUB 1.22fF $ **FLOATING
C7079 S.n6439 SUB 0.61fF $ **FLOATING
C7080 S.n6440 SUB 0.35fF $ **FLOATING
C7081 S.n6441 SUB 0.63fF $ **FLOATING
C7082 S.n6442 SUB 1.15fF $ **FLOATING
C7083 S.n6443 SUB 3.03fF $ **FLOATING
C7084 S.n6444 SUB 0.59fF $ **FLOATING
C7085 S.n6445 SUB 0.02fF $ **FLOATING
C7086 S.n6446 SUB 0.97fF $ **FLOATING
C7087 S.t125 SUB 21.38fF
C7088 S.n6447 SUB 20.25fF $ **FLOATING
C7089 S.n6449 SUB 0.38fF $ **FLOATING
C7090 S.n6450 SUB 0.23fF $ **FLOATING
C7091 S.n6451 SUB 2.90fF $ **FLOATING
C7092 S.n6452 SUB 2.46fF $ **FLOATING
C7093 S.n6453 SUB 1.96fF $ **FLOATING
C7094 S.n6454 SUB 3.94fF $ **FLOATING
C7095 S.n6455 SUB 0.25fF $ **FLOATING
C7096 S.n6456 SUB 0.01fF $ **FLOATING
C7097 S.t2271 SUB 0.02fF
C7098 S.n6457 SUB 0.25fF $ **FLOATING
C7099 S.t1498 SUB 0.02fF
C7100 S.n6458 SUB 0.95fF $ **FLOATING
C7101 S.n6459 SUB 0.70fF $ **FLOATING
C7102 S.n6460 SUB 0.78fF $ **FLOATING
C7103 S.n6461 SUB 1.93fF $ **FLOATING
C7104 S.n6462 SUB 1.88fF $ **FLOATING
C7105 S.n6463 SUB 0.12fF $ **FLOATING
C7106 S.t1415 SUB 0.02fF
C7107 S.n6464 SUB 0.14fF $ **FLOATING
C7108 S.t1654 SUB 0.02fF
C7109 S.n6466 SUB 0.24fF $ **FLOATING
C7110 S.n6467 SUB 0.36fF $ **FLOATING
C7111 S.n6468 SUB 0.61fF $ **FLOATING
C7112 S.n6469 SUB 1.52fF $ **FLOATING
C7113 S.n6470 SUB 2.99fF $ **FLOATING
C7114 S.t635 SUB 0.02fF
C7115 S.n6471 SUB 0.24fF $ **FLOATING
C7116 S.n6472 SUB 0.91fF $ **FLOATING
C7117 S.n6473 SUB 0.05fF $ **FLOATING
C7118 S.t2057 SUB 0.02fF
C7119 S.n6474 SUB 0.12fF $ **FLOATING
C7120 S.n6475 SUB 0.14fF $ **FLOATING
C7121 S.n6477 SUB 1.89fF $ **FLOATING
C7122 S.n6478 SUB 1.88fF $ **FLOATING
C7123 S.t783 SUB 0.02fF
C7124 S.n6479 SUB 0.24fF $ **FLOATING
C7125 S.n6480 SUB 0.36fF $ **FLOATING
C7126 S.n6481 SUB 0.61fF $ **FLOATING
C7127 S.n6482 SUB 0.12fF $ **FLOATING
C7128 S.t551 SUB 0.02fF
C7129 S.n6483 SUB 0.14fF $ **FLOATING
C7130 S.n6485 SUB 1.16fF $ **FLOATING
C7131 S.n6486 SUB 0.22fF $ **FLOATING
C7132 S.n6487 SUB 0.25fF $ **FLOATING
C7133 S.n6488 SUB 0.09fF $ **FLOATING
C7134 S.n6489 SUB 1.88fF $ **FLOATING
C7135 S.t2288 SUB 0.02fF
C7136 S.n6490 SUB 0.24fF $ **FLOATING
C7137 S.n6491 SUB 0.91fF $ **FLOATING
C7138 S.n6492 SUB 0.05fF $ **FLOATING
C7139 S.t1195 SUB 0.02fF
C7140 S.n6493 SUB 0.12fF $ **FLOATING
C7141 S.n6494 SUB 0.14fF $ **FLOATING
C7142 S.n6496 SUB 0.78fF $ **FLOATING
C7143 S.n6497 SUB 1.94fF $ **FLOATING
C7144 S.n6498 SUB 1.88fF $ **FLOATING
C7145 S.n6499 SUB 0.12fF $ **FLOATING
C7146 S.t2190 SUB 0.02fF
C7147 S.n6500 SUB 0.14fF $ **FLOATING
C7148 S.t2436 SUB 0.02fF
C7149 S.n6502 SUB 0.24fF $ **FLOATING
C7150 S.n6503 SUB 0.36fF $ **FLOATING
C7151 S.n6504 SUB 0.61fF $ **FLOATING
C7152 S.n6505 SUB 1.84fF $ **FLOATING
C7153 S.n6506 SUB 2.99fF $ **FLOATING
C7154 S.t1435 SUB 0.02fF
C7155 S.n6507 SUB 0.24fF $ **FLOATING
C7156 S.n6508 SUB 0.91fF $ **FLOATING
C7157 S.n6509 SUB 0.05fF $ **FLOATING
C7158 S.t468 SUB 0.02fF
C7159 S.n6510 SUB 0.12fF $ **FLOATING
C7160 S.n6511 SUB 0.14fF $ **FLOATING
C7161 S.n6513 SUB 1.89fF $ **FLOATING
C7162 S.n6514 SUB 1.88fF $ **FLOATING
C7163 S.t1572 SUB 0.02fF
C7164 S.n6515 SUB 0.24fF $ **FLOATING
C7165 S.n6516 SUB 0.36fF $ **FLOATING
C7166 S.n6517 SUB 0.61fF $ **FLOATING
C7167 S.n6518 SUB 0.12fF $ **FLOATING
C7168 S.t1328 SUB 0.02fF
C7169 S.n6519 SUB 0.14fF $ **FLOATING
C7170 S.n6521 SUB 1.16fF $ **FLOATING
C7171 S.n6522 SUB 0.22fF $ **FLOATING
C7172 S.n6523 SUB 0.25fF $ **FLOATING
C7173 S.n6524 SUB 0.09fF $ **FLOATING
C7174 S.n6525 SUB 1.88fF $ **FLOATING
C7175 S.t572 SUB 0.02fF
C7176 S.n6526 SUB 0.24fF $ **FLOATING
C7177 S.n6527 SUB 0.91fF $ **FLOATING
C7178 S.n6528 SUB 0.05fF $ **FLOATING
C7179 S.t2117 SUB 0.02fF
C7180 S.n6529 SUB 0.12fF $ **FLOATING
C7181 S.n6530 SUB 0.14fF $ **FLOATING
C7182 S.n6532 SUB 0.78fF $ **FLOATING
C7183 S.n6533 SUB 1.94fF $ **FLOATING
C7184 S.n6534 SUB 1.88fF $ **FLOATING
C7185 S.n6535 SUB 0.12fF $ **FLOATING
C7186 S.t449 SUB 0.02fF
C7187 S.n6536 SUB 0.14fF $ **FLOATING
C7188 S.t701 SUB 0.02fF
C7189 S.n6538 SUB 0.24fF $ **FLOATING
C7190 S.n6539 SUB 0.36fF $ **FLOATING
C7191 S.n6540 SUB 0.61fF $ **FLOATING
C7192 S.n6541 SUB 1.84fF $ **FLOATING
C7193 S.n6542 SUB 2.99fF $ **FLOATING
C7194 S.t2217 SUB 0.02fF
C7195 S.n6543 SUB 0.24fF $ **FLOATING
C7196 S.n6544 SUB 0.91fF $ **FLOATING
C7197 S.n6545 SUB 0.05fF $ **FLOATING
C7198 S.t1246 SUB 0.02fF
C7199 S.n6546 SUB 0.12fF $ **FLOATING
C7200 S.n6547 SUB 0.14fF $ **FLOATING
C7201 S.n6549 SUB 1.89fF $ **FLOATING
C7202 S.n6550 SUB 1.75fF $ **FLOATING
C7203 S.t2360 SUB 0.02fF
C7204 S.n6551 SUB 0.24fF $ **FLOATING
C7205 S.n6552 SUB 0.36fF $ **FLOATING
C7206 S.n6553 SUB 0.61fF $ **FLOATING
C7207 S.n6554 SUB 0.12fF $ **FLOATING
C7208 S.t2092 SUB 0.02fF
C7209 S.n6555 SUB 0.14fF $ **FLOATING
C7210 S.n6557 SUB 1.16fF $ **FLOATING
C7211 S.n6558 SUB 0.22fF $ **FLOATING
C7212 S.n6559 SUB 0.25fF $ **FLOATING
C7213 S.n6560 SUB 0.09fF $ **FLOATING
C7214 S.n6561 SUB 2.44fF $ **FLOATING
C7215 S.t1357 SUB 0.02fF
C7216 S.n6562 SUB 0.24fF $ **FLOATING
C7217 S.n6563 SUB 0.91fF $ **FLOATING
C7218 S.n6564 SUB 0.05fF $ **FLOATING
C7219 S.t364 SUB 0.02fF
C7220 S.n6565 SUB 0.12fF $ **FLOATING
C7221 S.n6566 SUB 0.14fF $ **FLOATING
C7222 S.n6568 SUB 1.88fF $ **FLOATING
C7223 S.n6569 SUB 0.48fF $ **FLOATING
C7224 S.n6570 SUB 0.09fF $ **FLOATING
C7225 S.n6571 SUB 0.33fF $ **FLOATING
C7226 S.n6572 SUB 0.30fF $ **FLOATING
C7227 S.n6573 SUB 0.77fF $ **FLOATING
C7228 S.n6574 SUB 0.59fF $ **FLOATING
C7229 S.t1504 SUB 0.02fF
C7230 S.n6575 SUB 0.24fF $ **FLOATING
C7231 S.n6576 SUB 0.36fF $ **FLOATING
C7232 S.n6577 SUB 0.61fF $ **FLOATING
C7233 S.n6578 SUB 0.12fF $ **FLOATING
C7234 S.t1375 SUB 0.02fF
C7235 S.n6579 SUB 0.14fF $ **FLOATING
C7236 S.n6581 SUB 2.61fF $ **FLOATING
C7237 S.n6582 SUB 2.16fF $ **FLOATING
C7238 S.t479 SUB 0.02fF
C7239 S.n6583 SUB 0.24fF $ **FLOATING
C7240 S.n6584 SUB 0.91fF $ **FLOATING
C7241 S.n6585 SUB 0.05fF $ **FLOATING
C7242 S.t2016 SUB 0.02fF
C7243 S.n6586 SUB 0.12fF $ **FLOATING
C7244 S.n6587 SUB 0.14fF $ **FLOATING
C7245 S.n6589 SUB 0.78fF $ **FLOATING
C7246 S.n6590 SUB 2.30fF $ **FLOATING
C7247 S.n6591 SUB 1.88fF $ **FLOATING
C7248 S.n6592 SUB 0.12fF $ **FLOATING
C7249 S.t1962 SUB 0.02fF
C7250 S.n6593 SUB 0.14fF $ **FLOATING
C7251 S.t1218 SUB 0.02fF
C7252 S.n6595 SUB 0.24fF $ **FLOATING
C7253 S.n6596 SUB 0.36fF $ **FLOATING
C7254 S.n6597 SUB 0.61fF $ **FLOATING
C7255 S.n6598 SUB 1.39fF $ **FLOATING
C7256 S.n6599 SUB 0.71fF $ **FLOATING
C7257 S.n6600 SUB 1.14fF $ **FLOATING
C7258 S.n6601 SUB 0.35fF $ **FLOATING
C7259 S.n6602 SUB 2.03fF $ **FLOATING
C7260 S.t95 SUB 0.02fF
C7261 S.n6603 SUB 0.24fF $ **FLOATING
C7262 S.n6604 SUB 0.91fF $ **FLOATING
C7263 S.n6605 SUB 0.05fF $ **FLOATING
C7264 S.t1163 SUB 0.02fF
C7265 S.n6606 SUB 0.12fF $ **FLOATING
C7266 S.n6607 SUB 0.14fF $ **FLOATING
C7267 S.n6609 SUB 1.89fF $ **FLOATING
C7268 S.n6610 SUB 1.88fF $ **FLOATING
C7269 S.t336 SUB 0.02fF
C7270 S.n6611 SUB 0.24fF $ **FLOATING
C7271 S.n6612 SUB 0.36fF $ **FLOATING
C7272 S.n6613 SUB 0.61fF $ **FLOATING
C7273 S.n6614 SUB 0.12fF $ **FLOATING
C7274 S.t1104 SUB 0.02fF
C7275 S.n6615 SUB 0.14fF $ **FLOATING
C7276 S.n6617 SUB 1.16fF $ **FLOATING
C7277 S.n6618 SUB 0.22fF $ **FLOATING
C7278 S.n6619 SUB 0.25fF $ **FLOATING
C7279 S.n6620 SUB 0.09fF $ **FLOATING
C7280 S.n6621 SUB 1.88fF $ **FLOATING
C7281 S.t1770 SUB 0.02fF
C7282 S.n6622 SUB 0.24fF $ **FLOATING
C7283 S.n6623 SUB 0.91fF $ **FLOATING
C7284 S.n6624 SUB 0.05fF $ **FLOATING
C7285 S.t1769 SUB 0.02fF
C7286 S.n6625 SUB 0.12fF $ **FLOATING
C7287 S.n6626 SUB 0.14fF $ **FLOATING
C7288 S.n6628 SUB 20.78fF $ **FLOATING
C7289 S.n6629 SUB 1.88fF $ **FLOATING
C7290 S.n6630 SUB 2.67fF $ **FLOATING
C7291 S.t268 SUB 0.02fF
C7292 S.n6631 SUB 0.24fF $ **FLOATING
C7293 S.n6632 SUB 0.36fF $ **FLOATING
C7294 S.n6633 SUB 0.61fF $ **FLOATING
C7295 S.n6634 SUB 0.12fF $ **FLOATING
C7296 S.t1034 SUB 0.02fF
C7297 S.n6635 SUB 0.14fF $ **FLOATING
C7298 S.n6637 SUB 2.80fF $ **FLOATING
C7299 S.n6638 SUB 2.30fF $ **FLOATING
C7300 S.t1669 SUB 0.02fF
C7301 S.n6639 SUB 0.12fF $ **FLOATING
C7302 S.n6640 SUB 0.14fF $ **FLOATING
C7303 S.t1667 SUB 0.02fF
C7304 S.n6642 SUB 0.24fF $ **FLOATING
C7305 S.n6643 SUB 0.91fF $ **FLOATING
C7306 S.n6644 SUB 0.05fF $ **FLOATING
C7307 S.n6645 SUB 1.88fF $ **FLOATING
C7308 S.n6646 SUB 2.67fF $ **FLOATING
C7309 S.t1930 SUB 0.02fF
C7310 S.n6647 SUB 0.24fF $ **FLOATING
C7311 S.n6648 SUB 0.36fF $ **FLOATING
C7312 S.n6649 SUB 0.61fF $ **FLOATING
C7313 S.n6650 SUB 0.12fF $ **FLOATING
C7314 S.t137 SUB 0.02fF
C7315 S.n6651 SUB 0.14fF $ **FLOATING
C7316 S.n6653 SUB 2.80fF $ **FLOATING
C7317 S.n6654 SUB 2.30fF $ **FLOATING
C7318 S.t957 SUB 0.02fF
C7319 S.n6655 SUB 0.12fF $ **FLOATING
C7320 S.n6656 SUB 0.14fF $ **FLOATING
C7321 S.t793 SUB 0.02fF
C7322 S.n6658 SUB 0.24fF $ **FLOATING
C7323 S.n6659 SUB 0.91fF $ **FLOATING
C7324 S.n6660 SUB 0.05fF $ **FLOATING
C7325 S.n6661 SUB 1.88fF $ **FLOATING
C7326 S.n6662 SUB 2.67fF $ **FLOATING
C7327 S.t1071 SUB 0.02fF
C7328 S.n6663 SUB 0.24fF $ **FLOATING
C7329 S.n6664 SUB 0.36fF $ **FLOATING
C7330 S.n6665 SUB 0.61fF $ **FLOATING
C7331 S.n6666 SUB 0.12fF $ **FLOATING
C7332 S.t1808 SUB 0.02fF
C7333 S.n6667 SUB 0.14fF $ **FLOATING
C7334 S.n6669 SUB 2.80fF $ **FLOATING
C7335 S.n6670 SUB 2.30fF $ **FLOATING
C7336 S.t9 SUB 0.02fF
C7337 S.n6671 SUB 0.12fF $ **FLOATING
C7338 S.n6672 SUB 0.14fF $ **FLOATING
C7339 S.t2444 SUB 0.02fF
C7340 S.n6674 SUB 0.24fF $ **FLOATING
C7341 S.n6675 SUB 0.91fF $ **FLOATING
C7342 S.n6676 SUB 0.05fF $ **FLOATING
C7343 S.n6677 SUB 1.88fF $ **FLOATING
C7344 S.n6678 SUB 2.67fF $ **FLOATING
C7345 S.t192 SUB 0.02fF
C7346 S.n6679 SUB 0.24fF $ **FLOATING
C7347 S.n6680 SUB 0.36fF $ **FLOATING
C7348 S.n6681 SUB 0.61fF $ **FLOATING
C7349 S.n6682 SUB 0.12fF $ **FLOATING
C7350 S.t942 SUB 0.02fF
C7351 S.n6683 SUB 0.14fF $ **FLOATING
C7352 S.n6685 SUB 2.80fF $ **FLOATING
C7353 S.n6686 SUB 2.30fF $ **FLOATING
C7354 S.t1721 SUB 0.02fF
C7355 S.n6687 SUB 0.12fF $ **FLOATING
C7356 S.n6688 SUB 0.14fF $ **FLOATING
C7357 S.t1577 SUB 0.02fF
C7358 S.n6690 SUB 0.24fF $ **FLOATING
C7359 S.n6691 SUB 0.91fF $ **FLOATING
C7360 S.n6692 SUB 0.05fF $ **FLOATING
C7361 S.n6693 SUB 2.73fF $ **FLOATING
C7362 S.n6694 SUB 1.59fF $ **FLOATING
C7363 S.n6695 SUB 0.12fF $ **FLOATING
C7364 S.t2102 SUB 0.02fF
C7365 S.n6696 SUB 0.14fF $ **FLOATING
C7366 S.t1050 SUB 0.02fF
C7367 S.n6698 SUB 0.24fF $ **FLOATING
C7368 S.n6699 SUB 0.36fF $ **FLOATING
C7369 S.n6700 SUB 0.61fF $ **FLOATING
C7370 S.n6701 SUB 0.07fF $ **FLOATING
C7371 S.n6702 SUB 0.01fF $ **FLOATING
C7372 S.n6703 SUB 0.24fF $ **FLOATING
C7373 S.n6704 SUB 1.16fF $ **FLOATING
C7374 S.n6705 SUB 1.35fF $ **FLOATING
C7375 S.n6706 SUB 2.30fF $ **FLOATING
C7376 S.t317 SUB 0.02fF
C7377 S.n6707 SUB 0.12fF $ **FLOATING
C7378 S.n6708 SUB 0.14fF $ **FLOATING
C7379 S.t1141 SUB 0.02fF
C7380 S.n6710 SUB 0.24fF $ **FLOATING
C7381 S.n6711 SUB 0.91fF $ **FLOATING
C7382 S.n6712 SUB 0.05fF $ **FLOATING
C7383 S.t8 SUB 48.31fF
C7384 S.t709 SUB 0.02fF
C7385 S.n6713 SUB 0.24fF $ **FLOATING
C7386 S.n6714 SUB 0.91fF $ **FLOATING
C7387 S.n6715 SUB 0.05fF $ **FLOATING
C7388 S.t849 SUB 0.02fF
C7389 S.n6716 SUB 0.12fF $ **FLOATING
C7390 S.n6717 SUB 0.14fF $ **FLOATING
C7391 S.n6719 SUB 0.12fF $ **FLOATING
C7392 S.t2581 SUB 0.02fF
C7393 S.n6720 SUB 0.14fF $ **FLOATING
C7394 S.n6722 SUB 5.17fF $ **FLOATING
C7395 S.n6723 SUB 5.44fF $ **FLOATING
C7396 S.t2112 SUB 0.02fF
C7397 S.n6724 SUB 0.12fF $ **FLOATING
C7398 S.n6725 SUB 0.14fF $ **FLOATING
C7399 S.t518 SUB 0.02fF
C7400 S.n6727 SUB 0.24fF $ **FLOATING
C7401 S.n6728 SUB 0.91fF $ **FLOATING
C7402 S.n6729 SUB 0.05fF $ **FLOATING
C7403 S.t119 SUB 47.92fF
C7404 S.t2552 SUB 0.02fF
C7405 S.n6730 SUB 1.19fF $ **FLOATING
C7406 S.n6731 SUB 0.05fF $ **FLOATING
C7407 S.t1558 SUB 0.02fF
C7408 S.n6732 SUB 0.01fF $ **FLOATING
C7409 S.n6733 SUB 0.26fF $ **FLOATING
C7410 S.n6735 SUB 1.50fF $ **FLOATING
C7411 S.n6736 SUB 1.30fF $ **FLOATING
C7412 S.n6737 SUB 0.28fF $ **FLOATING
C7413 S.n6738 SUB 0.24fF $ **FLOATING
C7414 S.n6739 SUB 4.39fF $ **FLOATING
C7415 S.n6740 SUB 0.01fF $ **FLOATING
C7416 S.n6741 SUB 0.02fF $ **FLOATING
C7417 S.n6742 SUB 0.03fF $ **FLOATING
C7418 S.n6743 SUB 0.04fF $ **FLOATING
C7419 S.n6744 SUB 0.17fF $ **FLOATING
C7420 S.n6745 SUB 0.01fF $ **FLOATING
C7421 S.n6746 SUB 0.02fF $ **FLOATING
C7422 S.n6747 SUB 0.01fF $ **FLOATING
C7423 S.n6748 SUB 0.01fF $ **FLOATING
C7424 S.n6749 SUB 0.01fF $ **FLOATING
C7425 S.n6750 SUB 0.01fF $ **FLOATING
C7426 S.n6751 SUB 0.02fF $ **FLOATING
C7427 S.n6752 SUB 0.01fF $ **FLOATING
C7428 S.n6753 SUB 0.02fF $ **FLOATING
C7429 S.n6754 SUB 0.05fF $ **FLOATING
C7430 S.n6755 SUB 0.04fF $ **FLOATING
C7431 S.n6756 SUB 0.11fF $ **FLOATING
C7432 S.n6757 SUB 0.38fF $ **FLOATING
C7433 S.n6758 SUB 0.20fF $ **FLOATING
C7434 S.n6759 SUB 8.97fF $ **FLOATING
C7435 S.n6760 SUB 8.97fF $ **FLOATING
C7436 S.n6761 SUB 0.60fF $ **FLOATING
C7437 S.n6762 SUB 0.22fF $ **FLOATING
C7438 S.n6763 SUB 0.59fF $ **FLOATING
C7439 S.n6764 SUB 3.43fF $ **FLOATING
C7440 S.n6765 SUB 0.29fF $ **FLOATING
C7441 S.t42 SUB 21.38fF
C7442 S.n6766 SUB 21.67fF $ **FLOATING
C7443 S.n6767 SUB 0.77fF $ **FLOATING
C7444 S.n6768 SUB 0.28fF $ **FLOATING
C7445 S.n6769 SUB 4.00fF $ **FLOATING
C7446 S.n6770 SUB 1.35fF $ **FLOATING
C7447 S.t2204 SUB 0.02fF
C7448 S.n6771 SUB 0.64fF $ **FLOATING
C7449 S.n6772 SUB 0.61fF $ **FLOATING
C7450 S.n6773 SUB 1.89fF $ **FLOATING
C7451 S.n6774 SUB 0.06fF $ **FLOATING
C7452 S.n6775 SUB 0.03fF $ **FLOATING
C7453 S.n6776 SUB 0.04fF $ **FLOATING
C7454 S.n6777 SUB 0.99fF $ **FLOATING
C7455 S.n6778 SUB 0.02fF $ **FLOATING
C7456 S.n6779 SUB 0.01fF $ **FLOATING
C7457 S.n6780 SUB 0.02fF $ **FLOATING
C7458 S.n6781 SUB 0.08fF $ **FLOATING
C7459 S.n6782 SUB 0.36fF $ **FLOATING
C7460 S.n6783 SUB 1.85fF $ **FLOATING
C7461 S.t2554 SUB 0.02fF
C7462 S.n6784 SUB 0.24fF $ **FLOATING
C7463 S.n6785 SUB 0.36fF $ **FLOATING
C7464 S.n6786 SUB 0.61fF $ **FLOATING
C7465 S.n6787 SUB 0.12fF $ **FLOATING
C7466 S.t2020 SUB 0.02fF
C7467 S.n6788 SUB 0.14fF $ **FLOATING
C7468 S.n6790 SUB 0.70fF $ **FLOATING
C7469 S.n6791 SUB 0.23fF $ **FLOATING
C7470 S.n6792 SUB 0.23fF $ **FLOATING
C7471 S.n6793 SUB 0.70fF $ **FLOATING
C7472 S.n6794 SUB 1.16fF $ **FLOATING
C7473 S.n6795 SUB 0.22fF $ **FLOATING
C7474 S.n6796 SUB 0.25fF $ **FLOATING
C7475 S.n6797 SUB 0.09fF $ **FLOATING
C7476 S.n6798 SUB 1.88fF $ **FLOATING
C7477 S.t869 SUB 0.02fF
C7478 S.n6799 SUB 0.24fF $ **FLOATING
C7479 S.n6800 SUB 0.91fF $ **FLOATING
C7480 S.n6801 SUB 0.05fF $ **FLOATING
C7481 S.t2238 SUB 0.02fF
C7482 S.n6802 SUB 0.12fF $ **FLOATING
C7483 S.n6803 SUB 0.14fF $ **FLOATING
C7484 S.n6805 SUB 0.25fF $ **FLOATING
C7485 S.n6806 SUB 0.09fF $ **FLOATING
C7486 S.n6807 SUB 0.21fF $ **FLOATING
C7487 S.n6808 SUB 0.92fF $ **FLOATING
C7488 S.n6809 SUB 0.44fF $ **FLOATING
C7489 S.n6810 SUB 1.88fF $ **FLOATING
C7490 S.n6811 SUB 0.12fF $ **FLOATING
C7491 S.t1302 SUB 0.02fF
C7492 S.n6812 SUB 0.14fF $ **FLOATING
C7493 S.t1840 SUB 0.02fF
C7494 S.n6814 SUB 0.24fF $ **FLOATING
C7495 S.n6815 SUB 0.36fF $ **FLOATING
C7496 S.n6816 SUB 0.61fF $ **FLOATING
C7497 S.n6817 SUB 0.02fF $ **FLOATING
C7498 S.n6818 SUB 0.01fF $ **FLOATING
C7499 S.n6819 SUB 0.02fF $ **FLOATING
C7500 S.n6820 SUB 0.08fF $ **FLOATING
C7501 S.n6821 SUB 0.06fF $ **FLOATING
C7502 S.n6822 SUB 0.03fF $ **FLOATING
C7503 S.n6823 SUB 0.04fF $ **FLOATING
C7504 S.n6824 SUB 1.00fF $ **FLOATING
C7505 S.n6825 SUB 0.36fF $ **FLOATING
C7506 S.n6826 SUB 1.87fF $ **FLOATING
C7507 S.n6827 SUB 1.99fF $ **FLOATING
C7508 S.t126 SUB 0.02fF
C7509 S.n6828 SUB 0.24fF $ **FLOATING
C7510 S.n6829 SUB 0.91fF $ **FLOATING
C7511 S.n6830 SUB 0.05fF $ **FLOATING
C7512 S.t1379 SUB 0.02fF
C7513 S.n6831 SUB 0.12fF $ **FLOATING
C7514 S.n6832 SUB 0.14fF $ **FLOATING
C7515 S.n6834 SUB 1.89fF $ **FLOATING
C7516 S.n6835 SUB 0.06fF $ **FLOATING
C7517 S.n6836 SUB 0.03fF $ **FLOATING
C7518 S.n6837 SUB 0.04fF $ **FLOATING
C7519 S.n6838 SUB 0.99fF $ **FLOATING
C7520 S.n6839 SUB 0.02fF $ **FLOATING
C7521 S.n6840 SUB 0.01fF $ **FLOATING
C7522 S.n6841 SUB 0.02fF $ **FLOATING
C7523 S.n6842 SUB 0.08fF $ **FLOATING
C7524 S.n6843 SUB 0.36fF $ **FLOATING
C7525 S.n6844 SUB 1.85fF $ **FLOATING
C7526 S.t976 SUB 0.02fF
C7527 S.n6845 SUB 0.24fF $ **FLOATING
C7528 S.n6846 SUB 0.36fF $ **FLOATING
C7529 S.n6847 SUB 0.61fF $ **FLOATING
C7530 S.n6848 SUB 0.12fF $ **FLOATING
C7531 S.t418 SUB 0.02fF
C7532 S.n6849 SUB 0.14fF $ **FLOATING
C7533 S.n6851 SUB 0.70fF $ **FLOATING
C7534 S.n6852 SUB 0.23fF $ **FLOATING
C7535 S.n6853 SUB 0.23fF $ **FLOATING
C7536 S.n6854 SUB 0.70fF $ **FLOATING
C7537 S.n6855 SUB 1.16fF $ **FLOATING
C7538 S.n6856 SUB 0.22fF $ **FLOATING
C7539 S.n6857 SUB 0.25fF $ **FLOATING
C7540 S.n6858 SUB 0.09fF $ **FLOATING
C7541 S.n6859 SUB 1.88fF $ **FLOATING
C7542 S.t1796 SUB 0.02fF
C7543 S.n6860 SUB 0.24fF $ **FLOATING
C7544 S.n6861 SUB 0.91fF $ **FLOATING
C7545 S.n6862 SUB 0.05fF $ **FLOATING
C7546 S.t505 SUB 0.02fF
C7547 S.n6863 SUB 0.12fF $ **FLOATING
C7548 S.n6864 SUB 0.14fF $ **FLOATING
C7549 S.n6866 SUB 0.25fF $ **FLOATING
C7550 S.n6867 SUB 0.09fF $ **FLOATING
C7551 S.n6868 SUB 0.21fF $ **FLOATING
C7552 S.n6869 SUB 0.92fF $ **FLOATING
C7553 S.n6870 SUB 0.44fF $ **FLOATING
C7554 S.n6871 SUB 1.88fF $ **FLOATING
C7555 S.n6872 SUB 0.12fF $ **FLOATING
C7556 S.t2067 SUB 0.02fF
C7557 S.n6873 SUB 0.14fF $ **FLOATING
C7558 S.t43 SUB 0.02fF
C7559 S.n6875 SUB 0.24fF $ **FLOATING
C7560 S.n6876 SUB 0.36fF $ **FLOATING
C7561 S.n6877 SUB 0.61fF $ **FLOATING
C7562 S.n6878 SUB 0.02fF $ **FLOATING
C7563 S.n6879 SUB 0.01fF $ **FLOATING
C7564 S.n6880 SUB 0.02fF $ **FLOATING
C7565 S.n6881 SUB 0.08fF $ **FLOATING
C7566 S.n6882 SUB 0.06fF $ **FLOATING
C7567 S.n6883 SUB 0.03fF $ **FLOATING
C7568 S.n6884 SUB 0.04fF $ **FLOATING
C7569 S.n6885 SUB 1.00fF $ **FLOATING
C7570 S.n6886 SUB 0.36fF $ **FLOATING
C7571 S.n6887 SUB 1.87fF $ **FLOATING
C7572 S.n6888 SUB 1.99fF $ **FLOATING
C7573 S.t930 SUB 0.02fF
C7574 S.n6889 SUB 0.24fF $ **FLOATING
C7575 S.n6890 SUB 0.91fF $ **FLOATING
C7576 S.n6891 SUB 0.05fF $ **FLOATING
C7577 S.t2148 SUB 0.02fF
C7578 S.n6892 SUB 0.12fF $ **FLOATING
C7579 S.n6893 SUB 0.14fF $ **FLOATING
C7580 S.n6895 SUB 1.89fF $ **FLOATING
C7581 S.n6896 SUB 0.07fF $ **FLOATING
C7582 S.n6897 SUB 0.04fF $ **FLOATING
C7583 S.n6898 SUB 0.05fF $ **FLOATING
C7584 S.n6899 SUB 0.87fF $ **FLOATING
C7585 S.n6900 SUB 0.01fF $ **FLOATING
C7586 S.n6901 SUB 0.01fF $ **FLOATING
C7587 S.n6902 SUB 0.01fF $ **FLOATING
C7588 S.n6903 SUB 0.07fF $ **FLOATING
C7589 S.n6904 SUB 0.68fF $ **FLOATING
C7590 S.n6905 SUB 0.72fF $ **FLOATING
C7591 S.t1737 SUB 0.02fF
C7592 S.n6906 SUB 0.24fF $ **FLOATING
C7593 S.n6907 SUB 0.36fF $ **FLOATING
C7594 S.n6908 SUB 0.61fF $ **FLOATING
C7595 S.n6909 SUB 0.12fF $ **FLOATING
C7596 S.t1205 SUB 0.02fF
C7597 S.n6910 SUB 0.14fF $ **FLOATING
C7598 S.n6912 SUB 0.70fF $ **FLOATING
C7599 S.n6913 SUB 0.23fF $ **FLOATING
C7600 S.n6914 SUB 0.23fF $ **FLOATING
C7601 S.n6915 SUB 0.70fF $ **FLOATING
C7602 S.n6916 SUB 1.16fF $ **FLOATING
C7603 S.n6917 SUB 0.22fF $ **FLOATING
C7604 S.n6918 SUB 0.25fF $ **FLOATING
C7605 S.n6919 SUB 0.09fF $ **FLOATING
C7606 S.n6920 SUB 2.31fF $ **FLOATING
C7607 S.t2570 SUB 0.02fF
C7608 S.n6921 SUB 0.24fF $ **FLOATING
C7609 S.n6922 SUB 0.91fF $ **FLOATING
C7610 S.n6923 SUB 0.05fF $ **FLOATING
C7611 S.t1288 SUB 0.02fF
C7612 S.n6924 SUB 0.12fF $ **FLOATING
C7613 S.n6925 SUB 0.14fF $ **FLOATING
C7614 S.n6927 SUB 1.88fF $ **FLOATING
C7615 S.n6928 SUB 0.46fF $ **FLOATING
C7616 S.n6929 SUB 0.22fF $ **FLOATING
C7617 S.n6930 SUB 0.38fF $ **FLOATING
C7618 S.n6931 SUB 0.16fF $ **FLOATING
C7619 S.n6932 SUB 0.28fF $ **FLOATING
C7620 S.n6933 SUB 0.21fF $ **FLOATING
C7621 S.n6934 SUB 0.30fF $ **FLOATING
C7622 S.n6935 SUB 0.42fF $ **FLOATING
C7623 S.n6936 SUB 0.21fF $ **FLOATING
C7624 S.t862 SUB 0.02fF
C7625 S.n6937 SUB 0.24fF $ **FLOATING
C7626 S.n6938 SUB 0.36fF $ **FLOATING
C7627 S.n6939 SUB 0.61fF $ **FLOATING
C7628 S.n6940 SUB 0.12fF $ **FLOATING
C7629 S.t327 SUB 0.02fF
C7630 S.n6941 SUB 0.14fF $ **FLOATING
C7631 S.n6943 SUB 0.04fF $ **FLOATING
C7632 S.n6944 SUB 0.03fF $ **FLOATING
C7633 S.n6945 SUB 0.03fF $ **FLOATING
C7634 S.n6946 SUB 0.10fF $ **FLOATING
C7635 S.n6947 SUB 0.36fF $ **FLOATING
C7636 S.n6948 SUB 0.38fF $ **FLOATING
C7637 S.n6949 SUB 0.11fF $ **FLOATING
C7638 S.n6950 SUB 0.12fF $ **FLOATING
C7639 S.n6951 SUB 0.07fF $ **FLOATING
C7640 S.n6952 SUB 0.12fF $ **FLOATING
C7641 S.n6953 SUB 0.18fF $ **FLOATING
C7642 S.n6954 SUB 4.00fF $ **FLOATING
C7643 S.t1694 SUB 0.02fF
C7644 S.n6955 SUB 0.24fF $ **FLOATING
C7645 S.n6956 SUB 0.91fF $ **FLOATING
C7646 S.n6957 SUB 0.05fF $ **FLOATING
C7647 S.t405 SUB 0.02fF
C7648 S.n6958 SUB 0.12fF $ **FLOATING
C7649 S.n6959 SUB 0.14fF $ **FLOATING
C7650 S.n6961 SUB 0.25fF $ **FLOATING
C7651 S.n6962 SUB 0.09fF $ **FLOATING
C7652 S.n6963 SUB 0.21fF $ **FLOATING
C7653 S.n6964 SUB 1.28fF $ **FLOATING
C7654 S.n6965 SUB 0.53fF $ **FLOATING
C7655 S.n6966 SUB 1.88fF $ **FLOATING
C7656 S.n6967 SUB 0.12fF $ **FLOATING
C7657 S.t1986 SUB 0.02fF
C7658 S.n6968 SUB 0.14fF $ **FLOATING
C7659 S.t2507 SUB 0.02fF
C7660 S.n6970 SUB 0.24fF $ **FLOATING
C7661 S.n6971 SUB 0.36fF $ **FLOATING
C7662 S.n6972 SUB 0.61fF $ **FLOATING
C7663 S.n6973 SUB 1.58fF $ **FLOATING
C7664 S.n6974 SUB 2.45fF $ **FLOATING
C7665 S.t819 SUB 0.02fF
C7666 S.n6975 SUB 0.24fF $ **FLOATING
C7667 S.n6976 SUB 0.91fF $ **FLOATING
C7668 S.n6977 SUB 0.05fF $ **FLOATING
C7669 S.t2196 SUB 0.02fF
C7670 S.n6978 SUB 0.12fF $ **FLOATING
C7671 S.n6979 SUB 0.14fF $ **FLOATING
C7672 S.n6981 SUB 1.89fF $ **FLOATING
C7673 S.n6982 SUB 0.06fF $ **FLOATING
C7674 S.n6983 SUB 0.03fF $ **FLOATING
C7675 S.n6984 SUB 0.04fF $ **FLOATING
C7676 S.n6985 SUB 0.99fF $ **FLOATING
C7677 S.n6986 SUB 0.02fF $ **FLOATING
C7678 S.n6987 SUB 0.01fF $ **FLOATING
C7679 S.n6988 SUB 0.02fF $ **FLOATING
C7680 S.n6989 SUB 0.08fF $ **FLOATING
C7681 S.n6990 SUB 0.36fF $ **FLOATING
C7682 S.n6991 SUB 1.85fF $ **FLOATING
C7683 S.t533 SUB 0.02fF
C7684 S.n6992 SUB 0.24fF $ **FLOATING
C7685 S.n6993 SUB 0.36fF $ **FLOATING
C7686 S.n6994 SUB 0.61fF $ **FLOATING
C7687 S.n6995 SUB 0.12fF $ **FLOATING
C7688 S.t2468 SUB 0.02fF
C7689 S.n6996 SUB 0.14fF $ **FLOATING
C7690 S.n6998 SUB 0.70fF $ **FLOATING
C7691 S.n6999 SUB 0.23fF $ **FLOATING
C7692 S.n7000 SUB 0.23fF $ **FLOATING
C7693 S.n7001 SUB 0.70fF $ **FLOATING
C7694 S.n7002 SUB 1.16fF $ **FLOATING
C7695 S.n7003 SUB 0.22fF $ **FLOATING
C7696 S.n7004 SUB 0.25fF $ **FLOATING
C7697 S.n7005 SUB 0.09fF $ **FLOATING
C7698 S.n7006 SUB 1.88fF $ **FLOATING
C7699 S.t413 SUB 0.02fF
C7700 S.n7007 SUB 0.24fF $ **FLOATING
C7701 S.n7008 SUB 0.91fF $ **FLOATING
C7702 S.n7009 SUB 0.05fF $ **FLOATING
C7703 S.t173 SUB 0.02fF
C7704 S.n7010 SUB 0.12fF $ **FLOATING
C7705 S.n7011 SUB 0.14fF $ **FLOATING
C7706 S.n7013 SUB 20.78fF $ **FLOATING
C7707 S.n7014 SUB 0.06fF $ **FLOATING
C7708 S.n7015 SUB 0.20fF $ **FLOATING
C7709 S.n7016 SUB 0.09fF $ **FLOATING
C7710 S.n7017 SUB 0.21fF $ **FLOATING
C7711 S.n7018 SUB 0.10fF $ **FLOATING
C7712 S.n7019 SUB 0.30fF $ **FLOATING
C7713 S.n7020 SUB 0.69fF $ **FLOATING
C7714 S.n7021 SUB 0.45fF $ **FLOATING
C7715 S.n7022 SUB 2.33fF $ **FLOATING
C7716 S.n7023 SUB 0.12fF $ **FLOATING
C7717 S.t368 SUB 0.02fF
C7718 S.n7024 SUB 0.14fF $ **FLOATING
C7719 S.t913 SUB 0.02fF
C7720 S.n7026 SUB 0.24fF $ **FLOATING
C7721 S.n7027 SUB 0.36fF $ **FLOATING
C7722 S.n7028 SUB 0.61fF $ **FLOATING
C7723 S.n7029 SUB 1.90fF $ **FLOATING
C7724 S.n7030 SUB 0.17fF $ **FLOATING
C7725 S.n7031 SUB 0.76fF $ **FLOATING
C7726 S.n7032 SUB 0.32fF $ **FLOATING
C7727 S.n7033 SUB 0.25fF $ **FLOATING
C7728 S.n7034 SUB 0.30fF $ **FLOATING
C7729 S.n7035 SUB 0.47fF $ **FLOATING
C7730 S.n7036 SUB 0.16fF $ **FLOATING
C7731 S.n7037 SUB 1.93fF $ **FLOATING
C7732 S.t591 SUB 0.02fF
C7733 S.n7038 SUB 0.12fF $ **FLOATING
C7734 S.n7039 SUB 0.14fF $ **FLOATING
C7735 S.t1745 SUB 0.02fF
C7736 S.n7041 SUB 0.24fF $ **FLOATING
C7737 S.n7042 SUB 0.91fF $ **FLOATING
C7738 S.n7043 SUB 0.05fF $ **FLOATING
C7739 S.n7044 SUB 1.88fF $ **FLOATING
C7740 S.n7045 SUB 0.12fF $ **FLOATING
C7741 S.t253 SUB 0.02fF
C7742 S.n7046 SUB 0.14fF $ **FLOATING
C7743 S.t933 SUB 0.02fF
C7744 S.n7048 SUB 0.12fF $ **FLOATING
C7745 S.n7049 SUB 0.14fF $ **FLOATING
C7746 S.t452 SUB 0.02fF
C7747 S.n7051 SUB 0.24fF $ **FLOATING
C7748 S.n7052 SUB 0.91fF $ **FLOATING
C7749 S.n7053 SUB 0.05fF $ **FLOATING
C7750 S.t2017 SUB 0.02fF
C7751 S.n7054 SUB 0.24fF $ **FLOATING
C7752 S.n7055 SUB 0.36fF $ **FLOATING
C7753 S.n7056 SUB 0.61fF $ **FLOATING
C7754 S.n7057 SUB 0.32fF $ **FLOATING
C7755 S.n7058 SUB 1.09fF $ **FLOATING
C7756 S.n7059 SUB 0.15fF $ **FLOATING
C7757 S.n7060 SUB 2.10fF $ **FLOATING
C7758 S.n7061 SUB 2.94fF $ **FLOATING
C7759 S.n7062 SUB 1.88fF $ **FLOATING
C7760 S.n7063 SUB 0.12fF $ **FLOATING
C7761 S.t1598 SUB 0.02fF
C7762 S.n7064 SUB 0.14fF $ **FLOATING
C7763 S.t2176 SUB 0.02fF
C7764 S.n7066 SUB 0.24fF $ **FLOATING
C7765 S.n7067 SUB 0.36fF $ **FLOATING
C7766 S.n7068 SUB 0.61fF $ **FLOATING
C7767 S.n7069 SUB 0.92fF $ **FLOATING
C7768 S.n7070 SUB 0.32fF $ **FLOATING
C7769 S.n7071 SUB 0.92fF $ **FLOATING
C7770 S.n7072 SUB 1.09fF $ **FLOATING
C7771 S.n7073 SUB 0.15fF $ **FLOATING
C7772 S.n7074 SUB 4.96fF $ **FLOATING
C7773 S.t1836 SUB 0.02fF
C7774 S.n7075 SUB 0.12fF $ **FLOATING
C7775 S.n7076 SUB 0.14fF $ **FLOATING
C7776 S.t2062 SUB 0.02fF
C7777 S.n7078 SUB 0.24fF $ **FLOATING
C7778 S.n7079 SUB 0.91fF $ **FLOATING
C7779 S.n7080 SUB 0.05fF $ **FLOATING
C7780 S.n7081 SUB 1.88fF $ **FLOATING
C7781 S.n7082 SUB 2.67fF $ **FLOATING
C7782 S.t1312 SUB 0.02fF
C7783 S.n7083 SUB 0.24fF $ **FLOATING
C7784 S.n7084 SUB 0.36fF $ **FLOATING
C7785 S.n7085 SUB 0.61fF $ **FLOATING
C7786 S.n7086 SUB 0.12fF $ **FLOATING
C7787 S.t735 SUB 0.02fF
C7788 S.n7087 SUB 0.14fF $ **FLOATING
C7789 S.n7089 SUB 1.88fF $ **FLOATING
C7790 S.n7090 SUB 2.67fF $ **FLOATING
C7791 S.t1164 SUB 0.02fF
C7792 S.n7091 SUB 0.24fF $ **FLOATING
C7793 S.n7092 SUB 0.36fF $ **FLOATING
C7794 S.n7093 SUB 0.61fF $ **FLOATING
C7795 S.t2097 SUB 0.02fF
C7796 S.n7094 SUB 0.24fF $ **FLOATING
C7797 S.n7095 SUB 0.91fF $ **FLOATING
C7798 S.n7096 SUB 0.05fF $ **FLOATING
C7799 S.t2576 SUB 0.02fF
C7800 S.n7097 SUB 0.12fF $ **FLOATING
C7801 S.n7098 SUB 0.14fF $ **FLOATING
C7802 S.n7100 SUB 0.12fF $ **FLOATING
C7803 S.t1920 SUB 0.02fF
C7804 S.n7101 SUB 0.14fF $ **FLOATING
C7805 S.n7103 SUB 2.30fF $ **FLOATING
C7806 S.n7104 SUB 2.94fF $ **FLOATING
C7807 S.n7105 SUB 5.16fF $ **FLOATING
C7808 S.t970 SUB 0.02fF
C7809 S.n7106 SUB 0.12fF $ **FLOATING
C7810 S.n7107 SUB 0.14fF $ **FLOATING
C7811 S.t1200 SUB 0.02fF
C7812 S.n7109 SUB 0.24fF $ **FLOATING
C7813 S.n7110 SUB 0.91fF $ **FLOATING
C7814 S.n7111 SUB 0.05fF $ **FLOATING
C7815 S.n7112 SUB 1.88fF $ **FLOATING
C7816 S.n7113 SUB 2.67fF $ **FLOATING
C7817 S.t435 SUB 0.02fF
C7818 S.n7114 SUB 0.24fF $ **FLOATING
C7819 S.n7115 SUB 0.36fF $ **FLOATING
C7820 S.n7116 SUB 0.61fF $ **FLOATING
C7821 S.n7117 SUB 0.12fF $ **FLOATING
C7822 S.t2385 SUB 0.02fF
C7823 S.n7118 SUB 0.14fF $ **FLOATING
C7824 S.n7120 SUB 5.17fF $ **FLOATING
C7825 S.t38 SUB 0.02fF
C7826 S.n7121 SUB 0.12fF $ **FLOATING
C7827 S.n7122 SUB 0.14fF $ **FLOATING
C7828 S.t322 SUB 0.02fF
C7829 S.n7124 SUB 0.24fF $ **FLOATING
C7830 S.n7125 SUB 0.91fF $ **FLOATING
C7831 S.n7126 SUB 0.05fF $ **FLOATING
C7832 S.n7127 SUB 1.88fF $ **FLOATING
C7833 S.n7128 SUB 2.67fF $ **FLOATING
C7834 S.t2224 SUB 0.02fF
C7835 S.n7129 SUB 0.24fF $ **FLOATING
C7836 S.n7130 SUB 0.36fF $ **FLOATING
C7837 S.n7131 SUB 0.61fF $ **FLOATING
C7838 S.n7132 SUB 0.12fF $ **FLOATING
C7839 S.t1646 SUB 0.02fF
C7840 S.n7133 SUB 0.14fF $ **FLOATING
C7841 S.n7135 SUB 5.17fF $ **FLOATING
C7842 S.t1735 SUB 0.02fF
C7843 S.n7136 SUB 0.12fF $ **FLOATING
C7844 S.n7137 SUB 0.14fF $ **FLOATING
C7845 S.t2121 SUB 0.02fF
C7846 S.n7139 SUB 0.24fF $ **FLOATING
C7847 S.n7140 SUB 0.91fF $ **FLOATING
C7848 S.n7141 SUB 0.05fF $ **FLOATING
C7849 S.n7142 SUB 1.88fF $ **FLOATING
C7850 S.n7143 SUB 2.67fF $ **FLOATING
C7851 S.t1362 SUB 0.02fF
C7852 S.n7144 SUB 0.24fF $ **FLOATING
C7853 S.n7145 SUB 0.36fF $ **FLOATING
C7854 S.n7146 SUB 0.61fF $ **FLOATING
C7855 S.n7147 SUB 0.12fF $ **FLOATING
C7856 S.t777 SUB 0.02fF
C7857 S.n7148 SUB 0.14fF $ **FLOATING
C7858 S.n7150 SUB 5.17fF $ **FLOATING
C7859 S.t861 SUB 0.02fF
C7860 S.n7151 SUB 0.12fF $ **FLOATING
C7861 S.n7152 SUB 0.14fF $ **FLOATING
C7862 S.t1253 SUB 0.02fF
C7863 S.n7154 SUB 0.24fF $ **FLOATING
C7864 S.n7155 SUB 0.91fF $ **FLOATING
C7865 S.n7156 SUB 0.05fF $ **FLOATING
C7866 S.n7157 SUB 1.88fF $ **FLOATING
C7867 S.n7158 SUB 2.67fF $ **FLOATING
C7868 S.t489 SUB 0.02fF
C7869 S.n7159 SUB 0.24fF $ **FLOATING
C7870 S.n7160 SUB 0.36fF $ **FLOATING
C7871 S.n7161 SUB 0.61fF $ **FLOATING
C7872 S.n7162 SUB 0.12fF $ **FLOATING
C7873 S.t2429 SUB 0.02fF
C7874 S.n7163 SUB 0.14fF $ **FLOATING
C7875 S.n7165 SUB 5.17fF $ **FLOATING
C7876 S.t2506 SUB 0.02fF
C7877 S.n7166 SUB 0.12fF $ **FLOATING
C7878 S.n7167 SUB 0.14fF $ **FLOATING
C7879 S.t371 SUB 0.02fF
C7880 S.n7169 SUB 0.24fF $ **FLOATING
C7881 S.n7170 SUB 0.91fF $ **FLOATING
C7882 S.n7171 SUB 0.05fF $ **FLOATING
C7883 S.n7172 SUB 1.88fF $ **FLOATING
C7884 S.n7173 SUB 2.67fF $ **FLOATING
C7885 S.t2134 SUB 0.02fF
C7886 S.n7174 SUB 0.24fF $ **FLOATING
C7887 S.n7175 SUB 0.36fF $ **FLOATING
C7888 S.n7176 SUB 0.61fF $ **FLOATING
C7889 S.n7177 SUB 0.12fF $ **FLOATING
C7890 S.t1565 SUB 0.02fF
C7891 S.n7178 SUB 0.14fF $ **FLOATING
C7892 S.n7180 SUB 4.90fF $ **FLOATING
C7893 S.t1631 SUB 0.02fF
C7894 S.n7181 SUB 0.12fF $ **FLOATING
C7895 S.n7182 SUB 0.14fF $ **FLOATING
C7896 S.t2024 SUB 0.02fF
C7897 S.n7184 SUB 0.24fF $ **FLOATING
C7898 S.n7185 SUB 0.91fF $ **FLOATING
C7899 S.n7186 SUB 0.05fF $ **FLOATING
C7900 S.n7187 SUB 1.88fF $ **FLOATING
C7901 S.n7188 SUB 2.67fF $ **FLOATING
C7902 S.t2183 SUB 0.02fF
C7903 S.n7189 SUB 0.24fF $ **FLOATING
C7904 S.n7190 SUB 0.36fF $ **FLOATING
C7905 S.n7191 SUB 0.61fF $ **FLOATING
C7906 S.n7192 SUB 0.12fF $ **FLOATING
C7907 S.t898 SUB 0.02fF
C7908 S.n7193 SUB 0.14fF $ **FLOATING
C7909 S.n7195 SUB 1.88fF $ **FLOATING
C7910 S.n7196 SUB 2.68fF $ **FLOATING
C7911 S.t1022 SUB 0.02fF
C7912 S.n7197 SUB 0.24fF $ **FLOATING
C7913 S.n7198 SUB 0.36fF $ **FLOATING
C7914 S.n7199 SUB 0.61fF $ **FLOATING
C7915 S.t2269 SUB 0.02fF
C7916 S.n7200 SUB 1.22fF $ **FLOATING
C7917 S.n7201 SUB 0.36fF $ **FLOATING
C7918 S.n7202 SUB 1.22fF $ **FLOATING
C7919 S.n7203 SUB 0.61fF $ **FLOATING
C7920 S.n7204 SUB 0.35fF $ **FLOATING
C7921 S.n7205 SUB 0.63fF $ **FLOATING
C7922 S.n7206 SUB 1.15fF $ **FLOATING
C7923 S.n7207 SUB 3.03fF $ **FLOATING
C7924 S.n7208 SUB 0.59fF $ **FLOATING
C7925 S.n7209 SUB 0.02fF $ **FLOATING
C7926 S.n7210 SUB 0.97fF $ **FLOATING
C7927 S.t219 SUB 21.38fF
C7928 S.n7211 SUB 20.25fF $ **FLOATING
C7929 S.n7213 SUB 0.38fF $ **FLOATING
C7930 S.n7214 SUB 0.23fF $ **FLOATING
C7931 S.n7215 SUB 2.79fF $ **FLOATING
C7932 S.n7216 SUB 2.46fF $ **FLOATING
C7933 S.n7217 SUB 4.00fF $ **FLOATING
C7934 S.n7218 SUB 0.25fF $ **FLOATING
C7935 S.n7219 SUB 0.01fF $ **FLOATING
C7936 S.t1976 SUB 0.02fF
C7937 S.n7220 SUB 0.25fF $ **FLOATING
C7938 S.t1700 SUB 0.02fF
C7939 S.n7221 SUB 0.95fF $ **FLOATING
C7940 S.n7222 SUB 0.70fF $ **FLOATING
C7941 S.n7223 SUB 1.89fF $ **FLOATING
C7942 S.n7224 SUB 1.88fF $ **FLOATING
C7943 S.t1410 SUB 0.02fF
C7944 S.n7225 SUB 0.24fF $ **FLOATING
C7945 S.n7226 SUB 0.36fF $ **FLOATING
C7946 S.n7227 SUB 0.61fF $ **FLOATING
C7947 S.n7228 SUB 0.12fF $ **FLOATING
C7948 S.t1122 SUB 0.02fF
C7949 S.n7229 SUB 0.14fF $ **FLOATING
C7950 S.n7231 SUB 1.16fF $ **FLOATING
C7951 S.n7232 SUB 0.22fF $ **FLOATING
C7952 S.n7233 SUB 0.25fF $ **FLOATING
C7953 S.n7234 SUB 0.09fF $ **FLOATING
C7954 S.n7235 SUB 1.88fF $ **FLOATING
C7955 S.t826 SUB 0.02fF
C7956 S.n7236 SUB 0.24fF $ **FLOATING
C7957 S.n7237 SUB 0.91fF $ **FLOATING
C7958 S.n7238 SUB 0.05fF $ **FLOATING
C7959 S.t1786 SUB 0.02fF
C7960 S.n7239 SUB 0.12fF $ **FLOATING
C7961 S.n7240 SUB 0.14fF $ **FLOATING
C7962 S.n7242 SUB 0.78fF $ **FLOATING
C7963 S.n7243 SUB 1.94fF $ **FLOATING
C7964 S.n7244 SUB 1.88fF $ **FLOATING
C7965 S.n7245 SUB 0.12fF $ **FLOATING
C7966 S.t244 SUB 0.02fF
C7967 S.n7246 SUB 0.14fF $ **FLOATING
C7968 S.t545 SUB 0.02fF
C7969 S.n7248 SUB 0.24fF $ **FLOATING
C7970 S.n7249 SUB 0.36fF $ **FLOATING
C7971 S.n7250 SUB 0.61fF $ **FLOATING
C7972 S.n7251 SUB 1.84fF $ **FLOATING
C7973 S.n7252 SUB 2.99fF $ **FLOATING
C7974 S.t2470 SUB 0.02fF
C7975 S.n7253 SUB 0.24fF $ **FLOATING
C7976 S.n7254 SUB 0.91fF $ **FLOATING
C7977 S.n7255 SUB 0.05fF $ **FLOATING
C7978 S.t920 SUB 0.02fF
C7979 S.n7256 SUB 0.12fF $ **FLOATING
C7980 S.n7257 SUB 0.14fF $ **FLOATING
C7981 S.n7259 SUB 1.89fF $ **FLOATING
C7982 S.n7260 SUB 1.88fF $ **FLOATING
C7983 S.t2186 SUB 0.02fF
C7984 S.n7261 SUB 0.24fF $ **FLOATING
C7985 S.n7262 SUB 0.36fF $ **FLOATING
C7986 S.n7263 SUB 0.61fF $ **FLOATING
C7987 S.n7264 SUB 0.12fF $ **FLOATING
C7988 S.t1910 SUB 0.02fF
C7989 S.n7265 SUB 0.14fF $ **FLOATING
C7990 S.n7267 SUB 1.16fF $ **FLOATING
C7991 S.n7268 SUB 0.22fF $ **FLOATING
C7992 S.n7269 SUB 0.25fF $ **FLOATING
C7993 S.n7270 SUB 0.09fF $ **FLOATING
C7994 S.n7271 SUB 1.88fF $ **FLOATING
C7995 S.t1600 SUB 0.02fF
C7996 S.n7272 SUB 0.24fF $ **FLOATING
C7997 S.n7273 SUB 0.91fF $ **FLOATING
C7998 S.n7274 SUB 0.05fF $ **FLOATING
C7999 S.t178 SUB 0.02fF
C8000 S.n7275 SUB 0.12fF $ **FLOATING
C8001 S.n7276 SUB 0.14fF $ **FLOATING
C8002 S.n7278 SUB 0.78fF $ **FLOATING
C8003 S.n7279 SUB 1.94fF $ **FLOATING
C8004 S.n7280 SUB 1.88fF $ **FLOATING
C8005 S.n7281 SUB 0.12fF $ **FLOATING
C8006 S.t1051 SUB 0.02fF
C8007 S.n7282 SUB 0.14fF $ **FLOATING
C8008 S.t1323 SUB 0.02fF
C8009 S.n7284 SUB 0.24fF $ **FLOATING
C8010 S.n7285 SUB 0.36fF $ **FLOATING
C8011 S.n7286 SUB 0.61fF $ **FLOATING
C8012 S.n7287 SUB 1.84fF $ **FLOATING
C8013 S.n7288 SUB 2.99fF $ **FLOATING
C8014 S.t736 SUB 0.02fF
C8015 S.n7289 SUB 0.24fF $ **FLOATING
C8016 S.n7290 SUB 0.91fF $ **FLOATING
C8017 S.n7291 SUB 0.05fF $ **FLOATING
C8018 S.t1843 SUB 0.02fF
C8019 S.n7292 SUB 0.12fF $ **FLOATING
C8020 S.n7293 SUB 0.14fF $ **FLOATING
C8021 S.n7295 SUB 1.89fF $ **FLOATING
C8022 S.n7296 SUB 1.75fF $ **FLOATING
C8023 S.t443 SUB 0.02fF
C8024 S.n7297 SUB 0.24fF $ **FLOATING
C8025 S.n7298 SUB 0.36fF $ **FLOATING
C8026 S.n7299 SUB 0.61fF $ **FLOATING
C8027 S.n7300 SUB 0.12fF $ **FLOATING
C8028 S.t162 SUB 0.02fF
C8029 S.n7301 SUB 0.14fF $ **FLOATING
C8030 S.n7303 SUB 1.16fF $ **FLOATING
C8031 S.n7304 SUB 0.22fF $ **FLOATING
C8032 S.n7305 SUB 0.25fF $ **FLOATING
C8033 S.n7306 SUB 0.09fF $ **FLOATING
C8034 S.n7307 SUB 2.44fF $ **FLOATING
C8035 S.t2386 SUB 0.02fF
C8036 S.n7308 SUB 0.24fF $ **FLOATING
C8037 S.n7309 SUB 0.91fF $ **FLOATING
C8038 S.n7310 SUB 0.05fF $ **FLOATING
C8039 S.t981 SUB 0.02fF
C8040 S.n7311 SUB 0.12fF $ **FLOATING
C8041 S.n7312 SUB 0.14fF $ **FLOATING
C8042 S.n7314 SUB 1.88fF $ **FLOATING
C8043 S.n7315 SUB 0.48fF $ **FLOATING
C8044 S.n7316 SUB 0.09fF $ **FLOATING
C8045 S.n7317 SUB 0.33fF $ **FLOATING
C8046 S.n7318 SUB 0.30fF $ **FLOATING
C8047 S.n7319 SUB 0.77fF $ **FLOATING
C8048 S.n7320 SUB 0.59fF $ **FLOATING
C8049 S.t2087 SUB 0.02fF
C8050 S.n7321 SUB 0.24fF $ **FLOATING
C8051 S.n7322 SUB 0.36fF $ **FLOATING
C8052 S.n7323 SUB 0.61fF $ **FLOATING
C8053 S.n7324 SUB 0.12fF $ **FLOATING
C8054 S.t1823 SUB 0.02fF
C8055 S.n7325 SUB 0.14fF $ **FLOATING
C8056 S.n7327 SUB 2.61fF $ **FLOATING
C8057 S.n7328 SUB 2.16fF $ **FLOATING
C8058 S.t1530 SUB 0.02fF
C8059 S.n7329 SUB 0.24fF $ **FLOATING
C8060 S.n7330 SUB 0.91fF $ **FLOATING
C8061 S.n7331 SUB 0.05fF $ **FLOATING
C8062 S.t48 SUB 0.02fF
C8063 S.n7332 SUB 0.12fF $ **FLOATING
C8064 S.n7333 SUB 0.14fF $ **FLOATING
C8065 S.n7335 SUB 0.78fF $ **FLOATING
C8066 S.n7336 SUB 2.30fF $ **FLOATING
C8067 S.n7337 SUB 1.88fF $ **FLOATING
C8068 S.n7338 SUB 0.12fF $ **FLOATING
C8069 S.t1084 SUB 0.02fF
C8070 S.n7339 SUB 0.14fF $ **FLOATING
C8071 S.t1223 SUB 0.02fF
C8072 S.n7341 SUB 0.24fF $ **FLOATING
C8073 S.n7342 SUB 0.36fF $ **FLOATING
C8074 S.n7343 SUB 0.61fF $ **FLOATING
C8075 S.n7344 SUB 1.39fF $ **FLOATING
C8076 S.n7345 SUB 0.71fF $ **FLOATING
C8077 S.n7346 SUB 1.14fF $ **FLOATING
C8078 S.n7347 SUB 0.35fF $ **FLOATING
C8079 S.n7348 SUB 2.03fF $ **FLOATING
C8080 S.t670 SUB 0.02fF
C8081 S.n7349 SUB 0.24fF $ **FLOATING
C8082 S.n7350 SUB 0.91fF $ **FLOATING
C8083 S.n7351 SUB 0.05fF $ **FLOATING
C8084 S.t1741 SUB 0.02fF
C8085 S.n7352 SUB 0.12fF $ **FLOATING
C8086 S.n7353 SUB 0.14fF $ **FLOATING
C8087 S.n7355 SUB 1.89fF $ **FLOATING
C8088 S.n7356 SUB 1.88fF $ **FLOATING
C8089 S.t365 SUB 0.02fF
C8090 S.n7357 SUB 0.24fF $ **FLOATING
C8091 S.n7358 SUB 0.36fF $ **FLOATING
C8092 S.n7359 SUB 0.61fF $ **FLOATING
C8093 S.n7360 SUB 0.12fF $ **FLOATING
C8094 S.t1133 SUB 0.02fF
C8095 S.n7361 SUB 0.14fF $ **FLOATING
C8096 S.n7363 SUB 1.16fF $ **FLOATING
C8097 S.n7364 SUB 0.22fF $ **FLOATING
C8098 S.n7365 SUB 0.25fF $ **FLOATING
C8099 S.n7366 SUB 0.09fF $ **FLOATING
C8100 S.n7367 SUB 1.88fF $ **FLOATING
C8101 S.t1331 SUB 0.02fF
C8102 S.n7368 SUB 0.24fF $ **FLOATING
C8103 S.n7369 SUB 0.91fF $ **FLOATING
C8104 S.n7370 SUB 0.05fF $ **FLOATING
C8105 S.t865 SUB 0.02fF
C8106 S.n7371 SUB 0.12fF $ **FLOATING
C8107 S.n7372 SUB 0.14fF $ **FLOATING
C8108 S.n7374 SUB 20.78fF $ **FLOATING
C8109 S.n7375 SUB 1.88fF $ **FLOATING
C8110 S.n7376 SUB 2.67fF $ **FLOATING
C8111 S.t291 SUB 0.02fF
C8112 S.n7377 SUB 0.24fF $ **FLOATING
C8113 S.n7378 SUB 0.36fF $ **FLOATING
C8114 S.n7379 SUB 0.61fF $ **FLOATING
C8115 S.n7380 SUB 0.12fF $ **FLOATING
C8116 S.t1060 SUB 0.02fF
C8117 S.n7381 SUB 0.14fF $ **FLOATING
C8118 S.n7383 SUB 2.80fF $ **FLOATING
C8119 S.n7384 SUB 2.30fF $ **FLOATING
C8120 S.t1699 SUB 0.02fF
C8121 S.n7385 SUB 0.12fF $ **FLOATING
C8122 S.n7386 SUB 0.14fF $ **FLOATING
C8123 S.t1232 SUB 0.02fF
C8124 S.n7388 SUB 0.24fF $ **FLOATING
C8125 S.n7389 SUB 0.91fF $ **FLOATING
C8126 S.n7390 SUB 0.05fF $ **FLOATING
C8127 S.n7391 SUB 1.88fF $ **FLOATING
C8128 S.n7392 SUB 2.67fF $ **FLOATING
C8129 S.t1954 SUB 0.02fF
C8130 S.n7393 SUB 0.24fF $ **FLOATING
C8131 S.n7394 SUB 0.36fF $ **FLOATING
C8132 S.n7395 SUB 0.61fF $ **FLOATING
C8133 S.n7396 SUB 0.12fF $ **FLOATING
C8134 S.t175 SUB 0.02fF
C8135 S.n7397 SUB 0.14fF $ **FLOATING
C8136 S.n7399 SUB 2.80fF $ **FLOATING
C8137 S.n7400 SUB 2.30fF $ **FLOATING
C8138 S.t825 SUB 0.02fF
C8139 S.n7401 SUB 0.12fF $ **FLOATING
C8140 S.n7402 SUB 0.14fF $ **FLOATING
C8141 S.t349 SUB 0.02fF
C8142 S.n7404 SUB 0.24fF $ **FLOATING
C8143 S.n7405 SUB 0.91fF $ **FLOATING
C8144 S.n7406 SUB 0.05fF $ **FLOATING
C8145 S.n7407 SUB 1.88fF $ **FLOATING
C8146 S.n7408 SUB 2.67fF $ **FLOATING
C8147 S.t1094 SUB 0.02fF
C8148 S.n7409 SUB 0.24fF $ **FLOATING
C8149 S.n7410 SUB 0.36fF $ **FLOATING
C8150 S.n7411 SUB 0.61fF $ **FLOATING
C8151 S.n7412 SUB 0.12fF $ **FLOATING
C8152 S.t1839 SUB 0.02fF
C8153 S.n7413 SUB 0.14fF $ **FLOATING
C8154 S.n7415 SUB 2.80fF $ **FLOATING
C8155 S.n7416 SUB 2.30fF $ **FLOATING
C8156 S.t76 SUB 0.02fF
C8157 S.n7417 SUB 0.12fF $ **FLOATING
C8158 S.n7418 SUB 0.14fF $ **FLOATING
C8159 S.t2006 SUB 0.02fF
C8160 S.n7420 SUB 0.24fF $ **FLOATING
C8161 S.n7421 SUB 0.91fF $ **FLOATING
C8162 S.n7422 SUB 0.05fF $ **FLOATING
C8163 S.n7423 SUB 1.88fF $ **FLOATING
C8164 S.n7424 SUB 2.67fF $ **FLOATING
C8165 S.t220 SUB 0.02fF
C8166 S.n7425 SUB 0.24fF $ **FLOATING
C8167 S.n7426 SUB 0.36fF $ **FLOATING
C8168 S.n7427 SUB 0.61fF $ **FLOATING
C8169 S.n7428 SUB 0.12fF $ **FLOATING
C8170 S.t974 SUB 0.02fF
C8171 S.n7429 SUB 0.14fF $ **FLOATING
C8172 S.n7431 SUB 2.80fF $ **FLOATING
C8173 S.n7432 SUB 2.30fF $ **FLOATING
C8174 S.t1757 SUB 0.02fF
C8175 S.n7433 SUB 0.12fF $ **FLOATING
C8176 S.n7434 SUB 0.14fF $ **FLOATING
C8177 S.t1156 SUB 0.02fF
C8178 S.n7436 SUB 0.24fF $ **FLOATING
C8179 S.n7437 SUB 0.91fF $ **FLOATING
C8180 S.n7438 SUB 0.05fF $ **FLOATING
C8181 S.n7439 SUB 1.88fF $ **FLOATING
C8182 S.n7440 SUB 2.67fF $ **FLOATING
C8183 S.t1884 SUB 0.02fF
C8184 S.n7441 SUB 0.24fF $ **FLOATING
C8185 S.n7442 SUB 0.36fF $ **FLOATING
C8186 S.n7443 SUB 0.61fF $ **FLOATING
C8187 S.n7444 SUB 0.12fF $ **FLOATING
C8188 S.t41 SUB 0.02fF
C8189 S.n7445 SUB 0.14fF $ **FLOATING
C8190 S.n7447 SUB 2.80fF $ **FLOATING
C8191 S.n7448 SUB 2.30fF $ **FLOATING
C8192 S.t879 SUB 0.02fF
C8193 S.n7449 SUB 0.12fF $ **FLOATING
C8194 S.n7450 SUB 0.14fF $ **FLOATING
C8195 S.t282 SUB 0.02fF
C8196 S.n7452 SUB 0.24fF $ **FLOATING
C8197 S.n7453 SUB 0.91fF $ **FLOATING
C8198 S.n7454 SUB 0.05fF $ **FLOATING
C8199 S.n7455 SUB 2.73fF $ **FLOATING
C8200 S.n7456 SUB 1.59fF $ **FLOATING
C8201 S.n7457 SUB 0.12fF $ **FLOATING
C8202 S.t711 SUB 0.02fF
C8203 S.n7458 SUB 0.14fF $ **FLOATING
C8204 S.t2153 SUB 0.02fF
C8205 S.n7460 SUB 0.24fF $ **FLOATING
C8206 S.n7461 SUB 0.36fF $ **FLOATING
C8207 S.n7462 SUB 0.61fF $ **FLOATING
C8208 S.n7463 SUB 0.07fF $ **FLOATING
C8209 S.n7464 SUB 0.01fF $ **FLOATING
C8210 S.n7465 SUB 0.24fF $ **FLOATING
C8211 S.n7466 SUB 1.16fF $ **FLOATING
C8212 S.n7467 SUB 1.35fF $ **FLOATING
C8213 S.n7468 SUB 2.30fF $ **FLOATING
C8214 S.t1486 SUB 0.02fF
C8215 S.n7469 SUB 0.12fF $ **FLOATING
C8216 S.n7470 SUB 0.14fF $ **FLOATING
C8217 S.t2445 SUB 0.02fF
C8218 S.n7472 SUB 0.24fF $ **FLOATING
C8219 S.n7473 SUB 0.91fF $ **FLOATING
C8220 S.n7474 SUB 0.05fF $ **FLOATING
C8221 S.t40 SUB 48.31fF
C8222 S.t1941 SUB 0.02fF
C8223 S.n7475 SUB 0.24fF $ **FLOATING
C8224 S.n7476 SUB 0.91fF $ **FLOATING
C8225 S.n7477 SUB 0.05fF $ **FLOATING
C8226 S.t2524 SUB 0.02fF
C8227 S.n7478 SUB 0.12fF $ **FLOATING
C8228 S.n7479 SUB 0.14fF $ **FLOATING
C8229 S.n7481 SUB 0.12fF $ **FLOATING
C8230 S.t1736 SUB 0.02fF
C8231 S.n7482 SUB 0.14fF $ **FLOATING
C8232 S.n7484 SUB 5.17fF $ **FLOATING
C8233 S.n7485 SUB 5.44fF $ **FLOATING
C8234 S.t763 SUB 0.02fF
C8235 S.n7486 SUB 0.12fF $ **FLOATING
C8236 S.n7487 SUB 0.14fF $ **FLOATING
C8237 S.t971 SUB 0.02fF
C8238 S.n7489 SUB 0.24fF $ **FLOATING
C8239 S.n7490 SUB 0.91fF $ **FLOATING
C8240 S.n7491 SUB 0.05fF $ **FLOATING
C8241 S.t37 SUB 47.92fF
C8242 S.t2091 SUB 0.02fF
C8243 S.n7492 SUB 1.19fF $ **FLOATING
C8244 S.n7493 SUB 0.05fF $ **FLOATING
C8245 S.t150 SUB 0.02fF
C8246 S.n7494 SUB 0.01fF $ **FLOATING
C8247 S.n7495 SUB 0.26fF $ **FLOATING
C8248 S.n7497 SUB 1.50fF $ **FLOATING
C8249 S.n7498 SUB 1.30fF $ **FLOATING
C8250 S.n7499 SUB 0.28fF $ **FLOATING
C8251 S.n7500 SUB 0.24fF $ **FLOATING
C8252 S.n7501 SUB 4.39fF $ **FLOATING
C8253 S.n7502 SUB 0.01fF $ **FLOATING
C8254 S.n7503 SUB 0.02fF $ **FLOATING
C8255 S.n7504 SUB 0.03fF $ **FLOATING
C8256 S.n7505 SUB 0.04fF $ **FLOATING
C8257 S.n7506 SUB 0.17fF $ **FLOATING
C8258 S.n7507 SUB 0.01fF $ **FLOATING
C8259 S.n7508 SUB 0.02fF $ **FLOATING
C8260 S.n7509 SUB 0.01fF $ **FLOATING
C8261 S.n7510 SUB 0.01fF $ **FLOATING
C8262 S.n7511 SUB 0.01fF $ **FLOATING
C8263 S.n7512 SUB 0.01fF $ **FLOATING
C8264 S.n7513 SUB 0.02fF $ **FLOATING
C8265 S.n7514 SUB 0.01fF $ **FLOATING
C8266 S.n7515 SUB 0.02fF $ **FLOATING
C8267 S.n7516 SUB 0.05fF $ **FLOATING
C8268 S.n7517 SUB 0.04fF $ **FLOATING
C8269 S.n7518 SUB 0.11fF $ **FLOATING
C8270 S.n7519 SUB 0.38fF $ **FLOATING
C8271 S.n7520 SUB 0.20fF $ **FLOATING
C8272 S.n7521 SUB 8.97fF $ **FLOATING
C8273 S.n7522 SUB 8.97fF $ **FLOATING
C8274 S.n7523 SUB 0.60fF $ **FLOATING
C8275 S.n7524 SUB 0.22fF $ **FLOATING
C8276 S.n7525 SUB 0.59fF $ **FLOATING
C8277 S.n7526 SUB 3.43fF $ **FLOATING
C8278 S.n7527 SUB 0.29fF $ **FLOATING
C8279 S.t299 SUB 21.38fF
C8280 S.n7528 SUB 21.67fF $ **FLOATING
C8281 S.n7529 SUB 0.77fF $ **FLOATING
C8282 S.n7530 SUB 0.28fF $ **FLOATING
C8283 S.n7531 SUB 4.00fF $ **FLOATING
C8284 S.n7532 SUB 1.35fF $ **FLOATING
C8285 S.t1368 SUB 0.02fF
C8286 S.n7533 SUB 0.64fF $ **FLOATING
C8287 S.n7534 SUB 0.61fF $ **FLOATING
C8288 S.n7535 SUB 0.25fF $ **FLOATING
C8289 S.n7536 SUB 0.09fF $ **FLOATING
C8290 S.n7537 SUB 0.21fF $ **FLOATING
C8291 S.n7538 SUB 0.92fF $ **FLOATING
C8292 S.n7539 SUB 0.44fF $ **FLOATING
C8293 S.n7540 SUB 1.88fF $ **FLOATING
C8294 S.n7541 SUB 0.12fF $ **FLOATING
C8295 S.t1747 SUB 0.02fF
C8296 S.n7542 SUB 0.14fF $ **FLOATING
C8297 S.t2285 SUB 0.02fF
C8298 S.n7544 SUB 0.24fF $ **FLOATING
C8299 S.n7545 SUB 0.36fF $ **FLOATING
C8300 S.n7546 SUB 0.61fF $ **FLOATING
C8301 S.n7547 SUB 0.02fF $ **FLOATING
C8302 S.n7548 SUB 0.01fF $ **FLOATING
C8303 S.n7549 SUB 0.02fF $ **FLOATING
C8304 S.n7550 SUB 0.08fF $ **FLOATING
C8305 S.n7551 SUB 0.06fF $ **FLOATING
C8306 S.n7552 SUB 0.03fF $ **FLOATING
C8307 S.n7553 SUB 0.04fF $ **FLOATING
C8308 S.n7554 SUB 1.00fF $ **FLOATING
C8309 S.n7555 SUB 0.36fF $ **FLOATING
C8310 S.n7556 SUB 1.87fF $ **FLOATING
C8311 S.n7557 SUB 1.99fF $ **FLOATING
C8312 S.t604 SUB 0.02fF
C8313 S.n7558 SUB 0.24fF $ **FLOATING
C8314 S.n7559 SUB 0.91fF $ **FLOATING
C8315 S.n7560 SUB 0.05fF $ **FLOATING
C8316 S.t1948 SUB 0.02fF
C8317 S.n7561 SUB 0.12fF $ **FLOATING
C8318 S.n7562 SUB 0.14fF $ **FLOATING
C8319 S.n7564 SUB 1.89fF $ **FLOATING
C8320 S.n7565 SUB 0.06fF $ **FLOATING
C8321 S.n7566 SUB 0.03fF $ **FLOATING
C8322 S.n7567 SUB 0.04fF $ **FLOATING
C8323 S.n7568 SUB 0.99fF $ **FLOATING
C8324 S.n7569 SUB 0.02fF $ **FLOATING
C8325 S.n7570 SUB 0.01fF $ **FLOATING
C8326 S.n7571 SUB 0.02fF $ **FLOATING
C8327 S.n7572 SUB 0.08fF $ **FLOATING
C8328 S.n7573 SUB 0.36fF $ **FLOATING
C8329 S.n7574 SUB 1.85fF $ **FLOATING
C8330 S.t1525 SUB 0.02fF
C8331 S.n7575 SUB 0.24fF $ **FLOATING
C8332 S.n7576 SUB 0.36fF $ **FLOATING
C8333 S.n7577 SUB 0.61fF $ **FLOATING
C8334 S.n7578 SUB 0.12fF $ **FLOATING
C8335 S.t1029 SUB 0.02fF
C8336 S.n7579 SUB 0.14fF $ **FLOATING
C8337 S.n7581 SUB 0.70fF $ **FLOATING
C8338 S.n7582 SUB 0.23fF $ **FLOATING
C8339 S.n7583 SUB 0.23fF $ **FLOATING
C8340 S.n7584 SUB 0.70fF $ **FLOATING
C8341 S.n7585 SUB 1.16fF $ **FLOATING
C8342 S.n7586 SUB 0.22fF $ **FLOATING
C8343 S.n7587 SUB 0.25fF $ **FLOATING
C8344 S.n7588 SUB 0.09fF $ **FLOATING
C8345 S.n7589 SUB 1.88fF $ **FLOATING
C8346 S.t2355 SUB 0.02fF
C8347 S.n7590 SUB 0.24fF $ **FLOATING
C8348 S.n7591 SUB 0.91fF $ **FLOATING
C8349 S.n7592 SUB 0.05fF $ **FLOATING
C8350 S.t1090 SUB 0.02fF
C8351 S.n7593 SUB 0.12fF $ **FLOATING
C8352 S.n7594 SUB 0.14fF $ **FLOATING
C8353 S.n7596 SUB 0.25fF $ **FLOATING
C8354 S.n7597 SUB 0.09fF $ **FLOATING
C8355 S.n7598 SUB 0.21fF $ **FLOATING
C8356 S.n7599 SUB 0.92fF $ **FLOATING
C8357 S.n7600 SUB 0.44fF $ **FLOATING
C8358 S.n7601 SUB 1.88fF $ **FLOATING
C8359 S.n7602 SUB 0.12fF $ **FLOATING
C8360 S.t133 SUB 0.02fF
C8361 S.n7603 SUB 0.14fF $ **FLOATING
C8362 S.t665 SUB 0.02fF
C8363 S.n7605 SUB 0.24fF $ **FLOATING
C8364 S.n7606 SUB 0.36fF $ **FLOATING
C8365 S.n7607 SUB 0.61fF $ **FLOATING
C8366 S.n7608 SUB 0.02fF $ **FLOATING
C8367 S.n7609 SUB 0.01fF $ **FLOATING
C8368 S.n7610 SUB 0.02fF $ **FLOATING
C8369 S.n7611 SUB 0.08fF $ **FLOATING
C8370 S.n7612 SUB 0.06fF $ **FLOATING
C8371 S.n7613 SUB 0.03fF $ **FLOATING
C8372 S.n7614 SUB 0.04fF $ **FLOATING
C8373 S.n7615 SUB 1.00fF $ **FLOATING
C8374 S.n7616 SUB 0.36fF $ **FLOATING
C8375 S.n7617 SUB 1.87fF $ **FLOATING
C8376 S.n7618 SUB 1.99fF $ **FLOATING
C8377 S.t1497 SUB 0.02fF
C8378 S.n7619 SUB 0.24fF $ **FLOATING
C8379 S.n7620 SUB 0.91fF $ **FLOATING
C8380 S.n7621 SUB 0.05fF $ **FLOATING
C8381 S.t211 SUB 0.02fF
C8382 S.n7622 SUB 0.12fF $ **FLOATING
C8383 S.n7623 SUB 0.14fF $ **FLOATING
C8384 S.n7625 SUB 1.89fF $ **FLOATING
C8385 S.n7626 SUB 0.07fF $ **FLOATING
C8386 S.n7627 SUB 0.04fF $ **FLOATING
C8387 S.n7628 SUB 0.05fF $ **FLOATING
C8388 S.n7629 SUB 0.87fF $ **FLOATING
C8389 S.n7630 SUB 0.01fF $ **FLOATING
C8390 S.n7631 SUB 0.01fF $ **FLOATING
C8391 S.n7632 SUB 0.01fF $ **FLOATING
C8392 S.n7633 SUB 0.07fF $ **FLOATING
C8393 S.n7634 SUB 0.68fF $ **FLOATING
C8394 S.n7635 SUB 0.72fF $ **FLOATING
C8395 S.t2319 SUB 0.02fF
C8396 S.n7636 SUB 0.24fF $ **FLOATING
C8397 S.n7637 SUB 0.36fF $ **FLOATING
C8398 S.n7638 SUB 0.61fF $ **FLOATING
C8399 S.n7639 SUB 0.12fF $ **FLOATING
C8400 S.t1802 SUB 0.02fF
C8401 S.n7640 SUB 0.14fF $ **FLOATING
C8402 S.n7642 SUB 0.70fF $ **FLOATING
C8403 S.n7643 SUB 0.23fF $ **FLOATING
C8404 S.n7644 SUB 0.23fF $ **FLOATING
C8405 S.n7645 SUB 0.70fF $ **FLOATING
C8406 S.n7646 SUB 1.16fF $ **FLOATING
C8407 S.n7647 SUB 0.22fF $ **FLOATING
C8408 S.n7648 SUB 0.25fF $ **FLOATING
C8409 S.n7649 SUB 0.09fF $ **FLOATING
C8410 S.n7650 SUB 2.31fF $ **FLOATING
C8411 S.t634 SUB 0.02fF
C8412 S.n7651 SUB 0.24fF $ **FLOATING
C8413 S.n7652 SUB 0.91fF $ **FLOATING
C8414 S.n7653 SUB 0.05fF $ **FLOATING
C8415 S.t1879 SUB 0.02fF
C8416 S.n7654 SUB 0.12fF $ **FLOATING
C8417 S.n7655 SUB 0.14fF $ **FLOATING
C8418 S.n7657 SUB 1.88fF $ **FLOATING
C8419 S.n7658 SUB 0.46fF $ **FLOATING
C8420 S.n7659 SUB 0.22fF $ **FLOATING
C8421 S.n7660 SUB 0.38fF $ **FLOATING
C8422 S.n7661 SUB 0.16fF $ **FLOATING
C8423 S.n7662 SUB 0.28fF $ **FLOATING
C8424 S.n7663 SUB 0.21fF $ **FLOATING
C8425 S.n7664 SUB 0.30fF $ **FLOATING
C8426 S.n7665 SUB 0.42fF $ **FLOATING
C8427 S.n7666 SUB 0.21fF $ **FLOATING
C8428 S.t1458 SUB 0.02fF
C8429 S.n7667 SUB 0.24fF $ **FLOATING
C8430 S.n7668 SUB 0.36fF $ **FLOATING
C8431 S.n7669 SUB 0.61fF $ **FLOATING
C8432 S.n7670 SUB 0.12fF $ **FLOATING
C8433 S.t932 SUB 0.02fF
C8434 S.n7671 SUB 0.14fF $ **FLOATING
C8435 S.n7673 SUB 0.04fF $ **FLOATING
C8436 S.n7674 SUB 0.03fF $ **FLOATING
C8437 S.n7675 SUB 0.03fF $ **FLOATING
C8438 S.n7676 SUB 0.10fF $ **FLOATING
C8439 S.n7677 SUB 0.36fF $ **FLOATING
C8440 S.n7678 SUB 0.38fF $ **FLOATING
C8441 S.n7679 SUB 0.11fF $ **FLOATING
C8442 S.n7680 SUB 0.12fF $ **FLOATING
C8443 S.n7681 SUB 0.07fF $ **FLOATING
C8444 S.n7682 SUB 0.12fF $ **FLOATING
C8445 S.n7683 SUB 0.18fF $ **FLOATING
C8446 S.n7684 SUB 4.00fF $ **FLOATING
C8447 S.t2290 SUB 0.02fF
C8448 S.n7685 SUB 0.24fF $ **FLOATING
C8449 S.n7686 SUB 0.91fF $ **FLOATING
C8450 S.n7687 SUB 0.05fF $ **FLOATING
C8451 S.t1015 SUB 0.02fF
C8452 S.n7688 SUB 0.12fF $ **FLOATING
C8453 S.n7689 SUB 0.14fF $ **FLOATING
C8454 S.n7691 SUB 0.25fF $ **FLOATING
C8455 S.n7692 SUB 0.09fF $ **FLOATING
C8456 S.n7693 SUB 0.21fF $ **FLOATING
C8457 S.n7694 SUB 1.28fF $ **FLOATING
C8458 S.n7695 SUB 0.53fF $ **FLOATING
C8459 S.n7696 SUB 1.88fF $ **FLOATING
C8460 S.n7697 SUB 0.12fF $ **FLOATING
C8461 S.t2573 SUB 0.02fF
C8462 S.n7698 SUB 0.14fF $ **FLOATING
C8463 S.t600 SUB 0.02fF
C8464 S.n7700 SUB 0.24fF $ **FLOATING
C8465 S.n7701 SUB 0.36fF $ **FLOATING
C8466 S.n7702 SUB 0.61fF $ **FLOATING
C8467 S.n7703 SUB 1.58fF $ **FLOATING
C8468 S.n7704 SUB 2.45fF $ **FLOATING
C8469 S.t1436 SUB 0.02fF
C8470 S.n7705 SUB 0.24fF $ **FLOATING
C8471 S.n7706 SUB 0.91fF $ **FLOATING
C8472 S.n7707 SUB 0.05fF $ **FLOATING
C8473 S.t111 SUB 0.02fF
C8474 S.n7708 SUB 0.12fF $ **FLOATING
C8475 S.n7709 SUB 0.14fF $ **FLOATING
C8476 S.n7711 SUB 1.89fF $ **FLOATING
C8477 S.n7712 SUB 0.06fF $ **FLOATING
C8478 S.n7713 SUB 0.03fF $ **FLOATING
C8479 S.n7714 SUB 0.04fF $ **FLOATING
C8480 S.n7715 SUB 0.99fF $ **FLOATING
C8481 S.n7716 SUB 0.02fF $ **FLOATING
C8482 S.n7717 SUB 0.01fF $ **FLOATING
C8483 S.n7718 SUB 0.02fF $ **FLOATING
C8484 S.n7719 SUB 0.08fF $ **FLOATING
C8485 S.n7720 SUB 0.36fF $ **FLOATING
C8486 S.n7721 SUB 1.85fF $ **FLOATING
C8487 S.t2251 SUB 0.02fF
C8488 S.n7722 SUB 0.24fF $ **FLOATING
C8489 S.n7723 SUB 0.36fF $ **FLOATING
C8490 S.n7724 SUB 0.61fF $ **FLOATING
C8491 S.n7725 SUB 0.12fF $ **FLOATING
C8492 S.t1696 SUB 0.02fF
C8493 S.n7726 SUB 0.14fF $ **FLOATING
C8494 S.n7728 SUB 0.70fF $ **FLOATING
C8495 S.n7729 SUB 0.23fF $ **FLOATING
C8496 S.n7730 SUB 0.23fF $ **FLOATING
C8497 S.n7731 SUB 0.70fF $ **FLOATING
C8498 S.n7732 SUB 1.16fF $ **FLOATING
C8499 S.n7733 SUB 0.22fF $ **FLOATING
C8500 S.n7734 SUB 0.25fF $ **FLOATING
C8501 S.n7735 SUB 0.09fF $ **FLOATING
C8502 S.n7736 SUB 1.88fF $ **FLOATING
C8503 S.t573 SUB 0.02fF
C8504 S.n7737 SUB 0.24fF $ **FLOATING
C8505 S.n7738 SUB 0.91fF $ **FLOATING
C8506 S.n7739 SUB 0.05fF $ **FLOATING
C8507 S.t1918 SUB 0.02fF
C8508 S.n7740 SUB 0.12fF $ **FLOATING
C8509 S.n7741 SUB 0.14fF $ **FLOATING
C8510 S.n7743 SUB 20.78fF $ **FLOATING
C8511 S.n7744 SUB 1.72fF $ **FLOATING
C8512 S.n7745 SUB 3.05fF $ **FLOATING
C8513 S.t626 SUB 0.02fF
C8514 S.n7746 SUB 0.24fF $ **FLOATING
C8515 S.n7747 SUB 0.36fF $ **FLOATING
C8516 S.n7748 SUB 0.61fF $ **FLOATING
C8517 S.n7749 SUB 0.12fF $ **FLOATING
C8518 S.t60 SUB 0.02fF
C8519 S.n7750 SUB 0.14fF $ **FLOATING
C8520 S.n7752 SUB 0.31fF $ **FLOATING
C8521 S.n7753 SUB 0.23fF $ **FLOATING
C8522 S.n7754 SUB 0.66fF $ **FLOATING
C8523 S.n7755 SUB 0.95fF $ **FLOATING
C8524 S.n7756 SUB 0.23fF $ **FLOATING
C8525 S.n7757 SUB 0.21fF $ **FLOATING
C8526 S.n7758 SUB 0.20fF $ **FLOATING
C8527 S.n7759 SUB 0.06fF $ **FLOATING
C8528 S.n7760 SUB 0.09fF $ **FLOATING
C8529 S.n7761 SUB 0.10fF $ **FLOATING
C8530 S.n7762 SUB 1.99fF $ **FLOATING
C8531 S.t285 SUB 0.02fF
C8532 S.n7763 SUB 0.12fF $ **FLOATING
C8533 S.n7764 SUB 0.14fF $ **FLOATING
C8534 S.t1463 SUB 0.02fF
C8535 S.n7766 SUB 0.24fF $ **FLOATING
C8536 S.n7767 SUB 0.91fF $ **FLOATING
C8537 S.n7768 SUB 0.05fF $ **FLOATING
C8538 S.n7769 SUB 1.88fF $ **FLOATING
C8539 S.n7770 SUB 0.12fF $ **FLOATING
C8540 S.t273 SUB 0.02fF
C8541 S.n7771 SUB 0.14fF $ **FLOATING
C8542 S.t1974 SUB 0.02fF
C8543 S.n7773 SUB 1.22fF $ **FLOATING
C8544 S.n7774 SUB 0.61fF $ **FLOATING
C8545 S.n7775 SUB 0.35fF $ **FLOATING
C8546 S.n7776 SUB 0.63fF $ **FLOATING
C8547 S.n7777 SUB 1.15fF $ **FLOATING
C8548 S.n7778 SUB 3.03fF $ **FLOATING
C8549 S.n7779 SUB 0.59fF $ **FLOATING
C8550 S.n7780 SUB 0.02fF $ **FLOATING
C8551 S.n7781 SUB 0.97fF $ **FLOATING
C8552 S.t156 SUB 21.38fF
C8553 S.n7782 SUB 20.25fF $ **FLOATING
C8554 S.n7784 SUB 0.38fF $ **FLOATING
C8555 S.n7785 SUB 0.23fF $ **FLOATING
C8556 S.n7786 SUB 2.90fF $ **FLOATING
C8557 S.n7787 SUB 2.46fF $ **FLOATING
C8558 S.n7788 SUB 1.96fF $ **FLOATING
C8559 S.n7789 SUB 3.94fF $ **FLOATING
C8560 S.n7790 SUB 0.25fF $ **FLOATING
C8561 S.n7791 SUB 0.01fF $ **FLOATING
C8562 S.t1677 SUB 0.02fF
C8563 S.n7792 SUB 0.25fF $ **FLOATING
C8564 S.t1439 SUB 0.02fF
C8565 S.n7793 SUB 0.95fF $ **FLOATING
C8566 S.n7794 SUB 0.70fF $ **FLOATING
C8567 S.n7795 SUB 0.78fF $ **FLOATING
C8568 S.n7796 SUB 1.93fF $ **FLOATING
C8569 S.n7797 SUB 1.88fF $ **FLOATING
C8570 S.n7798 SUB 0.12fF $ **FLOATING
C8571 S.t802 SUB 0.02fF
C8572 S.n7799 SUB 0.14fF $ **FLOATING
C8573 S.t1119 SUB 0.02fF
C8574 S.n7801 SUB 0.24fF $ **FLOATING
C8575 S.n7802 SUB 0.36fF $ **FLOATING
C8576 S.n7803 SUB 0.61fF $ **FLOATING
C8577 S.n7804 SUB 1.52fF $ **FLOATING
C8578 S.n7805 SUB 2.99fF $ **FLOATING
C8579 S.t576 SUB 0.02fF
C8580 S.n7806 SUB 0.24fF $ **FLOATING
C8581 S.n7807 SUB 0.91fF $ **FLOATING
C8582 S.n7808 SUB 0.05fF $ **FLOATING
C8583 S.t1492 SUB 0.02fF
C8584 S.n7809 SUB 0.12fF $ **FLOATING
C8585 S.n7810 SUB 0.14fF $ **FLOATING
C8586 S.n7812 SUB 1.89fF $ **FLOATING
C8587 S.n7813 SUB 1.88fF $ **FLOATING
C8588 S.t239 SUB 0.02fF
C8589 S.n7814 SUB 0.24fF $ **FLOATING
C8590 S.n7815 SUB 0.36fF $ **FLOATING
C8591 S.n7816 SUB 0.61fF $ **FLOATING
C8592 S.n7817 SUB 0.12fF $ **FLOATING
C8593 S.t2452 SUB 0.02fF
C8594 S.n7818 SUB 0.14fF $ **FLOATING
C8595 S.n7820 SUB 1.16fF $ **FLOATING
C8596 S.n7821 SUB 0.22fF $ **FLOATING
C8597 S.n7822 SUB 0.25fF $ **FLOATING
C8598 S.n7823 SUB 0.09fF $ **FLOATING
C8599 S.n7824 SUB 1.88fF $ **FLOATING
C8600 S.t2221 SUB 0.02fF
C8601 S.n7825 SUB 0.24fF $ **FLOATING
C8602 S.n7826 SUB 0.91fF $ **FLOATING
C8603 S.n7827 SUB 0.05fF $ **FLOATING
C8604 S.t629 SUB 0.02fF
C8605 S.n7828 SUB 0.12fF $ **FLOATING
C8606 S.n7829 SUB 0.14fF $ **FLOATING
C8607 S.n7831 SUB 0.78fF $ **FLOATING
C8608 S.n7832 SUB 1.94fF $ **FLOATING
C8609 S.n7833 SUB 1.88fF $ **FLOATING
C8610 S.n7834 SUB 0.12fF $ **FLOATING
C8611 S.t1584 SUB 0.02fF
C8612 S.n7835 SUB 0.14fF $ **FLOATING
C8613 S.t1906 SUB 0.02fF
C8614 S.n7837 SUB 0.24fF $ **FLOATING
C8615 S.n7838 SUB 0.36fF $ **FLOATING
C8616 S.n7839 SUB 0.61fF $ **FLOATING
C8617 S.n7840 SUB 1.84fF $ **FLOATING
C8618 S.n7841 SUB 2.99fF $ **FLOATING
C8619 S.t1360 SUB 0.02fF
C8620 S.n7842 SUB 0.24fF $ **FLOATING
C8621 S.n7843 SUB 0.91fF $ **FLOATING
C8622 S.n7844 SUB 0.05fF $ **FLOATING
C8623 S.t2381 SUB 0.02fF
C8624 S.n7845 SUB 0.12fF $ **FLOATING
C8625 S.n7846 SUB 0.14fF $ **FLOATING
C8626 S.n7848 SUB 1.89fF $ **FLOATING
C8627 S.n7849 SUB 1.75fF $ **FLOATING
C8628 S.t1047 SUB 0.02fF
C8629 S.n7850 SUB 0.24fF $ **FLOATING
C8630 S.n7851 SUB 0.36fF $ **FLOATING
C8631 S.n7852 SUB 0.61fF $ **FLOATING
C8632 S.n7853 SUB 0.12fF $ **FLOATING
C8633 S.t717 SUB 0.02fF
C8634 S.n7854 SUB 0.14fF $ **FLOATING
C8635 S.n7856 SUB 1.16fF $ **FLOATING
C8636 S.n7857 SUB 0.22fF $ **FLOATING
C8637 S.n7858 SUB 0.25fF $ **FLOATING
C8638 S.n7859 SUB 0.09fF $ **FLOATING
C8639 S.n7860 SUB 2.44fF $ **FLOATING
C8640 S.t487 SUB 0.02fF
C8641 S.n7861 SUB 0.24fF $ **FLOATING
C8642 S.n7862 SUB 0.91fF $ **FLOATING
C8643 S.n7863 SUB 0.05fF $ **FLOATING
C8644 S.t1527 SUB 0.02fF
C8645 S.n7864 SUB 0.12fF $ **FLOATING
C8646 S.n7865 SUB 0.14fF $ **FLOATING
C8647 S.n7867 SUB 1.88fF $ **FLOATING
C8648 S.n7868 SUB 0.48fF $ **FLOATING
C8649 S.n7869 SUB 0.09fF $ **FLOATING
C8650 S.n7870 SUB 0.33fF $ **FLOATING
C8651 S.n7871 SUB 0.30fF $ **FLOATING
C8652 S.n7872 SUB 0.77fF $ **FLOATING
C8653 S.n7873 SUB 0.59fF $ **FLOATING
C8654 S.t157 SUB 0.02fF
C8655 S.n7874 SUB 0.24fF $ **FLOATING
C8656 S.n7875 SUB 0.36fF $ **FLOATING
C8657 S.n7876 SUB 0.61fF $ **FLOATING
C8658 S.n7877 SUB 0.12fF $ **FLOATING
C8659 S.t2372 SUB 0.02fF
C8660 S.n7878 SUB 0.14fF $ **FLOATING
C8661 S.n7880 SUB 2.61fF $ **FLOATING
C8662 S.n7881 SUB 2.16fF $ **FLOATING
C8663 S.t2132 SUB 0.02fF
C8664 S.n7882 SUB 0.24fF $ **FLOATING
C8665 S.n7883 SUB 0.91fF $ **FLOATING
C8666 S.n7884 SUB 0.05fF $ **FLOATING
C8667 S.t666 SUB 0.02fF
C8668 S.n7885 SUB 0.12fF $ **FLOATING
C8669 S.n7886 SUB 0.14fF $ **FLOATING
C8670 S.n7888 SUB 0.78fF $ **FLOATING
C8671 S.n7889 SUB 2.30fF $ **FLOATING
C8672 S.n7890 SUB 1.88fF $ **FLOATING
C8673 S.n7891 SUB 0.12fF $ **FLOATING
C8674 S.t1515 SUB 0.02fF
C8675 S.n7892 SUB 0.14fF $ **FLOATING
C8676 S.t1820 SUB 0.02fF
C8677 S.n7894 SUB 0.24fF $ **FLOATING
C8678 S.n7895 SUB 0.36fF $ **FLOATING
C8679 S.n7896 SUB 0.61fF $ **FLOATING
C8680 S.n7897 SUB 1.39fF $ **FLOATING
C8681 S.n7898 SUB 0.71fF $ **FLOATING
C8682 S.n7899 SUB 1.14fF $ **FLOATING
C8683 S.n7900 SUB 0.35fF $ **FLOATING
C8684 S.n7901 SUB 2.03fF $ **FLOATING
C8685 S.t1267 SUB 0.02fF
C8686 S.n7902 SUB 0.24fF $ **FLOATING
C8687 S.n7903 SUB 0.91fF $ **FLOATING
C8688 S.n7904 SUB 0.05fF $ **FLOATING
C8689 S.t2320 SUB 0.02fF
C8690 S.n7905 SUB 0.12fF $ **FLOATING
C8691 S.n7906 SUB 0.14fF $ **FLOATING
C8692 S.n7908 SUB 1.89fF $ **FLOATING
C8693 S.n7909 SUB 1.88fF $ **FLOATING
C8694 S.t954 SUB 0.02fF
C8695 S.n7910 SUB 0.24fF $ **FLOATING
C8696 S.n7911 SUB 0.36fF $ **FLOATING
C8697 S.n7912 SUB 0.61fF $ **FLOATING
C8698 S.n7913 SUB 0.12fF $ **FLOATING
C8699 S.t756 SUB 0.02fF
C8700 S.n7914 SUB 0.14fF $ **FLOATING
C8701 S.n7916 SUB 1.16fF $ **FLOATING
C8702 S.n7917 SUB 0.22fF $ **FLOATING
C8703 S.n7918 SUB 0.25fF $ **FLOATING
C8704 S.n7919 SUB 0.09fF $ **FLOATING
C8705 S.n7920 SUB 1.88fF $ **FLOATING
C8706 S.t384 SUB 0.02fF
C8707 S.n7921 SUB 0.24fF $ **FLOATING
C8708 S.n7922 SUB 0.91fF $ **FLOATING
C8709 S.n7923 SUB 0.05fF $ **FLOATING
C8710 S.t1462 SUB 0.02fF
C8711 S.n7924 SUB 0.12fF $ **FLOATING
C8712 S.n7925 SUB 0.14fF $ **FLOATING
C8713 S.n7927 SUB 20.78fF $ **FLOATING
C8714 S.n7928 SUB 1.88fF $ **FLOATING
C8715 S.n7929 SUB 2.67fF $ **FLOATING
C8716 S.t312 SUB 0.02fF
C8717 S.n7930 SUB 0.24fF $ **FLOATING
C8718 S.n7931 SUB 0.36fF $ **FLOATING
C8719 S.n7932 SUB 0.61fF $ **FLOATING
C8720 S.n7933 SUB 0.12fF $ **FLOATING
C8721 S.t1078 SUB 0.02fF
C8722 S.n7934 SUB 0.14fF $ **FLOATING
C8723 S.n7936 SUB 2.80fF $ **FLOATING
C8724 S.n7937 SUB 2.30fF $ **FLOATING
C8725 S.t1731 SUB 0.02fF
C8726 S.n7938 SUB 0.12fF $ **FLOATING
C8727 S.n7939 SUB 0.14fF $ **FLOATING
C8728 S.t1265 SUB 0.02fF
C8729 S.n7941 SUB 0.24fF $ **FLOATING
C8730 S.n7942 SUB 0.91fF $ **FLOATING
C8731 S.n7943 SUB 0.05fF $ **FLOATING
C8732 S.n7944 SUB 1.88fF $ **FLOATING
C8733 S.n7945 SUB 2.67fF $ **FLOATING
C8734 S.t1975 SUB 0.02fF
C8735 S.n7946 SUB 0.24fF $ **FLOATING
C8736 S.n7947 SUB 0.36fF $ **FLOATING
C8737 S.n7948 SUB 0.61fF $ **FLOATING
C8738 S.n7949 SUB 0.12fF $ **FLOATING
C8739 S.t203 SUB 0.02fF
C8740 S.n7950 SUB 0.14fF $ **FLOATING
C8741 S.n7952 SUB 2.80fF $ **FLOATING
C8742 S.n7953 SUB 2.30fF $ **FLOATING
C8743 S.t857 SUB 0.02fF
C8744 S.n7954 SUB 0.12fF $ **FLOATING
C8745 S.n7955 SUB 0.14fF $ **FLOATING
C8746 S.t382 SUB 0.02fF
C8747 S.n7957 SUB 0.24fF $ **FLOATING
C8748 S.n7958 SUB 0.91fF $ **FLOATING
C8749 S.n7959 SUB 0.05fF $ **FLOATING
C8750 S.n7960 SUB 1.88fF $ **FLOATING
C8751 S.n7961 SUB 2.67fF $ **FLOATING
C8752 S.t1120 SUB 0.02fF
C8753 S.n7962 SUB 0.24fF $ **FLOATING
C8754 S.n7963 SUB 0.36fF $ **FLOATING
C8755 S.n7964 SUB 0.61fF $ **FLOATING
C8756 S.n7965 SUB 0.12fF $ **FLOATING
C8757 S.t1870 SUB 0.02fF
C8758 S.n7966 SUB 0.14fF $ **FLOATING
C8759 S.n7968 SUB 2.80fF $ **FLOATING
C8760 S.n7969 SUB 2.30fF $ **FLOATING
C8761 S.t2501 SUB 0.02fF
C8762 S.n7970 SUB 0.12fF $ **FLOATING
C8763 S.n7971 SUB 0.14fF $ **FLOATING
C8764 S.t2033 SUB 0.02fF
C8765 S.n7973 SUB 0.24fF $ **FLOATING
C8766 S.n7974 SUB 0.91fF $ **FLOATING
C8767 S.n7975 SUB 0.05fF $ **FLOATING
C8768 S.n7976 SUB 1.88fF $ **FLOATING
C8769 S.n7977 SUB 2.67fF $ **FLOATING
C8770 S.t243 SUB 0.02fF
C8771 S.n7978 SUB 0.24fF $ **FLOATING
C8772 S.n7979 SUB 0.36fF $ **FLOATING
C8773 S.n7980 SUB 0.61fF $ **FLOATING
C8774 S.n7981 SUB 0.12fF $ **FLOATING
C8775 S.t1001 SUB 0.02fF
C8776 S.n7982 SUB 0.14fF $ **FLOATING
C8777 S.n7984 SUB 2.80fF $ **FLOATING
C8778 S.n7985 SUB 2.30fF $ **FLOATING
C8779 S.t1785 SUB 0.02fF
C8780 S.n7986 SUB 0.12fF $ **FLOATING
C8781 S.n7987 SUB 0.14fF $ **FLOATING
C8782 S.t1177 SUB 0.02fF
C8783 S.n7989 SUB 0.24fF $ **FLOATING
C8784 S.n7990 SUB 0.91fF $ **FLOATING
C8785 S.n7991 SUB 0.05fF $ **FLOATING
C8786 S.n7992 SUB 1.88fF $ **FLOATING
C8787 S.n7993 SUB 2.67fF $ **FLOATING
C8788 S.t1909 SUB 0.02fF
C8789 S.n7994 SUB 0.24fF $ **FLOATING
C8790 S.n7995 SUB 0.36fF $ **FLOATING
C8791 S.n7996 SUB 0.61fF $ **FLOATING
C8792 S.n7997 SUB 0.12fF $ **FLOATING
C8793 S.t96 SUB 0.02fF
C8794 S.n7998 SUB 0.14fF $ **FLOATING
C8795 S.n8000 SUB 2.80fF $ **FLOATING
C8796 S.n8001 SUB 2.30fF $ **FLOATING
C8797 S.t916 SUB 0.02fF
C8798 S.n8002 SUB 0.12fF $ **FLOATING
C8799 S.n8003 SUB 0.14fF $ **FLOATING
C8800 S.t300 SUB 0.02fF
C8801 S.n8005 SUB 0.24fF $ **FLOATING
C8802 S.n8006 SUB 0.91fF $ **FLOATING
C8803 S.n8007 SUB 0.05fF $ **FLOATING
C8804 S.n8008 SUB 1.88fF $ **FLOATING
C8805 S.n8009 SUB 2.67fF $ **FLOATING
C8806 S.t1049 SUB 0.02fF
C8807 S.n8010 SUB 0.24fF $ **FLOATING
C8808 S.n8011 SUB 0.36fF $ **FLOATING
C8809 S.n8012 SUB 0.61fF $ **FLOATING
C8810 S.n8013 SUB 0.12fF $ **FLOATING
C8811 S.t1772 SUB 0.02fF
C8812 S.n8014 SUB 0.14fF $ **FLOATING
C8813 S.n8016 SUB 2.80fF $ **FLOATING
C8814 S.n8017 SUB 2.30fF $ **FLOATING
C8815 S.t2557 SUB 0.02fF
C8816 S.n8018 SUB 0.12fF $ **FLOATING
C8817 S.n8019 SUB 0.14fF $ **FLOATING
C8818 S.t1964 SUB 0.02fF
C8819 S.n8021 SUB 0.24fF $ **FLOATING
C8820 S.n8022 SUB 0.91fF $ **FLOATING
C8821 S.n8023 SUB 0.05fF $ **FLOATING
C8822 S.n8024 SUB 1.88fF $ **FLOATING
C8823 S.n8025 SUB 2.68fF $ **FLOATING
C8824 S.t159 SUB 0.02fF
C8825 S.n8026 SUB 0.24fF $ **FLOATING
C8826 S.n8027 SUB 0.36fF $ **FLOATING
C8827 S.n8028 SUB 0.61fF $ **FLOATING
C8828 S.n8029 SUB 0.12fF $ **FLOATING
C8829 S.t900 SUB 0.02fF
C8830 S.n8030 SUB 0.14fF $ **FLOATING
C8831 S.n8032 SUB 5.17fF $ **FLOATING
C8832 S.t1684 SUB 0.02fF
C8833 S.n8033 SUB 0.12fF $ **FLOATING
C8834 S.n8034 SUB 0.14fF $ **FLOATING
C8835 S.t1109 SUB 0.02fF
C8836 S.n8036 SUB 0.24fF $ **FLOATING
C8837 S.n8037 SUB 0.91fF $ **FLOATING
C8838 S.n8038 SUB 0.05fF $ **FLOATING
C8839 S.n8039 SUB 2.73fF $ **FLOATING
C8840 S.n8040 SUB 1.59fF $ **FLOATING
C8841 S.n8041 SUB 0.12fF $ **FLOATING
C8842 S.t1907 SUB 0.02fF
C8843 S.n8042 SUB 0.14fF $ **FLOATING
C8844 S.t725 SUB 0.02fF
C8845 S.n8044 SUB 0.24fF $ **FLOATING
C8846 S.n8045 SUB 0.36fF $ **FLOATING
C8847 S.n8046 SUB 0.61fF $ **FLOATING
C8848 S.n8047 SUB 0.07fF $ **FLOATING
C8849 S.n8048 SUB 0.01fF $ **FLOATING
C8850 S.n8049 SUB 0.24fF $ **FLOATING
C8851 S.n8050 SUB 1.16fF $ **FLOATING
C8852 S.n8051 SUB 1.35fF $ **FLOATING
C8853 S.n8052 SUB 2.30fF $ **FLOATING
C8854 S.t100 SUB 0.02fF
C8855 S.n8053 SUB 0.12fF $ **FLOATING
C8856 S.n8054 SUB 0.14fF $ **FLOATING
C8857 S.t1085 SUB 0.02fF
C8858 S.n8056 SUB 0.24fF $ **FLOATING
C8859 S.n8057 SUB 0.91fF $ **FLOATING
C8860 S.n8058 SUB 0.05fF $ **FLOATING
C8861 S.t22 SUB 48.31fF
C8862 S.t602 SUB 0.02fF
C8863 S.n8059 SUB 0.12fF $ **FLOATING
C8864 S.n8060 SUB 0.14fF $ **FLOATING
C8865 S.t481 SUB 0.02fF
C8866 S.n8062 SUB 0.24fF $ **FLOATING
C8867 S.n8063 SUB 0.91fF $ **FLOATING
C8868 S.n8064 SUB 0.05fF $ **FLOATING
C8869 S.t2043 SUB 0.02fF
C8870 S.n8065 SUB 0.24fF $ **FLOATING
C8871 S.n8066 SUB 0.36fF $ **FLOATING
C8872 S.n8067 SUB 0.61fF $ **FLOATING
C8873 S.n8068 SUB 0.32fF $ **FLOATING
C8874 S.n8069 SUB 1.09fF $ **FLOATING
C8875 S.n8070 SUB 0.15fF $ **FLOATING
C8876 S.n8071 SUB 2.10fF $ **FLOATING
C8877 S.n8072 SUB 2.94fF $ **FLOATING
C8878 S.n8073 SUB 1.88fF $ **FLOATING
C8879 S.n8074 SUB 0.12fF $ **FLOATING
C8880 S.t1623 SUB 0.02fF
C8881 S.n8075 SUB 0.14fF $ **FLOATING
C8882 S.t2205 SUB 0.02fF
C8883 S.n8077 SUB 0.24fF $ **FLOATING
C8884 S.n8078 SUB 0.36fF $ **FLOATING
C8885 S.n8079 SUB 0.61fF $ **FLOATING
C8886 S.n8080 SUB 0.92fF $ **FLOATING
C8887 S.n8081 SUB 0.32fF $ **FLOATING
C8888 S.n8082 SUB 0.92fF $ **FLOATING
C8889 S.n8083 SUB 1.09fF $ **FLOATING
C8890 S.n8084 SUB 0.15fF $ **FLOATING
C8891 S.n8085 SUB 4.96fF $ **FLOATING
C8892 S.t1868 SUB 0.02fF
C8893 S.n8086 SUB 0.12fF $ **FLOATING
C8894 S.n8087 SUB 0.14fF $ **FLOATING
C8895 S.t2094 SUB 0.02fF
C8896 S.n8089 SUB 0.24fF $ **FLOATING
C8897 S.n8090 SUB 0.91fF $ **FLOATING
C8898 S.n8091 SUB 0.05fF $ **FLOATING
C8899 S.n8092 SUB 1.88fF $ **FLOATING
C8900 S.n8093 SUB 2.67fF $ **FLOATING
C8901 S.t1346 SUB 0.02fF
C8902 S.n8094 SUB 0.24fF $ **FLOATING
C8903 S.n8095 SUB 0.36fF $ **FLOATING
C8904 S.n8096 SUB 0.61fF $ **FLOATING
C8905 S.n8097 SUB 0.12fF $ **FLOATING
C8906 S.t758 SUB 0.02fF
C8907 S.n8098 SUB 0.14fF $ **FLOATING
C8908 S.n8100 SUB 1.88fF $ **FLOATING
C8909 S.n8101 SUB 2.67fF $ **FLOATING
C8910 S.t1187 SUB 0.02fF
C8911 S.n8102 SUB 0.24fF $ **FLOATING
C8912 S.n8103 SUB 0.36fF $ **FLOATING
C8913 S.n8104 SUB 0.61fF $ **FLOATING
C8914 S.t2129 SUB 0.02fF
C8915 S.n8105 SUB 0.24fF $ **FLOATING
C8916 S.n8106 SUB 0.91fF $ **FLOATING
C8917 S.n8107 SUB 0.05fF $ **FLOATING
C8918 S.t23 SUB 0.02fF
C8919 S.n8108 SUB 0.12fF $ **FLOATING
C8920 S.n8109 SUB 0.14fF $ **FLOATING
C8921 S.n8111 SUB 0.12fF $ **FLOATING
C8922 S.t1936 SUB 0.02fF
C8923 S.n8112 SUB 0.14fF $ **FLOATING
C8924 S.n8114 SUB 2.30fF $ **FLOATING
C8925 S.n8115 SUB 2.94fF $ **FLOATING
C8926 S.n8116 SUB 5.16fF $ **FLOATING
C8927 S.t1000 SUB 0.02fF
C8928 S.n8117 SUB 0.12fF $ **FLOATING
C8929 S.n8118 SUB 0.14fF $ **FLOATING
C8930 S.t1229 SUB 0.02fF
C8931 S.n8120 SUB 0.24fF $ **FLOATING
C8932 S.n8121 SUB 0.91fF $ **FLOATING
C8933 S.n8122 SUB 0.05fF $ **FLOATING
C8934 S.n8123 SUB 1.88fF $ **FLOATING
C8935 S.n8124 SUB 2.67fF $ **FLOATING
C8936 S.t469 SUB 0.02fF
C8937 S.n8125 SUB 0.24fF $ **FLOATING
C8938 S.n8126 SUB 0.36fF $ **FLOATING
C8939 S.n8127 SUB 0.61fF $ **FLOATING
C8940 S.n8128 SUB 0.12fF $ **FLOATING
C8941 S.t2412 SUB 0.02fF
C8942 S.n8129 SUB 0.14fF $ **FLOATING
C8943 S.n8131 SUB 5.17fF $ **FLOATING
C8944 S.t94 SUB 0.02fF
C8945 S.n8132 SUB 0.12fF $ **FLOATING
C8946 S.n8133 SUB 0.14fF $ **FLOATING
C8947 S.t347 SUB 0.02fF
C8948 S.n8135 SUB 0.24fF $ **FLOATING
C8949 S.n8136 SUB 0.91fF $ **FLOATING
C8950 S.n8137 SUB 0.05fF $ **FLOATING
C8951 S.n8138 SUB 1.88fF $ **FLOATING
C8952 S.n8139 SUB 2.67fF $ **FLOATING
C8953 S.t2118 SUB 0.02fF
C8954 S.n8140 SUB 0.24fF $ **FLOATING
C8955 S.n8141 SUB 0.36fF $ **FLOATING
C8956 S.n8142 SUB 0.61fF $ **FLOATING
C8957 S.n8143 SUB 0.12fF $ **FLOATING
C8958 S.t1548 SUB 0.02fF
C8959 S.n8144 SUB 0.14fF $ **FLOATING
C8960 S.n8146 SUB 5.17fF $ **FLOATING
C8961 S.t1771 SUB 0.02fF
C8962 S.n8147 SUB 0.12fF $ **FLOATING
C8963 S.n8148 SUB 0.14fF $ **FLOATING
C8964 S.t2005 SUB 0.02fF
C8965 S.n8150 SUB 0.24fF $ **FLOATING
C8966 S.n8151 SUB 0.91fF $ **FLOATING
C8967 S.n8152 SUB 0.05fF $ **FLOATING
C8968 S.n8153 SUB 1.88fF $ **FLOATING
C8969 S.n8154 SUB 2.67fF $ **FLOATING
C8970 S.t1392 SUB 0.02fF
C8971 S.n8155 SUB 0.24fF $ **FLOATING
C8972 S.n8156 SUB 0.36fF $ **FLOATING
C8973 S.n8157 SUB 0.61fF $ **FLOATING
C8974 S.n8158 SUB 0.12fF $ **FLOATING
C8975 S.t808 SUB 0.02fF
C8976 S.n8159 SUB 0.14fF $ **FLOATING
C8977 S.n8161 SUB 5.17fF $ **FLOATING
C8978 S.t897 SUB 0.02fF
C8979 S.n8162 SUB 0.12fF $ **FLOATING
C8980 S.n8163 SUB 0.14fF $ **FLOATING
C8981 S.t1286 SUB 0.02fF
C8982 S.n8165 SUB 0.24fF $ **FLOATING
C8983 S.n8166 SUB 0.91fF $ **FLOATING
C8984 S.n8167 SUB 0.05fF $ **FLOATING
C8985 S.n8168 SUB 1.88fF $ **FLOATING
C8986 S.n8169 SUB 2.67fF $ **FLOATING
C8987 S.t520 SUB 0.02fF
C8988 S.n8170 SUB 0.24fF $ **FLOATING
C8989 S.n8171 SUB 0.36fF $ **FLOATING
C8990 S.n8172 SUB 0.61fF $ **FLOATING
C8991 S.n8173 SUB 0.12fF $ **FLOATING
C8992 S.t2458 SUB 0.02fF
C8993 S.n8174 SUB 0.14fF $ **FLOATING
C8994 S.n8176 SUB 5.17fF $ **FLOATING
C8995 S.t2539 SUB 0.02fF
C8996 S.n8177 SUB 0.12fF $ **FLOATING
C8997 S.n8178 SUB 0.14fF $ **FLOATING
C8998 S.t398 SUB 0.02fF
C8999 S.n8180 SUB 0.24fF $ **FLOATING
C9000 S.n8181 SUB 0.91fF $ **FLOATING
C9001 S.n8182 SUB 0.05fF $ **FLOATING
C9002 S.n8183 SUB 1.88fF $ **FLOATING
C9003 S.n8184 SUB 2.67fF $ **FLOATING
C9004 S.t2165 SUB 0.02fF
C9005 S.n8185 SUB 0.24fF $ **FLOATING
C9006 S.n8186 SUB 0.36fF $ **FLOATING
C9007 S.n8187 SUB 0.61fF $ **FLOATING
C9008 S.n8188 SUB 0.12fF $ **FLOATING
C9009 S.t1590 SUB 0.02fF
C9010 S.n8189 SUB 0.14fF $ **FLOATING
C9011 S.n8191 SUB 5.17fF $ **FLOATING
C9012 S.t1668 SUB 0.02fF
C9013 S.n8192 SUB 0.12fF $ **FLOATING
C9014 S.n8193 SUB 0.14fF $ **FLOATING
C9015 S.t2050 SUB 0.02fF
C9016 S.n8195 SUB 0.24fF $ **FLOATING
C9017 S.n8196 SUB 0.91fF $ **FLOATING
C9018 S.n8197 SUB 0.05fF $ **FLOATING
C9019 S.n8198 SUB 1.88fF $ **FLOATING
C9020 S.n8199 SUB 2.67fF $ **FLOATING
C9021 S.t1300 SUB 0.02fF
C9022 S.n8200 SUB 0.24fF $ **FLOATING
C9023 S.n8201 SUB 0.36fF $ **FLOATING
C9024 S.n8202 SUB 0.61fF $ **FLOATING
C9025 S.n8203 SUB 0.12fF $ **FLOATING
C9026 S.t726 SUB 0.02fF
C9027 S.n8204 SUB 0.14fF $ **FLOATING
C9028 S.n8206 SUB 4.90fF $ **FLOATING
C9029 S.t794 SUB 0.02fF
C9030 S.n8207 SUB 0.12fF $ **FLOATING
C9031 S.n8208 SUB 0.14fF $ **FLOATING
C9032 S.t1192 SUB 0.02fF
C9033 S.n8210 SUB 0.24fF $ **FLOATING
C9034 S.n8211 SUB 0.91fF $ **FLOATING
C9035 S.n8212 SUB 0.05fF $ **FLOATING
C9036 S.n8213 SUB 1.88fF $ **FLOATING
C9037 S.n8214 SUB 2.67fF $ **FLOATING
C9038 S.t782 SUB 0.02fF
C9039 S.n8215 SUB 0.24fF $ **FLOATING
C9040 S.n8216 SUB 0.36fF $ **FLOATING
C9041 S.n8217 SUB 0.61fF $ **FLOATING
C9042 S.n8218 SUB 0.12fF $ **FLOATING
C9043 S.t2042 SUB 0.02fF
C9044 S.n8219 SUB 0.14fF $ **FLOATING
C9045 S.n8221 SUB 5.44fF $ **FLOATING
C9046 S.t2442 SUB 0.02fF
C9047 S.n8222 SUB 0.12fF $ **FLOATING
C9048 S.n8223 SUB 0.14fF $ **FLOATING
C9049 S.t2111 SUB 0.02fF
C9050 S.n8225 SUB 0.24fF $ **FLOATING
C9051 S.n8226 SUB 0.91fF $ **FLOATING
C9052 S.n8227 SUB 0.05fF $ **FLOATING
C9053 S.t59 SUB 47.92fF
C9054 S.t1262 SUB 0.02fF
C9055 S.n8228 SUB 1.19fF $ **FLOATING
C9056 S.n8229 SUB 0.05fF $ **FLOATING
C9057 S.t1319 SUB 0.02fF
C9058 S.n8230 SUB 0.01fF $ **FLOATING
C9059 S.n8231 SUB 0.26fF $ **FLOATING
C9060 S.n8233 SUB 1.50fF $ **FLOATING
C9061 S.n8234 SUB 1.30fF $ **FLOATING
C9062 S.n8235 SUB 0.28fF $ **FLOATING
C9063 S.n8236 SUB 0.24fF $ **FLOATING
C9064 S.n8237 SUB 4.39fF $ **FLOATING
C9065 S.n8238 SUB 0.01fF $ **FLOATING
C9066 S.n8239 SUB 0.02fF $ **FLOATING
C9067 S.n8240 SUB 0.03fF $ **FLOATING
C9068 S.n8241 SUB 0.04fF $ **FLOATING
C9069 S.n8242 SUB 0.17fF $ **FLOATING
C9070 S.n8243 SUB 0.01fF $ **FLOATING
C9071 S.n8244 SUB 0.02fF $ **FLOATING
C9072 S.n8245 SUB 0.01fF $ **FLOATING
C9073 S.n8246 SUB 0.01fF $ **FLOATING
C9074 S.n8247 SUB 0.01fF $ **FLOATING
C9075 S.n8248 SUB 0.01fF $ **FLOATING
C9076 S.n8249 SUB 0.02fF $ **FLOATING
C9077 S.n8250 SUB 0.01fF $ **FLOATING
C9078 S.n8251 SUB 0.02fF $ **FLOATING
C9079 S.n8252 SUB 0.05fF $ **FLOATING
C9080 S.n8253 SUB 0.04fF $ **FLOATING
C9081 S.n8254 SUB 0.11fF $ **FLOATING
C9082 S.n8255 SUB 0.38fF $ **FLOATING
C9083 S.n8256 SUB 0.20fF $ **FLOATING
C9084 S.n8257 SUB 8.97fF $ **FLOATING
C9085 S.n8258 SUB 8.97fF $ **FLOATING
C9086 S.n8259 SUB 0.60fF $ **FLOATING
C9087 S.n8260 SUB 0.22fF $ **FLOATING
C9088 S.n8261 SUB 0.59fF $ **FLOATING
C9089 S.n8262 SUB 3.43fF $ **FLOATING
C9090 S.n8263 SUB 0.29fF $ **FLOATING
C9091 S.t84 SUB 21.38fF
C9092 S.n8264 SUB 21.67fF $ **FLOATING
C9093 S.n8265 SUB 0.77fF $ **FLOATING
C9094 S.n8266 SUB 0.28fF $ **FLOATING
C9095 S.n8267 SUB 4.00fF $ **FLOATING
C9096 S.n8268 SUB 1.35fF $ **FLOATING
C9097 S.t524 SUB 0.02fF
C9098 S.n8269 SUB 0.64fF $ **FLOATING
C9099 S.n8270 SUB 0.61fF $ **FLOATING
C9100 S.n8271 SUB 1.89fF $ **FLOATING
C9101 S.n8272 SUB 0.06fF $ **FLOATING
C9102 S.n8273 SUB 0.03fF $ **FLOATING
C9103 S.n8274 SUB 0.04fF $ **FLOATING
C9104 S.n8275 SUB 0.99fF $ **FLOATING
C9105 S.n8276 SUB 0.02fF $ **FLOATING
C9106 S.n8277 SUB 0.01fF $ **FLOATING
C9107 S.n8278 SUB 0.02fF $ **FLOATING
C9108 S.n8279 SUB 0.08fF $ **FLOATING
C9109 S.n8280 SUB 0.36fF $ **FLOATING
C9110 S.n8281 SUB 1.85fF $ **FLOATING
C9111 S.t1985 SUB 0.02fF
C9112 S.n8282 SUB 0.24fF $ **FLOATING
C9113 S.n8283 SUB 0.36fF $ **FLOATING
C9114 S.n8284 SUB 0.61fF $ **FLOATING
C9115 S.n8285 SUB 0.12fF $ **FLOATING
C9116 S.t1467 SUB 0.02fF
C9117 S.n8286 SUB 0.14fF $ **FLOATING
C9118 S.n8288 SUB 0.70fF $ **FLOATING
C9119 S.n8289 SUB 0.23fF $ **FLOATING
C9120 S.n8290 SUB 0.23fF $ **FLOATING
C9121 S.n8291 SUB 0.70fF $ **FLOATING
C9122 S.n8292 SUB 1.16fF $ **FLOATING
C9123 S.n8293 SUB 0.22fF $ **FLOATING
C9124 S.n8294 SUB 0.25fF $ **FLOATING
C9125 S.n8295 SUB 0.09fF $ **FLOATING
C9126 S.n8296 SUB 1.88fF $ **FLOATING
C9127 S.t297 SUB 0.02fF
C9128 S.n8297 SUB 0.24fF $ **FLOATING
C9129 S.n8298 SUB 0.91fF $ **FLOATING
C9130 S.n8299 SUB 0.05fF $ **FLOATING
C9131 S.t1628 SUB 0.02fF
C9132 S.n8300 SUB 0.12fF $ **FLOATING
C9133 S.n8301 SUB 0.14fF $ **FLOATING
C9134 S.n8303 SUB 0.25fF $ **FLOATING
C9135 S.n8304 SUB 0.09fF $ **FLOATING
C9136 S.n8305 SUB 0.21fF $ **FLOATING
C9137 S.n8306 SUB 0.92fF $ **FLOATING
C9138 S.n8307 SUB 0.44fF $ **FLOATING
C9139 S.n8308 SUB 1.88fF $ **FLOATING
C9140 S.n8309 SUB 0.12fF $ **FLOATING
C9141 S.t697 SUB 0.02fF
C9142 S.n8310 SUB 0.14fF $ **FLOATING
C9143 S.t1256 SUB 0.02fF
C9144 S.n8312 SUB 0.24fF $ **FLOATING
C9145 S.n8313 SUB 0.36fF $ **FLOATING
C9146 S.n8314 SUB 0.61fF $ **FLOATING
C9147 S.n8315 SUB 0.02fF $ **FLOATING
C9148 S.n8316 SUB 0.01fF $ **FLOATING
C9149 S.n8317 SUB 0.02fF $ **FLOATING
C9150 S.n8318 SUB 0.08fF $ **FLOATING
C9151 S.n8319 SUB 0.06fF $ **FLOATING
C9152 S.n8320 SUB 0.03fF $ **FLOATING
C9153 S.n8321 SUB 0.04fF $ **FLOATING
C9154 S.n8322 SUB 1.00fF $ **FLOATING
C9155 S.n8323 SUB 0.36fF $ **FLOATING
C9156 S.n8324 SUB 1.87fF $ **FLOATING
C9157 S.n8325 SUB 1.99fF $ **FLOATING
C9158 S.t2078 SUB 0.02fF
C9159 S.n8326 SUB 0.24fF $ **FLOATING
C9160 S.n8327 SUB 0.91fF $ **FLOATING
C9161 S.n8328 SUB 0.05fF $ **FLOATING
C9162 S.t761 SUB 0.02fF
C9163 S.n8329 SUB 0.12fF $ **FLOATING
C9164 S.n8330 SUB 0.14fF $ **FLOATING
C9165 S.n8332 SUB 1.89fF $ **FLOATING
C9166 S.n8333 SUB 0.07fF $ **FLOATING
C9167 S.n8334 SUB 0.04fF $ **FLOATING
C9168 S.n8335 SUB 0.05fF $ **FLOATING
C9169 S.n8336 SUB 0.87fF $ **FLOATING
C9170 S.n8337 SUB 0.01fF $ **FLOATING
C9171 S.n8338 SUB 0.01fF $ **FLOATING
C9172 S.n8339 SUB 0.01fF $ **FLOATING
C9173 S.n8340 SUB 0.07fF $ **FLOATING
C9174 S.n8341 SUB 0.68fF $ **FLOATING
C9175 S.n8342 SUB 0.72fF $ **FLOATING
C9176 S.t374 SUB 0.02fF
C9177 S.n8343 SUB 0.24fF $ **FLOATING
C9178 S.n8344 SUB 0.36fF $ **FLOATING
C9179 S.n8345 SUB 0.61fF $ **FLOATING
C9180 S.n8346 SUB 0.12fF $ **FLOATING
C9181 S.t2356 SUB 0.02fF
C9182 S.n8347 SUB 0.14fF $ **FLOATING
C9183 S.n8349 SUB 0.70fF $ **FLOATING
C9184 S.n8350 SUB 0.23fF $ **FLOATING
C9185 S.n8351 SUB 0.23fF $ **FLOATING
C9186 S.n8352 SUB 0.70fF $ **FLOATING
C9187 S.n8353 SUB 1.16fF $ **FLOATING
C9188 S.n8354 SUB 0.22fF $ **FLOATING
C9189 S.n8355 SUB 0.25fF $ **FLOATING
C9190 S.n8356 SUB 0.09fF $ **FLOATING
C9191 S.n8357 SUB 2.31fF $ **FLOATING
C9192 S.t1216 SUB 0.02fF
C9193 S.n8358 SUB 0.24fF $ **FLOATING
C9194 S.n8359 SUB 0.91fF $ **FLOATING
C9195 S.n8360 SUB 0.05fF $ **FLOATING
C9196 S.t2414 SUB 0.02fF
C9197 S.n8361 SUB 0.12fF $ **FLOATING
C9198 S.n8362 SUB 0.14fF $ **FLOATING
C9199 S.n8364 SUB 1.88fF $ **FLOATING
C9200 S.n8365 SUB 0.46fF $ **FLOATING
C9201 S.n8366 SUB 0.22fF $ **FLOATING
C9202 S.n8367 SUB 0.38fF $ **FLOATING
C9203 S.n8368 SUB 0.16fF $ **FLOATING
C9204 S.n8369 SUB 0.28fF $ **FLOATING
C9205 S.n8370 SUB 0.21fF $ **FLOATING
C9206 S.n8371 SUB 0.30fF $ **FLOATING
C9207 S.n8372 SUB 0.42fF $ **FLOATING
C9208 S.n8373 SUB 0.21fF $ **FLOATING
C9209 S.t2025 SUB 0.02fF
C9210 S.n8374 SUB 0.24fF $ **FLOATING
C9211 S.n8375 SUB 0.36fF $ **FLOATING
C9212 S.n8376 SUB 0.61fF $ **FLOATING
C9213 S.n8377 SUB 0.12fF $ **FLOATING
C9214 S.t1500 SUB 0.02fF
C9215 S.n8378 SUB 0.14fF $ **FLOATING
C9216 S.n8380 SUB 0.04fF $ **FLOATING
C9217 S.n8381 SUB 0.03fF $ **FLOATING
C9218 S.n8382 SUB 0.03fF $ **FLOATING
C9219 S.n8383 SUB 0.10fF $ **FLOATING
C9220 S.n8384 SUB 0.36fF $ **FLOATING
C9221 S.n8385 SUB 0.38fF $ **FLOATING
C9222 S.n8386 SUB 0.11fF $ **FLOATING
C9223 S.n8387 SUB 0.12fF $ **FLOATING
C9224 S.n8388 SUB 0.07fF $ **FLOATING
C9225 S.n8389 SUB 0.12fF $ **FLOATING
C9226 S.n8390 SUB 0.18fF $ **FLOATING
C9227 S.n8391 SUB 4.00fF $ **FLOATING
C9228 S.t335 SUB 0.02fF
C9229 S.n8392 SUB 0.24fF $ **FLOATING
C9230 S.n8393 SUB 0.91fF $ **FLOATING
C9231 S.n8394 SUB 0.05fF $ **FLOATING
C9232 S.t1550 SUB 0.02fF
C9233 S.n8395 SUB 0.12fF $ **FLOATING
C9234 S.n8396 SUB 0.14fF $ **FLOATING
C9235 S.n8398 SUB 0.25fF $ **FLOATING
C9236 S.n8399 SUB 0.09fF $ **FLOATING
C9237 S.n8400 SUB 0.21fF $ **FLOATING
C9238 S.n8401 SUB 1.28fF $ **FLOATING
C9239 S.n8402 SUB 0.53fF $ **FLOATING
C9240 S.n8403 SUB 1.88fF $ **FLOATING
C9241 S.n8404 SUB 0.12fF $ **FLOATING
C9242 S.t637 SUB 0.02fF
C9243 S.n8405 SUB 0.14fF $ **FLOATING
C9244 S.t1168 SUB 0.02fF
C9245 S.n8407 SUB 0.24fF $ **FLOATING
C9246 S.n8408 SUB 0.36fF $ **FLOATING
C9247 S.n8409 SUB 0.61fF $ **FLOATING
C9248 S.n8410 SUB 1.58fF $ **FLOATING
C9249 S.n8411 SUB 2.45fF $ **FLOATING
C9250 S.t1992 SUB 0.02fF
C9251 S.n8412 SUB 0.24fF $ **FLOATING
C9252 S.n8413 SUB 0.91fF $ **FLOATING
C9253 S.n8414 SUB 0.05fF $ **FLOATING
C9254 S.t688 SUB 0.02fF
C9255 S.n8415 SUB 0.12fF $ **FLOATING
C9256 S.n8416 SUB 0.14fF $ **FLOATING
C9257 S.n8418 SUB 1.89fF $ **FLOATING
C9258 S.n8419 SUB 0.06fF $ **FLOATING
C9259 S.n8420 SUB 0.03fF $ **FLOATING
C9260 S.n8421 SUB 0.04fF $ **FLOATING
C9261 S.n8422 SUB 0.99fF $ **FLOATING
C9262 S.n8423 SUB 0.02fF $ **FLOATING
C9263 S.n8424 SUB 0.01fF $ **FLOATING
C9264 S.n8425 SUB 0.02fF $ **FLOATING
C9265 S.n8426 SUB 0.08fF $ **FLOATING
C9266 S.n8427 SUB 0.36fF $ **FLOATING
C9267 S.n8428 SUB 1.85fF $ **FLOATING
C9268 S.t293 SUB 0.02fF
C9269 S.n8429 SUB 0.24fF $ **FLOATING
C9270 S.n8430 SUB 0.36fF $ **FLOATING
C9271 S.n8431 SUB 0.61fF $ **FLOATING
C9272 S.n8432 SUB 0.12fF $ **FLOATING
C9273 S.t2292 SUB 0.02fF
C9274 S.n8433 SUB 0.14fF $ **FLOATING
C9275 S.n8435 SUB 0.70fF $ **FLOATING
C9276 S.n8436 SUB 0.23fF $ **FLOATING
C9277 S.n8437 SUB 0.23fF $ **FLOATING
C9278 S.n8438 SUB 0.70fF $ **FLOATING
C9279 S.n8439 SUB 1.16fF $ **FLOATING
C9280 S.n8440 SUB 0.22fF $ **FLOATING
C9281 S.n8441 SUB 0.25fF $ **FLOATING
C9282 S.n8442 SUB 0.09fF $ **FLOATING
C9283 S.n8443 SUB 1.88fF $ **FLOATING
C9284 S.t1143 SUB 0.02fF
C9285 S.n8444 SUB 0.24fF $ **FLOATING
C9286 S.n8445 SUB 0.91fF $ **FLOATING
C9287 S.n8446 SUB 0.05fF $ **FLOATING
C9288 S.t2347 SUB 0.02fF
C9289 S.n8447 SUB 0.12fF $ **FLOATING
C9290 S.n8448 SUB 0.14fF $ **FLOATING
C9291 S.n8450 SUB 20.78fF $ **FLOATING
C9292 S.n8451 SUB 0.06fF $ **FLOATING
C9293 S.n8452 SUB 0.20fF $ **FLOATING
C9294 S.n8453 SUB 0.09fF $ **FLOATING
C9295 S.n8454 SUB 0.21fF $ **FLOATING
C9296 S.n8455 SUB 0.10fF $ **FLOATING
C9297 S.n8456 SUB 0.30fF $ **FLOATING
C9298 S.n8457 SUB 0.69fF $ **FLOATING
C9299 S.n8458 SUB 0.45fF $ **FLOATING
C9300 S.n8459 SUB 2.33fF $ **FLOATING
C9301 S.n8460 SUB 0.12fF $ **FLOATING
C9302 S.t2325 SUB 0.02fF
C9303 S.n8461 SUB 0.14fF $ **FLOATING
C9304 S.t325 SUB 0.02fF
C9305 S.n8463 SUB 0.24fF $ **FLOATING
C9306 S.n8464 SUB 0.36fF $ **FLOATING
C9307 S.n8465 SUB 0.61fF $ **FLOATING
C9308 S.n8466 SUB 1.90fF $ **FLOATING
C9309 S.n8467 SUB 0.17fF $ **FLOATING
C9310 S.n8468 SUB 0.76fF $ **FLOATING
C9311 S.n8469 SUB 0.32fF $ **FLOATING
C9312 S.n8470 SUB 0.25fF $ **FLOATING
C9313 S.n8471 SUB 0.30fF $ **FLOATING
C9314 S.n8472 SUB 0.47fF $ **FLOATING
C9315 S.n8473 SUB 0.16fF $ **FLOATING
C9316 S.n8474 SUB 1.93fF $ **FLOATING
C9317 S.t2503 SUB 0.02fF
C9318 S.n8475 SUB 0.12fF $ **FLOATING
C9319 S.n8476 SUB 0.14fF $ **FLOATING
C9320 S.t1173 SUB 0.02fF
C9321 S.n8478 SUB 0.24fF $ **FLOATING
C9322 S.n8479 SUB 0.91fF $ **FLOATING
C9323 S.n8480 SUB 0.05fF $ **FLOATING
C9324 S.n8481 SUB 1.88fF $ **FLOATING
C9325 S.n8482 SUB 0.12fF $ **FLOATING
C9326 S.t513 SUB 0.02fF
C9327 S.n8483 SUB 0.14fF $ **FLOATING
C9328 S.t1671 SUB 0.02fF
C9329 S.n8485 SUB 1.22fF $ **FLOATING
C9330 S.n8486 SUB 0.36fF $ **FLOATING
C9331 S.n8487 SUB 1.22fF $ **FLOATING
C9332 S.n8488 SUB 0.61fF $ **FLOATING
C9333 S.n8489 SUB 0.35fF $ **FLOATING
C9334 S.n8490 SUB 0.63fF $ **FLOATING
C9335 S.n8491 SUB 1.15fF $ **FLOATING
C9336 S.n8492 SUB 3.03fF $ **FLOATING
C9337 S.n8493 SUB 0.59fF $ **FLOATING
C9338 S.n8494 SUB 0.02fF $ **FLOATING
C9339 S.n8495 SUB 0.97fF $ **FLOATING
C9340 S.t188 SUB 21.38fF
C9341 S.n8496 SUB 20.25fF $ **FLOATING
C9342 S.n8498 SUB 0.38fF $ **FLOATING
C9343 S.n8499 SUB 0.23fF $ **FLOATING
C9344 S.n8500 SUB 2.79fF $ **FLOATING
C9345 S.n8501 SUB 2.46fF $ **FLOATING
C9346 S.n8502 SUB 4.00fF $ **FLOATING
C9347 S.n8503 SUB 0.25fF $ **FLOATING
C9348 S.n8504 SUB 0.01fF $ **FLOATING
C9349 S.t1427 SUB 0.02fF
C9350 S.n8505 SUB 0.25fF $ **FLOATING
C9351 S.t1147 SUB 0.02fF
C9352 S.n8506 SUB 0.95fF $ **FLOATING
C9353 S.n8507 SUB 0.70fF $ **FLOATING
C9354 S.n8508 SUB 1.89fF $ **FLOATING
C9355 S.n8509 SUB 1.88fF $ **FLOATING
C9356 S.t799 SUB 0.02fF
C9357 S.n8510 SUB 0.24fF $ **FLOATING
C9358 S.n8511 SUB 0.36fF $ **FLOATING
C9359 S.n8512 SUB 0.61fF $ **FLOATING
C9360 S.n8513 SUB 0.12fF $ **FLOATING
C9361 S.t560 SUB 0.02fF
C9362 S.n8514 SUB 0.14fF $ **FLOATING
C9363 S.n8516 SUB 1.16fF $ **FLOATING
C9364 S.n8517 SUB 0.22fF $ **FLOATING
C9365 S.n8518 SUB 0.25fF $ **FLOATING
C9366 S.n8519 SUB 0.09fF $ **FLOATING
C9367 S.n8520 SUB 1.88fF $ **FLOATING
C9368 S.t269 SUB 0.02fF
C9369 S.n8521 SUB 0.24fF $ **FLOATING
C9370 S.n8522 SUB 0.91fF $ **FLOATING
C9371 S.n8523 SUB 0.05fF $ **FLOATING
C9372 S.t1208 SUB 0.02fF
C9373 S.n8524 SUB 0.12fF $ **FLOATING
C9374 S.n8525 SUB 0.14fF $ **FLOATING
C9375 S.n8527 SUB 0.78fF $ **FLOATING
C9376 S.n8528 SUB 1.94fF $ **FLOATING
C9377 S.n8529 SUB 1.88fF $ **FLOATING
C9378 S.n8530 SUB 0.12fF $ **FLOATING
C9379 S.t2199 SUB 0.02fF
C9380 S.n8531 SUB 0.14fF $ **FLOATING
C9381 S.t2448 SUB 0.02fF
C9382 S.n8533 SUB 0.24fF $ **FLOATING
C9383 S.n8534 SUB 0.36fF $ **FLOATING
C9384 S.n8535 SUB 0.61fF $ **FLOATING
C9385 S.n8536 SUB 1.84fF $ **FLOATING
C9386 S.n8537 SUB 2.99fF $ **FLOATING
C9387 S.t1932 SUB 0.02fF
C9388 S.n8538 SUB 0.24fF $ **FLOATING
C9389 S.n8539 SUB 0.91fF $ **FLOATING
C9390 S.n8540 SUB 0.05fF $ **FLOATING
C9391 S.t330 SUB 0.02fF
C9392 S.n8541 SUB 0.12fF $ **FLOATING
C9393 S.n8542 SUB 0.14fF $ **FLOATING
C9394 S.n8544 SUB 1.89fF $ **FLOATING
C9395 S.n8545 SUB 1.75fF $ **FLOATING
C9396 S.t1580 SUB 0.02fF
C9397 S.n8546 SUB 0.24fF $ **FLOATING
C9398 S.n8547 SUB 0.36fF $ **FLOATING
C9399 S.n8548 SUB 0.61fF $ **FLOATING
C9400 S.n8549 SUB 0.12fF $ **FLOATING
C9401 S.t1341 SUB 0.02fF
C9402 S.n8550 SUB 0.14fF $ **FLOATING
C9403 S.n8552 SUB 1.16fF $ **FLOATING
C9404 S.n8553 SUB 0.22fF $ **FLOATING
C9405 S.n8554 SUB 0.25fF $ **FLOATING
C9406 S.n8555 SUB 0.09fF $ **FLOATING
C9407 S.n8556 SUB 2.44fF $ **FLOATING
C9408 S.t1072 SUB 0.02fF
C9409 S.n8557 SUB 0.24fF $ **FLOATING
C9410 S.n8558 SUB 0.91fF $ **FLOATING
C9411 S.n8559 SUB 0.05fF $ **FLOATING
C9412 S.t2126 SUB 0.02fF
C9413 S.n8560 SUB 0.12fF $ **FLOATING
C9414 S.n8561 SUB 0.14fF $ **FLOATING
C9415 S.n8563 SUB 1.88fF $ **FLOATING
C9416 S.n8564 SUB 0.48fF $ **FLOATING
C9417 S.n8565 SUB 0.09fF $ **FLOATING
C9418 S.n8566 SUB 0.33fF $ **FLOATING
C9419 S.n8567 SUB 0.30fF $ **FLOATING
C9420 S.n8568 SUB 0.77fF $ **FLOATING
C9421 S.n8569 SUB 0.59fF $ **FLOATING
C9422 S.t713 SUB 0.02fF
C9423 S.n8570 SUB 0.24fF $ **FLOATING
C9424 S.n8571 SUB 0.36fF $ **FLOATING
C9425 S.n8572 SUB 0.61fF $ **FLOATING
C9426 S.n8573 SUB 0.12fF $ **FLOATING
C9427 S.t462 SUB 0.02fF
C9428 S.n8574 SUB 0.14fF $ **FLOATING
C9429 S.n8576 SUB 2.61fF $ **FLOATING
C9430 S.n8577 SUB 2.16fF $ **FLOATING
C9431 S.t195 SUB 0.02fF
C9432 S.n8578 SUB 0.24fF $ **FLOATING
C9433 S.n8579 SUB 0.91fF $ **FLOATING
C9434 S.n8580 SUB 0.05fF $ **FLOATING
C9435 S.t1260 SUB 0.02fF
C9436 S.n8581 SUB 0.12fF $ **FLOATING
C9437 S.n8582 SUB 0.14fF $ **FLOATING
C9438 S.n8584 SUB 0.78fF $ **FLOATING
C9439 S.n8585 SUB 2.30fF $ **FLOATING
C9440 S.n8586 SUB 1.88fF $ **FLOATING
C9441 S.n8587 SUB 0.12fF $ **FLOATING
C9442 S.t2113 SUB 0.02fF
C9443 S.n8588 SUB 0.14fF $ **FLOATING
C9444 S.t2368 SUB 0.02fF
C9445 S.n8590 SUB 0.24fF $ **FLOATING
C9446 S.n8591 SUB 0.36fF $ **FLOATING
C9447 S.n8592 SUB 0.61fF $ **FLOATING
C9448 S.n8593 SUB 1.39fF $ **FLOATING
C9449 S.n8594 SUB 0.71fF $ **FLOATING
C9450 S.n8595 SUB 1.14fF $ **FLOATING
C9451 S.n8596 SUB 0.35fF $ **FLOATING
C9452 S.n8597 SUB 2.03fF $ **FLOATING
C9453 S.t1863 SUB 0.02fF
C9454 S.n8598 SUB 0.24fF $ **FLOATING
C9455 S.n8599 SUB 0.91fF $ **FLOATING
C9456 S.n8600 SUB 0.05fF $ **FLOATING
C9457 S.t377 SUB 0.02fF
C9458 S.n8601 SUB 0.12fF $ **FLOATING
C9459 S.n8602 SUB 0.14fF $ **FLOATING
C9460 S.n8604 SUB 1.89fF $ **FLOATING
C9461 S.n8605 SUB 1.88fF $ **FLOATING
C9462 S.t1512 SUB 0.02fF
C9463 S.n8606 SUB 0.24fF $ **FLOATING
C9464 S.n8607 SUB 0.36fF $ **FLOATING
C9465 S.n8608 SUB 0.61fF $ **FLOATING
C9466 S.n8609 SUB 0.12fF $ **FLOATING
C9467 S.t1242 SUB 0.02fF
C9468 S.n8610 SUB 0.14fF $ **FLOATING
C9469 S.n8612 SUB 1.16fF $ **FLOATING
C9470 S.n8613 SUB 0.22fF $ **FLOATING
C9471 S.n8614 SUB 0.25fF $ **FLOATING
C9472 S.n8615 SUB 0.09fF $ **FLOATING
C9473 S.n8616 SUB 1.88fF $ **FLOATING
C9474 S.t994 SUB 0.02fF
C9475 S.n8617 SUB 0.24fF $ **FLOATING
C9476 S.n8618 SUB 0.91fF $ **FLOATING
C9477 S.n8619 SUB 0.05fF $ **FLOATING
C9478 S.t2028 SUB 0.02fF
C9479 S.n8620 SUB 0.12fF $ **FLOATING
C9480 S.n8621 SUB 0.14fF $ **FLOATING
C9481 S.n8623 SUB 20.78fF $ **FLOATING
C9482 S.n8624 SUB 1.88fF $ **FLOATING
C9483 S.n8625 SUB 2.67fF $ **FLOATING
C9484 S.t333 SUB 0.02fF
C9485 S.n8626 SUB 0.24fF $ **FLOATING
C9486 S.n8627 SUB 0.36fF $ **FLOATING
C9487 S.n8628 SUB 0.61fF $ **FLOATING
C9488 S.n8629 SUB 0.12fF $ **FLOATING
C9489 S.t1100 SUB 0.02fF
C9490 S.n8630 SUB 0.14fF $ **FLOATING
C9491 S.n8632 SUB 2.80fF $ **FLOATING
C9492 S.n8633 SUB 2.30fF $ **FLOATING
C9493 S.t1763 SUB 0.02fF
C9494 S.n8634 SUB 0.12fF $ **FLOATING
C9495 S.n8635 SUB 0.14fF $ **FLOATING
C9496 S.t1295 SUB 0.02fF
C9497 S.n8637 SUB 0.24fF $ **FLOATING
C9498 S.n8638 SUB 0.91fF $ **FLOATING
C9499 S.n8639 SUB 0.05fF $ **FLOATING
C9500 S.n8640 SUB 1.88fF $ **FLOATING
C9501 S.n8641 SUB 2.67fF $ **FLOATING
C9502 S.t1990 SUB 0.02fF
C9503 S.n8642 SUB 0.24fF $ **FLOATING
C9504 S.n8643 SUB 0.36fF $ **FLOATING
C9505 S.n8644 SUB 0.61fF $ **FLOATING
C9506 S.n8645 SUB 0.12fF $ **FLOATING
C9507 S.t225 SUB 0.02fF
C9508 S.n8646 SUB 0.14fF $ **FLOATING
C9509 S.n8648 SUB 2.80fF $ **FLOATING
C9510 S.n8649 SUB 2.30fF $ **FLOATING
C9511 S.t890 SUB 0.02fF
C9512 S.n8650 SUB 0.12fF $ **FLOATING
C9513 S.n8651 SUB 0.14fF $ **FLOATING
C9514 S.t411 SUB 0.02fF
C9515 S.n8653 SUB 0.24fF $ **FLOATING
C9516 S.n8654 SUB 0.91fF $ **FLOATING
C9517 S.n8655 SUB 0.05fF $ **FLOATING
C9518 S.n8656 SUB 1.88fF $ **FLOATING
C9519 S.n8657 SUB 2.67fF $ **FLOATING
C9520 S.t1140 SUB 0.02fF
C9521 S.n8658 SUB 0.24fF $ **FLOATING
C9522 S.n8659 SUB 0.36fF $ **FLOATING
C9523 S.n8660 SUB 0.61fF $ **FLOATING
C9524 S.n8661 SUB 0.12fF $ **FLOATING
C9525 S.t1892 SUB 0.02fF
C9526 S.n8662 SUB 0.14fF $ **FLOATING
C9527 S.n8664 SUB 2.80fF $ **FLOATING
C9528 S.n8665 SUB 2.30fF $ **FLOATING
C9529 S.t2533 SUB 0.02fF
C9530 S.n8666 SUB 0.12fF $ **FLOATING
C9531 S.n8667 SUB 0.14fF $ **FLOATING
C9532 S.t2059 SUB 0.02fF
C9533 S.n8669 SUB 0.24fF $ **FLOATING
C9534 S.n8670 SUB 0.91fF $ **FLOATING
C9535 S.n8671 SUB 0.05fF $ **FLOATING
C9536 S.n8672 SUB 1.88fF $ **FLOATING
C9537 S.n8673 SUB 2.67fF $ **FLOATING
C9538 S.t265 SUB 0.02fF
C9539 S.n8674 SUB 0.24fF $ **FLOATING
C9540 S.n8675 SUB 0.36fF $ **FLOATING
C9541 S.n8676 SUB 0.61fF $ **FLOATING
C9542 S.n8677 SUB 0.12fF $ **FLOATING
C9543 S.t1031 SUB 0.02fF
C9544 S.n8678 SUB 0.14fF $ **FLOATING
C9545 S.n8680 SUB 2.80fF $ **FLOATING
C9546 S.n8681 SUB 2.30fF $ **FLOATING
C9547 S.t1660 SUB 0.02fF
C9548 S.n8682 SUB 0.12fF $ **FLOATING
C9549 S.n8683 SUB 0.14fF $ **FLOATING
C9550 S.t1199 SUB 0.02fF
C9551 S.n8685 SUB 0.24fF $ **FLOATING
C9552 S.n8686 SUB 0.91fF $ **FLOATING
C9553 S.n8687 SUB 0.05fF $ **FLOATING
C9554 S.n8688 SUB 1.88fF $ **FLOATING
C9555 S.n8689 SUB 2.67fF $ **FLOATING
C9556 S.t1928 SUB 0.02fF
C9557 S.n8690 SUB 0.24fF $ **FLOATING
C9558 S.n8691 SUB 0.36fF $ **FLOATING
C9559 S.n8692 SUB 0.61fF $ **FLOATING
C9560 S.n8693 SUB 0.12fF $ **FLOATING
C9561 S.t134 SUB 0.02fF
C9562 S.n8694 SUB 0.14fF $ **FLOATING
C9563 S.n8696 SUB 2.80fF $ **FLOATING
C9564 S.n8697 SUB 2.30fF $ **FLOATING
C9565 S.t952 SUB 0.02fF
C9566 S.n8698 SUB 0.12fF $ **FLOATING
C9567 S.n8699 SUB 0.14fF $ **FLOATING
C9568 S.t319 SUB 0.02fF
C9569 S.n8701 SUB 0.24fF $ **FLOATING
C9570 S.n8702 SUB 0.91fF $ **FLOATING
C9571 S.n8703 SUB 0.05fF $ **FLOATING
C9572 S.n8704 SUB 1.88fF $ **FLOATING
C9573 S.n8705 SUB 2.67fF $ **FLOATING
C9574 S.t1068 SUB 0.02fF
C9575 S.n8706 SUB 0.24fF $ **FLOATING
C9576 S.n8707 SUB 0.36fF $ **FLOATING
C9577 S.n8708 SUB 0.61fF $ **FLOATING
C9578 S.n8709 SUB 0.12fF $ **FLOATING
C9579 S.t1803 SUB 0.02fF
C9580 S.n8710 SUB 0.14fF $ **FLOATING
C9581 S.n8712 SUB 2.80fF $ **FLOATING
C9582 S.n8713 SUB 2.30fF $ **FLOATING
C9583 S.t1 SUB 0.02fF
C9584 S.n8714 SUB 0.12fF $ **FLOATING
C9585 S.n8715 SUB 0.14fF $ **FLOATING
C9586 S.t1982 SUB 0.02fF
C9587 S.n8717 SUB 0.24fF $ **FLOATING
C9588 S.n8718 SUB 0.91fF $ **FLOATING
C9589 S.n8719 SUB 0.05fF $ **FLOATING
C9590 S.n8720 SUB 1.88fF $ **FLOATING
C9591 S.n8721 SUB 2.67fF $ **FLOATING
C9592 S.t189 SUB 0.02fF
C9593 S.n8722 SUB 0.24fF $ **FLOATING
C9594 S.n8723 SUB 0.36fF $ **FLOATING
C9595 S.n8724 SUB 0.61fF $ **FLOATING
C9596 S.n8725 SUB 0.12fF $ **FLOATING
C9597 S.t935 SUB 0.02fF
C9598 S.n8726 SUB 0.14fF $ **FLOATING
C9599 S.n8728 SUB 2.80fF $ **FLOATING
C9600 S.n8729 SUB 2.30fF $ **FLOATING
C9601 S.t1716 SUB 0.02fF
C9602 S.n8730 SUB 0.12fF $ **FLOATING
C9603 S.n8731 SUB 0.14fF $ **FLOATING
C9604 S.t1134 SUB 0.02fF
C9605 S.n8733 SUB 0.24fF $ **FLOATING
C9606 S.n8734 SUB 0.91fF $ **FLOATING
C9607 S.n8735 SUB 0.05fF $ **FLOATING
C9608 S.n8736 SUB 1.88fF $ **FLOATING
C9609 S.n8737 SUB 2.68fF $ **FLOATING
C9610 S.t1856 SUB 0.02fF
C9611 S.n8738 SUB 0.24fF $ **FLOATING
C9612 S.n8739 SUB 0.36fF $ **FLOATING
C9613 S.n8740 SUB 0.61fF $ **FLOATING
C9614 S.n8741 SUB 0.12fF $ **FLOATING
C9615 S.t2577 SUB 0.02fF
C9616 S.n8742 SUB 0.14fF $ **FLOATING
C9617 S.n8744 SUB 5.17fF $ **FLOATING
C9618 S.t845 SUB 0.02fF
C9619 S.n8745 SUB 0.12fF $ **FLOATING
C9620 S.n8746 SUB 0.14fF $ **FLOATING
C9621 S.t255 SUB 0.02fF
C9622 S.n8748 SUB 0.24fF $ **FLOATING
C9623 S.n8749 SUB 0.91fF $ **FLOATING
C9624 S.n8750 SUB 0.05fF $ **FLOATING
C9625 S.n8751 SUB 2.73fF $ **FLOATING
C9626 S.n8752 SUB 1.59fF $ **FLOATING
C9627 S.n8753 SUB 0.12fF $ **FLOATING
C9628 S.t548 SUB 0.02fF
C9629 S.n8754 SUB 0.14fF $ **FLOATING
C9630 S.t1890 SUB 0.02fF
C9631 S.n8756 SUB 0.24fF $ **FLOATING
C9632 S.n8757 SUB 0.36fF $ **FLOATING
C9633 S.n8758 SUB 0.61fF $ **FLOATING
C9634 S.n8759 SUB 0.07fF $ **FLOATING
C9635 S.n8760 SUB 0.01fF $ **FLOATING
C9636 S.n8761 SUB 0.24fF $ **FLOATING
C9637 S.n8762 SUB 1.16fF $ **FLOATING
C9638 S.n8763 SUB 1.35fF $ **FLOATING
C9639 S.n8764 SUB 2.30fF $ **FLOATING
C9640 S.t1282 SUB 0.02fF
C9641 S.n8765 SUB 0.12fF $ **FLOATING
C9642 S.n8766 SUB 0.14fF $ **FLOATING
C9643 S.t2203 SUB 0.02fF
C9644 S.n8768 SUB 0.24fF $ **FLOATING
C9645 S.n8769 SUB 0.91fF $ **FLOATING
C9646 S.n8770 SUB 0.05fF $ **FLOATING
C9647 S.t0 SUB 48.31fF
C9648 S.t1170 SUB 0.02fF
C9649 S.n8771 SUB 0.12fF $ **FLOATING
C9650 S.n8772 SUB 0.14fF $ **FLOATING
C9651 S.t85 SUB 0.02fF
C9652 S.n8774 SUB 0.24fF $ **FLOATING
C9653 S.n8775 SUB 0.91fF $ **FLOATING
C9654 S.n8776 SUB 0.05fF $ **FLOATING
C9655 S.t651 SUB 0.02fF
C9656 S.n8777 SUB 0.24fF $ **FLOATING
C9657 S.n8778 SUB 0.36fF $ **FLOATING
C9658 S.n8779 SUB 0.61fF $ **FLOATING
C9659 S.n8780 SUB 0.32fF $ **FLOATING
C9660 S.n8781 SUB 1.09fF $ **FLOATING
C9661 S.n8782 SUB 0.15fF $ **FLOATING
C9662 S.n8783 SUB 2.10fF $ **FLOATING
C9663 S.n8784 SUB 2.94fF $ **FLOATING
C9664 S.n8785 SUB 1.88fF $ **FLOATING
C9665 S.n8786 SUB 0.12fF $ **FLOATING
C9666 S.t1437 SUB 0.02fF
C9667 S.n8787 SUB 0.14fF $ **FLOATING
C9668 S.t1958 SUB 0.02fF
C9669 S.n8789 SUB 0.24fF $ **FLOATING
C9670 S.n8790 SUB 0.36fF $ **FLOATING
C9671 S.n8791 SUB 0.61fF $ **FLOATING
C9672 S.n8792 SUB 0.92fF $ **FLOATING
C9673 S.n8793 SUB 0.32fF $ **FLOATING
C9674 S.n8794 SUB 0.92fF $ **FLOATING
C9675 S.n8795 SUB 1.09fF $ **FLOATING
C9676 S.n8796 SUB 0.15fF $ **FLOATING
C9677 S.n8797 SUB 4.96fF $ **FLOATING
C9678 S.t1591 SUB 0.02fF
C9679 S.n8798 SUB 0.12fF $ **FLOATING
C9680 S.n8799 SUB 0.14fF $ **FLOATING
C9681 S.t267 SUB 0.02fF
C9682 S.n8801 SUB 0.24fF $ **FLOATING
C9683 S.n8802 SUB 0.91fF $ **FLOATING
C9684 S.n8803 SUB 0.05fF $ **FLOATING
C9685 S.n8804 SUB 1.88fF $ **FLOATING
C9686 S.n8805 SUB 2.67fF $ **FLOATING
C9687 S.t1369 SUB 0.02fF
C9688 S.n8806 SUB 0.24fF $ **FLOATING
C9689 S.n8807 SUB 0.36fF $ **FLOATING
C9690 S.n8808 SUB 0.61fF $ **FLOATING
C9691 S.n8809 SUB 0.12fF $ **FLOATING
C9692 S.t787 SUB 0.02fF
C9693 S.n8810 SUB 0.14fF $ **FLOATING
C9694 S.n8812 SUB 1.88fF $ **FLOATING
C9695 S.n8813 SUB 2.67fF $ **FLOATING
C9696 S.t1212 SUB 0.02fF
C9697 S.n8814 SUB 0.24fF $ **FLOATING
C9698 S.n8815 SUB 0.36fF $ **FLOATING
C9699 S.n8816 SUB 0.61fF $ **FLOATING
C9700 S.t2158 SUB 0.02fF
C9701 S.n8817 SUB 0.24fF $ **FLOATING
C9702 S.n8818 SUB 0.91fF $ **FLOATING
C9703 S.n8819 SUB 0.05fF $ **FLOATING
C9704 S.t295 SUB 0.02fF
C9705 S.n8820 SUB 0.12fF $ **FLOATING
C9706 S.n8821 SUB 0.14fF $ **FLOATING
C9707 S.n8823 SUB 0.12fF $ **FLOATING
C9708 S.t1959 SUB 0.02fF
C9709 S.n8824 SUB 0.14fF $ **FLOATING
C9710 S.n8826 SUB 2.30fF $ **FLOATING
C9711 S.n8827 SUB 2.94fF $ **FLOATING
C9712 S.n8828 SUB 5.16fF $ **FLOATING
C9713 S.t1030 SUB 0.02fF
C9714 S.n8829 SUB 0.12fF $ **FLOATING
C9715 S.n8830 SUB 0.14fF $ **FLOATING
C9716 S.t1263 SUB 0.02fF
C9717 S.n8832 SUB 0.24fF $ **FLOATING
C9718 S.n8833 SUB 0.91fF $ **FLOATING
C9719 S.n8834 SUB 0.05fF $ **FLOATING
C9720 S.n8835 SUB 1.88fF $ **FLOATING
C9721 S.n8836 SUB 2.67fF $ **FLOATING
C9722 S.t496 SUB 0.02fF
C9723 S.n8837 SUB 0.24fF $ **FLOATING
C9724 S.n8838 SUB 0.36fF $ **FLOATING
C9725 S.n8839 SUB 0.61fF $ **FLOATING
C9726 S.n8840 SUB 0.12fF $ **FLOATING
C9727 S.t2438 SUB 0.02fF
C9728 S.n8841 SUB 0.14fF $ **FLOATING
C9729 S.n8843 SUB 5.17fF $ **FLOATING
C9730 S.t132 SUB 0.02fF
C9731 S.n8844 SUB 0.12fF $ **FLOATING
C9732 S.n8845 SUB 0.14fF $ **FLOATING
C9733 S.t379 SUB 0.02fF
C9734 S.n8847 SUB 0.24fF $ **FLOATING
C9735 S.n8848 SUB 0.91fF $ **FLOATING
C9736 S.n8849 SUB 0.05fF $ **FLOATING
C9737 S.n8850 SUB 1.88fF $ **FLOATING
C9738 S.n8851 SUB 2.67fF $ **FLOATING
C9739 S.t2142 SUB 0.02fF
C9740 S.n8852 SUB 0.24fF $ **FLOATING
C9741 S.n8853 SUB 0.36fF $ **FLOATING
C9742 S.n8854 SUB 0.61fF $ **FLOATING
C9743 S.n8855 SUB 0.12fF $ **FLOATING
C9744 S.t1574 SUB 0.02fF
C9745 S.n8856 SUB 0.14fF $ **FLOATING
C9746 S.n8858 SUB 5.17fF $ **FLOATING
C9747 S.t1801 SUB 0.02fF
C9748 S.n8859 SUB 0.12fF $ **FLOATING
C9749 S.n8860 SUB 0.14fF $ **FLOATING
C9750 S.t2031 SUB 0.02fF
C9751 S.n8862 SUB 0.24fF $ **FLOATING
C9752 S.n8863 SUB 0.91fF $ **FLOATING
C9753 S.n8864 SUB 0.05fF $ **FLOATING
C9754 S.n8865 SUB 1.88fF $ **FLOATING
C9755 S.n8866 SUB 2.67fF $ **FLOATING
C9756 S.t1280 SUB 0.02fF
C9757 S.n8867 SUB 0.24fF $ **FLOATING
C9758 S.n8868 SUB 0.36fF $ **FLOATING
C9759 S.n8869 SUB 0.61fF $ **FLOATING
C9760 S.n8870 SUB 0.12fF $ **FLOATING
C9761 S.t704 SUB 0.02fF
C9762 S.n8871 SUB 0.14fF $ **FLOATING
C9763 S.n8873 SUB 5.17fF $ **FLOATING
C9764 S.t934 SUB 0.02fF
C9765 S.n8874 SUB 0.12fF $ **FLOATING
C9766 S.n8875 SUB 0.14fF $ **FLOATING
C9767 S.t1176 SUB 0.02fF
C9768 S.n8877 SUB 0.24fF $ **FLOATING
C9769 S.n8878 SUB 0.91fF $ **FLOATING
C9770 S.n8879 SUB 0.05fF $ **FLOATING
C9771 S.n8880 SUB 1.88fF $ **FLOATING
C9772 S.n8881 SUB 2.67fF $ **FLOATING
C9773 S.t552 SUB 0.02fF
C9774 S.n8882 SUB 0.24fF $ **FLOATING
C9775 S.n8883 SUB 0.36fF $ **FLOATING
C9776 S.n8884 SUB 0.61fF $ **FLOATING
C9777 S.n8885 SUB 0.12fF $ **FLOATING
C9778 S.t2486 SUB 0.02fF
C9779 S.n8886 SUB 0.14fF $ **FLOATING
C9780 S.n8888 SUB 5.17fF $ **FLOATING
C9781 S.t2574 SUB 0.02fF
C9782 S.n8889 SUB 0.12fF $ **FLOATING
C9783 S.n8890 SUB 0.14fF $ **FLOATING
C9784 S.t432 SUB 0.02fF
C9785 S.n8892 SUB 0.24fF $ **FLOATING
C9786 S.n8893 SUB 0.91fF $ **FLOATING
C9787 S.n8894 SUB 0.05fF $ **FLOATING
C9788 S.n8895 SUB 1.88fF $ **FLOATING
C9789 S.n8896 SUB 2.67fF $ **FLOATING
C9790 S.t2191 SUB 0.02fF
C9791 S.n8897 SUB 0.24fF $ **FLOATING
C9792 S.n8898 SUB 0.36fF $ **FLOATING
C9793 S.n8899 SUB 0.61fF $ **FLOATING
C9794 S.n8900 SUB 0.12fF $ **FLOATING
C9795 S.t1614 SUB 0.02fF
C9796 S.n8901 SUB 0.14fF $ **FLOATING
C9797 S.n8903 SUB 5.17fF $ **FLOATING
C9798 S.t1698 SUB 0.02fF
C9799 S.n8904 SUB 0.12fF $ **FLOATING
C9800 S.n8905 SUB 0.14fF $ **FLOATING
C9801 S.t2079 SUB 0.02fF
C9802 S.n8907 SUB 0.24fF $ **FLOATING
C9803 S.n8908 SUB 0.91fF $ **FLOATING
C9804 S.n8909 SUB 0.05fF $ **FLOATING
C9805 S.n8910 SUB 1.88fF $ **FLOATING
C9806 S.n8911 SUB 2.67fF $ **FLOATING
C9807 S.t1334 SUB 0.02fF
C9808 S.n8912 SUB 0.24fF $ **FLOATING
C9809 S.n8913 SUB 0.36fF $ **FLOATING
C9810 S.n8914 SUB 0.61fF $ **FLOATING
C9811 S.n8915 SUB 0.12fF $ **FLOATING
C9812 S.t749 SUB 0.02fF
C9813 S.n8916 SUB 0.14fF $ **FLOATING
C9814 S.n8918 SUB 5.17fF $ **FLOATING
C9815 S.t824 SUB 0.02fF
C9816 S.n8919 SUB 0.12fF $ **FLOATING
C9817 S.n8920 SUB 0.14fF $ **FLOATING
C9818 S.t1219 SUB 0.02fF
C9819 S.n8922 SUB 0.24fF $ **FLOATING
C9820 S.n8923 SUB 0.91fF $ **FLOATING
C9821 S.n8924 SUB 0.05fF $ **FLOATING
C9822 S.n8925 SUB 1.88fF $ **FLOATING
C9823 S.n8926 SUB 2.67fF $ **FLOATING
C9824 S.t454 SUB 0.02fF
C9825 S.n8927 SUB 0.24fF $ **FLOATING
C9826 S.n8928 SUB 0.36fF $ **FLOATING
C9827 S.n8929 SUB 0.61fF $ **FLOATING
C9828 S.n8930 SUB 0.12fF $ **FLOATING
C9829 S.t2401 SUB 0.02fF
C9830 S.n8931 SUB 0.14fF $ **FLOATING
C9831 S.n8933 SUB 4.90fF $ **FLOATING
C9832 S.t2469 SUB 0.02fF
C9833 S.n8934 SUB 0.12fF $ **FLOATING
C9834 S.n8935 SUB 0.14fF $ **FLOATING
C9835 S.t337 SUB 0.02fF
C9836 S.n8937 SUB 0.24fF $ **FLOATING
C9837 S.n8938 SUB 0.91fF $ **FLOATING
C9838 S.n8939 SUB 0.05fF $ **FLOATING
C9839 S.n8940 SUB 1.88fF $ **FLOATING
C9840 S.n8941 SUB 2.67fF $ **FLOATING
C9841 S.t1963 SUB 0.02fF
C9842 S.n8942 SUB 0.24fF $ **FLOATING
C9843 S.n8943 SUB 0.36fF $ **FLOATING
C9844 S.n8944 SUB 0.61fF $ **FLOATING
C9845 S.n8945 SUB 0.12fF $ **FLOATING
C9846 S.t674 SUB 0.02fF
C9847 S.n8946 SUB 0.14fF $ **FLOATING
C9848 S.n8948 SUB 5.44fF $ **FLOATING
C9849 S.t1599 SUB 0.02fF
C9850 S.n8949 SUB 0.12fF $ **FLOATING
C9851 S.n8950 SUB 0.14fF $ **FLOATING
C9852 S.t718 SUB 0.02fF
C9853 S.n8952 SUB 0.24fF $ **FLOATING
C9854 S.n8953 SUB 0.91fF $ **FLOATING
C9855 S.n8954 SUB 0.05fF $ **FLOATING
C9856 S.t131 SUB 47.92fF
C9857 S.t407 SUB 0.02fF
C9858 S.n8955 SUB 1.19fF $ **FLOATING
C9859 S.n8956 SUB 0.05fF $ **FLOATING
C9860 S.t2430 SUB 0.02fF
C9861 S.n8957 SUB 0.01fF $ **FLOATING
C9862 S.n8958 SUB 0.26fF $ **FLOATING
C9863 S.n8960 SUB 1.50fF $ **FLOATING
C9864 S.n8961 SUB 1.30fF $ **FLOATING
C9865 S.n8962 SUB 0.28fF $ **FLOATING
C9866 S.n8963 SUB 0.24fF $ **FLOATING
C9867 S.n8964 SUB 4.39fF $ **FLOATING
C9868 S.n8965 SUB 0.01fF $ **FLOATING
C9869 S.n8966 SUB 0.02fF $ **FLOATING
C9870 S.n8967 SUB 0.03fF $ **FLOATING
C9871 S.n8968 SUB 0.04fF $ **FLOATING
C9872 S.n8969 SUB 0.17fF $ **FLOATING
C9873 S.n8970 SUB 0.01fF $ **FLOATING
C9874 S.n8971 SUB 0.02fF $ **FLOATING
C9875 S.n8972 SUB 0.01fF $ **FLOATING
C9876 S.n8973 SUB 0.01fF $ **FLOATING
C9877 S.n8974 SUB 0.01fF $ **FLOATING
C9878 S.n8975 SUB 0.01fF $ **FLOATING
C9879 S.n8976 SUB 0.02fF $ **FLOATING
C9880 S.n8977 SUB 0.01fF $ **FLOATING
C9881 S.n8978 SUB 0.02fF $ **FLOATING
C9882 S.n8979 SUB 0.05fF $ **FLOATING
C9883 S.n8980 SUB 0.04fF $ **FLOATING
C9884 S.n8981 SUB 0.11fF $ **FLOATING
C9885 S.n8982 SUB 0.38fF $ **FLOATING
C9886 S.n8983 SUB 0.20fF $ **FLOATING
C9887 S.n8984 SUB 8.97fF $ **FLOATING
C9888 S.n8985 SUB 8.97fF $ **FLOATING
C9889 S.n8986 SUB 0.60fF $ **FLOATING
C9890 S.n8987 SUB 0.22fF $ **FLOATING
C9891 S.n8988 SUB 0.59fF $ **FLOATING
C9892 S.n8989 SUB 3.43fF $ **FLOATING
C9893 S.n8990 SUB 0.29fF $ **FLOATING
C9894 S.t67 SUB 21.38fF
C9895 S.n8991 SUB 21.67fF $ **FLOATING
C9896 S.n8992 SUB 0.77fF $ **FLOATING
C9897 S.n8993 SUB 0.28fF $ **FLOATING
C9898 S.n8994 SUB 4.00fF $ **FLOATING
C9899 S.n8995 SUB 1.35fF $ **FLOATING
C9900 S.t2197 SUB 0.02fF
C9901 S.n8996 SUB 0.64fF $ **FLOATING
C9902 S.n8997 SUB 0.61fF $ **FLOATING
C9903 S.n8998 SUB 0.25fF $ **FLOATING
C9904 S.n8999 SUB 0.09fF $ **FLOATING
C9905 S.n9000 SUB 0.21fF $ **FLOATING
C9906 S.n9001 SUB 0.92fF $ **FLOATING
C9907 S.n9002 SUB 0.44fF $ **FLOATING
C9908 S.n9003 SUB 1.88fF $ **FLOATING
C9909 S.n9004 SUB 0.12fF $ **FLOATING
C9910 S.t1175 SUB 0.02fF
C9911 S.n9005 SUB 0.14fF $ **FLOATING
C9912 S.t1695 SUB 0.02fF
C9913 S.n9007 SUB 0.24fF $ **FLOATING
C9914 S.n9008 SUB 0.36fF $ **FLOATING
C9915 S.n9009 SUB 0.61fF $ **FLOATING
C9916 S.n9010 SUB 0.02fF $ **FLOATING
C9917 S.n9011 SUB 0.01fF $ **FLOATING
C9918 S.n9012 SUB 0.02fF $ **FLOATING
C9919 S.n9013 SUB 0.08fF $ **FLOATING
C9920 S.n9014 SUB 0.06fF $ **FLOATING
C9921 S.n9015 SUB 0.03fF $ **FLOATING
C9922 S.n9016 SUB 0.04fF $ **FLOATING
C9923 S.n9017 SUB 1.00fF $ **FLOATING
C9924 S.n9018 SUB 0.36fF $ **FLOATING
C9925 S.n9019 SUB 1.87fF $ **FLOATING
C9926 S.n9020 SUB 1.99fF $ **FLOATING
C9927 S.t2525 SUB 0.02fF
C9928 S.n9021 SUB 0.24fF $ **FLOATING
C9929 S.n9022 SUB 0.91fF $ **FLOATING
C9930 S.n9023 SUB 0.05fF $ **FLOATING
C9931 S.t1390 SUB 0.02fF
C9932 S.n9024 SUB 0.12fF $ **FLOATING
C9933 S.n9025 SUB 0.14fF $ **FLOATING
C9934 S.n9027 SUB 1.89fF $ **FLOATING
C9935 S.n9028 SUB 0.07fF $ **FLOATING
C9936 S.n9029 SUB 0.04fF $ **FLOATING
C9937 S.n9030 SUB 0.05fF $ **FLOATING
C9938 S.n9031 SUB 0.87fF $ **FLOATING
C9939 S.n9032 SUB 0.01fF $ **FLOATING
C9940 S.n9033 SUB 0.01fF $ **FLOATING
C9941 S.n9034 SUB 0.01fF $ **FLOATING
C9942 S.n9035 SUB 0.07fF $ **FLOATING
C9943 S.n9036 SUB 0.68fF $ **FLOATING
C9944 S.n9037 SUB 0.72fF $ **FLOATING
C9945 S.t987 SUB 0.02fF
C9946 S.n9038 SUB 0.24fF $ **FLOATING
C9947 S.n9039 SUB 0.36fF $ **FLOATING
C9948 S.n9040 SUB 0.61fF $ **FLOATING
C9949 S.n9041 SUB 0.12fF $ **FLOATING
C9950 S.t433 SUB 0.02fF
C9951 S.n9042 SUB 0.14fF $ **FLOATING
C9952 S.n9044 SUB 0.70fF $ **FLOATING
C9953 S.n9045 SUB 0.23fF $ **FLOATING
C9954 S.n9046 SUB 0.23fF $ **FLOATING
C9955 S.n9047 SUB 0.70fF $ **FLOATING
C9956 S.n9048 SUB 1.16fF $ **FLOATING
C9957 S.n9049 SUB 0.22fF $ **FLOATING
C9958 S.n9050 SUB 0.25fF $ **FLOATING
C9959 S.n9051 SUB 0.09fF $ **FLOATING
C9960 S.n9052 SUB 2.31fF $ **FLOATING
C9961 S.t1813 SUB 0.02fF
C9962 S.n9053 SUB 0.24fF $ **FLOATING
C9963 S.n9054 SUB 0.91fF $ **FLOATING
C9964 S.n9055 SUB 0.05fF $ **FLOATING
C9965 S.t517 SUB 0.02fF
C9966 S.n9056 SUB 0.12fF $ **FLOATING
C9967 S.n9057 SUB 0.14fF $ **FLOATING
C9968 S.n9059 SUB 1.88fF $ **FLOATING
C9969 S.n9060 SUB 0.46fF $ **FLOATING
C9970 S.n9061 SUB 0.22fF $ **FLOATING
C9971 S.n9062 SUB 0.38fF $ **FLOATING
C9972 S.n9063 SUB 0.16fF $ **FLOATING
C9973 S.n9064 SUB 0.28fF $ **FLOATING
C9974 S.n9065 SUB 0.21fF $ **FLOATING
C9975 S.n9066 SUB 0.30fF $ **FLOATING
C9976 S.n9067 SUB 0.42fF $ **FLOATING
C9977 S.n9068 SUB 0.21fF $ **FLOATING
C9978 S.t68 SUB 0.02fF
C9979 S.n9069 SUB 0.24fF $ **FLOATING
C9980 S.n9070 SUB 0.36fF $ **FLOATING
C9981 S.n9071 SUB 0.61fF $ **FLOATING
C9982 S.n9072 SUB 0.12fF $ **FLOATING
C9983 S.t2080 SUB 0.02fF
C9984 S.n9073 SUB 0.14fF $ **FLOATING
C9985 S.n9075 SUB 0.04fF $ **FLOATING
C9986 S.n9076 SUB 0.03fF $ **FLOATING
C9987 S.n9077 SUB 0.03fF $ **FLOATING
C9988 S.n9078 SUB 0.10fF $ **FLOATING
C9989 S.n9079 SUB 0.36fF $ **FLOATING
C9990 S.n9080 SUB 0.38fF $ **FLOATING
C9991 S.n9081 SUB 0.11fF $ **FLOATING
C9992 S.n9082 SUB 0.12fF $ **FLOATING
C9993 S.n9083 SUB 0.07fF $ **FLOATING
C9994 S.n9084 SUB 0.12fF $ **FLOATING
C9995 S.n9085 SUB 0.18fF $ **FLOATING
C9996 S.n9086 SUB 4.00fF $ **FLOATING
C9997 S.t946 SUB 0.02fF
C9998 S.n9087 SUB 0.24fF $ **FLOATING
C9999 S.n9088 SUB 0.91fF $ **FLOATING
C10000 S.n9089 SUB 0.05fF $ **FLOATING
C10001 S.t2162 SUB 0.02fF
C10002 S.n9090 SUB 0.12fF $ **FLOATING
C10003 S.n9091 SUB 0.14fF $ **FLOATING
C10004 S.n9093 SUB 0.25fF $ **FLOATING
C10005 S.n9094 SUB 0.09fF $ **FLOATING
C10006 S.n9095 SUB 0.21fF $ **FLOATING
C10007 S.n9096 SUB 1.28fF $ **FLOATING
C10008 S.n9097 SUB 0.53fF $ **FLOATING
C10009 S.n9098 SUB 1.88fF $ **FLOATING
C10010 S.n9099 SUB 0.12fF $ **FLOATING
C10011 S.t1217 SUB 0.02fF
C10012 S.n9100 SUB 0.14fF $ **FLOATING
C10013 S.t1752 SUB 0.02fF
C10014 S.n9102 SUB 0.24fF $ **FLOATING
C10015 S.n9103 SUB 0.36fF $ **FLOATING
C10016 S.n9104 SUB 0.61fF $ **FLOATING
C10017 S.n9105 SUB 1.58fF $ **FLOATING
C10018 S.n9106 SUB 2.45fF $ **FLOATING
C10019 S.t2583 SUB 0.02fF
C10020 S.n9107 SUB 0.24fF $ **FLOATING
C10021 S.n9108 SUB 0.91fF $ **FLOATING
C10022 S.n9109 SUB 0.05fF $ **FLOATING
C10023 S.t1298 SUB 0.02fF
C10024 S.n9110 SUB 0.12fF $ **FLOATING
C10025 S.n9111 SUB 0.14fF $ **FLOATING
C10026 S.n9113 SUB 1.89fF $ **FLOATING
C10027 S.n9114 SUB 0.06fF $ **FLOATING
C10028 S.n9115 SUB 0.03fF $ **FLOATING
C10029 S.n9116 SUB 0.04fF $ **FLOATING
C10030 S.n9117 SUB 0.99fF $ **FLOATING
C10031 S.n9118 SUB 0.02fF $ **FLOATING
C10032 S.n9119 SUB 0.01fF $ **FLOATING
C10033 S.n9120 SUB 0.02fF $ **FLOATING
C10034 S.n9121 SUB 0.08fF $ **FLOATING
C10035 S.n9122 SUB 0.36fF $ **FLOATING
C10036 S.n9123 SUB 1.85fF $ **FLOATING
C10037 S.t875 SUB 0.02fF
C10038 S.n9124 SUB 0.24fF $ **FLOATING
C10039 S.n9125 SUB 0.36fF $ **FLOATING
C10040 S.n9126 SUB 0.61fF $ **FLOATING
C10041 S.n9127 SUB 0.12fF $ **FLOATING
C10042 S.t338 SUB 0.02fF
C10043 S.n9128 SUB 0.14fF $ **FLOATING
C10044 S.n9130 SUB 0.70fF $ **FLOATING
C10045 S.n9131 SUB 0.23fF $ **FLOATING
C10046 S.n9132 SUB 0.23fF $ **FLOATING
C10047 S.n9133 SUB 0.70fF $ **FLOATING
C10048 S.n9134 SUB 1.16fF $ **FLOATING
C10049 S.n9135 SUB 0.22fF $ **FLOATING
C10050 S.n9136 SUB 0.25fF $ **FLOATING
C10051 S.n9137 SUB 0.09fF $ **FLOATING
C10052 S.n9138 SUB 1.88fF $ **FLOATING
C10053 S.t1705 SUB 0.02fF
C10054 S.n9139 SUB 0.24fF $ **FLOATING
C10055 S.n9140 SUB 0.91fF $ **FLOATING
C10056 S.n9141 SUB 0.05fF $ **FLOATING
C10057 S.t415 SUB 0.02fF
C10058 S.n9142 SUB 0.12fF $ **FLOATING
C10059 S.n9143 SUB 0.14fF $ **FLOATING
C10060 S.n9145 SUB 20.78fF $ **FLOATING
C10061 S.n9146 SUB 1.72fF $ **FLOATING
C10062 S.n9147 SUB 3.05fF $ **FLOATING
C10063 S.t2568 SUB 0.02fF
C10064 S.n9148 SUB 0.24fF $ **FLOATING
C10065 S.n9149 SUB 0.36fF $ **FLOATING
C10066 S.n9150 SUB 0.61fF $ **FLOATING
C10067 S.n9151 SUB 0.12fF $ **FLOATING
C10068 S.t2030 SUB 0.02fF
C10069 S.n9152 SUB 0.14fF $ **FLOATING
C10070 S.n9154 SUB 0.31fF $ **FLOATING
C10071 S.n9155 SUB 0.23fF $ **FLOATING
C10072 S.n9156 SUB 0.66fF $ **FLOATING
C10073 S.n9157 SUB 0.95fF $ **FLOATING
C10074 S.n9158 SUB 0.23fF $ **FLOATING
C10075 S.n9159 SUB 0.21fF $ **FLOATING
C10076 S.n9160 SUB 0.20fF $ **FLOATING
C10077 S.n9161 SUB 0.06fF $ **FLOATING
C10078 S.n9162 SUB 0.09fF $ **FLOATING
C10079 S.n9163 SUB 0.10fF $ **FLOATING
C10080 S.n9164 SUB 1.99fF $ **FLOATING
C10081 S.t2248 SUB 0.02fF
C10082 S.n9165 SUB 0.12fF $ **FLOATING
C10083 S.n9166 SUB 0.14fF $ **FLOATING
C10084 S.t880 SUB 0.02fF
C10085 S.n9168 SUB 0.24fF $ **FLOATING
C10086 S.n9169 SUB 0.91fF $ **FLOATING
C10087 S.n9170 SUB 0.05fF $ **FLOATING
C10088 S.n9171 SUB 1.88fF $ **FLOATING
C10089 S.n9172 SUB 0.12fF $ **FLOATING
C10090 S.t975 SUB 0.02fF
C10091 S.n9173 SUB 0.14fF $ **FLOATING
C10092 S.t1756 SUB 0.02fF
C10093 S.n9175 SUB 0.12fF $ **FLOATING
C10094 S.n9176 SUB 0.14fF $ **FLOATING
C10095 S.t677 SUB 0.02fF
C10096 S.n9178 SUB 0.24fF $ **FLOATING
C10097 S.n9179 SUB 0.91fF $ **FLOATING
C10098 S.n9180 SUB 0.05fF $ **FLOATING
C10099 S.t1238 SUB 0.02fF
C10100 S.n9181 SUB 0.24fF $ **FLOATING
C10101 S.n9182 SUB 0.36fF $ **FLOATING
C10102 S.n9183 SUB 0.61fF $ **FLOATING
C10103 S.n9184 SUB 0.32fF $ **FLOATING
C10104 S.n9185 SUB 1.09fF $ **FLOATING
C10105 S.n9186 SUB 0.15fF $ **FLOATING
C10106 S.n9187 SUB 2.10fF $ **FLOATING
C10107 S.n9188 SUB 2.94fF $ **FLOATING
C10108 S.n9189 SUB 1.88fF $ **FLOATING
C10109 S.n9190 SUB 0.12fF $ **FLOATING
C10110 S.t1996 SUB 0.02fF
C10111 S.n9191 SUB 0.14fF $ **FLOATING
C10112 S.t2521 SUB 0.02fF
C10113 S.n9193 SUB 0.24fF $ **FLOATING
C10114 S.n9194 SUB 0.36fF $ **FLOATING
C10115 S.n9195 SUB 0.61fF $ **FLOATING
C10116 S.n9196 SUB 0.92fF $ **FLOATING
C10117 S.n9197 SUB 0.32fF $ **FLOATING
C10118 S.n9198 SUB 0.92fF $ **FLOATING
C10119 S.n9199 SUB 1.09fF $ **FLOATING
C10120 S.n9200 SUB 0.15fF $ **FLOATING
C10121 S.n9201 SUB 4.96fF $ **FLOATING
C10122 S.t2063 SUB 0.02fF
C10123 S.n9202 SUB 0.12fF $ **FLOATING
C10124 S.n9203 SUB 0.14fF $ **FLOATING
C10125 S.t833 SUB 0.02fF
C10126 S.n9205 SUB 0.24fF $ **FLOATING
C10127 S.n9206 SUB 0.91fF $ **FLOATING
C10128 S.n9207 SUB 0.05fF $ **FLOATING
C10129 S.n9208 SUB 1.88fF $ **FLOATING
C10130 S.n9209 SUB 2.67fF $ **FLOATING
C10131 S.t1643 SUB 0.02fF
C10132 S.n9210 SUB 0.24fF $ **FLOATING
C10133 S.n9211 SUB 0.36fF $ **FLOATING
C10134 S.n9212 SUB 0.61fF $ **FLOATING
C10135 S.n9213 SUB 0.12fF $ **FLOATING
C10136 S.t1145 SUB 0.02fF
C10137 S.n9214 SUB 0.14fF $ **FLOATING
C10138 S.n9216 SUB 1.88fF $ **FLOATING
C10139 S.n9217 SUB 2.67fF $ **FLOATING
C10140 S.t353 SUB 0.02fF
C10141 S.n9218 SUB 0.24fF $ **FLOATING
C10142 S.n9219 SUB 0.36fF $ **FLOATING
C10143 S.n9220 SUB 0.61fF $ **FLOATING
C10144 S.t2334 SUB 0.02fF
C10145 S.n9221 SUB 0.24fF $ **FLOATING
C10146 S.n9222 SUB 0.91fF $ **FLOATING
C10147 S.n9223 SUB 0.05fF $ **FLOATING
C10148 S.t878 SUB 0.02fF
C10149 S.n9224 SUB 0.12fF $ **FLOATING
C10150 S.n9225 SUB 0.14fF $ **FLOATING
C10151 S.n9227 SUB 0.12fF $ **FLOATING
C10152 S.t218 SUB 0.02fF
C10153 S.n9228 SUB 0.14fF $ **FLOATING
C10154 S.n9230 SUB 2.30fF $ **FLOATING
C10155 S.n9231 SUB 2.94fF $ **FLOATING
C10156 S.n9232 SUB 5.16fF $ **FLOATING
C10157 S.t1351 SUB 0.02fF
C10158 S.n9233 SUB 0.12fF $ **FLOATING
C10159 S.n9234 SUB 0.14fF $ **FLOATING
C10160 S.t2478 SUB 0.02fF
C10161 S.n9236 SUB 0.24fF $ **FLOATING
C10162 S.n9237 SUB 0.91fF $ **FLOATING
C10163 S.n9238 SUB 0.05fF $ **FLOATING
C10164 S.n9239 SUB 1.88fF $ **FLOATING
C10165 S.n9240 SUB 2.67fF $ **FLOATING
C10166 S.t525 SUB 0.02fF
C10167 S.n9241 SUB 0.24fF $ **FLOATING
C10168 S.n9242 SUB 0.36fF $ **FLOATING
C10169 S.n9243 SUB 0.61fF $ **FLOATING
C10170 S.n9244 SUB 0.12fF $ **FLOATING
C10171 S.t2462 SUB 0.02fF
C10172 S.n9245 SUB 0.14fF $ **FLOATING
C10173 S.n9247 SUB 5.17fF $ **FLOATING
C10174 S.t166 SUB 0.02fF
C10175 S.n9248 SUB 0.12fF $ **FLOATING
C10176 S.n9249 SUB 0.14fF $ **FLOATING
C10177 S.t408 SUB 0.02fF
C10178 S.n9251 SUB 0.24fF $ **FLOATING
C10179 S.n9252 SUB 0.91fF $ **FLOATING
C10180 S.n9253 SUB 0.05fF $ **FLOATING
C10181 S.n9254 SUB 1.88fF $ **FLOATING
C10182 S.n9255 SUB 2.67fF $ **FLOATING
C10183 S.t2169 SUB 0.02fF
C10184 S.n9256 SUB 0.24fF $ **FLOATING
C10185 S.n9257 SUB 0.36fF $ **FLOATING
C10186 S.n9258 SUB 0.61fF $ **FLOATING
C10187 S.n9259 SUB 0.12fF $ **FLOATING
C10188 S.t1593 SUB 0.02fF
C10189 S.n9260 SUB 0.14fF $ **FLOATING
C10190 S.n9262 SUB 5.17fF $ **FLOATING
C10191 S.t1829 SUB 0.02fF
C10192 S.n9263 SUB 0.12fF $ **FLOATING
C10193 S.n9264 SUB 0.14fF $ **FLOATING
C10194 S.t2055 SUB 0.02fF
C10195 S.n9266 SUB 0.24fF $ **FLOATING
C10196 S.n9267 SUB 0.91fF $ **FLOATING
C10197 S.n9268 SUB 0.05fF $ **FLOATING
C10198 S.n9269 SUB 1.88fF $ **FLOATING
C10199 S.n9270 SUB 2.67fF $ **FLOATING
C10200 S.t1306 SUB 0.02fF
C10201 S.n9271 SUB 0.24fF $ **FLOATING
C10202 S.n9272 SUB 0.36fF $ **FLOATING
C10203 S.n9273 SUB 0.61fF $ **FLOATING
C10204 S.n9274 SUB 0.12fF $ **FLOATING
C10205 S.t730 SUB 0.02fF
C10206 S.n9275 SUB 0.14fF $ **FLOATING
C10207 S.n9277 SUB 5.17fF $ **FLOATING
C10208 S.t963 SUB 0.02fF
C10209 S.n9278 SUB 0.12fF $ **FLOATING
C10210 S.n9279 SUB 0.14fF $ **FLOATING
C10211 S.t1198 SUB 0.02fF
C10212 S.n9281 SUB 0.24fF $ **FLOATING
C10213 S.n9282 SUB 0.91fF $ **FLOATING
C10214 S.n9283 SUB 0.05fF $ **FLOATING
C10215 S.n9284 SUB 1.88fF $ **FLOATING
C10216 S.n9285 SUB 2.67fF $ **FLOATING
C10217 S.t424 SUB 0.02fF
C10218 S.n9286 SUB 0.24fF $ **FLOATING
C10219 S.n9287 SUB 0.36fF $ **FLOATING
C10220 S.n9288 SUB 0.61fF $ **FLOATING
C10221 S.n9289 SUB 0.12fF $ **FLOATING
C10222 S.t2383 SUB 0.02fF
C10223 S.n9290 SUB 0.14fF $ **FLOATING
C10224 S.n9292 SUB 5.17fF $ **FLOATING
C10225 S.t25 SUB 0.02fF
C10226 S.n9293 SUB 0.12fF $ **FLOATING
C10227 S.n9294 SUB 0.14fF $ **FLOATING
C10228 S.t318 SUB 0.02fF
C10229 S.n9296 SUB 0.24fF $ **FLOATING
C10230 S.n9297 SUB 0.91fF $ **FLOATING
C10231 S.n9298 SUB 0.05fF $ **FLOATING
C10232 S.n9299 SUB 1.88fF $ **FLOATING
C10233 S.n9300 SUB 2.67fF $ **FLOATING
C10234 S.t2218 SUB 0.02fF
C10235 S.n9301 SUB 0.24fF $ **FLOATING
C10236 S.n9302 SUB 0.36fF $ **FLOATING
C10237 S.n9303 SUB 0.61fF $ **FLOATING
C10238 S.n9304 SUB 0.12fF $ **FLOATING
C10239 S.t1641 SUB 0.02fF
C10240 S.n9305 SUB 0.14fF $ **FLOATING
C10241 S.n9307 SUB 5.17fF $ **FLOATING
C10242 S.t1729 SUB 0.02fF
C10243 S.n9308 SUB 0.12fF $ **FLOATING
C10244 S.n9309 SUB 0.14fF $ **FLOATING
C10245 S.t2115 SUB 0.02fF
C10246 S.n9311 SUB 0.24fF $ **FLOATING
C10247 S.n9312 SUB 0.91fF $ **FLOATING
C10248 S.n9313 SUB 0.05fF $ **FLOATING
C10249 S.n9314 SUB 1.88fF $ **FLOATING
C10250 S.n9315 SUB 2.67fF $ **FLOATING
C10251 S.t1358 SUB 0.02fF
C10252 S.n9316 SUB 0.24fF $ **FLOATING
C10253 S.n9317 SUB 0.36fF $ **FLOATING
C10254 S.n9318 SUB 0.61fF $ **FLOATING
C10255 S.n9319 SUB 0.12fF $ **FLOATING
C10256 S.t773 SUB 0.02fF
C10257 S.n9320 SUB 0.14fF $ **FLOATING
C10258 S.n9322 SUB 5.17fF $ **FLOATING
C10259 S.t856 SUB 0.02fF
C10260 S.n9323 SUB 0.12fF $ **FLOATING
C10261 S.n9324 SUB 0.14fF $ **FLOATING
C10262 S.t1247 SUB 0.02fF
C10263 S.n9326 SUB 0.24fF $ **FLOATING
C10264 S.n9327 SUB 0.91fF $ **FLOATING
C10265 S.n9328 SUB 0.05fF $ **FLOATING
C10266 S.n9329 SUB 1.88fF $ **FLOATING
C10267 S.n9330 SUB 2.67fF $ **FLOATING
C10268 S.t484 SUB 0.02fF
C10269 S.n9331 SUB 0.24fF $ **FLOATING
C10270 S.n9332 SUB 0.36fF $ **FLOATING
C10271 S.n9333 SUB 0.61fF $ **FLOATING
C10272 S.n9334 SUB 0.12fF $ **FLOATING
C10273 S.t2424 SUB 0.02fF
C10274 S.n9335 SUB 0.14fF $ **FLOATING
C10275 S.n9337 SUB 5.17fF $ **FLOATING
C10276 S.t2500 SUB 0.02fF
C10277 S.n9338 SUB 0.12fF $ **FLOATING
C10278 S.n9339 SUB 0.14fF $ **FLOATING
C10279 S.t366 SUB 0.02fF
C10280 S.n9341 SUB 0.24fF $ **FLOATING
C10281 S.n9342 SUB 0.91fF $ **FLOATING
C10282 S.n9343 SUB 0.05fF $ **FLOATING
C10283 S.n9344 SUB 1.88fF $ **FLOATING
C10284 S.n9345 SUB 2.67fF $ **FLOATING
C10285 S.t2131 SUB 0.02fF
C10286 S.n9346 SUB 0.24fF $ **FLOATING
C10287 S.n9347 SUB 0.36fF $ **FLOATING
C10288 S.n9348 SUB 0.61fF $ **FLOATING
C10289 S.n9349 SUB 0.12fF $ **FLOATING
C10290 S.t1559 SUB 0.02fF
C10291 S.n9350 SUB 0.14fF $ **FLOATING
C10292 S.n9352 SUB 4.90fF $ **FLOATING
C10293 S.t1625 SUB 0.02fF
C10294 S.n9353 SUB 0.12fF $ **FLOATING
C10295 S.n9354 SUB 0.14fF $ **FLOATING
C10296 S.t2018 SUB 0.02fF
C10297 S.n9356 SUB 0.24fF $ **FLOATING
C10298 S.n9357 SUB 0.91fF $ **FLOATING
C10299 S.n9358 SUB 0.05fF $ **FLOATING
C10300 S.n9359 SUB 1.88fF $ **FLOATING
C10301 S.n9360 SUB 2.67fF $ **FLOATING
C10302 S.t607 SUB 0.02fF
C10303 S.n9361 SUB 0.24fF $ **FLOATING
C10304 S.n9362 SUB 0.36fF $ **FLOATING
C10305 S.n9363 SUB 0.61fF $ **FLOATING
C10306 S.n9364 SUB 0.12fF $ **FLOATING
C10307 S.t1860 SUB 0.02fF
C10308 S.n9365 SUB 0.14fF $ **FLOATING
C10309 S.n9367 SUB 1.88fF $ **FLOATING
C10310 S.n9368 SUB 2.68fF $ **FLOATING
C10311 S.t1018 SUB 0.02fF
C10312 S.n9369 SUB 0.24fF $ **FLOATING
C10313 S.n9370 SUB 0.36fF $ **FLOATING
C10314 S.n9371 SUB 0.61fF $ **FLOATING
C10315 S.t1423 SUB 0.02fF
C10316 S.n9372 SUB 1.22fF $ **FLOATING
C10317 S.n9373 SUB 0.61fF $ **FLOATING
C10318 S.n9374 SUB 0.35fF $ **FLOATING
C10319 S.n9375 SUB 0.63fF $ **FLOATING
C10320 S.n9376 SUB 1.15fF $ **FLOATING
C10321 S.n9377 SUB 3.03fF $ **FLOATING
C10322 S.n9378 SUB 0.59fF $ **FLOATING
C10323 S.n9379 SUB 0.02fF $ **FLOATING
C10324 S.n9380 SUB 0.97fF $ **FLOATING
C10325 S.t212 SUB 21.38fF
C10326 S.n9381 SUB 20.25fF $ **FLOATING
C10327 S.n9383 SUB 0.38fF $ **FLOATING
C10328 S.n9384 SUB 0.23fF $ **FLOATING
C10329 S.n9385 SUB 2.90fF $ **FLOATING
C10330 S.n9386 SUB 2.46fF $ **FLOATING
C10331 S.n9387 SUB 1.96fF $ **FLOATING
C10332 S.n9388 SUB 3.94fF $ **FLOATING
C10333 S.n9389 SUB 0.25fF $ **FLOATING
C10334 S.n9390 SUB 0.01fF $ **FLOATING
C10335 S.t1132 SUB 0.02fF
C10336 S.n9391 SUB 0.25fF $ **FLOATING
C10337 S.t841 SUB 0.02fF
C10338 S.n9392 SUB 0.95fF $ **FLOATING
C10339 S.n9393 SUB 0.70fF $ **FLOATING
C10340 S.n9394 SUB 0.78fF $ **FLOATING
C10341 S.n9395 SUB 1.93fF $ **FLOATING
C10342 S.n9396 SUB 1.88fF $ **FLOATING
C10343 S.n9397 SUB 0.12fF $ **FLOATING
C10344 S.t254 SUB 0.02fF
C10345 S.n9398 SUB 0.14fF $ **FLOATING
C10346 S.t556 SUB 0.02fF
C10347 S.n9400 SUB 0.24fF $ **FLOATING
C10348 S.n9401 SUB 0.36fF $ **FLOATING
C10349 S.n9402 SUB 0.61fF $ **FLOATING
C10350 S.n9403 SUB 1.52fF $ **FLOATING
C10351 S.n9404 SUB 2.99fF $ **FLOATING
C10352 S.t2484 SUB 0.02fF
C10353 S.n9405 SUB 0.24fF $ **FLOATING
C10354 S.n9406 SUB 0.91fF $ **FLOATING
C10355 S.n9407 SUB 0.05fF $ **FLOATING
C10356 S.t936 SUB 0.02fF
C10357 S.n9408 SUB 0.12fF $ **FLOATING
C10358 S.n9409 SUB 0.14fF $ **FLOATING
C10359 S.n9411 SUB 1.89fF $ **FLOATING
C10360 S.n9412 SUB 1.75fF $ **FLOATING
C10361 S.t2195 SUB 0.02fF
C10362 S.n9413 SUB 0.24fF $ **FLOATING
C10363 S.n9414 SUB 0.36fF $ **FLOATING
C10364 S.n9415 SUB 0.61fF $ **FLOATING
C10365 S.n9416 SUB 0.12fF $ **FLOATING
C10366 S.t1921 SUB 0.02fF
C10367 S.n9417 SUB 0.14fF $ **FLOATING
C10368 S.n9419 SUB 1.16fF $ **FLOATING
C10369 S.n9420 SUB 0.22fF $ **FLOATING
C10370 S.n9421 SUB 0.25fF $ **FLOATING
C10371 S.n9422 SUB 0.09fF $ **FLOATING
C10372 S.n9423 SUB 2.44fF $ **FLOATING
C10373 S.t1610 SUB 0.02fF
C10374 S.n9424 SUB 0.24fF $ **FLOATING
C10375 S.n9425 SUB 0.91fF $ **FLOATING
C10376 S.n9426 SUB 0.05fF $ **FLOATING
C10377 S.t2575 SUB 0.02fF
C10378 S.n9427 SUB 0.12fF $ **FLOATING
C10379 S.n9428 SUB 0.14fF $ **FLOATING
C10380 S.n9430 SUB 1.88fF $ **FLOATING
C10381 S.n9431 SUB 0.48fF $ **FLOATING
C10382 S.n9432 SUB 0.09fF $ **FLOATING
C10383 S.n9433 SUB 0.33fF $ **FLOATING
C10384 S.n9434 SUB 0.30fF $ **FLOATING
C10385 S.n9435 SUB 0.77fF $ **FLOATING
C10386 S.n9436 SUB 0.59fF $ **FLOATING
C10387 S.t1339 SUB 0.02fF
C10388 S.n9437 SUB 0.24fF $ **FLOATING
C10389 S.n9438 SUB 0.36fF $ **FLOATING
C10390 S.n9439 SUB 0.61fF $ **FLOATING
C10391 S.n9440 SUB 0.12fF $ **FLOATING
C10392 S.t1059 SUB 0.02fF
C10393 S.n9441 SUB 0.14fF $ **FLOATING
C10394 S.n9443 SUB 2.61fF $ **FLOATING
C10395 S.n9444 SUB 2.16fF $ **FLOATING
C10396 S.t746 SUB 0.02fF
C10397 S.n9445 SUB 0.24fF $ **FLOATING
C10398 S.n9446 SUB 0.91fF $ **FLOATING
C10399 S.n9447 SUB 0.05fF $ **FLOATING
C10400 S.t1857 SUB 0.02fF
C10401 S.n9448 SUB 0.12fF $ **FLOATING
C10402 S.n9449 SUB 0.14fF $ **FLOATING
C10403 S.n9451 SUB 0.78fF $ **FLOATING
C10404 S.n9452 SUB 2.30fF $ **FLOATING
C10405 S.n9453 SUB 1.88fF $ **FLOATING
C10406 S.n9454 SUB 0.12fF $ **FLOATING
C10407 S.t174 SUB 0.02fF
C10408 S.n9455 SUB 0.14fF $ **FLOATING
C10409 S.t458 SUB 0.02fF
C10410 S.n9457 SUB 0.24fF $ **FLOATING
C10411 S.n9458 SUB 0.36fF $ **FLOATING
C10412 S.n9459 SUB 0.61fF $ **FLOATING
C10413 S.n9460 SUB 1.39fF $ **FLOATING
C10414 S.n9461 SUB 0.71fF $ **FLOATING
C10415 S.n9462 SUB 1.14fF $ **FLOATING
C10416 S.n9463 SUB 0.35fF $ **FLOATING
C10417 S.n9464 SUB 2.03fF $ **FLOATING
C10418 S.t2399 SUB 0.02fF
C10419 S.n9465 SUB 0.24fF $ **FLOATING
C10420 S.n9466 SUB 0.91fF $ **FLOATING
C10421 S.n9467 SUB 0.05fF $ **FLOATING
C10422 S.t990 SUB 0.02fF
C10423 S.n9468 SUB 0.12fF $ **FLOATING
C10424 S.n9469 SUB 0.14fF $ **FLOATING
C10425 S.n9471 SUB 1.89fF $ **FLOATING
C10426 S.n9472 SUB 1.88fF $ **FLOATING
C10427 S.t2104 SUB 0.02fF
C10428 S.n9473 SUB 0.24fF $ **FLOATING
C10429 S.n9474 SUB 0.36fF $ **FLOATING
C10430 S.n9475 SUB 0.61fF $ **FLOATING
C10431 S.n9476 SUB 0.12fF $ **FLOATING
C10432 S.t1837 SUB 0.02fF
C10433 S.n9477 SUB 0.14fF $ **FLOATING
C10434 S.n9479 SUB 1.16fF $ **FLOATING
C10435 S.n9480 SUB 0.22fF $ **FLOATING
C10436 S.n9481 SUB 0.25fF $ **FLOATING
C10437 S.n9482 SUB 0.09fF $ **FLOATING
C10438 S.n9483 SUB 1.88fF $ **FLOATING
C10439 S.t1538 SUB 0.02fF
C10440 S.n9484 SUB 0.24fF $ **FLOATING
C10441 S.n9485 SUB 0.91fF $ **FLOATING
C10442 S.n9486 SUB 0.05fF $ **FLOATING
C10443 S.t77 SUB 0.02fF
C10444 S.n9487 SUB 0.12fF $ **FLOATING
C10445 S.n9488 SUB 0.14fF $ **FLOATING
C10446 S.n9490 SUB 20.78fF $ **FLOATING
C10447 S.n9491 SUB 1.88fF $ **FLOATING
C10448 S.n9492 SUB 2.67fF $ **FLOATING
C10449 S.t358 SUB 0.02fF
C10450 S.n9493 SUB 0.24fF $ **FLOATING
C10451 S.n9494 SUB 0.36fF $ **FLOATING
C10452 S.n9495 SUB 0.61fF $ **FLOATING
C10453 S.n9496 SUB 0.12fF $ **FLOATING
C10454 S.t1126 SUB 0.02fF
C10455 S.n9497 SUB 0.14fF $ **FLOATING
C10456 S.n9499 SUB 2.80fF $ **FLOATING
C10457 S.n9500 SUB 2.30fF $ **FLOATING
C10458 S.t2522 SUB 0.02fF
C10459 S.n9501 SUB 0.12fF $ **FLOATING
C10460 S.n9502 SUB 0.14fF $ **FLOATING
C10461 S.t1324 SUB 0.02fF
C10462 S.n9504 SUB 0.24fF $ **FLOATING
C10463 S.n9505 SUB 0.91fF $ **FLOATING
C10464 S.n9506 SUB 0.05fF $ **FLOATING
C10465 S.n9507 SUB 1.88fF $ **FLOATING
C10466 S.n9508 SUB 2.67fF $ **FLOATING
C10467 S.t2012 SUB 0.02fF
C10468 S.n9509 SUB 0.24fF $ **FLOATING
C10469 S.n9510 SUB 0.36fF $ **FLOATING
C10470 S.n9511 SUB 0.61fF $ **FLOATING
C10471 S.n9512 SUB 0.12fF $ **FLOATING
C10472 S.t247 SUB 0.02fF
C10473 S.n9513 SUB 0.14fF $ **FLOATING
C10474 S.n9515 SUB 2.80fF $ **FLOATING
C10475 S.n9516 SUB 2.30fF $ **FLOATING
C10476 S.t924 SUB 0.02fF
C10477 S.n9517 SUB 0.12fF $ **FLOATING
C10478 S.n9518 SUB 0.14fF $ **FLOATING
C10479 S.t446 SUB 0.02fF
C10480 S.n9520 SUB 0.24fF $ **FLOATING
C10481 S.n9521 SUB 0.91fF $ **FLOATING
C10482 S.n9522 SUB 0.05fF $ **FLOATING
C10483 S.n9523 SUB 1.88fF $ **FLOATING
C10484 S.n9524 SUB 2.67fF $ **FLOATING
C10485 S.t1160 SUB 0.02fF
C10486 S.n9525 SUB 0.24fF $ **FLOATING
C10487 S.n9526 SUB 0.36fF $ **FLOATING
C10488 S.n9527 SUB 0.61fF $ **FLOATING
C10489 S.n9528 SUB 0.12fF $ **FLOATING
C10490 S.t1914 SUB 0.02fF
C10491 S.n9529 SUB 0.14fF $ **FLOATING
C10492 S.n9531 SUB 2.80fF $ **FLOATING
C10493 S.n9532 SUB 2.30fF $ **FLOATING
C10494 S.t2564 SUB 0.02fF
C10495 S.n9533 SUB 0.12fF $ **FLOATING
C10496 S.n9534 SUB 0.14fF $ **FLOATING
C10497 S.t2089 SUB 0.02fF
C10498 S.n9536 SUB 0.24fF $ **FLOATING
C10499 S.n9537 SUB 0.91fF $ **FLOATING
C10500 S.n9538 SUB 0.05fF $ **FLOATING
C10501 S.n9539 SUB 1.88fF $ **FLOATING
C10502 S.n9540 SUB 2.67fF $ **FLOATING
C10503 S.t288 SUB 0.02fF
C10504 S.n9541 SUB 0.24fF $ **FLOATING
C10505 S.n9542 SUB 0.36fF $ **FLOATING
C10506 S.n9543 SUB 0.61fF $ **FLOATING
C10507 S.n9544 SUB 0.12fF $ **FLOATING
C10508 S.t1054 SUB 0.02fF
C10509 S.n9545 SUB 0.14fF $ **FLOATING
C10510 S.n9547 SUB 2.80fF $ **FLOATING
C10511 S.n9548 SUB 2.30fF $ **FLOATING
C10512 S.t1690 SUB 0.02fF
C10513 S.n9549 SUB 0.12fF $ **FLOATING
C10514 S.n9550 SUB 0.14fF $ **FLOATING
C10515 S.t1227 SUB 0.02fF
C10516 S.n9552 SUB 0.24fF $ **FLOATING
C10517 S.n9553 SUB 0.91fF $ **FLOATING
C10518 S.n9554 SUB 0.05fF $ **FLOATING
C10519 S.n9555 SUB 1.88fF $ **FLOATING
C10520 S.n9556 SUB 2.67fF $ **FLOATING
C10521 S.t1949 SUB 0.02fF
C10522 S.n9557 SUB 0.24fF $ **FLOATING
C10523 S.n9558 SUB 0.36fF $ **FLOATING
C10524 S.n9559 SUB 0.61fF $ **FLOATING
C10525 S.n9560 SUB 0.12fF $ **FLOATING
C10526 S.t167 SUB 0.02fF
C10527 S.n9561 SUB 0.14fF $ **FLOATING
C10528 S.n9563 SUB 2.80fF $ **FLOATING
C10529 S.n9564 SUB 2.30fF $ **FLOATING
C10530 S.t816 SUB 0.02fF
C10531 S.n9565 SUB 0.12fF $ **FLOATING
C10532 S.n9566 SUB 0.14fF $ **FLOATING
C10533 S.t344 SUB 0.02fF
C10534 S.n9568 SUB 0.24fF $ **FLOATING
C10535 S.n9569 SUB 0.91fF $ **FLOATING
C10536 S.n9570 SUB 0.05fF $ **FLOATING
C10537 S.n9571 SUB 1.88fF $ **FLOATING
C10538 S.n9572 SUB 2.67fF $ **FLOATING
C10539 S.t1091 SUB 0.02fF
C10540 S.n9573 SUB 0.24fF $ **FLOATING
C10541 S.n9574 SUB 0.36fF $ **FLOATING
C10542 S.n9575 SUB 0.61fF $ **FLOATING
C10543 S.n9576 SUB 0.12fF $ **FLOATING
C10544 S.t1830 SUB 0.02fF
C10545 S.n9577 SUB 0.14fF $ **FLOATING
C10546 S.n9579 SUB 2.80fF $ **FLOATING
C10547 S.n9580 SUB 2.30fF $ **FLOATING
C10548 S.t65 SUB 0.02fF
C10549 S.n9581 SUB 0.12fF $ **FLOATING
C10550 S.n9582 SUB 0.14fF $ **FLOATING
C10551 S.t2003 SUB 0.02fF
C10552 S.n9584 SUB 0.24fF $ **FLOATING
C10553 S.n9585 SUB 0.91fF $ **FLOATING
C10554 S.n9586 SUB 0.05fF $ **FLOATING
C10555 S.n9587 SUB 1.88fF $ **FLOATING
C10556 S.n9588 SUB 2.67fF $ **FLOATING
C10557 S.t213 SUB 0.02fF
C10558 S.n9589 SUB 0.24fF $ **FLOATING
C10559 S.n9590 SUB 0.36fF $ **FLOATING
C10560 S.n9591 SUB 0.61fF $ **FLOATING
C10561 S.n9592 SUB 0.12fF $ **FLOATING
C10562 S.t964 SUB 0.02fF
C10563 S.n9593 SUB 0.14fF $ **FLOATING
C10564 S.n9595 SUB 2.80fF $ **FLOATING
C10565 S.n9596 SUB 2.30fF $ **FLOATING
C10566 S.t1751 SUB 0.02fF
C10567 S.n9597 SUB 0.12fF $ **FLOATING
C10568 S.n9598 SUB 0.14fF $ **FLOATING
C10569 S.t1151 SUB 0.02fF
C10570 S.n9600 SUB 0.24fF $ **FLOATING
C10571 S.n9601 SUB 0.91fF $ **FLOATING
C10572 S.n9602 SUB 0.05fF $ **FLOATING
C10573 S.n9603 SUB 1.88fF $ **FLOATING
C10574 S.n9604 SUB 2.67fF $ **FLOATING
C10575 S.t1880 SUB 0.02fF
C10576 S.n9605 SUB 0.24fF $ **FLOATING
C10577 S.n9606 SUB 0.36fF $ **FLOATING
C10578 S.n9607 SUB 0.61fF $ **FLOATING
C10579 S.n9608 SUB 0.12fF $ **FLOATING
C10580 S.t27 SUB 0.02fF
C10581 S.n9609 SUB 0.14fF $ **FLOATING
C10582 S.n9611 SUB 2.80fF $ **FLOATING
C10583 S.n9612 SUB 2.30fF $ **FLOATING
C10584 S.t873 SUB 0.02fF
C10585 S.n9613 SUB 0.12fF $ **FLOATING
C10586 S.n9614 SUB 0.14fF $ **FLOATING
C10587 S.t275 SUB 0.02fF
C10588 S.n9616 SUB 0.24fF $ **FLOATING
C10589 S.n9617 SUB 0.91fF $ **FLOATING
C10590 S.n9618 SUB 0.05fF $ **FLOATING
C10591 S.n9619 SUB 2.73fF $ **FLOATING
C10592 S.n9620 SUB 1.59fF $ **FLOATING
C10593 S.n9621 SUB 0.12fF $ **FLOATING
C10594 S.t1659 SUB 0.02fF
C10595 S.n9622 SUB 0.14fF $ **FLOATING
C10596 S.t480 SUB 0.02fF
C10597 S.n9624 SUB 0.24fF $ **FLOATING
C10598 S.n9625 SUB 0.36fF $ **FLOATING
C10599 S.n9626 SUB 0.61fF $ **FLOATING
C10600 S.n9627 SUB 0.07fF $ **FLOATING
C10601 S.n9628 SUB 0.01fF $ **FLOATING
C10602 S.n9629 SUB 0.24fF $ **FLOATING
C10603 S.n9630 SUB 1.16fF $ **FLOATING
C10604 S.n9631 SUB 1.35fF $ **FLOATING
C10605 S.n9632 SUB 2.30fF $ **FLOATING
C10606 S.t2400 SUB 0.02fF
C10607 S.n9633 SUB 0.12fF $ **FLOATING
C10608 S.n9634 SUB 0.14fF $ **FLOATING
C10609 S.t766 SUB 0.02fF
C10610 S.n9636 SUB 0.24fF $ **FLOATING
C10611 S.n9637 SUB 0.91fF $ **FLOATING
C10612 S.n9638 SUB 0.05fF $ **FLOATING
C10613 S.t26 SUB 48.31fF
C10614 S.t1938 SUB 0.02fF
C10615 S.n9639 SUB 0.24fF $ **FLOATING
C10616 S.n9640 SUB 0.91fF $ **FLOATING
C10617 S.n9641 SUB 0.05fF $ **FLOATING
C10618 S.t2518 SUB 0.02fF
C10619 S.n9642 SUB 0.12fF $ **FLOATING
C10620 S.n9643 SUB 0.14fF $ **FLOATING
C10621 S.n9645 SUB 0.12fF $ **FLOATING
C10622 S.t1732 SUB 0.02fF
C10623 S.n9646 SUB 0.14fF $ **FLOATING
C10624 S.n9648 SUB 5.17fF $ **FLOATING
C10625 S.n9649 SUB 5.44fF $ **FLOATING
C10626 S.t759 SUB 0.02fF
C10627 S.n9650 SUB 0.12fF $ **FLOATING
C10628 S.n9651 SUB 0.14fF $ **FLOATING
C10629 S.t1912 SUB 0.02fF
C10630 S.n9653 SUB 0.24fF $ **FLOATING
C10631 S.n9654 SUB 0.91fF $ **FLOATING
C10632 S.n9655 SUB 0.05fF $ **FLOATING
C10633 S.t24 SUB 47.92fF
C10634 S.t2084 SUB 0.02fF
C10635 S.n9656 SUB 1.19fF $ **FLOATING
C10636 S.n9657 SUB 0.05fF $ **FLOATING
C10637 S.t1103 SUB 0.02fF
C10638 S.n9658 SUB 0.01fF $ **FLOATING
C10639 S.n9659 SUB 0.26fF $ **FLOATING
C10640 S.n9661 SUB 1.50fF $ **FLOATING
C10641 S.n9662 SUB 1.30fF $ **FLOATING
C10642 S.n9663 SUB 0.28fF $ **FLOATING
C10643 S.n9664 SUB 0.24fF $ **FLOATING
C10644 S.n9665 SUB 4.39fF $ **FLOATING
C10645 S.n9666 SUB 0.01fF $ **FLOATING
C10646 S.n9667 SUB 0.02fF $ **FLOATING
C10647 S.n9668 SUB 0.03fF $ **FLOATING
C10648 S.n9669 SUB 0.04fF $ **FLOATING
C10649 S.n9670 SUB 0.17fF $ **FLOATING
C10650 S.n9671 SUB 0.01fF $ **FLOATING
C10651 S.n9672 SUB 0.02fF $ **FLOATING
C10652 S.n9673 SUB 0.01fF $ **FLOATING
C10653 S.n9674 SUB 0.01fF $ **FLOATING
C10654 S.n9675 SUB 0.01fF $ **FLOATING
C10655 S.n9676 SUB 0.01fF $ **FLOATING
C10656 S.n9677 SUB 0.02fF $ **FLOATING
C10657 S.n9678 SUB 0.01fF $ **FLOATING
C10658 S.n9679 SUB 0.02fF $ **FLOATING
C10659 S.n9680 SUB 0.05fF $ **FLOATING
C10660 S.n9681 SUB 0.04fF $ **FLOATING
C10661 S.n9682 SUB 0.11fF $ **FLOATING
C10662 S.n9683 SUB 0.38fF $ **FLOATING
C10663 S.n9684 SUB 0.20fF $ **FLOATING
C10664 S.n9685 SUB 8.97fF $ **FLOATING
C10665 S.n9686 SUB 8.97fF $ **FLOATING
C10666 S.n9687 SUB 0.60fF $ **FLOATING
C10667 S.n9688 SUB 0.22fF $ **FLOATING
C10668 S.n9689 SUB 0.59fF $ **FLOATING
C10669 S.n9690 SUB 3.43fF $ **FLOATING
C10670 S.n9691 SUB 0.29fF $ **FLOATING
C10671 S.t101 SUB 21.38fF
C10672 S.n9692 SUB 21.67fF $ **FLOATING
C10673 S.n9693 SUB 0.77fF $ **FLOATING
C10674 S.n9694 SUB 0.28fF $ **FLOATING
C10675 S.n9695 SUB 4.00fF $ **FLOATING
C10676 S.n9696 SUB 1.35fF $ **FLOATING
C10677 S.t2212 SUB 0.02fF
C10678 S.n9697 SUB 0.64fF $ **FLOATING
C10679 S.n9698 SUB 0.61fF $ **FLOATING
C10680 S.n9699 SUB 1.89fF $ **FLOATING
C10681 S.n9700 SUB 0.07fF $ **FLOATING
C10682 S.n9701 SUB 0.04fF $ **FLOATING
C10683 S.n9702 SUB 0.05fF $ **FLOATING
C10684 S.n9703 SUB 0.87fF $ **FLOATING
C10685 S.n9704 SUB 0.01fF $ **FLOATING
C10686 S.n9705 SUB 0.01fF $ **FLOATING
C10687 S.n9706 SUB 0.01fF $ **FLOATING
C10688 S.n9707 SUB 0.07fF $ **FLOATING
C10689 S.n9708 SUB 0.68fF $ **FLOATING
C10690 S.n9709 SUB 0.72fF $ **FLOATING
C10691 S.t1144 SUB 0.02fF
C10692 S.n9710 SUB 0.24fF $ **FLOATING
C10693 S.n9711 SUB 0.36fF $ **FLOATING
C10694 S.n9712 SUB 0.61fF $ **FLOATING
C10695 S.n9713 SUB 0.12fF $ **FLOATING
C10696 S.t883 SUB 0.02fF
C10697 S.n9714 SUB 0.14fF $ **FLOATING
C10698 S.n9716 SUB 0.70fF $ **FLOATING
C10699 S.n9717 SUB 0.23fF $ **FLOATING
C10700 S.n9718 SUB 0.23fF $ **FLOATING
C10701 S.n9719 SUB 0.70fF $ **FLOATING
C10702 S.n9720 SUB 1.16fF $ **FLOATING
C10703 S.n9721 SUB 0.22fF $ **FLOATING
C10704 S.n9722 SUB 0.25fF $ **FLOATING
C10705 S.n9723 SUB 0.09fF $ **FLOATING
C10706 S.n9724 SUB 2.31fF $ **FLOATING
C10707 S.t2265 SUB 0.02fF
C10708 S.n9725 SUB 0.24fF $ **FLOATING
C10709 S.n9726 SUB 0.91fF $ **FLOATING
C10710 S.n9727 SUB 0.05fF $ **FLOATING
C10711 S.t1097 SUB 0.02fF
C10712 S.n9728 SUB 0.12fF $ **FLOATING
C10713 S.n9729 SUB 0.14fF $ **FLOATING
C10714 S.n9731 SUB 1.88fF $ **FLOATING
C10715 S.n9732 SUB 0.46fF $ **FLOATING
C10716 S.n9733 SUB 0.22fF $ **FLOATING
C10717 S.n9734 SUB 0.38fF $ **FLOATING
C10718 S.n9735 SUB 0.16fF $ **FLOATING
C10719 S.n9736 SUB 0.28fF $ **FLOATING
C10720 S.n9737 SUB 0.21fF $ **FLOATING
C10721 S.n9738 SUB 0.30fF $ **FLOATING
C10722 S.n9739 SUB 0.42fF $ **FLOATING
C10723 S.n9740 SUB 0.21fF $ **FLOATING
C10724 S.t385 SUB 0.02fF
C10725 S.n9741 SUB 0.24fF $ **FLOATING
C10726 S.n9742 SUB 0.36fF $ **FLOATING
C10727 S.n9743 SUB 0.61fF $ **FLOATING
C10728 S.n9744 SUB 0.12fF $ **FLOATING
C10729 S.t147 SUB 0.02fF
C10730 S.n9745 SUB 0.14fF $ **FLOATING
C10731 S.n9747 SUB 0.04fF $ **FLOATING
C10732 S.n9748 SUB 0.03fF $ **FLOATING
C10733 S.n9749 SUB 0.03fF $ **FLOATING
C10734 S.n9750 SUB 0.10fF $ **FLOATING
C10735 S.n9751 SUB 0.36fF $ **FLOATING
C10736 S.n9752 SUB 0.38fF $ **FLOATING
C10737 S.n9753 SUB 0.11fF $ **FLOATING
C10738 S.n9754 SUB 0.12fF $ **FLOATING
C10739 S.n9755 SUB 0.07fF $ **FLOATING
C10740 S.n9756 SUB 0.12fF $ **FLOATING
C10741 S.n9757 SUB 0.18fF $ **FLOATING
C10742 S.n9758 SUB 4.00fF $ **FLOATING
C10743 S.t1506 SUB 0.02fF
C10744 S.n9759 SUB 0.24fF $ **FLOATING
C10745 S.n9760 SUB 0.91fF $ **FLOATING
C10746 S.n9761 SUB 0.05fF $ **FLOATING
C10747 S.t222 SUB 0.02fF
C10748 S.n9762 SUB 0.12fF $ **FLOATING
C10749 S.n9763 SUB 0.14fF $ **FLOATING
C10750 S.n9765 SUB 0.25fF $ **FLOATING
C10751 S.n9766 SUB 0.09fF $ **FLOATING
C10752 S.n9767 SUB 0.21fF $ **FLOATING
C10753 S.n9768 SUB 1.28fF $ **FLOATING
C10754 S.n9769 SUB 0.53fF $ **FLOATING
C10755 S.n9770 SUB 1.88fF $ **FLOATING
C10756 S.n9771 SUB 0.12fF $ **FLOATING
C10757 S.t1816 SUB 0.02fF
C10758 S.n9772 SUB 0.14fF $ **FLOATING
C10759 S.t2035 SUB 0.02fF
C10760 S.n9774 SUB 0.24fF $ **FLOATING
C10761 S.n9775 SUB 0.36fF $ **FLOATING
C10762 S.n9776 SUB 0.61fF $ **FLOATING
C10763 S.n9777 SUB 1.58fF $ **FLOATING
C10764 S.n9778 SUB 2.45fF $ **FLOATING
C10765 S.t645 SUB 0.02fF
C10766 S.n9779 SUB 0.24fF $ **FLOATING
C10767 S.n9780 SUB 0.91fF $ **FLOATING
C10768 S.n9781 SUB 0.05fF $ **FLOATING
C10769 S.t1887 SUB 0.02fF
C10770 S.n9782 SUB 0.12fF $ **FLOATING
C10771 S.n9783 SUB 0.14fF $ **FLOATING
C10772 S.n9785 SUB 1.89fF $ **FLOATING
C10773 S.n9786 SUB 0.06fF $ **FLOATING
C10774 S.n9787 SUB 0.03fF $ **FLOATING
C10775 S.n9788 SUB 0.04fF $ **FLOATING
C10776 S.n9789 SUB 0.99fF $ **FLOATING
C10777 S.n9790 SUB 0.02fF $ **FLOATING
C10778 S.n9791 SUB 0.01fF $ **FLOATING
C10779 S.n9792 SUB 0.02fF $ **FLOATING
C10780 S.n9793 SUB 0.08fF $ **FLOATING
C10781 S.n9794 SUB 0.36fF $ **FLOATING
C10782 S.n9795 SUB 1.85fF $ **FLOATING
C10783 S.t1180 SUB 0.02fF
C10784 S.n9796 SUB 0.24fF $ **FLOATING
C10785 S.n9797 SUB 0.36fF $ **FLOATING
C10786 S.n9798 SUB 0.61fF $ **FLOATING
C10787 S.n9799 SUB 0.12fF $ **FLOATING
C10788 S.t949 SUB 0.02fF
C10789 S.n9800 SUB 0.14fF $ **FLOATING
C10790 S.n9802 SUB 0.70fF $ **FLOATING
C10791 S.n9803 SUB 0.23fF $ **FLOATING
C10792 S.n9804 SUB 0.23fF $ **FLOATING
C10793 S.n9805 SUB 0.70fF $ **FLOATING
C10794 S.n9806 SUB 1.16fF $ **FLOATING
C10795 S.n9807 SUB 0.22fF $ **FLOATING
C10796 S.n9808 SUB 0.25fF $ **FLOATING
C10797 S.n9809 SUB 0.09fF $ **FLOATING
C10798 S.n9810 SUB 1.88fF $ **FLOATING
C10799 S.t2301 SUB 0.02fF
C10800 S.n9811 SUB 0.24fF $ **FLOATING
C10801 S.n9812 SUB 0.91fF $ **FLOATING
C10802 S.n9813 SUB 0.05fF $ **FLOATING
C10803 S.t1024 SUB 0.02fF
C10804 S.n9814 SUB 0.12fF $ **FLOATING
C10805 S.n9815 SUB 0.14fF $ **FLOATING
C10806 S.n9817 SUB 20.78fF $ **FLOATING
C10807 S.n9818 SUB 0.06fF $ **FLOATING
C10808 S.n9819 SUB 0.20fF $ **FLOATING
C10809 S.n9820 SUB 0.09fF $ **FLOATING
C10810 S.n9821 SUB 0.21fF $ **FLOATING
C10811 S.n9822 SUB 0.10fF $ **FLOATING
C10812 S.n9823 SUB 0.30fF $ **FLOATING
C10813 S.n9824 SUB 0.69fF $ **FLOATING
C10814 S.n9825 SUB 0.45fF $ **FLOATING
C10815 S.n9826 SUB 2.33fF $ **FLOATING
C10816 S.n9827 SUB 0.12fF $ **FLOATING
C10817 S.t1760 SUB 0.02fF
C10818 S.n9828 SUB 0.14fF $ **FLOATING
C10819 S.t1994 SUB 0.02fF
C10820 S.n9830 SUB 0.24fF $ **FLOATING
C10821 S.n9831 SUB 0.36fF $ **FLOATING
C10822 S.n9832 SUB 0.61fF $ **FLOATING
C10823 S.n9833 SUB 1.90fF $ **FLOATING
C10824 S.n9834 SUB 0.17fF $ **FLOATING
C10825 S.n9835 SUB 0.76fF $ **FLOATING
C10826 S.n9836 SUB 0.25fF $ **FLOATING
C10827 S.n9837 SUB 0.30fF $ **FLOATING
C10828 S.n9838 SUB 0.32fF $ **FLOATING
C10829 S.n9839 SUB 0.47fF $ **FLOATING
C10830 S.n9840 SUB 0.16fF $ **FLOATING
C10831 S.n9841 SUB 1.93fF $ **FLOATING
C10832 S.t1957 SUB 0.02fF
C10833 S.n9842 SUB 0.12fF $ **FLOATING
C10834 S.n9843 SUB 0.14fF $ **FLOATING
C10835 S.t611 SUB 0.02fF
C10836 S.n9845 SUB 0.24fF $ **FLOATING
C10837 S.n9846 SUB 0.91fF $ **FLOATING
C10838 S.n9847 SUB 0.05fF $ **FLOATING
C10839 S.n9848 SUB 1.88fF $ **FLOATING
C10840 S.n9849 SUB 0.12fF $ **FLOATING
C10841 S.t1524 SUB 0.02fF
C10842 S.n9850 SUB 0.14fF $ **FLOATING
C10843 S.t2330 SUB 0.02fF
C10844 S.n9852 SUB 0.12fF $ **FLOATING
C10845 S.n9853 SUB 0.14fF $ **FLOATING
C10846 S.t1006 SUB 0.02fF
C10847 S.n9855 SUB 0.24fF $ **FLOATING
C10848 S.n9856 SUB 0.91fF $ **FLOATING
C10849 S.n9857 SUB 0.05fF $ **FLOATING
C10850 S.t1834 SUB 0.02fF
C10851 S.n9858 SUB 0.24fF $ **FLOATING
C10852 S.n9859 SUB 0.36fF $ **FLOATING
C10853 S.n9860 SUB 0.61fF $ **FLOATING
C10854 S.n9861 SUB 0.32fF $ **FLOATING
C10855 S.n9862 SUB 1.09fF $ **FLOATING
C10856 S.n9863 SUB 0.15fF $ **FLOATING
C10857 S.n9864 SUB 2.10fF $ **FLOATING
C10858 S.n9865 SUB 2.94fF $ **FLOATING
C10859 S.n9866 SUB 1.88fF $ **FLOATING
C10860 S.n9867 SUB 0.12fF $ **FLOATING
C10861 S.t2585 SUB 0.02fF
C10862 S.n9868 SUB 0.14fF $ **FLOATING
C10863 S.t303 SUB 0.02fF
C10864 S.n9870 SUB 0.24fF $ **FLOATING
C10865 S.n9871 SUB 0.36fF $ **FLOATING
C10866 S.n9872 SUB 0.61fF $ **FLOATING
C10867 S.n9873 SUB 0.92fF $ **FLOATING
C10868 S.n9874 SUB 0.32fF $ **FLOATING
C10869 S.n9875 SUB 0.92fF $ **FLOATING
C10870 S.n9876 SUB 1.09fF $ **FLOATING
C10871 S.n9877 SUB 0.15fF $ **FLOATING
C10872 S.n9878 SUB 4.96fF $ **FLOATING
C10873 S.t124 SUB 0.02fF
C10874 S.n9879 SUB 0.12fF $ **FLOATING
C10875 S.n9880 SUB 0.14fF $ **FLOATING
C10876 S.t1444 SUB 0.02fF
C10877 S.n9882 SUB 0.24fF $ **FLOATING
C10878 S.n9883 SUB 0.91fF $ **FLOATING
C10879 S.n9884 SUB 0.05fF $ **FLOATING
C10880 S.n9885 SUB 1.88fF $ **FLOATING
C10881 S.n9886 SUB 2.67fF $ **FLOATING
C10882 S.t1967 SUB 0.02fF
C10883 S.n9887 SUB 0.24fF $ **FLOATING
C10884 S.n9888 SUB 0.36fF $ **FLOATING
C10885 S.n9889 SUB 0.61fF $ **FLOATING
C10886 S.n9890 SUB 0.12fF $ **FLOATING
C10887 S.t1711 SUB 0.02fF
C10888 S.n9891 SUB 0.14fF $ **FLOATING
C10889 S.n9893 SUB 1.88fF $ **FLOATING
C10890 S.n9894 SUB 2.67fF $ **FLOATING
C10891 S.t968 SUB 0.02fF
C10892 S.n9895 SUB 0.24fF $ **FLOATING
C10893 S.n9896 SUB 0.36fF $ **FLOATING
C10894 S.n9897 SUB 0.61fF $ **FLOATING
C10895 S.t102 SUB 0.02fF
C10896 S.n9898 SUB 0.24fF $ **FLOATING
C10897 S.n9899 SUB 0.91fF $ **FLOATING
C10898 S.n9900 SUB 0.05fF $ **FLOATING
C10899 S.t1471 SUB 0.02fF
C10900 S.n9901 SUB 0.12fF $ **FLOATING
C10901 S.n9902 SUB 0.14fF $ **FLOATING
C10902 S.n9904 SUB 0.12fF $ **FLOATING
C10903 S.t663 SUB 0.02fF
C10904 S.n9905 SUB 0.14fF $ **FLOATING
C10905 S.n9907 SUB 2.30fF $ **FLOATING
C10906 S.n9908 SUB 2.94fF $ **FLOATING
C10907 S.n9909 SUB 5.16fF $ **FLOATING
C10908 S.t1794 SUB 0.02fF
C10909 S.n9910 SUB 0.12fF $ **FLOATING
C10910 S.n9911 SUB 0.14fF $ **FLOATING
C10911 S.t583 SUB 0.02fF
C10912 S.n9913 SUB 0.24fF $ **FLOATING
C10913 S.n9914 SUB 0.91fF $ **FLOATING
C10914 S.n9915 SUB 0.05fF $ **FLOATING
C10915 S.n9916 SUB 1.88fF $ **FLOATING
C10916 S.n9917 SUB 2.67fF $ **FLOATING
C10917 S.t1113 SUB 0.02fF
C10918 S.n9918 SUB 0.24fF $ **FLOATING
C10919 S.n9919 SUB 0.36fF $ **FLOATING
C10920 S.n9920 SUB 0.61fF $ **FLOATING
C10921 S.n9921 SUB 0.12fF $ **FLOATING
C10922 S.t838 SUB 0.02fF
C10923 S.n9922 SUB 0.14fF $ **FLOATING
C10924 S.n9924 SUB 5.17fF $ **FLOATING
C10925 S.t1064 SUB 0.02fF
C10926 S.n9925 SUB 0.12fF $ **FLOATING
C10927 S.n9926 SUB 0.14fF $ **FLOATING
C10928 S.t2230 SUB 0.02fF
C10929 S.n9928 SUB 0.24fF $ **FLOATING
C10930 S.n9929 SUB 0.91fF $ **FLOATING
C10931 S.n9930 SUB 0.05fF $ **FLOATING
C10932 S.n9931 SUB 1.88fF $ **FLOATING
C10933 S.n9932 SUB 2.67fF $ **FLOATING
C10934 S.t542 SUB 0.02fF
C10935 S.n9933 SUB 0.24fF $ **FLOATING
C10936 S.n9934 SUB 0.36fF $ **FLOATING
C10937 S.n9935 SUB 0.61fF $ **FLOATING
C10938 S.n9936 SUB 0.12fF $ **FLOATING
C10939 S.t1617 SUB 0.02fF
C10940 S.n9937 SUB 0.14fF $ **FLOATING
C10941 S.n9939 SUB 5.17fF $ **FLOATING
C10942 S.t1862 SUB 0.02fF
C10943 S.n9940 SUB 0.12fF $ **FLOATING
C10944 S.n9941 SUB 0.14fF $ **FLOATING
C10945 S.t2085 SUB 0.02fF
C10946 S.n9943 SUB 0.24fF $ **FLOATING
C10947 S.n9944 SUB 0.91fF $ **FLOATING
C10948 S.n9945 SUB 0.05fF $ **FLOATING
C10949 S.n9946 SUB 1.88fF $ **FLOATING
C10950 S.n9947 SUB 2.67fF $ **FLOATING
C10951 S.t2187 SUB 0.02fF
C10952 S.n9948 SUB 0.24fF $ **FLOATING
C10953 S.n9949 SUB 0.36fF $ **FLOATING
C10954 S.n9950 SUB 0.61fF $ **FLOATING
C10955 S.n9951 SUB 0.12fF $ **FLOATING
C10956 S.t751 SUB 0.02fF
C10957 S.n9952 SUB 0.14fF $ **FLOATING
C10958 S.n9954 SUB 5.17fF $ **FLOATING
C10959 S.t993 SUB 0.02fF
C10960 S.n9955 SUB 0.12fF $ **FLOATING
C10961 S.n9956 SUB 0.14fF $ **FLOATING
C10962 S.t1225 SUB 0.02fF
C10963 S.n9958 SUB 0.24fF $ **FLOATING
C10964 S.n9959 SUB 0.91fF $ **FLOATING
C10965 S.n9960 SUB 0.05fF $ **FLOATING
C10966 S.n9961 SUB 1.88fF $ **FLOATING
C10967 S.n9962 SUB 2.67fF $ **FLOATING
C10968 S.t1322 SUB 0.02fF
C10969 S.n9963 SUB 0.24fF $ **FLOATING
C10970 S.n9964 SUB 0.36fF $ **FLOATING
C10971 S.n9965 SUB 0.61fF $ **FLOATING
C10972 S.n9966 SUB 0.12fF $ **FLOATING
C10973 S.t2407 SUB 0.02fF
C10974 S.n9967 SUB 0.14fF $ **FLOATING
C10975 S.n9969 SUB 5.17fF $ **FLOATING
C10976 S.t87 SUB 0.02fF
C10977 S.n9970 SUB 0.12fF $ **FLOATING
C10978 S.n9971 SUB 0.14fF $ **FLOATING
C10979 S.t342 SUB 0.02fF
C10980 S.n9973 SUB 0.24fF $ **FLOATING
C10981 S.n9974 SUB 0.91fF $ **FLOATING
C10982 S.n9975 SUB 0.05fF $ **FLOATING
C10983 S.n9976 SUB 1.88fF $ **FLOATING
C10984 S.n9977 SUB 2.67fF $ **FLOATING
C10985 S.t442 SUB 0.02fF
C10986 S.n9978 SUB 0.24fF $ **FLOATING
C10987 S.n9979 SUB 0.36fF $ **FLOATING
C10988 S.n9980 SUB 0.61fF $ **FLOATING
C10989 S.n9981 SUB 0.12fF $ **FLOATING
C10990 S.t1545 SUB 0.02fF
C10991 S.n9982 SUB 0.14fF $ **FLOATING
C10992 S.n9984 SUB 5.17fF $ **FLOATING
C10993 S.t1764 SUB 0.02fF
C10994 S.n9985 SUB 0.12fF $ **FLOATING
C10995 S.n9986 SUB 0.14fF $ **FLOATING
C10996 S.t2001 SUB 0.02fF
C10997 S.n9988 SUB 0.24fF $ **FLOATING
C10998 S.n9989 SUB 0.91fF $ **FLOATING
C10999 S.n9990 SUB 0.05fF $ **FLOATING
C11000 S.n9991 SUB 1.88fF $ **FLOATING
C11001 S.n9992 SUB 2.67fF $ **FLOATING
C11002 S.t2233 SUB 0.02fF
C11003 S.n9993 SUB 0.24fF $ **FLOATING
C11004 S.n9994 SUB 0.36fF $ **FLOATING
C11005 S.n9995 SUB 0.61fF $ **FLOATING
C11006 S.n9996 SUB 0.12fF $ **FLOATING
C11007 S.t806 SUB 0.02fF
C11008 S.n9997 SUB 0.14fF $ **FLOATING
C11009 S.n9999 SUB 5.17fF $ **FLOATING
C11010 S.t889 SUB 0.02fF
C11011 S.n10000 SUB 0.12fF $ **FLOATING
C11012 S.n10001 SUB 0.14fF $ **FLOATING
C11013 S.t1278 SUB 0.02fF
C11014 S.n10003 SUB 0.24fF $ **FLOATING
C11015 S.n10004 SUB 0.91fF $ **FLOATING
C11016 S.n10005 SUB 0.05fF $ **FLOATING
C11017 S.n10006 SUB 1.88fF $ **FLOATING
C11018 S.n10007 SUB 2.67fF $ **FLOATING
C11019 S.t1371 SUB 0.02fF
C11020 S.n10008 SUB 0.24fF $ **FLOATING
C11021 S.n10009 SUB 0.36fF $ **FLOATING
C11022 S.n10010 SUB 0.61fF $ **FLOATING
C11023 S.n10011 SUB 0.12fF $ **FLOATING
C11024 S.t2455 SUB 0.02fF
C11025 S.n10012 SUB 0.14fF $ **FLOATING
C11026 S.n10014 SUB 5.17fF $ **FLOATING
C11027 S.t2531 SUB 0.02fF
C11028 S.n10015 SUB 0.12fF $ **FLOATING
C11029 S.n10016 SUB 0.14fF $ **FLOATING
C11030 S.t394 SUB 0.02fF
C11031 S.n10018 SUB 0.24fF $ **FLOATING
C11032 S.n10019 SUB 0.91fF $ **FLOATING
C11033 S.n10020 SUB 0.05fF $ **FLOATING
C11034 S.n10021 SUB 1.88fF $ **FLOATING
C11035 S.n10022 SUB 2.67fF $ **FLOATING
C11036 S.t498 SUB 0.02fF
C11037 S.n10023 SUB 0.24fF $ **FLOATING
C11038 S.n10024 SUB 0.36fF $ **FLOATING
C11039 S.n10025 SUB 0.61fF $ **FLOATING
C11040 S.n10026 SUB 0.12fF $ **FLOATING
C11041 S.t1586 SUB 0.02fF
C11042 S.n10027 SUB 0.14fF $ **FLOATING
C11043 S.n10029 SUB 5.17fF $ **FLOATING
C11044 S.t1658 SUB 0.02fF
C11045 S.n10030 SUB 0.12fF $ **FLOATING
C11046 S.n10031 SUB 0.14fF $ **FLOATING
C11047 S.t2044 SUB 0.02fF
C11048 S.n10033 SUB 0.24fF $ **FLOATING
C11049 S.n10034 SUB 0.91fF $ **FLOATING
C11050 S.n10035 SUB 0.05fF $ **FLOATING
C11051 S.n10036 SUB 1.88fF $ **FLOATING
C11052 S.n10037 SUB 2.67fF $ **FLOATING
C11053 S.t2144 SUB 0.02fF
C11054 S.n10038 SUB 0.24fF $ **FLOATING
C11055 S.n10039 SUB 0.36fF $ **FLOATING
C11056 S.n10040 SUB 0.61fF $ **FLOATING
C11057 S.n10041 SUB 0.12fF $ **FLOATING
C11058 S.t721 SUB 0.02fF
C11059 S.n10042 SUB 0.14fF $ **FLOATING
C11060 S.n10044 SUB 4.90fF $ **FLOATING
C11061 S.t789 SUB 0.02fF
C11062 S.n10045 SUB 0.12fF $ **FLOATING
C11063 S.n10046 SUB 0.14fF $ **FLOATING
C11064 S.t1188 SUB 0.02fF
C11065 S.n10048 SUB 0.24fF $ **FLOATING
C11066 S.n10049 SUB 0.91fF $ **FLOATING
C11067 S.n10050 SUB 0.05fF $ **FLOATING
C11068 S.n10051 SUB 1.88fF $ **FLOATING
C11069 S.n10052 SUB 2.67fF $ **FLOATING
C11070 S.t1130 SUB 0.02fF
C11071 S.n10053 SUB 0.24fF $ **FLOATING
C11072 S.n10054 SUB 0.36fF $ **FLOATING
C11073 S.n10055 SUB 0.61fF $ **FLOATING
C11074 S.n10056 SUB 0.12fF $ **FLOATING
C11075 S.t485 SUB 0.02fF
C11076 S.n10057 SUB 0.14fF $ **FLOATING
C11077 S.n10059 SUB 1.88fF $ **FLOATING
C11078 S.n10060 SUB 2.68fF $ **FLOATING
C11079 S.t151 SUB 0.02fF
C11080 S.n10061 SUB 0.24fF $ **FLOATING
C11081 S.n10062 SUB 0.36fF $ **FLOATING
C11082 S.n10063 SUB 0.61fF $ **FLOATING
C11083 S.t1128 SUB 0.02fF
C11084 S.n10064 SUB 1.22fF $ **FLOATING
C11085 S.n10065 SUB 0.36fF $ **FLOATING
C11086 S.n10066 SUB 1.22fF $ **FLOATING
C11087 S.n10067 SUB 0.61fF $ **FLOATING
C11088 S.n10068 SUB 0.35fF $ **FLOATING
C11089 S.n10069 SUB 0.63fF $ **FLOATING
C11090 S.n10070 SUB 1.15fF $ **FLOATING
C11091 S.n10071 SUB 3.03fF $ **FLOATING
C11092 S.n10072 SUB 0.59fF $ **FLOATING
C11093 S.n10073 SUB 0.02fF $ **FLOATING
C11094 S.n10074 SUB 0.97fF $ **FLOATING
C11095 S.t30 SUB 21.38fF
C11096 S.n10075 SUB 20.25fF $ **FLOATING
C11097 S.n10077 SUB 0.38fF $ **FLOATING
C11098 S.n10078 SUB 0.23fF $ **FLOATING
C11099 S.n10079 SUB 2.79fF $ **FLOATING
C11100 S.n10080 SUB 2.46fF $ **FLOATING
C11101 S.n10081 SUB 4.00fF $ **FLOATING
C11102 S.n10082 SUB 0.25fF $ **FLOATING
C11103 S.n10083 SUB 0.01fF $ **FLOATING
C11104 S.t812 SUB 0.02fF
C11105 S.n10084 SUB 0.25fF $ **FLOATING
C11106 S.t281 SUB 0.02fF
C11107 S.n10085 SUB 0.95fF $ **FLOATING
C11108 S.n10086 SUB 0.70fF $ **FLOATING
C11109 S.n10087 SUB 1.89fF $ **FLOATING
C11110 S.n10088 SUB 1.73fF $ **FLOATING
C11111 S.t250 SUB 0.02fF
C11112 S.n10089 SUB 0.24fF $ **FLOATING
C11113 S.n10090 SUB 0.36fF $ **FLOATING
C11114 S.n10091 SUB 0.61fF $ **FLOATING
C11115 S.n10092 SUB 0.12fF $ **FLOATING
C11116 S.t2460 SUB 0.02fF
C11117 S.n10093 SUB 0.14fF $ **FLOATING
C11118 S.n10095 SUB 1.16fF $ **FLOATING
C11119 S.n10096 SUB 0.22fF $ **FLOATING
C11120 S.n10097 SUB 0.25fF $ **FLOATING
C11121 S.n10098 SUB 0.09fF $ **FLOATING
C11122 S.n10099 SUB 2.44fF $ **FLOATING
C11123 S.t1940 SUB 0.02fF
C11124 S.n10100 SUB 0.24fF $ **FLOATING
C11125 S.n10101 SUB 0.91fF $ **FLOATING
C11126 S.n10102 SUB 0.05fF $ **FLOATING
C11127 S.t638 SUB 0.02fF
C11128 S.n10103 SUB 0.12fF $ **FLOATING
C11129 S.n10104 SUB 0.14fF $ **FLOATING
C11130 S.n10106 SUB 1.88fF $ **FLOATING
C11131 S.n10107 SUB 0.48fF $ **FLOATING
C11132 S.n10108 SUB 0.09fF $ **FLOATING
C11133 S.n10109 SUB 0.33fF $ **FLOATING
C11134 S.n10110 SUB 0.30fF $ **FLOATING
C11135 S.n10111 SUB 0.77fF $ **FLOATING
C11136 S.n10112 SUB 0.59fF $ **FLOATING
C11137 S.t1916 SUB 0.02fF
C11138 S.n10113 SUB 0.24fF $ **FLOATING
C11139 S.n10114 SUB 0.36fF $ **FLOATING
C11140 S.n10115 SUB 0.61fF $ **FLOATING
C11141 S.n10116 SUB 0.12fF $ **FLOATING
C11142 S.t1592 SUB 0.02fF
C11143 S.n10117 SUB 0.14fF $ **FLOATING
C11144 S.n10119 SUB 2.61fF $ **FLOATING
C11145 S.n10120 SUB 2.16fF $ **FLOATING
C11146 S.t1080 SUB 0.02fF
C11147 S.n10121 SUB 0.24fF $ **FLOATING
C11148 S.n10122 SUB 0.91fF $ **FLOATING
C11149 S.n10123 SUB 0.05fF $ **FLOATING
C11150 S.t2295 SUB 0.02fF
C11151 S.n10124 SUB 0.12fF $ **FLOATING
C11152 S.n10125 SUB 0.14fF $ **FLOATING
C11153 S.n10127 SUB 0.78fF $ **FLOATING
C11154 S.n10128 SUB 2.30fF $ **FLOATING
C11155 S.n10129 SUB 1.88fF $ **FLOATING
C11156 S.n10130 SUB 0.12fF $ **FLOATING
C11157 S.t728 SUB 0.02fF
C11158 S.n10131 SUB 0.14fF $ **FLOATING
C11159 S.t1056 SUB 0.02fF
C11160 S.n10133 SUB 0.24fF $ **FLOATING
C11161 S.n10134 SUB 0.36fF $ **FLOATING
C11162 S.n10135 SUB 0.61fF $ **FLOATING
C11163 S.n10136 SUB 1.39fF $ **FLOATING
C11164 S.n10137 SUB 0.71fF $ **FLOATING
C11165 S.n10138 SUB 1.14fF $ **FLOATING
C11166 S.n10139 SUB 0.35fF $ **FLOATING
C11167 S.n10140 SUB 2.03fF $ **FLOATING
C11168 S.t204 SUB 0.02fF
C11169 S.n10141 SUB 0.24fF $ **FLOATING
C11170 S.n10142 SUB 0.91fF $ **FLOATING
C11171 S.n10143 SUB 0.05fF $ **FLOATING
C11172 S.t1533 SUB 0.02fF
C11173 S.n10144 SUB 0.12fF $ **FLOATING
C11174 S.n10145 SUB 0.14fF $ **FLOATING
C11175 S.n10147 SUB 1.89fF $ **FLOATING
C11176 S.n10148 SUB 1.88fF $ **FLOATING
C11177 S.t170 SUB 0.02fF
C11178 S.n10149 SUB 0.24fF $ **FLOATING
C11179 S.n10150 SUB 0.36fF $ **FLOATING
C11180 S.n10151 SUB 0.61fF $ **FLOATING
C11181 S.n10152 SUB 0.12fF $ **FLOATING
C11182 S.t2380 SUB 0.02fF
C11183 S.n10153 SUB 0.14fF $ **FLOATING
C11184 S.n10155 SUB 1.16fF $ **FLOATING
C11185 S.n10156 SUB 0.22fF $ **FLOATING
C11186 S.n10157 SUB 0.25fF $ **FLOATING
C11187 S.n10158 SUB 0.09fF $ **FLOATING
C11188 S.n10159 SUB 1.88fF $ **FLOATING
C11189 S.t1872 SUB 0.02fF
C11190 S.n10160 SUB 0.24fF $ **FLOATING
C11191 S.n10161 SUB 0.91fF $ **FLOATING
C11192 S.n10162 SUB 0.05fF $ **FLOATING
C11193 S.t673 SUB 0.02fF
C11194 S.n10163 SUB 0.12fF $ **FLOATING
C11195 S.n10164 SUB 0.14fF $ **FLOATING
C11196 S.n10166 SUB 20.78fF $ **FLOATING
C11197 S.n10167 SUB 1.88fF $ **FLOATING
C11198 S.n10168 SUB 2.67fF $ **FLOATING
C11199 S.t31 SUB 0.02fF
C11200 S.n10169 SUB 0.24fF $ **FLOATING
C11201 S.n10170 SUB 0.36fF $ **FLOATING
C11202 S.n10171 SUB 0.61fF $ **FLOATING
C11203 S.n10172 SUB 0.12fF $ **FLOATING
C11204 S.t2419 SUB 0.02fF
C11205 S.n10173 SUB 0.14fF $ **FLOATING
C11206 S.n10175 SUB 2.80fF $ **FLOATING
C11207 S.n10176 SUB 2.30fF $ **FLOATING
C11208 S.t609 SUB 0.02fF
C11209 S.n10177 SUB 0.12fF $ **FLOATING
C11210 S.n10178 SUB 0.14fF $ **FLOATING
C11211 S.t1777 SUB 0.02fF
C11212 S.n10180 SUB 0.24fF $ **FLOATING
C11213 S.n10181 SUB 0.91fF $ **FLOATING
C11214 S.n10182 SUB 0.05fF $ **FLOATING
C11215 S.n10183 SUB 1.88fF $ **FLOATING
C11216 S.n10184 SUB 2.67fF $ **FLOATING
C11217 S.t2037 SUB 0.02fF
C11218 S.n10185 SUB 0.24fF $ **FLOATING
C11219 S.n10186 SUB 0.36fF $ **FLOATING
C11220 S.n10187 SUB 0.61fF $ **FLOATING
C11221 S.n10188 SUB 0.12fF $ **FLOATING
C11222 S.t270 SUB 0.02fF
C11223 S.n10189 SUB 0.14fF $ **FLOATING
C11224 S.n10191 SUB 2.80fF $ **FLOATING
C11225 S.n10192 SUB 2.30fF $ **FLOATING
C11226 S.t2262 SUB 0.02fF
C11227 S.n10193 SUB 0.12fF $ **FLOATING
C11228 S.n10194 SUB 0.14fF $ **FLOATING
C11229 S.t1342 SUB 0.02fF
C11230 S.n10196 SUB 0.24fF $ **FLOATING
C11231 S.n10197 SUB 0.91fF $ **FLOATING
C11232 S.n10198 SUB 0.05fF $ **FLOATING
C11233 S.n10199 SUB 1.88fF $ **FLOATING
C11234 S.n10200 SUB 2.67fF $ **FLOATING
C11235 S.t1182 SUB 0.02fF
C11236 S.n10201 SUB 0.24fF $ **FLOATING
C11237 S.n10202 SUB 0.36fF $ **FLOATING
C11238 S.n10203 SUB 0.61fF $ **FLOATING
C11239 S.n10204 SUB 0.12fF $ **FLOATING
C11240 S.t1931 SUB 0.02fF
C11241 S.n10205 SUB 0.14fF $ **FLOATING
C11242 S.n10207 SUB 2.80fF $ **FLOATING
C11243 S.n10208 SUB 2.30fF $ **FLOATING
C11244 S.t17 SUB 0.02fF
C11245 S.n10209 SUB 0.12fF $ **FLOATING
C11246 S.n10210 SUB 0.14fF $ **FLOATING
C11247 S.t464 SUB 0.02fF
C11248 S.n10212 SUB 0.24fF $ **FLOATING
C11249 S.n10213 SUB 0.91fF $ **FLOATING
C11250 S.n10214 SUB 0.05fF $ **FLOATING
C11251 S.n10215 SUB 1.88fF $ **FLOATING
C11252 S.n10216 SUB 2.67fF $ **FLOATING
C11253 S.t306 SUB 0.02fF
C11254 S.n10217 SUB 0.24fF $ **FLOATING
C11255 S.n10218 SUB 0.36fF $ **FLOATING
C11256 S.n10219 SUB 0.61fF $ **FLOATING
C11257 S.n10220 SUB 0.12fF $ **FLOATING
C11258 S.t1073 SUB 0.02fF
C11259 S.n10221 SUB 0.14fF $ **FLOATING
C11260 S.n10223 SUB 2.80fF $ **FLOATING
C11261 S.n10224 SUB 2.30fF $ **FLOATING
C11262 S.t1725 SUB 0.02fF
C11263 S.n10225 SUB 0.12fF $ **FLOATING
C11264 S.n10226 SUB 0.14fF $ **FLOATING
C11265 S.t2109 SUB 0.02fF
C11266 S.n10228 SUB 0.24fF $ **FLOATING
C11267 S.n10229 SUB 0.91fF $ **FLOATING
C11268 S.n10230 SUB 0.05fF $ **FLOATING
C11269 S.n10231 SUB 1.88fF $ **FLOATING
C11270 S.n10232 SUB 2.67fF $ **FLOATING
C11271 S.t1969 SUB 0.02fF
C11272 S.n10233 SUB 0.24fF $ **FLOATING
C11273 S.n10234 SUB 0.36fF $ **FLOATING
C11274 S.n10235 SUB 0.61fF $ **FLOATING
C11275 S.n10236 SUB 0.12fF $ **FLOATING
C11276 S.t196 SUB 0.02fF
C11277 S.n10237 SUB 0.14fF $ **FLOATING
C11278 S.n10239 SUB 2.80fF $ **FLOATING
C11279 S.n10240 SUB 2.30fF $ **FLOATING
C11280 S.t853 SUB 0.02fF
C11281 S.n10241 SUB 0.12fF $ **FLOATING
C11282 S.n10242 SUB 0.14fF $ **FLOATING
C11283 S.t1244 SUB 0.02fF
C11284 S.n10244 SUB 0.24fF $ **FLOATING
C11285 S.n10245 SUB 0.91fF $ **FLOATING
C11286 S.n10246 SUB 0.05fF $ **FLOATING
C11287 S.n10247 SUB 1.88fF $ **FLOATING
C11288 S.n10248 SUB 2.67fF $ **FLOATING
C11289 S.t1114 SUB 0.02fF
C11290 S.n10249 SUB 0.24fF $ **FLOATING
C11291 S.n10250 SUB 0.36fF $ **FLOATING
C11292 S.n10251 SUB 0.61fF $ **FLOATING
C11293 S.n10252 SUB 0.12fF $ **FLOATING
C11294 S.t1864 SUB 0.02fF
C11295 S.n10253 SUB 0.14fF $ **FLOATING
C11296 S.n10255 SUB 2.80fF $ **FLOATING
C11297 S.n10256 SUB 2.30fF $ **FLOATING
C11298 S.t2495 SUB 0.02fF
C11299 S.n10257 SUB 0.12fF $ **FLOATING
C11300 S.n10258 SUB 0.14fF $ **FLOATING
C11301 S.t362 SUB 0.02fF
C11302 S.n10260 SUB 0.24fF $ **FLOATING
C11303 S.n10261 SUB 0.91fF $ **FLOATING
C11304 S.n10262 SUB 0.05fF $ **FLOATING
C11305 S.n10263 SUB 1.88fF $ **FLOATING
C11306 S.n10264 SUB 2.67fF $ **FLOATING
C11307 S.t236 SUB 0.02fF
C11308 S.n10265 SUB 0.24fF $ **FLOATING
C11309 S.n10266 SUB 0.36fF $ **FLOATING
C11310 S.n10267 SUB 0.61fF $ **FLOATING
C11311 S.n10268 SUB 0.12fF $ **FLOATING
C11312 S.t995 SUB 0.02fF
C11313 S.n10269 SUB 0.14fF $ **FLOATING
C11314 S.n10271 SUB 2.80fF $ **FLOATING
C11315 S.n10272 SUB 2.30fF $ **FLOATING
C11316 S.t1782 SUB 0.02fF
C11317 S.n10273 SUB 0.12fF $ **FLOATING
C11318 S.n10274 SUB 0.14fF $ **FLOATING
C11319 S.t2014 SUB 0.02fF
C11320 S.n10276 SUB 0.24fF $ **FLOATING
C11321 S.n10277 SUB 0.91fF $ **FLOATING
C11322 S.n10278 SUB 0.05fF $ **FLOATING
C11323 S.n10279 SUB 1.88fF $ **FLOATING
C11324 S.n10280 SUB 2.67fF $ **FLOATING
C11325 S.t1903 SUB 0.02fF
C11326 S.n10281 SUB 0.24fF $ **FLOATING
C11327 S.n10282 SUB 0.36fF $ **FLOATING
C11328 S.n10283 SUB 0.61fF $ **FLOATING
C11329 S.n10284 SUB 0.12fF $ **FLOATING
C11330 S.t88 SUB 0.02fF
C11331 S.n10285 SUB 0.14fF $ **FLOATING
C11332 S.n10287 SUB 2.80fF $ **FLOATING
C11333 S.n10288 SUB 2.30fF $ **FLOATING
C11334 S.t910 SUB 0.02fF
C11335 S.n10289 SUB 0.12fF $ **FLOATING
C11336 S.n10290 SUB 0.14fF $ **FLOATING
C11337 S.t1161 SUB 0.02fF
C11338 S.n10292 SUB 0.24fF $ **FLOATING
C11339 S.n10293 SUB 0.91fF $ **FLOATING
C11340 S.n10294 SUB 0.05fF $ **FLOATING
C11341 S.n10295 SUB 1.88fF $ **FLOATING
C11342 S.n10296 SUB 2.67fF $ **FLOATING
C11343 S.t1044 SUB 0.02fF
C11344 S.n10297 SUB 0.24fF $ **FLOATING
C11345 S.n10298 SUB 0.36fF $ **FLOATING
C11346 S.n10299 SUB 0.61fF $ **FLOATING
C11347 S.n10300 SUB 0.12fF $ **FLOATING
C11348 S.t1766 SUB 0.02fF
C11349 S.n10301 SUB 0.14fF $ **FLOATING
C11350 S.n10303 SUB 2.80fF $ **FLOATING
C11351 S.n10304 SUB 2.30fF $ **FLOATING
C11352 S.t2551 SUB 0.02fF
C11353 S.n10305 SUB 0.12fF $ **FLOATING
C11354 S.n10306 SUB 0.14fF $ **FLOATING
C11355 S.t289 SUB 0.02fF
C11356 S.n10308 SUB 0.24fF $ **FLOATING
C11357 S.n10309 SUB 0.91fF $ **FLOATING
C11358 S.n10310 SUB 0.05fF $ **FLOATING
C11359 S.n10311 SUB 2.73fF $ **FLOATING
C11360 S.n10312 SUB 1.59fF $ **FLOATING
C11361 S.n10313 SUB 0.12fF $ **FLOATING
C11362 S.t302 SUB 0.02fF
C11363 S.n10314 SUB 0.14fF $ **FLOATING
C11364 S.t1568 SUB 0.02fF
C11365 S.n10316 SUB 0.24fF $ **FLOATING
C11366 S.n10317 SUB 0.36fF $ **FLOATING
C11367 S.n10318 SUB 0.61fF $ **FLOATING
C11368 S.n10319 SUB 0.07fF $ **FLOATING
C11369 S.n10320 SUB 0.01fF $ **FLOATING
C11370 S.n10321 SUB 0.24fF $ **FLOATING
C11371 S.n10322 SUB 1.16fF $ **FLOATING
C11372 S.n10323 SUB 1.35fF $ **FLOATING
C11373 S.n10324 SUB 2.30fF $ **FLOATING
C11374 S.t1076 SUB 0.02fF
C11375 S.n10325 SUB 0.12fF $ **FLOATING
C11376 S.n10326 SUB 0.14fF $ **FLOATING
C11377 S.t2560 SUB 0.02fF
C11378 S.n10328 SUB 0.24fF $ **FLOATING
C11379 S.n10329 SUB 0.91fF $ **FLOATING
C11380 S.n10330 SUB 0.05fF $ **FLOATING
C11381 S.t16 SUB 48.31fF
C11382 S.t1950 SUB 0.02fF
C11383 S.n10331 SUB 0.24fF $ **FLOATING
C11384 S.n10332 SUB 0.91fF $ **FLOATING
C11385 S.n10333 SUB 0.05fF $ **FLOATING
C11386 S.t1681 SUB 0.02fF
C11387 S.n10334 SUB 0.12fF $ **FLOATING
C11388 S.n10335 SUB 0.14fF $ **FLOATING
C11389 S.n10337 SUB 0.12fF $ **FLOATING
C11390 S.t892 SUB 0.02fF
C11391 S.n10338 SUB 0.14fF $ **FLOATING
C11392 S.n10340 SUB 5.17fF $ **FLOATING
C11393 S.n10341 SUB 5.44fF $ **FLOATING
C11394 S.t2439 SUB 0.02fF
C11395 S.n10342 SUB 0.12fF $ **FLOATING
C11396 S.n10343 SUB 0.14fF $ **FLOATING
C11397 S.t553 SUB 0.02fF
C11398 S.n10345 SUB 0.24fF $ **FLOATING
C11399 S.n10346 SUB 0.91fF $ **FLOATING
C11400 S.n10347 SUB 0.05fF $ **FLOATING
C11401 S.t86 SUB 47.92fF
C11402 S.t1254 SUB 0.02fF
C11403 S.n10348 SUB 1.19fF $ **FLOATING
C11404 S.n10349 SUB 0.05fF $ **FLOATING
C11405 S.t2255 SUB 0.02fF
C11406 S.n10350 SUB 0.01fF $ **FLOATING
C11407 S.n10351 SUB 0.26fF $ **FLOATING
C11408 S.n10353 SUB 1.50fF $ **FLOATING
C11409 S.n10354 SUB 1.30fF $ **FLOATING
C11410 S.n10355 SUB 0.28fF $ **FLOATING
C11411 S.n10356 SUB 0.24fF $ **FLOATING
C11412 S.n10357 SUB 4.39fF $ **FLOATING
C11413 S.n10358 SUB 0.01fF $ **FLOATING
C11414 S.n10359 SUB 0.02fF $ **FLOATING
C11415 S.n10360 SUB 0.03fF $ **FLOATING
C11416 S.n10361 SUB 0.04fF $ **FLOATING
C11417 S.n10362 SUB 0.17fF $ **FLOATING
C11418 S.n10363 SUB 0.01fF $ **FLOATING
C11419 S.n10364 SUB 0.02fF $ **FLOATING
C11420 S.n10365 SUB 0.01fF $ **FLOATING
C11421 S.n10366 SUB 0.01fF $ **FLOATING
C11422 S.n10367 SUB 0.01fF $ **FLOATING
C11423 S.n10368 SUB 0.01fF $ **FLOATING
C11424 S.n10369 SUB 0.02fF $ **FLOATING
C11425 S.n10370 SUB 0.01fF $ **FLOATING
C11426 S.n10371 SUB 0.02fF $ **FLOATING
C11427 S.n10372 SUB 0.05fF $ **FLOATING
C11428 S.n10373 SUB 0.04fF $ **FLOATING
C11429 S.n10374 SUB 0.11fF $ **FLOATING
C11430 S.n10375 SUB 0.38fF $ **FLOATING
C11431 S.n10376 SUB 0.20fF $ **FLOATING
C11432 S.n10377 SUB 8.97fF $ **FLOATING
C11433 S.n10378 SUB 8.97fF $ **FLOATING
C11434 S.n10379 SUB 0.60fF $ **FLOATING
C11435 S.n10380 SUB 0.22fF $ **FLOATING
C11436 S.n10381 SUB 0.59fF $ **FLOATING
C11437 S.n10382 SUB 3.43fF $ **FLOATING
C11438 S.n10383 SUB 0.29fF $ **FLOATING
C11439 S.t91 SUB 21.38fF
C11440 S.n10384 SUB 21.67fF $ **FLOATING
C11441 S.n10385 SUB 0.77fF $ **FLOATING
C11442 S.n10386 SUB 0.28fF $ **FLOATING
C11443 S.n10387 SUB 4.00fF $ **FLOATING
C11444 S.n10388 SUB 1.35fF $ **FLOATING
C11445 S.t1377 SUB 0.02fF
C11446 S.n10389 SUB 0.64fF $ **FLOATING
C11447 S.n10390 SUB 0.61fF $ **FLOATING
C11448 S.n10391 SUB 1.88fF $ **FLOATING
C11449 S.n10392 SUB 0.46fF $ **FLOATING
C11450 S.n10393 SUB 0.22fF $ **FLOATING
C11451 S.n10394 SUB 0.38fF $ **FLOATING
C11452 S.n10395 SUB 0.16fF $ **FLOATING
C11453 S.n10396 SUB 0.28fF $ **FLOATING
C11454 S.n10397 SUB 0.21fF $ **FLOATING
C11455 S.n10398 SUB 0.30fF $ **FLOATING
C11456 S.n10399 SUB 0.42fF $ **FLOATING
C11457 S.n10400 SUB 0.21fF $ **FLOATING
C11458 S.t837 SUB 0.02fF
C11459 S.n10401 SUB 0.24fF $ **FLOATING
C11460 S.n10402 SUB 0.36fF $ **FLOATING
C11461 S.n10403 SUB 0.61fF $ **FLOATING
C11462 S.n10404 SUB 0.12fF $ **FLOATING
C11463 S.t311 SUB 0.02fF
C11464 S.n10405 SUB 0.14fF $ **FLOATING
C11465 S.n10407 SUB 0.04fF $ **FLOATING
C11466 S.n10408 SUB 0.03fF $ **FLOATING
C11467 S.n10409 SUB 0.03fF $ **FLOATING
C11468 S.n10410 SUB 0.10fF $ **FLOATING
C11469 S.n10411 SUB 0.36fF $ **FLOATING
C11470 S.n10412 SUB 0.38fF $ **FLOATING
C11471 S.n10413 SUB 0.11fF $ **FLOATING
C11472 S.n10414 SUB 0.12fF $ **FLOATING
C11473 S.n10415 SUB 0.07fF $ **FLOATING
C11474 S.n10416 SUB 0.12fF $ **FLOATING
C11475 S.n10417 SUB 0.18fF $ **FLOATING
C11476 S.n10418 SUB 4.00fF $ **FLOATING
C11477 S.t1970 SUB 0.02fF
C11478 S.n10419 SUB 0.24fF $ **FLOATING
C11479 S.n10420 SUB 0.91fF $ **FLOATING
C11480 S.n10421 SUB 0.05fF $ **FLOATING
C11481 S.t530 SUB 0.02fF
C11482 S.n10422 SUB 0.12fF $ **FLOATING
C11483 S.n10423 SUB 0.14fF $ **FLOATING
C11484 S.n10425 SUB 0.25fF $ **FLOATING
C11485 S.n10426 SUB 0.09fF $ **FLOATING
C11486 S.n10427 SUB 0.21fF $ **FLOATING
C11487 S.n10428 SUB 1.28fF $ **FLOATING
C11488 S.n10429 SUB 0.53fF $ **FLOATING
C11489 S.n10430 SUB 1.88fF $ **FLOATING
C11490 S.n10431 SUB 0.12fF $ **FLOATING
C11491 S.t2095 SUB 0.02fF
C11492 S.n10432 SUB 0.14fF $ **FLOATING
C11493 S.t92 SUB 0.02fF
C11494 S.n10434 SUB 0.24fF $ **FLOATING
C11495 S.n10435 SUB 0.36fF $ **FLOATING
C11496 S.n10436 SUB 0.61fF $ **FLOATING
C11497 S.n10437 SUB 1.58fF $ **FLOATING
C11498 S.n10438 SUB 2.45fF $ **FLOATING
C11499 S.t1226 SUB 0.02fF
C11500 S.n10439 SUB 0.24fF $ **FLOATING
C11501 S.n10440 SUB 0.91fF $ **FLOATING
C11502 S.n10441 SUB 0.05fF $ **FLOATING
C11503 S.t2173 SUB 0.02fF
C11504 S.n10442 SUB 0.12fF $ **FLOATING
C11505 S.n10443 SUB 0.14fF $ **FLOATING
C11506 S.n10445 SUB 1.89fF $ **FLOATING
C11507 S.n10446 SUB 0.06fF $ **FLOATING
C11508 S.n10447 SUB 0.03fF $ **FLOATING
C11509 S.n10448 SUB 0.04fF $ **FLOATING
C11510 S.n10449 SUB 0.99fF $ **FLOATING
C11511 S.n10450 SUB 0.02fF $ **FLOATING
C11512 S.n10451 SUB 0.01fF $ **FLOATING
C11513 S.n10452 SUB 0.02fF $ **FLOATING
C11514 S.n10453 SUB 0.08fF $ **FLOATING
C11515 S.n10454 SUB 0.36fF $ **FLOATING
C11516 S.n10455 SUB 1.85fF $ **FLOATING
C11517 S.t1767 SUB 0.02fF
C11518 S.n10456 SUB 0.24fF $ **FLOATING
C11519 S.n10457 SUB 0.36fF $ **FLOATING
C11520 S.n10458 SUB 0.61fF $ **FLOATING
C11521 S.n10459 SUB 0.12fF $ **FLOATING
C11522 S.t1230 SUB 0.02fF
C11523 S.n10460 SUB 0.14fF $ **FLOATING
C11524 S.n10462 SUB 0.70fF $ **FLOATING
C11525 S.n10463 SUB 0.23fF $ **FLOATING
C11526 S.n10464 SUB 0.23fF $ **FLOATING
C11527 S.n10465 SUB 0.70fF $ **FLOATING
C11528 S.n10466 SUB 1.16fF $ **FLOATING
C11529 S.n10467 SUB 0.22fF $ **FLOATING
C11530 S.n10468 SUB 0.25fF $ **FLOATING
C11531 S.n10469 SUB 0.09fF $ **FLOATING
C11532 S.n10470 SUB 1.88fF $ **FLOATING
C11533 S.t343 SUB 0.02fF
C11534 S.n10471 SUB 0.24fF $ **FLOATING
C11535 S.n10472 SUB 0.91fF $ **FLOATING
C11536 S.n10473 SUB 0.05fF $ **FLOATING
C11537 S.t1310 SUB 0.02fF
C11538 S.n10474 SUB 0.12fF $ **FLOATING
C11539 S.n10475 SUB 0.14fF $ **FLOATING
C11540 S.n10477 SUB 20.78fF $ **FLOATING
C11541 S.n10478 SUB 1.72fF $ **FLOATING
C11542 S.n10479 SUB 0.66fF $ **FLOATING
C11543 S.n10480 SUB 0.69fF $ **FLOATING
C11544 S.n10481 SUB 0.72fF $ **FLOATING
C11545 S.n10482 SUB 0.36fF $ **FLOATING
C11546 S.t1708 SUB 0.02fF
C11547 S.n10483 SUB 0.24fF $ **FLOATING
C11548 S.n10484 SUB 0.36fF $ **FLOATING
C11549 S.n10485 SUB 0.61fF $ **FLOATING
C11550 S.n10486 SUB 0.12fF $ **FLOATING
C11551 S.t1186 SUB 0.02fF
C11552 S.n10487 SUB 0.14fF $ **FLOATING
C11553 S.n10489 SUB 0.31fF $ **FLOATING
C11554 S.n10490 SUB 0.23fF $ **FLOATING
C11555 S.n10491 SUB 0.66fF $ **FLOATING
C11556 S.n10492 SUB 0.95fF $ **FLOATING
C11557 S.n10493 SUB 0.23fF $ **FLOATING
C11558 S.n10494 SUB 0.21fF $ **FLOATING
C11559 S.n10495 SUB 0.20fF $ **FLOATING
C11560 S.n10496 SUB 0.06fF $ **FLOATING
C11561 S.n10497 SUB 0.09fF $ **FLOATING
C11562 S.n10498 SUB 0.10fF $ **FLOATING
C11563 S.n10499 SUB 1.67fF $ **FLOATING
C11564 S.t1402 SUB 0.02fF
C11565 S.n10500 SUB 0.12fF $ **FLOATING
C11566 S.n10501 SUB 0.14fF $ **FLOATING
C11567 S.t305 SUB 0.02fF
C11568 S.n10503 SUB 0.24fF $ **FLOATING
C11569 S.n10504 SUB 0.91fF $ **FLOATING
C11570 S.n10505 SUB 0.05fF $ **FLOATING
C11571 S.n10506 SUB 1.88fF $ **FLOATING
C11572 S.n10507 SUB 0.12fF $ **FLOATING
C11573 S.t2122 SUB 0.02fF
C11574 S.n10508 SUB 0.14fF $ **FLOATING
C11575 S.t387 SUB 0.02fF
C11576 S.n10510 SUB 0.12fF $ **FLOATING
C11577 S.n10511 SUB 0.14fF $ **FLOATING
C11578 S.t1546 SUB 0.02fF
C11579 S.n10513 SUB 0.24fF $ **FLOATING
C11580 S.n10514 SUB 0.91fF $ **FLOATING
C11581 S.n10515 SUB 0.05fF $ **FLOATING
C11582 S.t2378 SUB 0.02fF
C11583 S.n10516 SUB 0.24fF $ **FLOATING
C11584 S.n10517 SUB 0.36fF $ **FLOATING
C11585 S.n10518 SUB 0.61fF $ **FLOATING
C11586 S.n10519 SUB 0.32fF $ **FLOATING
C11587 S.n10520 SUB 1.09fF $ **FLOATING
C11588 S.n10521 SUB 0.15fF $ **FLOATING
C11589 S.n10522 SUB 2.10fF $ **FLOATING
C11590 S.n10523 SUB 2.94fF $ **FLOATING
C11591 S.n10524 SUB 1.88fF $ **FLOATING
C11592 S.n10525 SUB 0.12fF $ **FLOATING
C11593 S.t346 SUB 0.02fF
C11594 S.n10526 SUB 0.14fF $ **FLOATING
C11595 S.t893 SUB 0.02fF
C11596 S.n10528 SUB 0.24fF $ **FLOATING
C11597 S.n10529 SUB 0.36fF $ **FLOATING
C11598 S.n10530 SUB 0.61fF $ **FLOATING
C11599 S.n10531 SUB 0.92fF $ **FLOATING
C11600 S.n10532 SUB 0.32fF $ **FLOATING
C11601 S.n10533 SUB 0.92fF $ **FLOATING
C11602 S.n10534 SUB 1.09fF $ **FLOATING
C11603 S.n10535 SUB 0.15fF $ **FLOATING
C11604 S.n10536 SUB 4.96fF $ **FLOATING
C11605 S.t428 SUB 0.02fF
C11606 S.n10537 SUB 0.12fF $ **FLOATING
C11607 S.n10538 SUB 0.14fF $ **FLOATING
C11608 S.t2002 SUB 0.02fF
C11609 S.n10540 SUB 0.24fF $ **FLOATING
C11610 S.n10541 SUB 0.91fF $ **FLOATING
C11611 S.n10542 SUB 0.05fF $ **FLOATING
C11612 S.n10543 SUB 1.88fF $ **FLOATING
C11613 S.n10544 SUB 2.67fF $ **FLOATING
C11614 S.t2535 SUB 0.02fF
C11615 S.n10545 SUB 0.24fF $ **FLOATING
C11616 S.n10546 SUB 0.36fF $ **FLOATING
C11617 S.n10547 SUB 0.61fF $ **FLOATING
C11618 S.n10548 SUB 0.12fF $ **FLOATING
C11619 S.t2004 SUB 0.02fF
C11620 S.n10549 SUB 0.14fF $ **FLOATING
C11621 S.n10551 SUB 1.88fF $ **FLOATING
C11622 S.n10552 SUB 2.67fF $ **FLOATING
C11623 S.t1522 SUB 0.02fF
C11624 S.n10553 SUB 0.24fF $ **FLOATING
C11625 S.n10554 SUB 0.36fF $ **FLOATING
C11626 S.n10555 SUB 0.61fF $ **FLOATING
C11627 S.t684 SUB 0.02fF
C11628 S.n10556 SUB 0.24fF $ **FLOATING
C11629 S.n10557 SUB 0.91fF $ **FLOATING
C11630 S.n10558 SUB 0.05fF $ **FLOATING
C11631 S.t2036 SUB 0.02fF
C11632 S.n10559 SUB 0.12fF $ **FLOATING
C11633 S.n10560 SUB 0.14fF $ **FLOATING
C11634 S.n10562 SUB 0.12fF $ **FLOATING
C11635 S.t1255 SUB 0.02fF
C11636 S.n10563 SUB 0.14fF $ **FLOATING
C11637 S.n10565 SUB 2.30fF $ **FLOATING
C11638 S.n10566 SUB 2.94fF $ **FLOATING
C11639 S.n10567 SUB 5.16fF $ **FLOATING
C11640 S.t2077 SUB 0.02fF
C11641 S.n10568 SUB 0.12fF $ **FLOATING
C11642 S.n10569 SUB 0.14fF $ **FLOATING
C11643 S.t1150 SUB 0.02fF
C11644 S.n10571 SUB 0.24fF $ **FLOATING
C11645 S.n10572 SUB 0.91fF $ **FLOATING
C11646 S.n10573 SUB 0.05fF $ **FLOATING
C11647 S.n10574 SUB 1.88fF $ **FLOATING
C11648 S.n10575 SUB 2.67fF $ **FLOATING
C11649 S.t1661 SUB 0.02fF
C11650 S.n10576 SUB 0.24fF $ **FLOATING
C11651 S.n10577 SUB 0.36fF $ **FLOATING
C11652 S.n10578 SUB 0.61fF $ **FLOATING
C11653 S.n10579 SUB 0.12fF $ **FLOATING
C11654 S.t1153 SUB 0.02fF
C11655 S.n10580 SUB 0.14fF $ **FLOATING
C11656 S.n10582 SUB 5.17fF $ **FLOATING
C11657 S.t1215 SUB 0.02fF
C11658 S.n10583 SUB 0.12fF $ **FLOATING
C11659 S.n10584 SUB 0.14fF $ **FLOATING
C11660 S.t274 SUB 0.02fF
C11661 S.n10586 SUB 0.24fF $ **FLOATING
C11662 S.n10587 SUB 0.91fF $ **FLOATING
C11663 S.n10588 SUB 0.05fF $ **FLOATING
C11664 S.n10589 SUB 1.88fF $ **FLOATING
C11665 S.n10590 SUB 2.67fF $ **FLOATING
C11666 S.t790 SUB 0.02fF
C11667 S.n10591 SUB 0.24fF $ **FLOATING
C11668 S.n10592 SUB 0.36fF $ **FLOATING
C11669 S.n10593 SUB 0.61fF $ **FLOATING
C11670 S.n10594 SUB 0.12fF $ **FLOATING
C11671 S.t277 SUB 0.02fF
C11672 S.n10595 SUB 0.14fF $ **FLOATING
C11673 S.n10597 SUB 5.17fF $ **FLOATING
C11674 S.t486 SUB 0.02fF
C11675 S.n10598 SUB 0.12fF $ **FLOATING
C11676 S.n10599 SUB 0.14fF $ **FLOATING
C11677 S.t1937 SUB 0.02fF
C11678 S.n10601 SUB 0.24fF $ **FLOATING
C11679 S.n10602 SUB 0.91fF $ **FLOATING
C11680 S.n10603 SUB 0.05fF $ **FLOATING
C11681 S.n10604 SUB 1.88fF $ **FLOATING
C11682 S.n10605 SUB 2.67fF $ **FLOATING
C11683 S.t2215 SUB 0.02fF
C11684 S.n10606 SUB 0.24fF $ **FLOATING
C11685 S.n10607 SUB 0.36fF $ **FLOATING
C11686 S.n10608 SUB 0.61fF $ **FLOATING
C11687 S.n10609 SUB 0.12fF $ **FLOATING
C11688 S.t1632 SUB 0.02fF
C11689 S.n10610 SUB 0.14fF $ **FLOATING
C11690 S.n10612 SUB 5.17fF $ **FLOATING
C11691 S.t1873 SUB 0.02fF
C11692 S.n10613 SUB 0.12fF $ **FLOATING
C11693 S.n10614 SUB 0.14fF $ **FLOATING
C11694 S.t1257 SUB 0.02fF
C11695 S.n10616 SUB 0.24fF $ **FLOATING
C11696 S.n10617 SUB 0.91fF $ **FLOATING
C11697 S.n10618 SUB 0.05fF $ **FLOATING
C11698 S.n10619 SUB 1.88fF $ **FLOATING
C11699 S.n10620 SUB 2.67fF $ **FLOATING
C11700 S.t1354 SUB 0.02fF
C11701 S.n10621 SUB 0.24fF $ **FLOATING
C11702 S.n10622 SUB 0.36fF $ **FLOATING
C11703 S.n10623 SUB 0.61fF $ **FLOATING
C11704 S.n10624 SUB 0.12fF $ **FLOATING
C11705 S.t765 SUB 0.02fF
C11706 S.n10625 SUB 0.14fF $ **FLOATING
C11707 S.n10627 SUB 5.17fF $ **FLOATING
C11708 S.t1008 SUB 0.02fF
C11709 S.n10628 SUB 0.12fF $ **FLOATING
C11710 S.n10629 SUB 0.14fF $ **FLOATING
C11711 S.t375 SUB 0.02fF
C11712 S.n10631 SUB 0.24fF $ **FLOATING
C11713 S.n10632 SUB 0.91fF $ **FLOATING
C11714 S.n10633 SUB 0.05fF $ **FLOATING
C11715 S.n10634 SUB 1.88fF $ **FLOATING
C11716 S.n10635 SUB 2.67fF $ **FLOATING
C11717 S.t474 SUB 0.02fF
C11718 S.n10636 SUB 0.24fF $ **FLOATING
C11719 S.n10637 SUB 0.36fF $ **FLOATING
C11720 S.n10638 SUB 0.61fF $ **FLOATING
C11721 S.n10639 SUB 0.12fF $ **FLOATING
C11722 S.t2418 SUB 0.02fF
C11723 S.n10640 SUB 0.14fF $ **FLOATING
C11724 S.n10642 SUB 5.17fF $ **FLOATING
C11725 S.t104 SUB 0.02fF
C11726 S.n10643 SUB 0.12fF $ **FLOATING
C11727 S.n10644 SUB 0.14fF $ **FLOATING
C11728 S.t2026 SUB 0.02fF
C11729 S.n10646 SUB 0.24fF $ **FLOATING
C11730 S.n10647 SUB 0.91fF $ **FLOATING
C11731 S.n10648 SUB 0.05fF $ **FLOATING
C11732 S.n10649 SUB 1.88fF $ **FLOATING
C11733 S.n10650 SUB 2.67fF $ **FLOATING
C11734 S.t2124 SUB 0.02fF
C11735 S.n10651 SUB 0.24fF $ **FLOATING
C11736 S.n10652 SUB 0.36fF $ **FLOATING
C11737 S.n10653 SUB 0.61fF $ **FLOATING
C11738 S.n10654 SUB 0.12fF $ **FLOATING
C11739 S.t1553 SUB 0.02fF
C11740 S.n10655 SUB 0.14fF $ **FLOATING
C11741 S.n10657 SUB 5.17fF $ **FLOATING
C11742 S.t1779 SUB 0.02fF
C11743 S.n10658 SUB 0.12fF $ **FLOATING
C11744 S.n10659 SUB 0.14fF $ **FLOATING
C11745 S.t1169 SUB 0.02fF
C11746 S.n10661 SUB 0.24fF $ **FLOATING
C11747 S.n10662 SUB 0.91fF $ **FLOATING
C11748 S.n10663 SUB 0.05fF $ **FLOATING
C11749 S.n10664 SUB 1.88fF $ **FLOATING
C11750 S.n10665 SUB 2.67fF $ **FLOATING
C11751 S.t1400 SUB 0.02fF
C11752 S.n10666 SUB 0.24fF $ **FLOATING
C11753 S.n10667 SUB 0.36fF $ **FLOATING
C11754 S.n10668 SUB 0.61fF $ **FLOATING
C11755 S.n10669 SUB 0.12fF $ **FLOATING
C11756 S.t817 SUB 0.02fF
C11757 S.n10670 SUB 0.14fF $ **FLOATING
C11758 S.n10672 SUB 5.17fF $ **FLOATING
C11759 S.t907 SUB 0.02fF
C11760 S.n10673 SUB 0.12fF $ **FLOATING
C11761 S.n10674 SUB 0.14fF $ **FLOATING
C11762 S.t422 SUB 0.02fF
C11763 S.n10676 SUB 0.24fF $ **FLOATING
C11764 S.n10677 SUB 0.91fF $ **FLOATING
C11765 S.n10678 SUB 0.05fF $ **FLOATING
C11766 S.n10679 SUB 1.88fF $ **FLOATING
C11767 S.n10680 SUB 2.67fF $ **FLOATING
C11768 S.t529 SUB 0.02fF
C11769 S.n10681 SUB 0.24fF $ **FLOATING
C11770 S.n10682 SUB 0.36fF $ **FLOATING
C11771 S.n10683 SUB 0.61fF $ **FLOATING
C11772 S.n10684 SUB 0.12fF $ **FLOATING
C11773 S.t2464 SUB 0.02fF
C11774 S.n10685 SUB 0.14fF $ **FLOATING
C11775 S.n10687 SUB 5.17fF $ **FLOATING
C11776 S.t2549 SUB 0.02fF
C11777 S.n10688 SUB 0.12fF $ **FLOATING
C11778 S.n10689 SUB 0.14fF $ **FLOATING
C11779 S.t2076 SUB 0.02fF
C11780 S.n10691 SUB 0.24fF $ **FLOATING
C11781 S.n10692 SUB 0.91fF $ **FLOATING
C11782 S.n10693 SUB 0.05fF $ **FLOATING
C11783 S.n10694 SUB 1.88fF $ **FLOATING
C11784 S.n10695 SUB 2.67fF $ **FLOATING
C11785 S.t2171 SUB 0.02fF
C11786 S.n10696 SUB 0.24fF $ **FLOATING
C11787 S.n10697 SUB 0.36fF $ **FLOATING
C11788 S.n10698 SUB 0.61fF $ **FLOATING
C11789 S.n10699 SUB 0.12fF $ **FLOATING
C11790 S.t1594 SUB 0.02fF
C11791 S.n10700 SUB 0.14fF $ **FLOATING
C11792 S.n10702 SUB 5.17fF $ **FLOATING
C11793 S.t1679 SUB 0.02fF
C11794 S.n10703 SUB 0.12fF $ **FLOATING
C11795 S.n10704 SUB 0.14fF $ **FLOATING
C11796 S.t1213 SUB 0.02fF
C11797 S.n10706 SUB 0.24fF $ **FLOATING
C11798 S.n10707 SUB 0.91fF $ **FLOATING
C11799 S.n10708 SUB 0.05fF $ **FLOATING
C11800 S.n10709 SUB 1.88fF $ **FLOATING
C11801 S.n10710 SUB 2.67fF $ **FLOATING
C11802 S.t1307 SUB 0.02fF
C11803 S.n10711 SUB 0.24fF $ **FLOATING
C11804 S.n10712 SUB 0.36fF $ **FLOATING
C11805 S.n10713 SUB 0.61fF $ **FLOATING
C11806 S.n10714 SUB 0.12fF $ **FLOATING
C11807 S.t731 SUB 0.02fF
C11808 S.n10715 SUB 0.14fF $ **FLOATING
C11809 S.n10717 SUB 4.90fF $ **FLOATING
C11810 S.t805 SUB 0.02fF
C11811 S.n10718 SUB 0.12fF $ **FLOATING
C11812 S.n10719 SUB 0.14fF $ **FLOATING
C11813 S.t334 SUB 0.02fF
C11814 S.n10721 SUB 0.24fF $ **FLOATING
C11815 S.n10722 SUB 0.91fF $ **FLOATING
C11816 S.n10723 SUB 0.05fF $ **FLOATING
C11817 S.n10724 SUB 1.88fF $ **FLOATING
C11818 S.n10725 SUB 2.67fF $ **FLOATING
C11819 S.t2281 SUB 0.02fF
C11820 S.n10726 SUB 0.24fF $ **FLOATING
C11821 S.n10727 SUB 0.36fF $ **FLOATING
C11822 S.n10728 SUB 0.61fF $ **FLOATING
C11823 S.n10729 SUB 0.12fF $ **FLOATING
C11824 S.t1017 SUB 0.02fF
C11825 S.n10730 SUB 0.14fF $ **FLOATING
C11826 S.n10732 SUB 1.88fF $ **FLOATING
C11827 S.n10733 SUB 2.68fF $ **FLOATING
C11828 S.t1848 SUB 0.02fF
C11829 S.n10734 SUB 0.24fF $ **FLOATING
C11830 S.n10735 SUB 0.36fF $ **FLOATING
C11831 S.n10736 SUB 0.61fF $ **FLOATING
C11832 S.t810 SUB 0.02fF
C11833 S.n10737 SUB 1.22fF $ **FLOATING
C11834 S.n10738 SUB 0.61fF $ **FLOATING
C11835 S.n10739 SUB 0.35fF $ **FLOATING
C11836 S.n10740 SUB 0.63fF $ **FLOATING
C11837 S.n10741 SUB 1.15fF $ **FLOATING
C11838 S.n10742 SUB 3.03fF $ **FLOATING
C11839 S.n10743 SUB 0.59fF $ **FLOATING
C11840 S.n10744 SUB 0.02fF $ **FLOATING
C11841 S.n10745 SUB 0.97fF $ **FLOATING
C11842 S.t6 SUB 21.38fF
C11843 S.n10746 SUB 20.25fF $ **FLOATING
C11844 S.n10748 SUB 0.38fF $ **FLOATING
C11845 S.n10749 SUB 0.23fF $ **FLOATING
C11846 S.n10750 SUB 2.89fF $ **FLOATING
C11847 S.n10751 SUB 2.46fF $ **FLOATING
C11848 S.n10752 SUB 2.53fF $ **FLOATING
C11849 S.n10753 SUB 3.94fF $ **FLOATING
C11850 S.n10754 SUB 0.25fF $ **FLOATING
C11851 S.n10755 SUB 0.01fF $ **FLOATING
C11852 S.t568 SUB 0.02fF
C11853 S.n10756 SUB 0.25fF $ **FLOATING
C11854 S.t2498 SUB 0.02fF
C11855 S.n10757 SUB 0.95fF $ **FLOATING
C11856 S.n10758 SUB 0.70fF $ **FLOATING
C11857 S.n10759 SUB 1.88fF $ **FLOATING
C11858 S.n10760 SUB 0.48fF $ **FLOATING
C11859 S.n10761 SUB 0.09fF $ **FLOATING
C11860 S.n10762 SUB 0.33fF $ **FLOATING
C11861 S.n10763 SUB 0.30fF $ **FLOATING
C11862 S.n10764 SUB 0.77fF $ **FLOATING
C11863 S.n10765 SUB 0.59fF $ **FLOATING
C11864 S.t2457 SUB 0.02fF
C11865 S.n10766 SUB 0.24fF $ **FLOATING
C11866 S.n10767 SUB 0.36fF $ **FLOATING
C11867 S.n10768 SUB 0.61fF $ **FLOATING
C11868 S.n10769 SUB 0.12fF $ **FLOATING
C11869 S.t2211 SUB 0.02fF
C11870 S.n10770 SUB 0.14fF $ **FLOATING
C11871 S.n10772 SUB 1.44fF $ **FLOATING
C11872 S.n10773 SUB 2.16fF $ **FLOATING
C11873 S.t1621 SUB 0.02fF
C11874 S.n10774 SUB 0.24fF $ **FLOATING
C11875 S.n10775 SUB 0.91fF $ **FLOATING
C11876 S.n10776 SUB 0.05fF $ **FLOATING
C11877 S.t339 SUB 0.02fF
C11878 S.n10777 SUB 0.12fF $ **FLOATING
C11879 S.n10778 SUB 0.14fF $ **FLOATING
C11880 S.n10780 SUB 0.78fF $ **FLOATING
C11881 S.n10781 SUB 2.30fF $ **FLOATING
C11882 S.n10782 SUB 1.88fF $ **FLOATING
C11883 S.n10783 SUB 0.12fF $ **FLOATING
C11884 S.t1352 SUB 0.02fF
C11885 S.n10784 SUB 0.14fF $ **FLOATING
C11886 S.t1589 SUB 0.02fF
C11887 S.n10786 SUB 0.24fF $ **FLOATING
C11888 S.n10787 SUB 0.36fF $ **FLOATING
C11889 S.n10788 SUB 0.61fF $ **FLOATING
C11890 S.n10789 SUB 1.39fF $ **FLOATING
C11891 S.n10790 SUB 0.71fF $ **FLOATING
C11892 S.n10791 SUB 1.14fF $ **FLOATING
C11893 S.n10792 SUB 0.35fF $ **FLOATING
C11894 S.n10793 SUB 2.03fF $ **FLOATING
C11895 S.t754 SUB 0.02fF
C11896 S.n10794 SUB 0.24fF $ **FLOATING
C11897 S.n10795 SUB 0.91fF $ **FLOATING
C11898 S.n10796 SUB 0.05fF $ **FLOATING
C11899 S.t1997 SUB 0.02fF
C11900 S.n10797 SUB 0.12fF $ **FLOATING
C11901 S.n10798 SUB 0.14fF $ **FLOATING
C11902 S.n10800 SUB 1.89fF $ **FLOATING
C11903 S.n10801 SUB 1.88fF $ **FLOATING
C11904 S.t724 SUB 0.02fF
C11905 S.n10802 SUB 0.24fF $ **FLOATING
C11906 S.n10803 SUB 0.36fF $ **FLOATING
C11907 S.n10804 SUB 0.61fF $ **FLOATING
C11908 S.n10805 SUB 0.12fF $ **FLOATING
C11909 S.t472 SUB 0.02fF
C11910 S.n10806 SUB 0.14fF $ **FLOATING
C11911 S.n10808 SUB 1.16fF $ **FLOATING
C11912 S.n10809 SUB 0.22fF $ **FLOATING
C11913 S.n10810 SUB 0.25fF $ **FLOATING
C11914 S.n10811 SUB 0.09fF $ **FLOATING
C11915 S.n10812 SUB 1.88fF $ **FLOATING
C11916 S.t2409 SUB 0.02fF
C11917 S.n10813 SUB 0.24fF $ **FLOATING
C11918 S.n10814 SUB 0.91fF $ **FLOATING
C11919 S.n10815 SUB 0.05fF $ **FLOATING
C11920 S.t1270 SUB 0.02fF
C11921 S.n10816 SUB 0.12fF $ **FLOATING
C11922 S.n10817 SUB 0.14fF $ **FLOATING
C11923 S.n10819 SUB 20.78fF $ **FLOATING
C11924 S.n10820 SUB 1.88fF $ **FLOATING
C11925 S.n10821 SUB 2.67fF $ **FLOATING
C11926 S.t661 SUB 0.02fF
C11927 S.n10822 SUB 0.24fF $ **FLOATING
C11928 S.n10823 SUB 0.36fF $ **FLOATING
C11929 S.n10824 SUB 0.61fF $ **FLOATING
C11930 S.n10825 SUB 0.12fF $ **FLOATING
C11931 S.t372 SUB 0.02fF
C11932 S.n10826 SUB 0.14fF $ **FLOATING
C11933 S.n10828 SUB 2.80fF $ **FLOATING
C11934 S.n10829 SUB 2.30fF $ **FLOATING
C11935 S.t1181 SUB 0.02fF
C11936 S.n10830 SUB 0.12fF $ **FLOATING
C11937 S.n10831 SUB 0.14fF $ **FLOATING
C11938 S.t2344 SUB 0.02fF
C11939 S.n10833 SUB 0.24fF $ **FLOATING
C11940 S.n10834 SUB 0.91fF $ **FLOATING
C11941 S.n10835 SUB 0.05fF $ **FLOATING
C11942 S.n10836 SUB 1.88fF $ **FLOATING
C11943 S.n10837 SUB 2.67fF $ **FLOATING
C11944 S.t2314 SUB 0.02fF
C11945 S.n10838 SUB 0.24fF $ **FLOATING
C11946 S.n10839 SUB 0.36fF $ **FLOATING
C11947 S.n10840 SUB 0.61fF $ **FLOATING
C11948 S.n10841 SUB 0.12fF $ **FLOATING
C11949 S.t2168 SUB 0.02fF
C11950 S.n10842 SUB 0.14fF $ **FLOATING
C11951 S.n10844 SUB 2.80fF $ **FLOATING
C11952 S.n10845 SUB 2.30fF $ **FLOATING
C11953 S.t304 SUB 0.02fF
C11954 S.n10846 SUB 0.12fF $ **FLOATING
C11955 S.n10847 SUB 0.14fF $ **FLOATING
C11956 S.t1484 SUB 0.02fF
C11957 S.n10849 SUB 0.24fF $ **FLOATING
C11958 S.n10850 SUB 0.91fF $ **FLOATING
C11959 S.n10851 SUB 0.05fF $ **FLOATING
C11960 S.n10852 SUB 1.88fF $ **FLOATING
C11961 S.n10853 SUB 2.67fF $ **FLOATING
C11962 S.t1206 SUB 0.02fF
C11963 S.n10854 SUB 0.24fF $ **FLOATING
C11964 S.n10855 SUB 0.36fF $ **FLOATING
C11965 S.n10856 SUB 0.61fF $ **FLOATING
C11966 S.n10857 SUB 0.12fF $ **FLOATING
C11967 S.t1956 SUB 0.02fF
C11968 S.n10858 SUB 0.14fF $ **FLOATING
C11969 S.n10860 SUB 2.80fF $ **FLOATING
C11970 S.n10861 SUB 2.30fF $ **FLOATING
C11971 S.t1968 SUB 0.02fF
C11972 S.n10862 SUB 0.12fF $ **FLOATING
C11973 S.n10863 SUB 0.14fF $ **FLOATING
C11974 S.t494 SUB 0.02fF
C11975 S.n10865 SUB 0.24fF $ **FLOATING
C11976 S.n10866 SUB 0.91fF $ **FLOATING
C11977 S.n10867 SUB 0.05fF $ **FLOATING
C11978 S.n10868 SUB 1.88fF $ **FLOATING
C11979 S.n10869 SUB 2.67fF $ **FLOATING
C11980 S.t328 SUB 0.02fF
C11981 S.n10870 SUB 0.24fF $ **FLOATING
C11982 S.n10871 SUB 0.36fF $ **FLOATING
C11983 S.n10872 SUB 0.61fF $ **FLOATING
C11984 S.n10873 SUB 0.12fF $ **FLOATING
C11985 S.t1098 SUB 0.02fF
C11986 S.n10874 SUB 0.14fF $ **FLOATING
C11987 S.n10876 SUB 2.80fF $ **FLOATING
C11988 S.n10877 SUB 2.30fF $ **FLOATING
C11989 S.t1761 SUB 0.02fF
C11990 S.n10878 SUB 0.12fF $ **FLOATING
C11991 S.n10879 SUB 0.14fF $ **FLOATING
C11992 S.t2140 SUB 0.02fF
C11993 S.n10881 SUB 0.24fF $ **FLOATING
C11994 S.n10882 SUB 0.91fF $ **FLOATING
C11995 S.n10883 SUB 0.05fF $ **FLOATING
C11996 S.n10884 SUB 1.88fF $ **FLOATING
C11997 S.n10885 SUB 2.67fF $ **FLOATING
C11998 S.t1987 SUB 0.02fF
C11999 S.n10886 SUB 0.24fF $ **FLOATING
C12000 S.n10887 SUB 0.36fF $ **FLOATING
C12001 S.n10888 SUB 0.61fF $ **FLOATING
C12002 S.n10889 SUB 0.12fF $ **FLOATING
C12003 S.t223 SUB 0.02fF
C12004 S.n10890 SUB 0.14fF $ **FLOATING
C12005 S.n10892 SUB 2.80fF $ **FLOATING
C12006 S.n10893 SUB 2.30fF $ **FLOATING
C12007 S.t884 SUB 0.02fF
C12008 S.n10894 SUB 0.12fF $ **FLOATING
C12009 S.n10895 SUB 0.14fF $ **FLOATING
C12010 S.t1274 SUB 0.02fF
C12011 S.n10897 SUB 0.24fF $ **FLOATING
C12012 S.n10898 SUB 0.91fF $ **FLOATING
C12013 S.n10899 SUB 0.05fF $ **FLOATING
C12014 S.n10900 SUB 1.88fF $ **FLOATING
C12015 S.n10901 SUB 2.67fF $ **FLOATING
C12016 S.t1137 SUB 0.02fF
C12017 S.n10902 SUB 0.24fF $ **FLOATING
C12018 S.n10903 SUB 0.36fF $ **FLOATING
C12019 S.n10904 SUB 0.61fF $ **FLOATING
C12020 S.n10905 SUB 0.12fF $ **FLOATING
C12021 S.t1888 SUB 0.02fF
C12022 S.n10906 SUB 0.14fF $ **FLOATING
C12023 S.n10908 SUB 2.80fF $ **FLOATING
C12024 S.n10909 SUB 2.30fF $ **FLOATING
C12025 S.t2528 SUB 0.02fF
C12026 S.n10910 SUB 0.12fF $ **FLOATING
C12027 S.n10911 SUB 0.14fF $ **FLOATING
C12028 S.t392 SUB 0.02fF
C12029 S.n10913 SUB 0.24fF $ **FLOATING
C12030 S.n10914 SUB 0.91fF $ **FLOATING
C12031 S.n10915 SUB 0.05fF $ **FLOATING
C12032 S.n10916 SUB 1.88fF $ **FLOATING
C12033 S.n10917 SUB 2.67fF $ **FLOATING
C12034 S.t259 SUB 0.02fF
C12035 S.n10918 SUB 0.24fF $ **FLOATING
C12036 S.n10919 SUB 0.36fF $ **FLOATING
C12037 S.n10920 SUB 0.61fF $ **FLOATING
C12038 S.n10921 SUB 0.12fF $ **FLOATING
C12039 S.t1026 SUB 0.02fF
C12040 S.n10922 SUB 0.14fF $ **FLOATING
C12041 S.n10924 SUB 2.80fF $ **FLOATING
C12042 S.n10925 SUB 2.30fF $ **FLOATING
C12043 S.t1652 SUB 0.02fF
C12044 S.n10926 SUB 0.12fF $ **FLOATING
C12045 S.n10927 SUB 0.14fF $ **FLOATING
C12046 S.t2041 SUB 0.02fF
C12047 S.n10929 SUB 0.24fF $ **FLOATING
C12048 S.n10930 SUB 0.91fF $ **FLOATING
C12049 S.n10931 SUB 0.05fF $ **FLOATING
C12050 S.n10932 SUB 1.88fF $ **FLOATING
C12051 S.n10933 SUB 2.67fF $ **FLOATING
C12052 S.t1925 SUB 0.02fF
C12053 S.n10934 SUB 0.24fF $ **FLOATING
C12054 S.n10935 SUB 0.36fF $ **FLOATING
C12055 S.n10936 SUB 0.61fF $ **FLOATING
C12056 S.n10937 SUB 0.12fF $ **FLOATING
C12057 S.t123 SUB 0.02fF
C12058 S.n10938 SUB 0.14fF $ **FLOATING
C12059 S.n10940 SUB 2.80fF $ **FLOATING
C12060 S.n10941 SUB 2.30fF $ **FLOATING
C12061 S.t950 SUB 0.02fF
C12062 S.n10942 SUB 0.12fF $ **FLOATING
C12063 S.n10943 SUB 0.14fF $ **FLOATING
C12064 S.t1184 SUB 0.02fF
C12065 S.n10945 SUB 0.24fF $ **FLOATING
C12066 S.n10946 SUB 0.91fF $ **FLOATING
C12067 S.n10947 SUB 0.05fF $ **FLOATING
C12068 S.n10948 SUB 1.88fF $ **FLOATING
C12069 S.n10949 SUB 2.67fF $ **FLOATING
C12070 S.t1065 SUB 0.02fF
C12071 S.n10950 SUB 0.24fF $ **FLOATING
C12072 S.n10951 SUB 0.36fF $ **FLOATING
C12073 S.n10952 SUB 0.61fF $ **FLOATING
C12074 S.n10953 SUB 0.12fF $ **FLOATING
C12075 S.t1793 SUB 0.02fF
C12076 S.n10954 SUB 0.14fF $ **FLOATING
C12077 S.n10956 SUB 2.80fF $ **FLOATING
C12078 S.n10957 SUB 2.30fF $ **FLOATING
C12079 S.t2587 SUB 0.02fF
C12080 S.n10958 SUB 0.12fF $ **FLOATING
C12081 S.n10959 SUB 0.14fF $ **FLOATING
C12082 S.t309 SUB 0.02fF
C12083 S.n10961 SUB 0.24fF $ **FLOATING
C12084 S.n10962 SUB 0.91fF $ **FLOATING
C12085 S.n10963 SUB 0.05fF $ **FLOATING
C12086 S.n10964 SUB 1.88fF $ **FLOATING
C12087 S.n10965 SUB 2.67fF $ **FLOATING
C12088 S.t184 SUB 0.02fF
C12089 S.n10966 SUB 0.24fF $ **FLOATING
C12090 S.n10967 SUB 0.36fF $ **FLOATING
C12091 S.n10968 SUB 0.61fF $ **FLOATING
C12092 S.n10969 SUB 0.12fF $ **FLOATING
C12093 S.t926 SUB 0.02fF
C12094 S.n10970 SUB 0.14fF $ **FLOATING
C12095 S.n10972 SUB 2.80fF $ **FLOATING
C12096 S.n10973 SUB 2.30fF $ **FLOATING
C12097 S.t1710 SUB 0.02fF
C12098 S.n10974 SUB 0.12fF $ **FLOATING
C12099 S.n10975 SUB 0.14fF $ **FLOATING
C12100 S.t1971 SUB 0.02fF
C12101 S.n10977 SUB 0.24fF $ **FLOATING
C12102 S.n10978 SUB 0.91fF $ **FLOATING
C12103 S.n10979 SUB 0.05fF $ **FLOATING
C12104 S.n10980 SUB 2.73fF $ **FLOATING
C12105 S.n10981 SUB 1.59fF $ **FLOATING
C12106 S.n10982 SUB 0.12fF $ **FLOATING
C12107 S.t1469 SUB 0.02fF
C12108 S.n10983 SUB 0.14fF $ **FLOATING
C12109 S.t199 SUB 0.02fF
C12110 S.n10985 SUB 0.24fF $ **FLOATING
C12111 S.n10986 SUB 0.36fF $ **FLOATING
C12112 S.n10987 SUB 0.61fF $ **FLOATING
C12113 S.n10988 SUB 0.07fF $ **FLOATING
C12114 S.n10989 SUB 0.01fF $ **FLOATING
C12115 S.n10990 SUB 0.24fF $ **FLOATING
C12116 S.n10991 SUB 1.16fF $ **FLOATING
C12117 S.n10992 SUB 1.35fF $ **FLOATING
C12118 S.n10993 SUB 2.30fF $ **FLOATING
C12119 S.t2229 SUB 0.02fF
C12120 S.n10994 SUB 0.12fF $ **FLOATING
C12121 S.n10995 SUB 0.14fF $ **FLOATING
C12122 S.t1167 SUB 0.02fF
C12123 S.n10997 SUB 0.24fF $ **FLOATING
C12124 S.n10998 SUB 0.91fF $ **FLOATING
C12125 S.n10999 SUB 0.05fF $ **FLOATING
C12126 S.t122 SUB 48.31fF
C12127 S.t1116 SUB 0.02fF
C12128 S.n11000 SUB 0.24fF $ **FLOATING
C12129 S.n11001 SUB 0.91fF $ **FLOATING
C12130 S.n11002 SUB 0.05fF $ **FLOATING
C12131 S.t840 SUB 0.02fF
C12132 S.n11003 SUB 0.12fF $ **FLOATING
C12133 S.n11004 SUB 0.14fF $ **FLOATING
C12134 S.n11006 SUB 0.12fF $ **FLOATING
C12135 S.t2566 SUB 0.02fF
C12136 S.n11007 SUB 0.14fF $ **FLOATING
C12137 S.n11009 SUB 5.17fF $ **FLOATING
C12138 S.n11010 SUB 5.44fF $ **FLOATING
C12139 S.t2454 SUB 0.02fF
C12140 S.n11011 SUB 0.12fF $ **FLOATING
C12141 S.n11012 SUB 0.14fF $ **FLOATING
C12142 S.t1665 SUB 0.02fF
C12143 S.n11014 SUB 0.24fF $ **FLOATING
C12144 S.n11015 SUB 0.91fF $ **FLOATING
C12145 S.n11016 SUB 0.05fF $ **FLOATING
C12146 S.t103 SUB 47.92fF
C12147 S.t401 SUB 0.02fF
C12148 S.n11017 SUB 1.19fF $ **FLOATING
C12149 S.n11018 SUB 0.05fF $ **FLOATING
C12150 S.t248 SUB 0.02fF
C12151 S.n11019 SUB 0.01fF $ **FLOATING
C12152 S.n11020 SUB 0.26fF $ **FLOATING
C12153 S.n11022 SUB 1.50fF $ **FLOATING
C12154 S.n11023 SUB 1.30fF $ **FLOATING
C12155 S.n11024 SUB 0.28fF $ **FLOATING
C12156 S.n11025 SUB 0.24fF $ **FLOATING
C12157 S.n11026 SUB 4.39fF $ **FLOATING
C12158 S.n11027 SUB 0.02fF $ **FLOATING
C12159 S.n11028 SUB 0.03fF $ **FLOATING
C12160 S.n11029 SUB 0.24fF $ **FLOATING
C12161 S.n11030 SUB 0.13fF $ **FLOATING
C12162 S.n11031 SUB 0.56fF $ **FLOATING
C12163 S.n11032 SUB 0.03fF $ **FLOATING
C12164 S.n11033 SUB 0.86fF $ **FLOATING
C12165 S.n11034 SUB 0.22fF $ **FLOATING
C12166 S.n11035 SUB 0.15fF $ **FLOATING
C12167 S.n11036 SUB 8.97fF $ **FLOATING
C12168 S.n11037 SUB 8.97fF $ **FLOATING
C12169 S.n11038 SUB 0.60fF $ **FLOATING
C12170 S.n11039 SUB 0.22fF $ **FLOATING
C12171 S.n11040 SUB 0.59fF $ **FLOATING
C12172 S.n11041 SUB 3.43fF $ **FLOATING
C12173 S.n11042 SUB 0.29fF $ **FLOATING
C12174 S.t261 SUB 21.38fF
C12175 S.n11043 SUB 21.67fF $ **FLOATING
C12176 S.n11044 SUB 0.77fF $ **FLOATING
C12177 S.n11045 SUB 0.28fF $ **FLOATING
C12178 S.n11046 SUB 4.00fF $ **FLOATING
C12179 S.n11047 SUB 1.14fF $ **FLOATING
C12180 S.t535 SUB 0.02fF
C12181 S.n11048 SUB 0.64fF $ **FLOATING
C12182 S.n11049 SUB 0.61fF $ **FLOATING
C12183 S.n11050 SUB 0.25fF $ **FLOATING
C12184 S.n11051 SUB 0.09fF $ **FLOATING
C12185 S.n11052 SUB 0.21fF $ **FLOATING
C12186 S.n11053 SUB 1.28fF $ **FLOATING
C12187 S.n11054 SUB 0.53fF $ **FLOATING
C12188 S.n11055 SUB 1.88fF $ **FLOATING
C12189 S.n11056 SUB 0.12fF $ **FLOATING
C12190 S.t2544 SUB 0.02fF
C12191 S.n11057 SUB 0.14fF $ **FLOATING
C12192 S.t584 SUB 0.02fF
C12193 S.n11059 SUB 0.24fF $ **FLOATING
C12194 S.n11060 SUB 0.36fF $ **FLOATING
C12195 S.n11061 SUB 0.61fF $ **FLOATING
C12196 S.n11062 SUB 1.58fF $ **FLOATING
C12197 S.n11063 SUB 2.45fF $ **FLOATING
C12198 S.t1666 SUB 0.02fF
C12199 S.n11064 SUB 0.24fF $ **FLOATING
C12200 S.n11065 SUB 0.91fF $ **FLOATING
C12201 S.n11066 SUB 0.05fF $ **FLOATING
C12202 S.t231 SUB 0.02fF
C12203 S.n11067 SUB 0.12fF $ **FLOATING
C12204 S.n11068 SUB 0.14fF $ **FLOATING
C12205 S.n11070 SUB 1.89fF $ **FLOATING
C12206 S.n11071 SUB 0.06fF $ **FLOATING
C12207 S.n11072 SUB 0.03fF $ **FLOATING
C12208 S.n11073 SUB 0.04fF $ **FLOATING
C12209 S.n11074 SUB 0.99fF $ **FLOATING
C12210 S.n11075 SUB 0.02fF $ **FLOATING
C12211 S.n11076 SUB 0.01fF $ **FLOATING
C12212 S.n11077 SUB 0.02fF $ **FLOATING
C12213 S.n11078 SUB 0.08fF $ **FLOATING
C12214 S.n11079 SUB 0.36fF $ **FLOATING
C12215 S.n11080 SUB 1.85fF $ **FLOATING
C12216 S.t2337 SUB 0.02fF
C12217 S.n11081 SUB 0.24fF $ **FLOATING
C12218 S.n11082 SUB 0.36fF $ **FLOATING
C12219 S.n11083 SUB 0.61fF $ **FLOATING
C12220 S.n11084 SUB 0.12fF $ **FLOATING
C12221 S.t1824 SUB 0.02fF
C12222 S.n11085 SUB 0.14fF $ **FLOATING
C12223 S.n11087 SUB 0.70fF $ **FLOATING
C12224 S.n11088 SUB 0.23fF $ **FLOATING
C12225 S.n11089 SUB 0.23fF $ **FLOATING
C12226 S.n11090 SUB 0.70fF $ **FLOATING
C12227 S.n11091 SUB 1.16fF $ **FLOATING
C12228 S.n11092 SUB 0.22fF $ **FLOATING
C12229 S.n11093 SUB 0.25fF $ **FLOATING
C12230 S.n11094 SUB 0.09fF $ **FLOATING
C12231 S.n11095 SUB 1.88fF $ **FLOATING
C12232 S.t956 SUB 0.02fF
C12233 S.n11096 SUB 0.24fF $ **FLOATING
C12234 S.n11097 SUB 0.91fF $ **FLOATING
C12235 S.n11098 SUB 0.05fF $ **FLOATING
C12236 S.t1897 SUB 0.02fF
C12237 S.n11099 SUB 0.12fF $ **FLOATING
C12238 S.n11100 SUB 0.14fF $ **FLOATING
C12239 S.n11102 SUB 20.78fF $ **FLOATING
C12240 S.n11103 SUB 2.38fF $ **FLOATING
C12241 S.n11104 SUB 0.46fF $ **FLOATING
C12242 S.n11105 SUB 0.22fF $ **FLOATING
C12243 S.n11106 SUB 0.38fF $ **FLOATING
C12244 S.n11107 SUB 0.16fF $ **FLOATING
C12245 S.n11108 SUB 0.28fF $ **FLOATING
C12246 S.n11109 SUB 0.21fF $ **FLOATING
C12247 S.n11110 SUB 0.30fF $ **FLOATING
C12248 S.n11111 SUB 0.21fF $ **FLOATING
C12249 S.t1446 SUB 0.02fF
C12250 S.n11112 SUB 0.24fF $ **FLOATING
C12251 S.n11113 SUB 0.36fF $ **FLOATING
C12252 S.n11114 SUB 0.61fF $ **FLOATING
C12253 S.n11115 SUB 0.12fF $ **FLOATING
C12254 S.t901 SUB 0.02fF
C12255 S.n11116 SUB 0.14fF $ **FLOATING
C12256 S.n11118 SUB 0.19fF $ **FLOATING
C12257 S.n11119 SUB 1.57fF $ **FLOATING
C12258 S.n11120 SUB 2.21fF $ **FLOATING
C12259 S.n11121 SUB 0.32fF $ **FLOATING
C12260 S.n11122 SUB 2.39fF $ **FLOATING
C12261 S.t1107 SUB 0.02fF
C12262 S.n11123 SUB 0.12fF $ **FLOATING
C12263 S.n11124 SUB 0.14fF $ **FLOATING
C12264 S.t2537 SUB 0.02fF
C12265 S.n11126 SUB 0.24fF $ **FLOATING
C12266 S.n11127 SUB 0.91fF $ **FLOATING
C12267 S.n11128 SUB 0.05fF $ **FLOATING
C12268 S.n11129 SUB 1.88fF $ **FLOATING
C12269 S.n11130 SUB 0.12fF $ **FLOATING
C12270 S.t185 SUB 0.02fF
C12271 S.n11131 SUB 0.14fF $ **FLOATING
C12272 S.t997 SUB 0.02fF
C12273 S.n11133 SUB 0.12fF $ **FLOATING
C12274 S.n11134 SUB 0.14fF $ **FLOATING
C12275 S.t2156 SUB 0.02fF
C12276 S.n11136 SUB 0.24fF $ **FLOATING
C12277 S.n11137 SUB 0.91fF $ **FLOATING
C12278 S.n11138 SUB 0.05fF $ **FLOATING
C12279 S.t471 SUB 0.02fF
C12280 S.n11139 SUB 0.24fF $ **FLOATING
C12281 S.n11140 SUB 0.36fF $ **FLOATING
C12282 S.n11141 SUB 0.61fF $ **FLOATING
C12283 S.n11142 SUB 0.32fF $ **FLOATING
C12284 S.n11143 SUB 1.09fF $ **FLOATING
C12285 S.n11144 SUB 0.15fF $ **FLOATING
C12286 S.n11145 SUB 2.10fF $ **FLOATING
C12287 S.n11146 SUB 2.94fF $ **FLOATING
C12288 S.n11147 SUB 1.88fF $ **FLOATING
C12289 S.n11148 SUB 0.12fF $ **FLOATING
C12290 S.t960 SUB 0.02fF
C12291 S.n11149 SUB 0.14fF $ **FLOATING
C12292 S.t1478 SUB 0.02fF
C12293 S.n11151 SUB 0.24fF $ **FLOATING
C12294 S.n11152 SUB 0.36fF $ **FLOATING
C12295 S.n11153 SUB 0.61fF $ **FLOATING
C12296 S.n11154 SUB 0.92fF $ **FLOATING
C12297 S.n11155 SUB 0.32fF $ **FLOATING
C12298 S.n11156 SUB 0.92fF $ **FLOATING
C12299 S.n11157 SUB 1.09fF $ **FLOATING
C12300 S.n11158 SUB 0.15fF $ **FLOATING
C12301 S.n11159 SUB 4.96fF $ **FLOATING
C12302 S.t1037 SUB 0.02fF
C12303 S.n11160 SUB 0.12fF $ **FLOATING
C12304 S.n11161 SUB 0.14fF $ **FLOATING
C12305 S.t7 SUB 0.02fF
C12306 S.n11163 SUB 0.24fF $ **FLOATING
C12307 S.n11164 SUB 0.91fF $ **FLOATING
C12308 S.n11165 SUB 0.05fF $ **FLOATING
C12309 S.n11166 SUB 1.88fF $ **FLOATING
C12310 S.n11167 SUB 2.67fF $ **FLOATING
C12311 S.t616 SUB 0.02fF
C12312 S.n11168 SUB 0.24fF $ **FLOATING
C12313 S.n11169 SUB 0.36fF $ **FLOATING
C12314 S.n11170 SUB 0.61fF $ **FLOATING
C12315 S.n11171 SUB 0.12fF $ **FLOATING
C12316 S.t13 SUB 0.02fF
C12317 S.n11172 SUB 0.14fF $ **FLOATING
C12318 S.n11174 SUB 1.88fF $ **FLOATING
C12319 S.n11175 SUB 2.67fF $ **FLOATING
C12320 S.t2120 SUB 0.02fF
C12321 S.n11176 SUB 0.24fF $ **FLOATING
C12322 S.n11177 SUB 0.36fF $ **FLOATING
C12323 S.n11178 SUB 0.61fF $ **FLOATING
C12324 S.t1293 SUB 0.02fF
C12325 S.n11179 SUB 0.24fF $ **FLOATING
C12326 S.n11180 SUB 0.91fF $ **FLOATING
C12327 S.n11181 SUB 0.05fF $ **FLOATING
C12328 S.t93 SUB 0.02fF
C12329 S.n11182 SUB 0.12fF $ **FLOATING
C12330 S.n11183 SUB 0.14fF $ **FLOATING
C12331 S.n11185 SUB 0.12fF $ **FLOATING
C12332 S.t1850 SUB 0.02fF
C12333 S.n11186 SUB 0.14fF $ **FLOATING
C12334 S.n11188 SUB 2.30fF $ **FLOATING
C12335 S.n11189 SUB 2.94fF $ **FLOATING
C12336 S.n11190 SUB 5.16fF $ **FLOATING
C12337 S.t140 SUB 0.02fF
C12338 S.n11191 SUB 0.12fF $ **FLOATING
C12339 S.n11192 SUB 0.14fF $ **FLOATING
C12340 S.t1719 SUB 0.02fF
C12341 S.n11194 SUB 0.24fF $ **FLOATING
C12342 S.n11195 SUB 0.91fF $ **FLOATING
C12343 S.n11196 SUB 0.05fF $ **FLOATING
C12344 S.n11197 SUB 1.88fF $ **FLOATING
C12345 S.n11198 SUB 2.67fF $ **FLOATING
C12346 S.t2272 SUB 0.02fF
C12347 S.n11199 SUB 0.24fF $ **FLOATING
C12348 S.n11200 SUB 0.36fF $ **FLOATING
C12349 S.n11201 SUB 0.61fF $ **FLOATING
C12350 S.n11202 SUB 0.12fF $ **FLOATING
C12351 S.t1723 SUB 0.02fF
C12352 S.n11203 SUB 0.14fF $ **FLOATING
C12353 S.n11205 SUB 5.17fF $ **FLOATING
C12354 S.t1810 SUB 0.02fF
C12355 S.n11206 SUB 0.12fF $ **FLOATING
C12356 S.n11207 SUB 0.14fF $ **FLOATING
C12357 S.t848 SUB 0.02fF
C12358 S.n11209 SUB 0.24fF $ **FLOATING
C12359 S.n11210 SUB 0.91fF $ **FLOATING
C12360 S.n11211 SUB 0.05fF $ **FLOATING
C12361 S.n11212 SUB 1.88fF $ **FLOATING
C12362 S.n11213 SUB 2.67fF $ **FLOATING
C12363 S.t1416 SUB 0.02fF
C12364 S.n11214 SUB 0.24fF $ **FLOATING
C12365 S.n11215 SUB 0.36fF $ **FLOATING
C12366 S.n11216 SUB 0.61fF $ **FLOATING
C12367 S.n11217 SUB 0.12fF $ **FLOATING
C12368 S.t851 SUB 0.02fF
C12369 S.n11218 SUB 0.14fF $ **FLOATING
C12370 S.n11220 SUB 5.17fF $ **FLOATING
C12371 S.t943 SUB 0.02fF
C12372 S.n11221 SUB 0.12fF $ **FLOATING
C12373 S.n11222 SUB 0.14fF $ **FLOATING
C12374 S.t2491 SUB 0.02fF
C12375 S.n11224 SUB 0.24fF $ **FLOATING
C12376 S.n11225 SUB 0.91fF $ **FLOATING
C12377 S.n11226 SUB 0.05fF $ **FLOATING
C12378 S.n11227 SUB 1.88fF $ **FLOATING
C12379 S.n11228 SUB 2.67fF $ **FLOATING
C12380 S.t550 SUB 0.02fF
C12381 S.n11229 SUB 0.24fF $ **FLOATING
C12382 S.n11230 SUB 0.36fF $ **FLOATING
C12383 S.n11231 SUB 0.61fF $ **FLOATING
C12384 S.n11232 SUB 0.12fF $ **FLOATING
C12385 S.t2493 SUB 0.02fF
C12386 S.n11233 SUB 0.14fF $ **FLOATING
C12387 S.n11235 SUB 5.17fF $ **FLOATING
C12388 S.t194 SUB 0.02fF
C12389 S.n11236 SUB 0.12fF $ **FLOATING
C12390 S.n11237 SUB 0.14fF $ **FLOATING
C12391 S.t1616 SUB 0.02fF
C12392 S.n11239 SUB 0.24fF $ **FLOATING
C12393 S.n11240 SUB 0.91fF $ **FLOATING
C12394 S.n11241 SUB 0.05fF $ **FLOATING
C12395 S.n11242 SUB 1.88fF $ **FLOATING
C12396 S.n11243 SUB 2.67fF $ **FLOATING
C12397 S.t1382 SUB 0.02fF
C12398 S.n11244 SUB 0.24fF $ **FLOATING
C12399 S.n11245 SUB 0.36fF $ **FLOATING
C12400 S.n11246 SUB 0.61fF $ **FLOATING
C12401 S.n11247 SUB 0.12fF $ **FLOATING
C12402 S.t796 SUB 0.02fF
C12403 S.n11248 SUB 0.14fF $ **FLOATING
C12404 S.n11250 SUB 5.17fF $ **FLOATING
C12405 S.t1036 SUB 0.02fF
C12406 S.n11251 SUB 0.12fF $ **FLOATING
C12407 S.n11252 SUB 0.14fF $ **FLOATING
C12408 S.t403 SUB 0.02fF
C12409 S.n11254 SUB 0.24fF $ **FLOATING
C12410 S.n11255 SUB 0.91fF $ **FLOATING
C12411 S.n11256 SUB 0.05fF $ **FLOATING
C12412 S.n11257 SUB 1.88fF $ **FLOATING
C12413 S.n11258 SUB 2.67fF $ **FLOATING
C12414 S.t507 SUB 0.02fF
C12415 S.n11259 SUB 0.24fF $ **FLOATING
C12416 S.n11260 SUB 0.36fF $ **FLOATING
C12417 S.n11261 SUB 0.61fF $ **FLOATING
C12418 S.n11262 SUB 0.12fF $ **FLOATING
C12419 S.t2447 SUB 0.02fF
C12420 S.n11263 SUB 0.14fF $ **FLOATING
C12421 S.n11265 SUB 5.17fF $ **FLOATING
C12422 S.t144 SUB 0.02fF
C12423 S.n11266 SUB 0.12fF $ **FLOATING
C12424 S.n11267 SUB 0.14fF $ **FLOATING
C12425 S.t2053 SUB 0.02fF
C12426 S.n11269 SUB 0.24fF $ **FLOATING
C12427 S.n11270 SUB 0.91fF $ **FLOATING
C12428 S.n11271 SUB 0.05fF $ **FLOATING
C12429 S.n11272 SUB 1.88fF $ **FLOATING
C12430 S.n11273 SUB 2.67fF $ **FLOATING
C12431 S.t2152 SUB 0.02fF
C12432 S.n11274 SUB 0.24fF $ **FLOATING
C12433 S.n11275 SUB 0.36fF $ **FLOATING
C12434 S.n11276 SUB 0.61fF $ **FLOATING
C12435 S.n11277 SUB 0.12fF $ **FLOATING
C12436 S.t1578 SUB 0.02fF
C12437 S.n11278 SUB 0.14fF $ **FLOATING
C12438 S.n11280 SUB 5.17fF $ **FLOATING
C12439 S.t1812 SUB 0.02fF
C12440 S.n11281 SUB 0.12fF $ **FLOATING
C12441 S.n11282 SUB 0.14fF $ **FLOATING
C12442 S.t1193 SUB 0.02fF
C12443 S.n11284 SUB 0.24fF $ **FLOATING
C12444 S.n11285 SUB 0.91fF $ **FLOATING
C12445 S.n11286 SUB 0.05fF $ **FLOATING
C12446 S.n11287 SUB 1.88fF $ **FLOATING
C12447 S.n11288 SUB 2.67fF $ **FLOATING
C12448 S.t1292 SUB 0.02fF
C12449 S.n11289 SUB 0.24fF $ **FLOATING
C12450 S.n11290 SUB 0.36fF $ **FLOATING
C12451 S.n11291 SUB 0.61fF $ **FLOATING
C12452 S.n11292 SUB 0.12fF $ **FLOATING
C12453 S.t710 SUB 0.02fF
C12454 S.n11293 SUB 0.14fF $ **FLOATING
C12455 S.n11295 SUB 5.17fF $ **FLOATING
C12456 S.t945 SUB 0.02fF
C12457 S.n11296 SUB 0.12fF $ **FLOATING
C12458 S.n11297 SUB 0.14fF $ **FLOATING
C12459 S.t314 SUB 0.02fF
C12460 S.n11299 SUB 0.24fF $ **FLOATING
C12461 S.n11300 SUB 0.91fF $ **FLOATING
C12462 S.n11301 SUB 0.05fF $ **FLOATING
C12463 S.n11302 SUB 1.88fF $ **FLOATING
C12464 S.n11303 SUB 2.67fF $ **FLOATING
C12465 S.t562 SUB 0.02fF
C12466 S.n11304 SUB 0.24fF $ **FLOATING
C12467 S.n11305 SUB 0.36fF $ **FLOATING
C12468 S.n11306 SUB 0.61fF $ **FLOATING
C12469 S.n11307 SUB 0.12fF $ **FLOATING
C12470 S.t2496 SUB 0.02fF
C12471 S.n11308 SUB 0.14fF $ **FLOATING
C12472 S.n11310 SUB 5.17fF $ **FLOATING
C12473 S.t2582 SUB 0.02fF
C12474 S.n11311 SUB 0.12fF $ **FLOATING
C12475 S.n11312 SUB 0.14fF $ **FLOATING
C12476 S.t2110 SUB 0.02fF
C12477 S.n11314 SUB 0.24fF $ **FLOATING
C12478 S.n11315 SUB 0.91fF $ **FLOATING
C12479 S.n11316 SUB 0.05fF $ **FLOATING
C12480 S.n11317 SUB 1.88fF $ **FLOATING
C12481 S.n11318 SUB 2.67fF $ **FLOATING
C12482 S.t2201 SUB 0.02fF
C12483 S.n11319 SUB 0.24fF $ **FLOATING
C12484 S.n11320 SUB 0.36fF $ **FLOATING
C12485 S.n11321 SUB 0.61fF $ **FLOATING
C12486 S.n11322 SUB 0.12fF $ **FLOATING
C12487 S.t1619 SUB 0.02fF
C12488 S.n11323 SUB 0.14fF $ **FLOATING
C12489 S.n11325 SUB 5.17fF $ **FLOATING
C12490 S.t1704 SUB 0.02fF
C12491 S.n11326 SUB 0.12fF $ **FLOATING
C12492 S.n11327 SUB 0.14fF $ **FLOATING
C12493 S.t1241 SUB 0.02fF
C12494 S.n11329 SUB 0.24fF $ **FLOATING
C12495 S.n11330 SUB 0.91fF $ **FLOATING
C12496 S.n11331 SUB 0.05fF $ **FLOATING
C12497 S.n11332 SUB 1.88fF $ **FLOATING
C12498 S.n11333 SUB 2.67fF $ **FLOATING
C12499 S.t1344 SUB 0.02fF
C12500 S.n11334 SUB 0.24fF $ **FLOATING
C12501 S.n11335 SUB 0.36fF $ **FLOATING
C12502 S.n11336 SUB 0.61fF $ **FLOATING
C12503 S.n11337 SUB 0.12fF $ **FLOATING
C12504 S.t752 SUB 0.02fF
C12505 S.n11338 SUB 0.14fF $ **FLOATING
C12506 S.n11340 SUB 5.17fF $ **FLOATING
C12507 S.t835 SUB 0.02fF
C12508 S.n11341 SUB 0.12fF $ **FLOATING
C12509 S.n11342 SUB 0.14fF $ **FLOATING
C12510 S.t359 SUB 0.02fF
C12511 S.n11344 SUB 0.24fF $ **FLOATING
C12512 S.n11345 SUB 0.91fF $ **FLOATING
C12513 S.n11346 SUB 0.05fF $ **FLOATING
C12514 S.n11347 SUB 1.88fF $ **FLOATING
C12515 S.n11348 SUB 2.67fF $ **FLOATING
C12516 S.t465 SUB 0.02fF
C12517 S.n11349 SUB 0.24fF $ **FLOATING
C12518 S.n11350 SUB 0.36fF $ **FLOATING
C12519 S.n11351 SUB 0.61fF $ **FLOATING
C12520 S.n11352 SUB 0.12fF $ **FLOATING
C12521 S.t2408 SUB 0.02fF
C12522 S.n11353 SUB 0.14fF $ **FLOATING
C12523 S.n11355 SUB 4.90fF $ **FLOATING
C12524 S.t2481 SUB 0.02fF
C12525 S.n11356 SUB 0.12fF $ **FLOATING
C12526 S.n11357 SUB 0.14fF $ **FLOATING
C12527 S.t2013 SUB 0.02fF
C12528 S.n11359 SUB 0.24fF $ **FLOATING
C12529 S.n11360 SUB 0.91fF $ **FLOATING
C12530 S.n11361 SUB 0.05fF $ **FLOATING
C12531 S.n11362 SUB 1.88fF $ **FLOATING
C12532 S.n11363 SUB 2.67fF $ **FLOATING
C12533 S.t906 SUB 0.02fF
C12534 S.n11364 SUB 0.24fF $ **FLOATING
C12535 S.n11365 SUB 0.36fF $ **FLOATING
C12536 S.n11366 SUB 0.61fF $ **FLOATING
C12537 S.n11367 SUB 0.12fF $ **FLOATING
C12538 S.t2155 SUB 0.02fF
C12539 S.n11368 SUB 0.14fF $ **FLOATING
C12540 S.n11370 SUB 1.88fF $ **FLOATING
C12541 S.n11371 SUB 2.68fF $ **FLOATING
C12542 S.t1012 SUB 0.02fF
C12543 S.n11372 SUB 0.24fF $ **FLOATING
C12544 S.n11373 SUB 0.36fF $ **FLOATING
C12545 S.n11374 SUB 0.61fF $ **FLOATING
C12546 S.t567 SUB 0.02fF
C12547 S.n11375 SUB 1.22fF $ **FLOATING
C12548 S.n11376 SUB 0.42fF $ **FLOATING
C12549 S.n11377 SUB 0.44fF $ **FLOATING
C12550 S.n11378 SUB 0.36fF $ **FLOATING
C12551 S.n11379 SUB 0.21fF $ **FLOATING
C12552 S.n11380 SUB 0.25fF $ **FLOATING
C12553 S.n11381 SUB 1.28fF $ **FLOATING
C12554 S.n11382 SUB 0.35fF $ **FLOATING
C12555 S.n11383 SUB 0.63fF $ **FLOATING
C12556 S.n11384 SUB 1.15fF $ **FLOATING
C12557 S.n11385 SUB 3.03fF $ **FLOATING
C12558 S.n11386 SUB 0.59fF $ **FLOATING
C12559 S.n11387 SUB 0.02fF $ **FLOATING
C12560 S.n11388 SUB 0.97fF $ **FLOATING
C12561 S.t208 SUB 21.38fF
C12562 S.n11389 SUB 20.25fF $ **FLOATING
C12563 S.n11391 SUB 0.38fF $ **FLOATING
C12564 S.n11392 SUB 0.23fF $ **FLOATING
C12565 S.n11393 SUB 2.82fF $ **FLOATING
C12566 S.n11394 SUB 2.00fF $ **FLOATING
C12567 S.n11395 SUB 4.08fF $ **FLOATING
C12568 S.n11396 SUB 0.25fF $ **FLOATING
C12569 S.n11397 SUB 0.01fF $ **FLOATING
C12570 S.t260 SUB 0.02fF
C12571 S.n11398 SUB 0.25fF $ **FLOATING
C12572 S.t2243 SUB 0.02fF
C12573 S.n11399 SUB 0.95fF $ **FLOATING
C12574 S.n11400 SUB 0.70fF $ **FLOATING
C12575 S.n11401 SUB 0.78fF $ **FLOATING
C12576 S.n11402 SUB 2.26fF $ **FLOATING
C12577 S.n11403 SUB 1.88fF $ **FLOATING
C12578 S.n11404 SUB 0.12fF $ **FLOATING
C12579 S.t1926 SUB 0.02fF
C12580 S.n11405 SUB 0.14fF $ **FLOATING
C12581 S.t2210 SUB 0.02fF
C12582 S.n11407 SUB 0.24fF $ **FLOATING
C12583 S.n11408 SUB 0.36fF $ **FLOATING
C12584 S.n11409 SUB 0.61fF $ **FLOATING
C12585 S.n11410 SUB 1.39fF $ **FLOATING
C12586 S.n11411 SUB 0.71fF $ **FLOATING
C12587 S.n11412 SUB 1.14fF $ **FLOATING
C12588 S.n11413 SUB 0.35fF $ **FLOATING
C12589 S.n11414 SUB 2.03fF $ **FLOATING
C12590 S.t1384 SUB 0.02fF
C12591 S.n11415 SUB 0.24fF $ **FLOATING
C12592 S.n11416 SUB 0.91fF $ **FLOATING
C12593 S.n11417 SUB 0.05fF $ **FLOATING
C12594 S.t2588 SUB 0.02fF
C12595 S.n11418 SUB 0.12fF $ **FLOATING
C12596 S.n11419 SUB 0.14fF $ **FLOATING
C12597 S.n11421 SUB 1.89fF $ **FLOATING
C12598 S.n11422 SUB 1.88fF $ **FLOATING
C12599 S.t1349 SUB 0.02fF
C12600 S.n11423 SUB 0.24fF $ **FLOATING
C12601 S.n11424 SUB 0.36fF $ **FLOATING
C12602 S.n11425 SUB 0.61fF $ **FLOATING
C12603 S.n11426 SUB 0.12fF $ **FLOATING
C12604 S.t1066 SUB 0.02fF
C12605 S.n11427 SUB 0.14fF $ **FLOATING
C12606 S.n11429 SUB 1.16fF $ **FLOATING
C12607 S.n11430 SUB 0.22fF $ **FLOATING
C12608 S.n11431 SUB 0.25fF $ **FLOATING
C12609 S.n11432 SUB 0.09fF $ **FLOATING
C12610 S.n11433 SUB 1.88fF $ **FLOATING
C12611 S.t512 SUB 0.02fF
C12612 S.n11434 SUB 0.24fF $ **FLOATING
C12613 S.n11435 SUB 0.91fF $ **FLOATING
C12614 S.n11436 SUB 0.05fF $ **FLOATING
C12615 S.t1712 SUB 0.02fF
C12616 S.n11437 SUB 0.12fF $ **FLOATING
C12617 S.n11438 SUB 0.14fF $ **FLOATING
C12618 S.n11440 SUB 20.78fF $ **FLOATING
C12619 S.n11441 SUB 1.88fF $ **FLOATING
C12620 S.n11442 SUB 2.67fF $ **FLOATING
C12621 S.t1252 SUB 0.02fF
C12622 S.n11443 SUB 0.24fF $ **FLOATING
C12623 S.n11444 SUB 0.36fF $ **FLOATING
C12624 S.n11445 SUB 0.61fF $ **FLOATING
C12625 S.n11446 SUB 0.12fF $ **FLOATING
C12626 S.t986 SUB 0.02fF
C12627 S.n11447 SUB 0.14fF $ **FLOATING
C12628 S.n11449 SUB 2.80fF $ **FLOATING
C12629 S.n11450 SUB 2.30fF $ **FLOATING
C12630 S.t1768 SUB 0.02fF
C12631 S.n11451 SUB 0.12fF $ **FLOATING
C12632 S.n11452 SUB 0.14fF $ **FLOATING
C12633 S.t409 SUB 0.02fF
C12634 S.n11454 SUB 0.24fF $ **FLOATING
C12635 S.n11455 SUB 0.91fF $ **FLOATING
C12636 S.n11456 SUB 0.05fF $ **FLOATING
C12637 S.n11457 SUB 1.88fF $ **FLOATING
C12638 S.n11458 SUB 2.67fF $ **FLOATING
C12639 S.t370 SUB 0.02fF
C12640 S.n11459 SUB 0.24fF $ **FLOATING
C12641 S.n11460 SUB 0.36fF $ **FLOATING
C12642 S.n11461 SUB 0.61fF $ **FLOATING
C12643 S.n11462 SUB 0.12fF $ **FLOATING
C12644 S.t66 SUB 0.02fF
C12645 S.n11463 SUB 0.14fF $ **FLOATING
C12646 S.n11465 SUB 2.80fF $ **FLOATING
C12647 S.n11466 SUB 2.30fF $ **FLOATING
C12648 S.t894 SUB 0.02fF
C12649 S.n11467 SUB 0.12fF $ **FLOATING
C12650 S.n11468 SUB 0.14fF $ **FLOATING
C12651 S.t2056 SUB 0.02fF
C12652 S.n11470 SUB 0.24fF $ **FLOATING
C12653 S.n11471 SUB 0.91fF $ **FLOATING
C12654 S.n11472 SUB 0.05fF $ **FLOATING
C12655 S.n11473 SUB 1.88fF $ **FLOATING
C12656 S.n11474 SUB 2.67fF $ **FLOATING
C12657 S.t2021 SUB 0.02fF
C12658 S.n11475 SUB 0.24fF $ **FLOATING
C12659 S.n11476 SUB 0.36fF $ **FLOATING
C12660 S.n11477 SUB 0.61fF $ **FLOATING
C12661 S.n11478 SUB 0.12fF $ **FLOATING
C12662 S.t1894 SUB 0.02fF
C12663 S.n11479 SUB 0.14fF $ **FLOATING
C12664 S.n11481 SUB 2.80fF $ **FLOATING
C12665 S.n11482 SUB 2.30fF $ **FLOATING
C12666 S.t2536 SUB 0.02fF
C12667 S.n11483 SUB 0.12fF $ **FLOATING
C12668 S.n11484 SUB 0.14fF $ **FLOATING
C12669 S.t1196 SUB 0.02fF
C12670 S.n11486 SUB 0.24fF $ **FLOATING
C12671 S.n11487 SUB 0.91fF $ **FLOATING
C12672 S.n11488 SUB 0.05fF $ **FLOATING
C12673 S.n11489 SUB 1.88fF $ **FLOATING
C12674 S.n11490 SUB 2.67fF $ **FLOATING
C12675 S.t352 SUB 0.02fF
C12676 S.n11491 SUB 0.24fF $ **FLOATING
C12677 S.n11492 SUB 0.36fF $ **FLOATING
C12678 S.n11493 SUB 0.61fF $ **FLOATING
C12679 S.n11494 SUB 0.12fF $ **FLOATING
C12680 S.t1123 SUB 0.02fF
C12681 S.n11495 SUB 0.14fF $ **FLOATING
C12682 S.n11497 SUB 2.80fF $ **FLOATING
C12683 S.n11498 SUB 2.30fF $ **FLOATING
C12684 S.t1663 SUB 0.02fF
C12685 S.n11499 SUB 0.12fF $ **FLOATING
C12686 S.n11500 SUB 0.14fF $ **FLOATING
C12687 S.t2166 SUB 0.02fF
C12688 S.n11502 SUB 0.24fF $ **FLOATING
C12689 S.n11503 SUB 0.91fF $ **FLOATING
C12690 S.n11504 SUB 0.05fF $ **FLOATING
C12691 S.n11505 SUB 1.88fF $ **FLOATING
C12692 S.n11506 SUB 2.67fF $ **FLOATING
C12693 S.t2009 SUB 0.02fF
C12694 S.n11507 SUB 0.24fF $ **FLOATING
C12695 S.n11508 SUB 0.36fF $ **FLOATING
C12696 S.n11509 SUB 0.61fF $ **FLOATING
C12697 S.n11510 SUB 0.12fF $ **FLOATING
C12698 S.t246 SUB 0.02fF
C12699 S.n11511 SUB 0.14fF $ **FLOATING
C12700 S.n11513 SUB 2.80fF $ **FLOATING
C12701 S.n11514 SUB 2.30fF $ **FLOATING
C12702 S.t922 SUB 0.02fF
C12703 S.n11515 SUB 0.12fF $ **FLOATING
C12704 S.n11516 SUB 0.14fF $ **FLOATING
C12705 S.t1304 SUB 0.02fF
C12706 S.n11518 SUB 0.24fF $ **FLOATING
C12707 S.n11519 SUB 0.91fF $ **FLOATING
C12708 S.n11520 SUB 0.05fF $ **FLOATING
C12709 S.n11521 SUB 1.88fF $ **FLOATING
C12710 S.n11522 SUB 2.67fF $ **FLOATING
C12711 S.t1157 SUB 0.02fF
C12712 S.n11523 SUB 0.24fF $ **FLOATING
C12713 S.n11524 SUB 0.36fF $ **FLOATING
C12714 S.n11525 SUB 0.61fF $ **FLOATING
C12715 S.n11526 SUB 0.12fF $ **FLOATING
C12716 S.t1911 SUB 0.02fF
C12717 S.n11527 SUB 0.14fF $ **FLOATING
C12718 S.n11529 SUB 2.80fF $ **FLOATING
C12719 S.n11530 SUB 2.30fF $ **FLOATING
C12720 S.t2559 SUB 0.02fF
C12721 S.n11531 SUB 0.12fF $ **FLOATING
C12722 S.n11532 SUB 0.14fF $ **FLOATING
C12723 S.t420 SUB 0.02fF
C12724 S.n11534 SUB 0.24fF $ **FLOATING
C12725 S.n11535 SUB 0.91fF $ **FLOATING
C12726 S.n11536 SUB 0.05fF $ **FLOATING
C12727 S.n11537 SUB 1.88fF $ **FLOATING
C12728 S.n11538 SUB 2.67fF $ **FLOATING
C12729 S.t283 SUB 0.02fF
C12730 S.n11539 SUB 0.24fF $ **FLOATING
C12731 S.n11540 SUB 0.36fF $ **FLOATING
C12732 S.n11541 SUB 0.61fF $ **FLOATING
C12733 S.n11542 SUB 0.12fF $ **FLOATING
C12734 S.t1052 SUB 0.02fF
C12735 S.n11543 SUB 0.14fF $ **FLOATING
C12736 S.n11545 SUB 2.80fF $ **FLOATING
C12737 S.n11546 SUB 2.30fF $ **FLOATING
C12738 S.t1686 SUB 0.02fF
C12739 S.n11547 SUB 0.12fF $ **FLOATING
C12740 S.n11548 SUB 0.14fF $ **FLOATING
C12741 S.t2071 SUB 0.02fF
C12742 S.n11550 SUB 0.24fF $ **FLOATING
C12743 S.n11551 SUB 0.91fF $ **FLOATING
C12744 S.n11552 SUB 0.05fF $ **FLOATING
C12745 S.n11553 SUB 1.88fF $ **FLOATING
C12746 S.n11554 SUB 2.67fF $ **FLOATING
C12747 S.t1944 SUB 0.02fF
C12748 S.n11555 SUB 0.24fF $ **FLOATING
C12749 S.n11556 SUB 0.36fF $ **FLOATING
C12750 S.n11557 SUB 0.61fF $ **FLOATING
C12751 S.n11558 SUB 0.12fF $ **FLOATING
C12752 S.t164 SUB 0.02fF
C12753 S.n11559 SUB 0.14fF $ **FLOATING
C12754 S.n11561 SUB 2.80fF $ **FLOATING
C12755 S.n11562 SUB 2.30fF $ **FLOATING
C12756 S.t813 SUB 0.02fF
C12757 S.n11563 SUB 0.12fF $ **FLOATING
C12758 S.n11564 SUB 0.14fF $ **FLOATING
C12759 S.t1210 SUB 0.02fF
C12760 S.n11566 SUB 0.24fF $ **FLOATING
C12761 S.n11567 SUB 0.91fF $ **FLOATING
C12762 S.n11568 SUB 0.05fF $ **FLOATING
C12763 S.n11569 SUB 1.88fF $ **FLOATING
C12764 S.n11570 SUB 2.67fF $ **FLOATING
C12765 S.t1087 SUB 0.02fF
C12766 S.n11571 SUB 0.24fF $ **FLOATING
C12767 S.n11572 SUB 0.36fF $ **FLOATING
C12768 S.n11573 SUB 0.61fF $ **FLOATING
C12769 S.n11574 SUB 0.12fF $ **FLOATING
C12770 S.t1827 SUB 0.02fF
C12771 S.n11575 SUB 0.14fF $ **FLOATING
C12772 S.n11577 SUB 2.80fF $ **FLOATING
C12773 S.n11578 SUB 2.30fF $ **FLOATING
C12774 S.t50 SUB 0.02fF
C12775 S.n11579 SUB 0.12fF $ **FLOATING
C12776 S.n11580 SUB 0.14fF $ **FLOATING
C12777 S.t331 SUB 0.02fF
C12778 S.n11582 SUB 0.24fF $ **FLOATING
C12779 S.n11583 SUB 0.91fF $ **FLOATING
C12780 S.n11584 SUB 0.05fF $ **FLOATING
C12781 S.n11585 SUB 1.88fF $ **FLOATING
C12782 S.n11586 SUB 2.67fF $ **FLOATING
C12783 S.t209 SUB 0.02fF
C12784 S.n11587 SUB 0.24fF $ **FLOATING
C12785 S.n11588 SUB 0.36fF $ **FLOATING
C12786 S.n11589 SUB 0.61fF $ **FLOATING
C12787 S.n11590 SUB 0.12fF $ **FLOATING
C12788 S.t959 SUB 0.02fF
C12789 S.n11591 SUB 0.14fF $ **FLOATING
C12790 S.n11593 SUB 2.80fF $ **FLOATING
C12791 S.n11594 SUB 2.30fF $ **FLOATING
C12792 S.t1744 SUB 0.02fF
C12793 S.n11595 SUB 0.12fF $ **FLOATING
C12794 S.n11596 SUB 0.14fF $ **FLOATING
C12795 S.t1988 SUB 0.02fF
C12796 S.n11598 SUB 0.24fF $ **FLOATING
C12797 S.n11599 SUB 0.91fF $ **FLOATING
C12798 S.n11600 SUB 0.05fF $ **FLOATING
C12799 S.n11601 SUB 1.88fF $ **FLOATING
C12800 S.n11602 SUB 2.67fF $ **FLOATING
C12801 S.t1877 SUB 0.02fF
C12802 S.n11603 SUB 0.24fF $ **FLOATING
C12803 S.n11604 SUB 0.36fF $ **FLOATING
C12804 S.n11605 SUB 0.61fF $ **FLOATING
C12805 S.n11606 SUB 0.12fF $ **FLOATING
C12806 S.t19 SUB 0.02fF
C12807 S.n11607 SUB 0.14fF $ **FLOATING
C12808 S.n11609 SUB 2.80fF $ **FLOATING
C12809 S.n11610 SUB 2.30fF $ **FLOATING
C12810 S.t868 SUB 0.02fF
C12811 S.n11611 SUB 0.12fF $ **FLOATING
C12812 S.n11612 SUB 0.14fF $ **FLOATING
C12813 S.t1138 SUB 0.02fF
C12814 S.n11614 SUB 0.24fF $ **FLOATING
C12815 S.n11615 SUB 0.91fF $ **FLOATING
C12816 S.n11616 SUB 0.05fF $ **FLOATING
C12817 S.n11617 SUB 0.12fF $ **FLOATING
C12818 S.t71 SUB 0.02fF
C12819 S.n11618 SUB 0.14fF $ **FLOATING
C12820 S.t1335 SUB 0.02fF
C12821 S.n11620 SUB 0.24fF $ **FLOATING
C12822 S.n11621 SUB 0.36fF $ **FLOATING
C12823 S.n11622 SUB 0.61fF $ **FLOATING
C12824 S.n11623 SUB 1.60fF $ **FLOATING
C12825 S.n11624 SUB 0.03fF $ **FLOATING
C12826 S.n11625 SUB 0.14fF $ **FLOATING
C12827 S.n11626 SUB 0.58fF $ **FLOATING
C12828 S.n11627 SUB 0.12fF $ **FLOATING
C12829 S.n11628 SUB 0.53fF $ **FLOATING
C12830 S.n11629 SUB 0.41fF $ **FLOATING
C12831 S.n11630 SUB 0.25fF $ **FLOATING
C12832 S.n11631 SUB 0.25fF $ **FLOATING
C12833 S.n11632 SUB 0.68fF $ **FLOATING
C12834 S.n11633 SUB 1.97fF $ **FLOATING
C12835 S.t832 SUB 0.02fF
C12836 S.n11634 SUB 0.12fF $ **FLOATING
C12837 S.n11635 SUB 0.14fF $ **FLOATING
C12838 S.t2294 SUB 0.02fF
C12839 S.n11637 SUB 0.24fF $ **FLOATING
C12840 S.n11638 SUB 0.91fF $ **FLOATING
C12841 S.n11639 SUB 0.05fF $ **FLOATING
C12842 S.t18 SUB 48.31fF
C12843 S.t262 SUB 0.02fF
C12844 S.n11640 SUB 0.24fF $ **FLOATING
C12845 S.n11641 SUB 0.91fF $ **FLOATING
C12846 S.n11642 SUB 0.05fF $ **FLOATING
C12847 S.t2513 SUB 0.02fF
C12848 S.n11643 SUB 0.12fF $ **FLOATING
C12849 S.n11644 SUB 0.14fF $ **FLOATING
C12850 S.n11646 SUB 0.12fF $ **FLOATING
C12851 S.t1726 SUB 0.02fF
C12852 S.n11647 SUB 0.14fF $ **FLOATING
C12853 S.n11649 SUB 5.17fF $ **FLOATING
C12854 S.n11650 SUB 5.44fF $ **FLOATING
C12855 S.t1607 SUB 0.02fF
C12856 S.n11651 SUB 0.12fF $ **FLOATING
C12857 S.n11652 SUB 0.14fF $ **FLOATING
C12858 S.t307 SUB 0.02fF
C12859 S.n11654 SUB 0.24fF $ **FLOATING
C12860 S.n11655 SUB 0.91fF $ **FLOATING
C12861 S.n11656 SUB 0.05fF $ **FLOATING
C12862 S.t12 SUB 47.92fF
C12863 S.t2081 SUB 0.02fF
C12864 S.n11657 SUB 1.19fF $ **FLOATING
C12865 S.n11658 SUB 0.05fF $ **FLOATING
C12866 S.t1422 SUB 0.02fF
C12867 S.n11659 SUB 0.01fF $ **FLOATING
C12868 S.n11660 SUB 0.26fF $ **FLOATING
C12869 S.n11662 SUB 1.50fF $ **FLOATING
C12870 S.n11663 SUB 1.26fF $ **FLOATING
C12871 S.n11664 SUB 0.28fF $ **FLOATING
C12872 S.n11665 SUB 0.24fF $ **FLOATING
C12873 S.n11666 SUB 4.38fF $ **FLOATING
C12874 S.n11667 SUB 1.89fF $ **FLOATING
C12875 S.n11668 SUB 0.06fF $ **FLOATING
C12876 S.n11669 SUB 0.03fF $ **FLOATING
C12877 S.n11670 SUB 0.04fF $ **FLOATING
C12878 S.n11671 SUB 0.99fF $ **FLOATING
C12879 S.n11672 SUB 0.02fF $ **FLOATING
C12880 S.n11673 SUB 0.01fF $ **FLOATING
C12881 S.n11674 SUB 0.02fF $ **FLOATING
C12882 S.n11675 SUB 0.08fF $ **FLOATING
C12883 S.n11676 SUB 0.36fF $ **FLOATING
C12884 S.n11677 SUB 1.85fF $ **FLOATING
C12885 S.t276 SUB 0.02fF
C12886 S.n11678 SUB 0.24fF $ **FLOATING
C12887 S.n11679 SUB 0.36fF $ **FLOATING
C12888 S.n11680 SUB 0.61fF $ **FLOATING
C12889 S.n11681 SUB 0.12fF $ **FLOATING
C12890 S.t2278 SUB 0.02fF
C12891 S.n11682 SUB 0.14fF $ **FLOATING
C12892 S.n11684 SUB 0.70fF $ **FLOATING
C12893 S.n11685 SUB 0.23fF $ **FLOATING
C12894 S.n11686 SUB 0.23fF $ **FLOATING
C12895 S.n11687 SUB 0.70fF $ **FLOATING
C12896 S.n11688 SUB 1.16fF $ **FLOATING
C12897 S.n11689 SUB 0.22fF $ **FLOATING
C12898 S.n11690 SUB 0.25fF $ **FLOATING
C12899 S.n11691 SUB 0.09fF $ **FLOATING
C12900 S.n11692 SUB 1.88fF $ **FLOATING
C12901 S.t1419 SUB 0.02fF
C12902 S.n11693 SUB 0.24fF $ **FLOATING
C12903 S.n11694 SUB 0.91fF $ **FLOATING
C12904 S.n11695 SUB 0.05fF $ **FLOATING
C12905 S.t2434 SUB 0.02fF
C12906 S.n11696 SUB 0.12fF $ **FLOATING
C12907 S.n11697 SUB 0.14fF $ **FLOATING
C12908 S.n11699 SUB 20.78fF $ **FLOATING
C12909 S.n11700 SUB 0.09fF $ **FLOATING
C12910 S.n11701 SUB 0.21fF $ **FLOATING
C12911 S.n11702 SUB 0.07fF $ **FLOATING
C12912 S.n11703 SUB 0.06fF $ **FLOATING
C12913 S.n11704 SUB 0.07fF $ **FLOATING
C12914 S.n11705 SUB 0.18fF $ **FLOATING
C12915 S.n11706 SUB 0.20fF $ **FLOATING
C12916 S.n11707 SUB 1.04fF $ **FLOATING
C12917 S.n11708 SUB 0.54fF $ **FLOATING
C12918 S.n11709 SUB 2.34fF $ **FLOATING
C12919 S.n11710 SUB 0.12fF $ **FLOATING
C12920 S.t620 SUB 0.02fF
C12921 S.n11711 SUB 0.14fF $ **FLOATING
C12922 S.t1152 SUB 0.02fF
C12923 S.n11713 SUB 0.24fF $ **FLOATING
C12924 S.n11714 SUB 0.36fF $ **FLOATING
C12925 S.n11715 SUB 0.61fF $ **FLOATING
C12926 S.n11716 SUB 1.73fF $ **FLOATING
C12927 S.n11717 SUB 2.44fF $ **FLOATING
C12928 S.t784 SUB 0.02fF
C12929 S.n11718 SUB 0.12fF $ **FLOATING
C12930 S.n11719 SUB 0.14fF $ **FLOATING
C12931 S.t2275 SUB 0.02fF
C12932 S.n11721 SUB 0.24fF $ **FLOATING
C12933 S.n11722 SUB 0.91fF $ **FLOATING
C12934 S.n11723 SUB 0.05fF $ **FLOATING
C12935 S.n11724 SUB 2.94fF $ **FLOATING
C12936 S.n11725 SUB 1.88fF $ **FLOATING
C12937 S.n11726 SUB 0.12fF $ **FLOATING
C12938 S.t1516 SUB 0.02fF
C12939 S.n11727 SUB 0.14fF $ **FLOATING
C12940 S.t2047 SUB 0.02fF
C12941 S.n11729 SUB 0.24fF $ **FLOATING
C12942 S.n11730 SUB 0.36fF $ **FLOATING
C12943 S.n11731 SUB 0.61fF $ **FLOATING
C12944 S.n11732 SUB 0.92fF $ **FLOATING
C12945 S.n11733 SUB 0.32fF $ **FLOATING
C12946 S.n11734 SUB 0.92fF $ **FLOATING
C12947 S.n11735 SUB 1.09fF $ **FLOATING
C12948 S.n11736 SUB 0.15fF $ **FLOATING
C12949 S.n11737 SUB 4.96fF $ **FLOATING
C12950 S.t1570 SUB 0.02fF
C12951 S.n11738 SUB 0.12fF $ **FLOATING
C12952 S.n11739 SUB 0.14fF $ **FLOATING
C12953 S.t653 SUB 0.02fF
C12954 S.n11741 SUB 0.24fF $ **FLOATING
C12955 S.n11742 SUB 0.91fF $ **FLOATING
C12956 S.n11743 SUB 0.05fF $ **FLOATING
C12957 S.n11744 SUB 1.88fF $ **FLOATING
C12958 S.n11745 SUB 2.67fF $ **FLOATING
C12959 S.t1189 SUB 0.02fF
C12960 S.n11746 SUB 0.24fF $ **FLOATING
C12961 S.n11747 SUB 0.36fF $ **FLOATING
C12962 S.n11748 SUB 0.61fF $ **FLOATING
C12963 S.n11749 SUB 0.12fF $ **FLOATING
C12964 S.t655 SUB 0.02fF
C12965 S.n11750 SUB 0.14fF $ **FLOATING
C12966 S.n11752 SUB 2.94fF $ **FLOATING
C12967 S.n11753 SUB 5.16fF $ **FLOATING
C12968 S.t702 SUB 0.02fF
C12969 S.n11754 SUB 0.12fF $ **FLOATING
C12970 S.n11755 SUB 0.14fF $ **FLOATING
C12971 S.t2307 SUB 0.02fF
C12972 S.n11757 SUB 0.24fF $ **FLOATING
C12973 S.n11758 SUB 0.91fF $ **FLOATING
C12974 S.n11759 SUB 0.05fF $ **FLOATING
C12975 S.n11760 SUB 1.88fF $ **FLOATING
C12976 S.n11761 SUB 2.67fF $ **FLOATING
C12977 S.t313 SUB 0.02fF
C12978 S.n11762 SUB 0.24fF $ **FLOATING
C12979 S.n11763 SUB 0.36fF $ **FLOATING
C12980 S.n11764 SUB 0.61fF $ **FLOATING
C12981 S.n11765 SUB 0.12fF $ **FLOATING
C12982 S.t2309 SUB 0.02fF
C12983 S.n11766 SUB 0.14fF $ **FLOATING
C12984 S.n11768 SUB 5.17fF $ **FLOATING
C12985 S.t2361 SUB 0.02fF
C12986 S.n11769 SUB 0.12fF $ **FLOATING
C12987 S.n11770 SUB 0.14fF $ **FLOATING
C12988 S.t1451 SUB 0.02fF
C12989 S.n11772 SUB 0.24fF $ **FLOATING
C12990 S.n11773 SUB 0.91fF $ **FLOATING
C12991 S.n11774 SUB 0.05fF $ **FLOATING
C12992 S.n11775 SUB 1.88fF $ **FLOATING
C12993 S.n11776 SUB 2.67fF $ **FLOATING
C12994 S.t1977 SUB 0.02fF
C12995 S.n11777 SUB 0.24fF $ **FLOATING
C12996 S.n11778 SUB 0.36fF $ **FLOATING
C12997 S.n11779 SUB 0.61fF $ **FLOATING
C12998 S.n11780 SUB 0.12fF $ **FLOATING
C12999 S.t1452 SUB 0.02fF
C13000 S.n11781 SUB 0.14fF $ **FLOATING
C13001 S.n11783 SUB 5.17fF $ **FLOATING
C13002 S.t1505 SUB 0.02fF
C13003 S.n11784 SUB 0.12fF $ **FLOATING
C13004 S.n11785 SUB 0.14fF $ **FLOATING
C13005 S.t590 SUB 0.02fF
C13006 S.n11787 SUB 0.24fF $ **FLOATING
C13007 S.n11788 SUB 0.91fF $ **FLOATING
C13008 S.n11789 SUB 0.05fF $ **FLOATING
C13009 S.n11790 SUB 1.88fF $ **FLOATING
C13010 S.n11791 SUB 2.67fF $ **FLOATING
C13011 S.t1124 SUB 0.02fF
C13012 S.n11792 SUB 0.24fF $ **FLOATING
C13013 S.n11793 SUB 0.36fF $ **FLOATING
C13014 S.n11794 SUB 0.61fF $ **FLOATING
C13015 S.n11795 SUB 0.12fF $ **FLOATING
C13016 S.t594 SUB 0.02fF
C13017 S.n11796 SUB 0.14fF $ **FLOATING
C13018 S.n11798 SUB 5.17fF $ **FLOATING
C13019 S.t644 SUB 0.02fF
C13020 S.n11799 SUB 0.12fF $ **FLOATING
C13021 S.n11800 SUB 0.14fF $ **FLOATING
C13022 S.t2240 SUB 0.02fF
C13023 S.n11802 SUB 0.24fF $ **FLOATING
C13024 S.n11803 SUB 0.91fF $ **FLOATING
C13025 S.n11804 SUB 0.05fF $ **FLOATING
C13026 S.n11805 SUB 1.88fF $ **FLOATING
C13027 S.n11806 SUB 2.67fF $ **FLOATING
C13028 S.t245 SUB 0.02fF
C13029 S.n11807 SUB 0.24fF $ **FLOATING
C13030 S.n11808 SUB 0.36fF $ **FLOATING
C13031 S.n11809 SUB 0.61fF $ **FLOATING
C13032 S.n11810 SUB 0.12fF $ **FLOATING
C13033 S.t2241 SUB 0.02fF
C13034 S.n11811 SUB 0.14fF $ **FLOATING
C13035 S.n11813 SUB 5.17fF $ **FLOATING
C13036 S.t2397 SUB 0.02fF
C13037 S.n11814 SUB 0.12fF $ **FLOATING
C13038 S.n11815 SUB 0.14fF $ **FLOATING
C13039 S.t1380 SUB 0.02fF
C13040 S.n11817 SUB 0.24fF $ **FLOATING
C13041 S.n11818 SUB 0.91fF $ **FLOATING
C13042 S.n11819 SUB 0.05fF $ **FLOATING
C13043 S.n11820 SUB 1.88fF $ **FLOATING
C13044 S.n11821 SUB 2.67fF $ **FLOATING
C13045 S.t538 SUB 0.02fF
C13046 S.n11822 SUB 0.24fF $ **FLOATING
C13047 S.n11823 SUB 0.36fF $ **FLOATING
C13048 S.n11824 SUB 0.61fF $ **FLOATING
C13049 S.n11825 SUB 0.12fF $ **FLOATING
C13050 S.t2472 SUB 0.02fF
C13051 S.n11826 SUB 0.14fF $ **FLOATING
C13052 S.n11828 SUB 5.17fF $ **FLOATING
C13053 S.t177 SUB 0.02fF
C13054 S.n11829 SUB 0.12fF $ **FLOATING
C13055 S.n11830 SUB 0.14fF $ **FLOATING
C13056 S.t2083 SUB 0.02fF
C13057 S.n11832 SUB 0.24fF $ **FLOATING
C13058 S.n11833 SUB 0.91fF $ **FLOATING
C13059 S.n11834 SUB 0.05fF $ **FLOATING
C13060 S.n11835 SUB 1.88fF $ **FLOATING
C13061 S.n11836 SUB 2.67fF $ **FLOATING
C13062 S.t2179 SUB 0.02fF
C13063 S.n11837 SUB 0.24fF $ **FLOATING
C13064 S.n11838 SUB 0.36fF $ **FLOATING
C13065 S.n11839 SUB 0.61fF $ **FLOATING
C13066 S.n11840 SUB 0.12fF $ **FLOATING
C13067 S.t1602 SUB 0.02fF
C13068 S.n11841 SUB 0.14fF $ **FLOATING
C13069 S.n11843 SUB 5.17fF $ **FLOATING
C13070 S.t1842 SUB 0.02fF
C13071 S.n11844 SUB 0.12fF $ **FLOATING
C13072 S.n11845 SUB 0.14fF $ **FLOATING
C13073 S.t1221 SUB 0.02fF
C13074 S.n11847 SUB 0.24fF $ **FLOATING
C13075 S.n11848 SUB 0.91fF $ **FLOATING
C13076 S.n11849 SUB 0.05fF $ **FLOATING
C13077 S.n11850 SUB 1.88fF $ **FLOATING
C13078 S.n11851 SUB 2.67fF $ **FLOATING
C13079 S.t1318 SUB 0.02fF
C13080 S.n11852 SUB 0.24fF $ **FLOATING
C13081 S.n11853 SUB 0.36fF $ **FLOATING
C13082 S.n11854 SUB 0.61fF $ **FLOATING
C13083 S.n11855 SUB 0.12fF $ **FLOATING
C13084 S.t738 SUB 0.02fF
C13085 S.n11856 SUB 0.14fF $ **FLOATING
C13086 S.n11858 SUB 5.17fF $ **FLOATING
C13087 S.t977 SUB 0.02fF
C13088 S.n11859 SUB 0.12fF $ **FLOATING
C13089 S.n11860 SUB 0.14fF $ **FLOATING
C13090 S.t340 SUB 0.02fF
C13091 S.n11862 SUB 0.24fF $ **FLOATING
C13092 S.n11863 SUB 0.91fF $ **FLOATING
C13093 S.n11864 SUB 0.05fF $ **FLOATING
C13094 S.n11865 SUB 1.88fF $ **FLOATING
C13095 S.n11866 SUB 2.67fF $ **FLOATING
C13096 S.t440 SUB 0.02fF
C13097 S.n11867 SUB 0.24fF $ **FLOATING
C13098 S.n11868 SUB 0.36fF $ **FLOATING
C13099 S.n11869 SUB 0.61fF $ **FLOATING
C13100 S.n11870 SUB 0.12fF $ **FLOATING
C13101 S.t2388 SUB 0.02fF
C13102 S.n11871 SUB 0.14fF $ **FLOATING
C13103 S.n11873 SUB 5.17fF $ **FLOATING
C13104 S.t45 SUB 0.02fF
C13105 S.n11874 SUB 0.12fF $ **FLOATING
C13106 S.n11875 SUB 0.14fF $ **FLOATING
C13107 S.t1998 SUB 0.02fF
C13108 S.n11877 SUB 0.24fF $ **FLOATING
C13109 S.n11878 SUB 0.91fF $ **FLOATING
C13110 S.n11879 SUB 0.05fF $ **FLOATING
C13111 S.n11880 SUB 1.88fF $ **FLOATING
C13112 S.n11881 SUB 2.67fF $ **FLOATING
C13113 S.t2231 SUB 0.02fF
C13114 S.n11882 SUB 0.24fF $ **FLOATING
C13115 S.n11883 SUB 0.36fF $ **FLOATING
C13116 S.n11884 SUB 0.61fF $ **FLOATING
C13117 S.n11885 SUB 0.12fF $ **FLOATING
C13118 S.t1653 SUB 0.02fF
C13119 S.n11886 SUB 0.14fF $ **FLOATING
C13120 S.n11888 SUB 5.17fF $ **FLOATING
C13121 S.t1738 SUB 0.02fF
C13122 S.n11889 SUB 0.12fF $ **FLOATING
C13123 S.n11890 SUB 0.14fF $ **FLOATING
C13124 S.t1275 SUB 0.02fF
C13125 S.n11892 SUB 0.24fF $ **FLOATING
C13126 S.n11893 SUB 0.91fF $ **FLOATING
C13127 S.n11894 SUB 0.05fF $ **FLOATING
C13128 S.n11895 SUB 1.88fF $ **FLOATING
C13129 S.n11896 SUB 2.67fF $ **FLOATING
C13130 S.t1367 SUB 0.02fF
C13131 S.n11897 SUB 0.24fF $ **FLOATING
C13132 S.n11898 SUB 0.36fF $ **FLOATING
C13133 S.n11899 SUB 0.61fF $ **FLOATING
C13134 S.n11900 SUB 0.12fF $ **FLOATING
C13135 S.t781 SUB 0.02fF
C13136 S.n11901 SUB 0.14fF $ **FLOATING
C13137 S.n11903 SUB 5.17fF $ **FLOATING
C13138 S.t863 SUB 0.02fF
C13139 S.n11904 SUB 0.12fF $ **FLOATING
C13140 S.n11905 SUB 0.14fF $ **FLOATING
C13141 S.t388 SUB 0.02fF
C13142 S.n11907 SUB 0.24fF $ **FLOATING
C13143 S.n11908 SUB 0.91fF $ **FLOATING
C13144 S.n11909 SUB 0.05fF $ **FLOATING
C13145 S.n11910 SUB 1.88fF $ **FLOATING
C13146 S.n11911 SUB 2.67fF $ **FLOATING
C13147 S.t495 SUB 0.02fF
C13148 S.n11912 SUB 0.24fF $ **FLOATING
C13149 S.n11913 SUB 0.36fF $ **FLOATING
C13150 S.n11914 SUB 0.61fF $ **FLOATING
C13151 S.n11915 SUB 0.12fF $ **FLOATING
C13152 S.t2432 SUB 0.02fF
C13153 S.n11916 SUB 0.14fF $ **FLOATING
C13154 S.n11918 SUB 5.17fF $ **FLOATING
C13155 S.t2510 SUB 0.02fF
C13156 S.n11919 SUB 0.12fF $ **FLOATING
C13157 S.n11920 SUB 0.14fF $ **FLOATING
C13158 S.t2038 SUB 0.02fF
C13159 S.n11922 SUB 0.24fF $ **FLOATING
C13160 S.n11923 SUB 0.91fF $ **FLOATING
C13161 S.n11924 SUB 0.05fF $ **FLOATING
C13162 S.n11925 SUB 1.88fF $ **FLOATING
C13163 S.n11926 SUB 2.67fF $ **FLOATING
C13164 S.t2141 SUB 0.02fF
C13165 S.n11927 SUB 0.24fF $ **FLOATING
C13166 S.n11928 SUB 0.36fF $ **FLOATING
C13167 S.n11929 SUB 0.61fF $ **FLOATING
C13168 S.n11930 SUB 0.12fF $ **FLOATING
C13169 S.t1569 SUB 0.02fF
C13170 S.n11931 SUB 0.14fF $ **FLOATING
C13171 S.n11933 SUB 4.90fF $ **FLOATING
C13172 S.t1635 SUB 0.02fF
C13173 S.n11934 SUB 0.12fF $ **FLOATING
C13174 S.n11935 SUB 0.14fF $ **FLOATING
C13175 S.t1183 SUB 0.02fF
C13176 S.n11937 SUB 0.24fF $ **FLOATING
C13177 S.n11938 SUB 0.91fF $ **FLOATING
C13178 S.n11939 SUB 0.05fF $ **FLOATING
C13179 S.n11940 SUB 0.11fF $ **FLOATING
C13180 S.n11941 SUB 0.12fF $ **FLOATING
C13181 S.n11942 SUB 0.09fF $ **FLOATING
C13182 S.n11943 SUB 0.12fF $ **FLOATING
C13183 S.n11944 SUB 0.18fF $ **FLOATING
C13184 S.n11945 SUB 1.88fF $ **FLOATING
C13185 S.n11946 SUB 0.12fF $ **FLOATING
C13186 S.t885 SUB 0.02fF
C13187 S.n11947 SUB 0.14fF $ **FLOATING
C13188 S.t258 SUB 0.02fF
C13189 S.n11949 SUB 1.22fF $ **FLOATING
C13190 S.n11950 SUB 0.06fF $ **FLOATING
C13191 S.n11951 SUB 0.10fF $ **FLOATING
C13192 S.n11952 SUB 0.60fF $ **FLOATING
C13193 S.n11953 SUB 0.35fF $ **FLOATING
C13194 S.n11954 SUB 0.63fF $ **FLOATING
C13195 S.n11955 SUB 1.15fF $ **FLOATING
C13196 S.n11956 SUB 3.03fF $ **FLOATING
C13197 S.n11957 SUB 0.59fF $ **FLOATING
C13198 S.n11958 SUB 0.02fF $ **FLOATING
C13199 S.n11959 SUB 0.97fF $ **FLOATING
C13200 S.t57 SUB 21.38fF
C13201 S.n11960 SUB 20.25fF $ **FLOATING
C13202 S.n11962 SUB 0.38fF $ **FLOATING
C13203 S.n11963 SUB 0.23fF $ **FLOATING
C13204 S.n11964 SUB 2.89fF $ **FLOATING
C13205 S.n11965 SUB 2.42fF $ **FLOATING
C13206 S.n11966 SUB 2.47fF $ **FLOATING
C13207 S.n11967 SUB 4.29fF $ **FLOATING
C13208 S.n11968 SUB 0.25fF $ **FLOATING
C13209 S.n11969 SUB 0.01fF $ **FLOATING
C13210 S.t2471 SUB 0.02fF
C13211 S.n11970 SUB 0.25fF $ **FLOATING
C13212 S.t1952 SUB 0.02fF
C13213 S.n11971 SUB 0.95fF $ **FLOATING
C13214 S.n11972 SUB 0.70fF $ **FLOATING
C13215 S.n11973 SUB 1.89fF $ **FLOATING
C13216 S.n11974 SUB 1.88fF $ **FLOATING
C13217 S.t1924 SUB 0.02fF
C13218 S.n11975 SUB 0.24fF $ **FLOATING
C13219 S.n11976 SUB 0.36fF $ **FLOATING
C13220 S.n11977 SUB 0.61fF $ **FLOATING
C13221 S.n11978 SUB 0.12fF $ **FLOATING
C13222 S.t1601 SUB 0.02fF
C13223 S.n11979 SUB 0.14fF $ **FLOATING
C13224 S.n11981 SUB 1.16fF $ **FLOATING
C13225 S.n11982 SUB 0.22fF $ **FLOATING
C13226 S.n11983 SUB 0.25fF $ **FLOATING
C13227 S.n11984 SUB 0.09fF $ **FLOATING
C13228 S.n11985 SUB 1.88fF $ **FLOATING
C13229 S.t1092 SUB 0.02fF
C13230 S.n11986 SUB 0.24fF $ **FLOATING
C13231 S.n11987 SUB 0.91fF $ **FLOATING
C13232 S.n11988 SUB 0.05fF $ **FLOATING
C13233 S.t2302 SUB 0.02fF
C13234 S.n11989 SUB 0.12fF $ **FLOATING
C13235 S.n11990 SUB 0.14fF $ **FLOATING
C13236 S.n11992 SUB 0.77fF $ **FLOATING
C13237 S.n11993 SUB 0.44fF $ **FLOATING
C13238 S.n11994 SUB 1.59fF $ **FLOATING
C13239 S.n11995 SUB 0.12fF $ **FLOATING
C13240 S.t1259 SUB 0.02fF
C13241 S.n11996 SUB 0.14fF $ **FLOATING
C13242 S.t2410 SUB 0.02fF
C13243 S.n11998 SUB 0.24fF $ **FLOATING
C13244 S.n11999 SUB 0.36fF $ **FLOATING
C13245 S.n12000 SUB 0.61fF $ **FLOATING
C13246 S.n12001 SUB 0.01fF $ **FLOATING
C13247 S.n12002 SUB 0.07fF $ **FLOATING
C13248 S.n12003 SUB 0.01fF $ **FLOATING
C13249 S.n12004 SUB 0.02fF $ **FLOATING
C13250 S.n12005 SUB 0.01fF $ **FLOATING
C13251 S.n12006 SUB 0.24fF $ **FLOATING
C13252 S.n12007 SUB 1.16fF $ **FLOATING
C13253 S.n12008 SUB 1.34fF $ **FLOATING
C13254 S.n12009 SUB 1.99fF $ **FLOATING
C13255 S.t887 SUB 0.02fF
C13256 S.n12010 SUB 0.24fF $ **FLOATING
C13257 S.n12011 SUB 0.91fF $ **FLOATING
C13258 S.n12012 SUB 0.05fF $ **FLOATING
C13259 S.t1991 SUB 0.02fF
C13260 S.n12013 SUB 0.12fF $ **FLOATING
C13261 S.n12014 SUB 0.14fF $ **FLOATING
C13262 S.n12016 SUB 20.78fF $ **FLOATING
C13263 S.n12017 SUB 1.88fF $ **FLOATING
C13264 S.n12018 SUB 0.12fF $ **FLOATING
C13265 S.t737 SUB 0.02fF
C13266 S.n12019 SUB 0.14fF $ **FLOATING
C13267 S.t1063 SUB 0.02fF
C13268 S.n12021 SUB 0.24fF $ **FLOATING
C13269 S.n12022 SUB 0.36fF $ **FLOATING
C13270 S.n12023 SUB 0.61fF $ **FLOATING
C13271 S.n12024 SUB 0.32fF $ **FLOATING
C13272 S.n12025 SUB 1.09fF $ **FLOATING
C13273 S.n12026 SUB 0.15fF $ **FLOATING
C13274 S.n12027 SUB 2.10fF $ **FLOATING
C13275 S.t1447 SUB 0.02fF
C13276 S.n12028 SUB 0.12fF $ **FLOATING
C13277 S.n12029 SUB 0.14fF $ **FLOATING
C13278 S.t214 SUB 0.02fF
C13279 S.n12031 SUB 0.24fF $ **FLOATING
C13280 S.n12032 SUB 0.91fF $ **FLOATING
C13281 S.n12033 SUB 0.05fF $ **FLOATING
C13282 S.n12034 SUB 1.88fF $ **FLOATING
C13283 S.n12035 SUB 2.67fF $ **FLOATING
C13284 S.t182 SUB 0.02fF
C13285 S.n12036 SUB 0.24fF $ **FLOATING
C13286 S.n12037 SUB 0.36fF $ **FLOATING
C13287 S.n12038 SUB 0.61fF $ **FLOATING
C13288 S.n12039 SUB 0.12fF $ **FLOATING
C13289 S.t2387 SUB 0.02fF
C13290 S.n12040 SUB 0.14fF $ **FLOATING
C13291 S.n12042 SUB 2.30fF $ **FLOATING
C13292 S.t679 SUB 0.02fF
C13293 S.n12043 SUB 0.12fF $ **FLOATING
C13294 S.n12044 SUB 0.14fF $ **FLOATING
C13295 S.t1883 SUB 0.02fF
C13296 S.n12046 SUB 0.24fF $ **FLOATING
C13297 S.n12047 SUB 0.91fF $ **FLOATING
C13298 S.n12048 SUB 0.05fF $ **FLOATING
C13299 S.n12049 SUB 1.88fF $ **FLOATING
C13300 S.n12050 SUB 2.67fF $ **FLOATING
C13301 S.t1845 SUB 0.02fF
C13302 S.n12051 SUB 0.24fF $ **FLOATING
C13303 S.n12052 SUB 0.36fF $ **FLOATING
C13304 S.n12053 SUB 0.61fF $ **FLOATING
C13305 S.n12054 SUB 0.12fF $ **FLOATING
C13306 S.t1529 SUB 0.02fF
C13307 S.n12055 SUB 0.14fF $ **FLOATING
C13308 S.n12057 SUB 2.80fF $ **FLOATING
C13309 S.n12058 SUB 2.30fF $ **FLOATING
C13310 S.t2339 SUB 0.02fF
C13311 S.n12059 SUB 0.12fF $ **FLOATING
C13312 S.n12060 SUB 0.14fF $ **FLOATING
C13313 S.t1020 SUB 0.02fF
C13314 S.n12062 SUB 0.24fF $ **FLOATING
C13315 S.n12063 SUB 0.91fF $ **FLOATING
C13316 S.n12064 SUB 0.05fF $ **FLOATING
C13317 S.n12065 SUB 1.88fF $ **FLOATING
C13318 S.n12066 SUB 2.67fF $ **FLOATING
C13319 S.t983 SUB 0.02fF
C13320 S.n12067 SUB 0.24fF $ **FLOATING
C13321 S.n12068 SUB 0.36fF $ **FLOATING
C13322 S.n12069 SUB 0.61fF $ **FLOATING
C13323 S.n12070 SUB 0.12fF $ **FLOATING
C13324 S.t671 SUB 0.02fF
C13325 S.n12071 SUB 0.14fF $ **FLOATING
C13326 S.n12073 SUB 2.80fF $ **FLOATING
C13327 S.n12074 SUB 2.30fF $ **FLOATING
C13328 S.t1479 SUB 0.02fF
C13329 S.n12075 SUB 0.12fF $ **FLOATING
C13330 S.n12076 SUB 0.14fF $ **FLOATING
C13331 S.t115 SUB 0.02fF
C13332 S.n12078 SUB 0.24fF $ **FLOATING
C13333 S.n12079 SUB 0.91fF $ **FLOATING
C13334 S.n12080 SUB 0.05fF $ **FLOATING
C13335 S.n12081 SUB 1.88fF $ **FLOATING
C13336 S.n12082 SUB 2.67fF $ **FLOATING
C13337 S.t58 SUB 0.02fF
C13338 S.n12083 SUB 0.24fF $ **FLOATING
C13339 S.n12084 SUB 0.36fF $ **FLOATING
C13340 S.n12085 SUB 0.61fF $ **FLOATING
C13341 S.n12086 SUB 0.12fF $ **FLOATING
C13342 S.t2326 SUB 0.02fF
C13343 S.n12087 SUB 0.14fF $ **FLOATING
C13344 S.n12089 SUB 2.80fF $ **FLOATING
C13345 S.n12090 SUB 2.30fF $ **FLOATING
C13346 S.t617 SUB 0.02fF
C13347 S.n12091 SUB 0.12fF $ **FLOATING
C13348 S.n12092 SUB 0.14fF $ **FLOATING
C13349 S.t1788 SUB 0.02fF
C13350 S.n12094 SUB 0.24fF $ **FLOATING
C13351 S.n12095 SUB 0.91fF $ **FLOATING
C13352 S.n12096 SUB 0.05fF $ **FLOATING
C13353 S.n12097 SUB 1.88fF $ **FLOATING
C13354 S.n12098 SUB 2.67fF $ **FLOATING
C13355 S.t1748 SUB 0.02fF
C13356 S.n12099 SUB 0.24fF $ **FLOATING
C13357 S.n12100 SUB 0.36fF $ **FLOATING
C13358 S.n12101 SUB 0.61fF $ **FLOATING
C13359 S.n12102 SUB 0.12fF $ **FLOATING
C13360 S.t1564 SUB 0.02fF
C13361 S.n12103 SUB 0.14fF $ **FLOATING
C13362 S.n12105 SUB 2.80fF $ **FLOATING
C13363 S.n12106 SUB 2.30fF $ **FLOATING
C13364 S.t2273 SUB 0.02fF
C13365 S.n12107 SUB 0.12fF $ **FLOATING
C13366 S.n12108 SUB 0.14fF $ **FLOATING
C13367 S.t917 SUB 0.02fF
C13368 S.n12110 SUB 0.24fF $ **FLOATING
C13369 S.n12111 SUB 0.91fF $ **FLOATING
C13370 S.n12112 SUB 0.05fF $ **FLOATING
C13371 S.n12113 SUB 1.88fF $ **FLOATING
C13372 S.n12114 SUB 2.67fF $ **FLOATING
C13373 S.t2034 SUB 0.02fF
C13374 S.n12115 SUB 0.24fF $ **FLOATING
C13375 S.n12116 SUB 0.36fF $ **FLOATING
C13376 S.n12117 SUB 0.61fF $ **FLOATING
C13377 S.n12118 SUB 0.12fF $ **FLOATING
C13378 S.t266 SUB 0.02fF
C13379 S.n12119 SUB 0.14fF $ **FLOATING
C13380 S.n12121 SUB 2.80fF $ **FLOATING
C13381 S.n12122 SUB 2.30fF $ **FLOATING
C13382 S.t1417 SUB 0.02fF
C13383 S.n12123 SUB 0.12fF $ **FLOATING
C13384 S.n12124 SUB 0.14fF $ **FLOATING
C13385 S.t1336 SUB 0.02fF
C13386 S.n12126 SUB 0.24fF $ **FLOATING
C13387 S.n12127 SUB 0.91fF $ **FLOATING
C13388 S.n12128 SUB 0.05fF $ **FLOATING
C13389 S.n12129 SUB 1.88fF $ **FLOATING
C13390 S.n12130 SUB 2.67fF $ **FLOATING
C13391 S.t1178 SUB 0.02fF
C13392 S.n12131 SUB 0.24fF $ **FLOATING
C13393 S.n12132 SUB 0.36fF $ **FLOATING
C13394 S.n12133 SUB 0.61fF $ **FLOATING
C13395 S.n12134 SUB 0.12fF $ **FLOATING
C13396 S.t1929 SUB 0.02fF
C13397 S.n12135 SUB 0.14fF $ **FLOATING
C13398 S.n12137 SUB 2.80fF $ **FLOATING
C13399 S.n12138 SUB 2.30fF $ **FLOATING
C13400 S.t3 SUB 0.02fF
C13401 S.n12139 SUB 0.12fF $ **FLOATING
C13402 S.n12140 SUB 0.14fF $ **FLOATING
C13403 S.t455 SUB 0.02fF
C13404 S.n12142 SUB 0.24fF $ **FLOATING
C13405 S.n12143 SUB 0.91fF $ **FLOATING
C13406 S.n12144 SUB 0.05fF $ **FLOATING
C13407 S.n12145 SUB 1.88fF $ **FLOATING
C13408 S.n12146 SUB 2.67fF $ **FLOATING
C13409 S.t301 SUB 0.02fF
C13410 S.n12147 SUB 0.24fF $ **FLOATING
C13411 S.n12148 SUB 0.36fF $ **FLOATING
C13412 S.n12149 SUB 0.61fF $ **FLOATING
C13413 S.n12150 SUB 0.12fF $ **FLOATING
C13414 S.t1070 SUB 0.02fF
C13415 S.n12151 SUB 0.14fF $ **FLOATING
C13416 S.n12153 SUB 2.80fF $ **FLOATING
C13417 S.n12154 SUB 2.30fF $ **FLOATING
C13418 S.t1718 SUB 0.02fF
C13419 S.n12155 SUB 0.12fF $ **FLOATING
C13420 S.n12156 SUB 0.14fF $ **FLOATING
C13421 S.t2100 SUB 0.02fF
C13422 S.n12158 SUB 0.24fF $ **FLOATING
C13423 S.n12159 SUB 0.91fF $ **FLOATING
C13424 S.n12160 SUB 0.05fF $ **FLOATING
C13425 S.n12161 SUB 1.88fF $ **FLOATING
C13426 S.n12162 SUB 2.67fF $ **FLOATING
C13427 S.t1966 SUB 0.02fF
C13428 S.n12163 SUB 0.24fF $ **FLOATING
C13429 S.n12164 SUB 0.36fF $ **FLOATING
C13430 S.n12165 SUB 0.61fF $ **FLOATING
C13431 S.n12166 SUB 0.12fF $ **FLOATING
C13432 S.t191 SUB 0.02fF
C13433 S.n12167 SUB 0.14fF $ **FLOATING
C13434 S.n12169 SUB 2.80fF $ **FLOATING
C13435 S.n12170 SUB 2.30fF $ **FLOATING
C13436 S.t847 SUB 0.02fF
C13437 S.n12171 SUB 0.12fF $ **FLOATING
C13438 S.n12172 SUB 0.14fF $ **FLOATING
C13439 S.t1235 SUB 0.02fF
C13440 S.n12174 SUB 0.24fF $ **FLOATING
C13441 S.n12175 SUB 0.91fF $ **FLOATING
C13442 S.n12176 SUB 0.05fF $ **FLOATING
C13443 S.n12177 SUB 1.88fF $ **FLOATING
C13444 S.n12178 SUB 2.67fF $ **FLOATING
C13445 S.t1112 SUB 0.02fF
C13446 S.n12179 SUB 0.24fF $ **FLOATING
C13447 S.n12180 SUB 0.36fF $ **FLOATING
C13448 S.n12181 SUB 0.61fF $ **FLOATING
C13449 S.n12182 SUB 0.12fF $ **FLOATING
C13450 S.t1859 SUB 0.02fF
C13451 S.n12183 SUB 0.14fF $ **FLOATING
C13452 S.n12185 SUB 2.80fF $ **FLOATING
C13453 S.n12186 SUB 2.30fF $ **FLOATING
C13454 S.t2490 SUB 0.02fF
C13455 S.n12187 SUB 0.12fF $ **FLOATING
C13456 S.n12188 SUB 0.14fF $ **FLOATING
C13457 S.t355 SUB 0.02fF
C13458 S.n12190 SUB 0.24fF $ **FLOATING
C13459 S.n12191 SUB 0.91fF $ **FLOATING
C13460 S.n12192 SUB 0.05fF $ **FLOATING
C13461 S.n12193 SUB 1.88fF $ **FLOATING
C13462 S.n12194 SUB 2.67fF $ **FLOATING
C13463 S.t234 SUB 0.02fF
C13464 S.n12195 SUB 0.24fF $ **FLOATING
C13465 S.n12196 SUB 0.36fF $ **FLOATING
C13466 S.n12197 SUB 0.61fF $ **FLOATING
C13467 S.n12198 SUB 0.12fF $ **FLOATING
C13468 S.t992 SUB 0.02fF
C13469 S.n12199 SUB 0.14fF $ **FLOATING
C13470 S.n12201 SUB 2.80fF $ **FLOATING
C13471 S.n12202 SUB 2.30fF $ **FLOATING
C13472 S.t1775 SUB 0.02fF
C13473 S.n12203 SUB 0.12fF $ **FLOATING
C13474 S.n12204 SUB 0.14fF $ **FLOATING
C13475 S.t2010 SUB 0.02fF
C13476 S.n12206 SUB 0.24fF $ **FLOATING
C13477 S.n12207 SUB 0.91fF $ **FLOATING
C13478 S.n12208 SUB 0.05fF $ **FLOATING
C13479 S.n12209 SUB 1.88fF $ **FLOATING
C13480 S.n12210 SUB 2.67fF $ **FLOATING
C13481 S.t1900 SUB 0.02fF
C13482 S.n12211 SUB 0.24fF $ **FLOATING
C13483 S.n12212 SUB 0.36fF $ **FLOATING
C13484 S.n12213 SUB 0.61fF $ **FLOATING
C13485 S.n12214 SUB 0.12fF $ **FLOATING
C13486 S.t83 SUB 0.02fF
C13487 S.n12215 SUB 0.14fF $ **FLOATING
C13488 S.n12217 SUB 2.80fF $ **FLOATING
C13489 S.n12218 SUB 2.30fF $ **FLOATING
C13490 S.t905 SUB 0.02fF
C13491 S.n12219 SUB 0.12fF $ **FLOATING
C13492 S.n12220 SUB 0.14fF $ **FLOATING
C13493 S.t1158 SUB 0.02fF
C13494 S.n12222 SUB 0.24fF $ **FLOATING
C13495 S.n12223 SUB 0.91fF $ **FLOATING
C13496 S.n12224 SUB 0.05fF $ **FLOATING
C13497 S.n12225 SUB 1.88fF $ **FLOATING
C13498 S.n12226 SUB 2.67fF $ **FLOATING
C13499 S.t1041 SUB 0.02fF
C13500 S.n12227 SUB 0.24fF $ **FLOATING
C13501 S.n12228 SUB 0.36fF $ **FLOATING
C13502 S.n12229 SUB 0.61fF $ **FLOATING
C13503 S.n12230 SUB 0.12fF $ **FLOATING
C13504 S.t1762 SUB 0.02fF
C13505 S.n12231 SUB 0.14fF $ **FLOATING
C13506 S.n12233 SUB 2.80fF $ **FLOATING
C13507 S.n12234 SUB 2.30fF $ **FLOATING
C13508 S.t2548 SUB 0.02fF
C13509 S.n12235 SUB 0.12fF $ **FLOATING
C13510 S.n12236 SUB 0.14fF $ **FLOATING
C13511 S.t284 SUB 0.02fF
C13512 S.n12238 SUB 0.24fF $ **FLOATING
C13513 S.n12239 SUB 0.91fF $ **FLOATING
C13514 S.n12240 SUB 0.05fF $ **FLOATING
C13515 S.t2 SUB 48.31fF
C13516 S.t1676 SUB 0.02fF
C13517 S.n12241 SUB 0.12fF $ **FLOATING
C13518 S.n12242 SUB 0.14fF $ **FLOATING
C13519 S.t1946 SUB 0.02fF
C13520 S.n12244 SUB 0.24fF $ **FLOATING
C13521 S.n12245 SUB 0.91fF $ **FLOATING
C13522 S.n12246 SUB 0.05fF $ **FLOATING
C13523 S.t149 SUB 0.02fF
C13524 S.n12247 SUB 0.24fF $ **FLOATING
C13525 S.n12248 SUB 0.36fF $ **FLOATING
C13526 S.n12249 SUB 0.61fF $ **FLOATING
C13527 S.n12250 SUB 2.66fF $ **FLOATING
C13528 S.n12251 SUB 3.28fF $ **FLOATING
C13529 S.n12252 SUB 0.11fF $ **FLOATING
C13530 S.n12253 SUB 0.36fF $ **FLOATING
C13531 S.n12254 SUB 0.47fF $ **FLOATING
C13532 S.n12255 SUB 1.14fF $ **FLOATING
C13533 S.n12256 SUB 1.87fF $ **FLOATING
C13534 S.n12257 SUB 0.12fF $ **FLOATING
C13535 S.t753 SUB 0.02fF
C13536 S.n12258 SUB 0.14fF $ **FLOATING
C13537 S.t2046 SUB 0.02fF
C13538 S.n12260 SUB 0.24fF $ **FLOATING
C13539 S.n12261 SUB 0.36fF $ **FLOATING
C13540 S.n12262 SUB 0.61fF $ **FLOATING
C13541 S.n12263 SUB 1.27fF $ **FLOATING
C13542 S.n12264 SUB 2.38fF $ **FLOATING
C13543 S.n12265 SUB 4.20fF $ **FLOATING
C13544 S.t767 SUB 0.02fF
C13545 S.n12266 SUB 0.12fF $ **FLOATING
C13546 S.n12267 SUB 0.14fF $ **FLOATING
C13547 S.t1474 SUB 0.02fF
C13548 S.n12269 SUB 0.24fF $ **FLOATING
C13549 S.n12270 SUB 0.91fF $ **FLOATING
C13550 S.n12271 SUB 0.05fF $ **FLOATING
C13551 S.t44 SUB 47.92fF
C13552 S.t2543 SUB 0.02fF
C13553 S.n12272 SUB 0.01fF $ **FLOATING
C13554 S.n12273 SUB 0.26fF $ **FLOATING
C13555 S.t1248 SUB 0.02fF
C13556 S.n12275 SUB 1.19fF $ **FLOATING
C13557 S.n12276 SUB 0.05fF $ **FLOATING
C13558 S.t2207 SUB 0.02fF
C13559 S.n12277 SUB 0.64fF $ **FLOATING
C13560 S.n12278 SUB 0.61fF $ **FLOATING
C13561 S.n12279 SUB 8.97fF $ **FLOATING
C13562 S.n12280 SUB 8.97fF $ **FLOATING
C13563 S.n12281 SUB 0.60fF $ **FLOATING
C13564 S.n12282 SUB 0.22fF $ **FLOATING
C13565 S.n12283 SUB 0.59fF $ **FLOATING
C13566 S.n12284 SUB 3.43fF $ **FLOATING
C13567 S.n12285 SUB 0.29fF $ **FLOATING
C13568 S.t114 SUB 21.38fF
C13569 S.n12286 SUB 21.67fF $ **FLOATING
C13570 S.n12287 SUB 0.77fF $ **FLOATING
C13571 S.n12288 SUB 0.28fF $ **FLOATING
C13572 S.n12289 SUB 4.26fF $ **FLOATING
C13573 S.n12290 SUB 2.81fF $ **FLOATING
C13574 S.n12291 SUB 1.50fF $ **FLOATING
C13575 S.n12292 SUB 0.02fF $ **FLOATING
C13576 S.n12293 SUB 0.01fF $ **FLOATING
C13577 S.n12294 SUB 0.01fF $ **FLOATING
C13578 S.n12295 SUB 0.01fF $ **FLOATING
C13579 S.n12296 SUB 0.01fF $ **FLOATING
C13580 S.n12297 SUB 0.02fF $ **FLOATING
C13581 S.n12298 SUB 0.03fF $ **FLOATING
C13582 S.n12299 SUB 0.04fF $ **FLOATING
C13583 S.n12300 SUB 0.16fF $ **FLOATING
C13584 S.n12301 SUB 0.10fF $ **FLOATING
C13585 S.n12302 SUB 0.17fF $ **FLOATING
C13586 S.n12303 SUB 0.15fF $ **FLOATING
C13587 S.n12304 SUB 0.28fF $ **FLOATING
C13588 S.n12305 SUB 0.24fF $ **FLOATING
C13589 S.n12306 SUB 4.68fF $ **FLOATING
C13590 S.n12307 SUB 21.10fF $ **FLOATING
C13591 S.n12308 SUB 1.73fF $ **FLOATING
C13592 S.n12309 SUB 31.46fF $ **FLOATING
C13593 S.n12311 SUB 2.40fF $ **FLOATING
C13594 S.n12312 SUB 0.77fF $ **FLOATING
C13595 S.n12313 SUB 0.52fF $ **FLOATING
C13596 S.n12314 SUB 11.63fF $ **FLOATING
C13597 S.n12315 SUB 2.52fF $ **FLOATING
C13598 S.n12316 SUB 0.03fF $ **FLOATING
C13599 S.n12317 SUB 0.02fF $ **FLOATING
C13600 S.n12318 SUB 0.03fF $ **FLOATING
C13601 S.n12319 SUB 0.03fF $ **FLOATING
C13602 S.n12320 SUB 0.02fF $ **FLOATING
C13603 S.n12321 SUB 0.02fF $ **FLOATING
C13604 S.n12322 SUB 0.62fF $ **FLOATING
C13605 S.n12323 SUB 0.24fF $ **FLOATING
C13606 S.n12324 SUB 0.15fF $ **FLOATING
C13607 S.n12325 SUB 0.18fF $ **FLOATING
C13608 S.n12326 SUB 3.95fF $ **FLOATING
C13609 S.n12327 SUB 2.78fF $ **FLOATING
C13610 S.n12328 SUB 2.43fF $ **FLOATING
C13611 S.n12329 SUB 0.96fF $ **FLOATING
C13612 S.n12330 SUB 3.60fF $ **FLOATING
C13613 S.n12331 SUB 2.80fF $ **FLOATING
C13614 S.n12332 SUB 0.96fF $ **FLOATING
C13615 S.n12333 SUB 3.60fF $ **FLOATING
C13616 S.n12334 SUB 2.79fF $ **FLOATING
C13617 S.n12335 SUB 2.43fF $ **FLOATING
C13618 S.n12336 SUB 0.96fF $ **FLOATING
C13619 S.n12337 SUB 3.60fF $ **FLOATING
C13620 S.n12338 SUB 2.79fF $ **FLOATING
C13621 S.n12339 SUB 2.43fF $ **FLOATING
C13622 S.n12340 SUB 0.96fF $ **FLOATING
C13623 S.n12341 SUB 3.60fF $ **FLOATING
C13624 S.n12342 SUB 2.79fF $ **FLOATING
C13625 S.n12343 SUB 2.43fF $ **FLOATING
C13626 S.n12344 SUB 0.96fF $ **FLOATING
C13627 S.n12345 SUB 3.60fF $ **FLOATING
C13628 S.n12346 SUB 2.79fF $ **FLOATING
C13629 S.n12347 SUB 2.43fF $ **FLOATING
C13630 S.n12348 SUB 0.96fF $ **FLOATING
C13631 S.n12349 SUB 3.60fF $ **FLOATING
C13632 S.n12350 SUB 2.79fF $ **FLOATING
C13633 S.n12351 SUB 2.43fF $ **FLOATING
C13634 S.n12352 SUB 0.96fF $ **FLOATING
C13635 S.n12353 SUB 3.60fF $ **FLOATING
C13636 S.n12354 SUB 2.79fF $ **FLOATING
C13637 S.n12355 SUB 2.43fF $ **FLOATING
C13638 S.n12356 SUB 0.96fF $ **FLOATING
C13639 S.n12357 SUB 3.60fF $ **FLOATING
C13640 S.n12358 SUB 2.79fF $ **FLOATING
C13641 S.n12359 SUB 2.43fF $ **FLOATING
C13642 S.n12360 SUB 0.96fF $ **FLOATING
C13643 S.n12361 SUB 3.60fF $ **FLOATING
C13644 S.n12362 SUB 2.79fF $ **FLOATING
C13645 S.n12363 SUB 2.43fF $ **FLOATING
C13646 S.n12364 SUB 0.96fF $ **FLOATING
C13647 S.n12365 SUB 3.60fF $ **FLOATING
C13648 S.n12366 SUB 2.79fF $ **FLOATING
C13649 S.n12367 SUB 2.43fF $ **FLOATING
C13650 S.n12368 SUB 0.96fF $ **FLOATING
C13651 S.n12369 SUB 3.60fF $ **FLOATING
C13652 S.n12370 SUB 2.79fF $ **FLOATING
C13653 S.n12371 SUB 2.43fF $ **FLOATING
C13654 S.n12372 SUB 0.96fF $ **FLOATING
C13655 S.n12373 SUB 3.60fF $ **FLOATING
C13656 S.n12374 SUB 2.79fF $ **FLOATING
C13657 S.n12375 SUB 2.43fF $ **FLOATING
C13658 S.n12376 SUB 0.96fF $ **FLOATING
C13659 S.n12377 SUB 3.60fF $ **FLOATING
C13660 S.n12378 SUB 2.79fF $ **FLOATING
C13661 S.n12379 SUB 2.43fF $ **FLOATING
C13662 S.n12380 SUB 3.85fF $ **FLOATING
C13663 S.n12381 SUB 2.79fF $ **FLOATING
C13664 S.n12382 SUB 0.21fF $ **FLOATING
C13665 S.n12383 SUB 2.19fF $ **FLOATING
C13666 S.n12384 SUB 1.27fF $ **FLOATING
C13667 S.n12385 SUB 0.31fF $ **FLOATING
C13668 S.n12386 SUB 0.31fF $ **FLOATING
C13669 S.n12387 SUB 1.19fF $ **FLOATING
C13670 S.n12388 SUB 0.33fF $ **FLOATING
C13671 S.n12389 SUB 0.93fF $ **FLOATING
C13672 S.n12390 SUB 4.08fF $ **FLOATING
C13673 S.n12391 SUB 1.85fF $ **FLOATING
C13674 S.n12392 SUB 2.08fF $ **FLOATING
C13675 S.n12393 SUB 1.23fF $ **FLOATING
C13676 S.n12394 SUB 0.24fF $ **FLOATING
C13677 S.n12395 SUB 1.23fF $ **FLOATING
C13678 S.n12396 SUB 0.24fF $ **FLOATING
C13679 S.n12397 SUB 1.23fF $ **FLOATING
C13680 S.n12398 SUB 0.24fF $ **FLOATING
C13681 S.n12399 SUB 1.23fF $ **FLOATING
C13682 S.n12400 SUB 0.24fF $ **FLOATING
C13683 S.n12401 SUB 1.23fF $ **FLOATING
C13684 S.n12402 SUB 0.24fF $ **FLOATING
C13685 S.n12403 SUB 1.23fF $ **FLOATING
C13686 S.n12404 SUB 0.24fF $ **FLOATING
C13687 S.n12405 SUB 1.23fF $ **FLOATING
C13688 S.n12406 SUB 0.24fF $ **FLOATING
C13689 S.n12407 SUB 1.23fF $ **FLOATING
C13690 S.n12408 SUB 0.24fF $ **FLOATING
C13691 S.n12409 SUB 1.23fF $ **FLOATING
C13692 S.n12410 SUB 0.24fF $ **FLOATING
C13693 S.n12411 SUB 1.23fF $ **FLOATING
C13694 S.n12412 SUB 0.24fF $ **FLOATING
C13695 S.n12413 SUB 1.23fF $ **FLOATING
C13696 S.n12414 SUB 0.24fF $ **FLOATING
C13697 S.n12415 SUB 1.23fF $ **FLOATING
C13698 S.n12416 SUB 0.24fF $ **FLOATING
C13699 S.n12417 SUB 1.23fF $ **FLOATING
C13700 S.n12418 SUB 0.24fF $ **FLOATING
C13701 S.n12419 SUB 1.23fF $ **FLOATING
C13702 S.n12420 SUB 0.23fF $ **FLOATING
C13703 S.n12422 SUB 1.46fF $ **FLOATING
C13704 S.n12423 SUB 0.39fF $ **FLOATING
C13705 S.n12425 SUB 1.46fF $ **FLOATING
C13706 S.n12426 SUB 0.39fF $ **FLOATING
C13707 S.n12428 SUB 1.46fF $ **FLOATING
C13708 S.n12429 SUB 0.39fF $ **FLOATING
C13709 S.n12431 SUB 1.46fF $ **FLOATING
C13710 S.n12432 SUB 0.39fF $ **FLOATING
C13711 S.n12434 SUB 1.46fF $ **FLOATING
C13712 S.n12435 SUB 0.39fF $ **FLOATING
C13713 S.n12437 SUB 1.46fF $ **FLOATING
C13714 S.n12438 SUB 0.39fF $ **FLOATING
C13715 S.n12440 SUB 1.46fF $ **FLOATING
C13716 S.n12441 SUB 0.39fF $ **FLOATING
C13717 S.n12443 SUB 1.46fF $ **FLOATING
C13718 S.n12444 SUB 0.39fF $ **FLOATING
C13719 S.n12446 SUB 1.46fF $ **FLOATING
C13720 S.n12447 SUB 0.39fF $ **FLOATING
C13721 S.n12449 SUB 1.46fF $ **FLOATING
C13722 S.n12450 SUB 0.39fF $ **FLOATING
C13723 S.n12452 SUB 1.46fF $ **FLOATING
C13724 S.n12453 SUB 0.39fF $ **FLOATING
C13725 S.n12455 SUB 1.46fF $ **FLOATING
C13726 S.n12456 SUB 0.39fF $ **FLOATING
C13727 S.n12458 SUB 1.46fF $ **FLOATING
C13728 S.n12459 SUB 0.39fF $ **FLOATING
C13729 S.n12461 SUB 1.68fF $ **FLOATING
C13730 S.n12462 SUB 0.39fF $ **FLOATING
C13731 S.n12463 SUB 124.41fF $ **FLOATING
C13732 S.n12464 SUB 4.69fF $ **FLOATING
C13733 S.n12465 SUB 0.03fF $ **FLOATING
C13734 S.n12466 SUB 0.02fF $ **FLOATING
C13735 S.n12467 SUB 0.03fF $ **FLOATING
C13736 S.n12468 SUB 0.03fF $ **FLOATING
C13737 S.n12469 SUB 0.02fF $ **FLOATING
C13738 S.n12470 SUB 0.02fF $ **FLOATING
C13739 S.n12471 SUB 0.62fF $ **FLOATING
C13740 S.n12472 SUB 0.24fF $ **FLOATING
C13741 S.n12473 SUB 0.15fF $ **FLOATING
C13742 S.n12474 SUB 0.18fF $ **FLOATING
C13743 S.t2392 SUB 0.02fF
C13744 S.n12475 SUB 0.89fF $ **FLOATING
C13745 S.t2300 SUB 0.02fF
C13746 S.n12476 SUB 0.89fF $ **FLOATING
C13747 S.t499 SUB 0.02fF
C13748 S.n12477 SUB 0.02fF $ **FLOATING
C13749 S.n12478 SUB 0.37fF $ **FLOATING
C13750 S.n12479 SUB 20.78fF $ **FLOATING
C13751 S.t1973 SUB 0.02fF
C13752 S.n12480 SUB 0.89fF $ **FLOATING
C13753 S.t1440 SUB 0.02fF
C13754 S.n12481 SUB 0.02fF $ **FLOATING
C13755 S.n12482 SUB 0.37fF $ **FLOATING
C13756 S.t1783 SUB 0.02fF
C13757 S.n12483 SUB 0.89fF $ **FLOATING
C13758 S.t1118 SUB 0.02fF
C13759 S.n12484 SUB 0.89fF $ **FLOATING
C13760 S.t578 SUB 0.02fF
C13761 S.n12485 SUB 0.02fF $ **FLOATING
C13762 S.n12486 SUB 0.37fF $ **FLOATING
C13763 S.t911 SUB 0.02fF
C13764 S.n12487 SUB 0.89fF $ **FLOATING
C13765 S.t237 SUB 0.02fF
C13766 S.n12488 SUB 0.89fF $ **FLOATING
C13767 S.t2331 SUB 0.02fF
C13768 S.n12489 SUB 0.02fF $ **FLOATING
C13769 S.n12490 SUB 0.37fF $ **FLOATING
C13770 S.t172 SUB 0.02fF
C13771 S.n12491 SUB 0.89fF $ **FLOATING
C13772 S.t1904 SUB 0.02fF
C13773 S.n12492 SUB 0.89fF $ **FLOATING
C13774 S.t1473 SUB 0.02fF
C13775 S.n12493 SUB 0.02fF $ **FLOATING
C13776 S.n12494 SUB 0.37fF $ **FLOATING
C13777 S.t1835 SUB 0.02fF
C13778 S.n12495 SUB 0.89fF $ **FLOATING
C13779 S.t1045 SUB 0.02fF
C13780 S.n12496 SUB 0.89fF $ **FLOATING
C13781 S.t613 SUB 0.02fF
C13782 S.n12497 SUB 0.02fF $ **FLOATING
C13783 S.n12498 SUB 0.37fF $ **FLOATING
C13784 S.t969 SUB 0.02fF
C13785 S.n12499 SUB 0.89fF $ **FLOATING
C13786 S.t153 SUB 0.02fF
C13787 S.n12500 SUB 0.89fF $ **FLOATING
C13788 S.t2266 SUB 0.02fF
C13789 S.n12501 SUB 0.02fF $ **FLOATING
C13790 S.n12502 SUB 0.37fF $ **FLOATING
C13791 S.t36 SUB 0.02fF
C13792 S.n12503 SUB 0.89fF $ **FLOATING
C13793 S.t1817 SUB 0.02fF
C13794 S.n12504 SUB 0.89fF $ **FLOATING
C13795 S.t1407 SUB 0.02fF
C13796 S.n12505 SUB 0.02fF $ **FLOATING
C13797 S.n12506 SUB 0.37fF $ **FLOATING
C13798 S.t1733 SUB 0.02fF
C13799 S.n12507 SUB 0.89fF $ **FLOATING
C13800 S.t1079 SUB 0.02fF
C13801 S.n12508 SUB 0.89fF $ **FLOATING
C13802 S.t540 SUB 0.02fF
C13803 S.n12509 SUB 0.02fF $ **FLOATING
C13804 S.n12510 SUB 0.37fF $ **FLOATING
C13805 S.t859 SUB 0.02fF
C13806 S.n12511 SUB 0.89fF $ **FLOATING
C13807 S.t1649 SUB 0.02fF
C13808 S.n12512 SUB 0.89fF $ **FLOATING
C13809 S.t1943 SUB 0.02fF
C13810 S.n12513 SUB 0.02fF $ **FLOATING
C13811 S.n12514 SUB 0.37fF $ **FLOATING
C13812 S.t1480 SUB 0.02fF
C13813 S.n12515 SUB 0.89fF $ **FLOATING
C13814 S.t778 SUB 0.02fF
C13815 S.n12516 SUB 0.89fF $ **FLOATING
C13816 S.t1086 SUB 0.02fF
C13817 S.n12517 SUB 0.02fF $ **FLOATING
C13818 S.n12518 SUB 0.37fF $ **FLOATING
C13819 S.t618 SUB 0.02fF
C13820 S.n12519 SUB 0.89fF $ **FLOATING
C13821 S.t2431 SUB 0.02fF
C13822 S.n12520 SUB 0.89fF $ **FLOATING
C13823 S.t207 SUB 0.02fF
C13824 S.n12521 SUB 0.02fF $ **FLOATING
C13825 S.n12522 SUB 0.37fF $ **FLOATING
C13826 S.t2274 SUB 0.02fF
C13827 S.n12523 SUB 0.89fF $ **FLOATING
C13828 S.t1567 SUB 0.02fF
C13829 S.n12524 SUB 0.89fF $ **FLOATING
C13830 S.t1875 SUB 0.02fF
C13831 S.n12525 SUB 0.02fF $ **FLOATING
C13832 S.n12526 SUB 0.37fF $ **FLOATING
C13833 S.t1418 SUB 0.02fF
C13834 S.n12527 SUB 0.89fF $ **FLOATING
C13835 S.t699 SUB 0.02fF
C13836 S.n12528 SUB 0.89fF $ **FLOATING
C13837 S.t1129 SUB 0.02fF
C13838 S.n12529 SUB 0.02fF $ **FLOATING
C13839 S.n12530 SUB 0.37fF $ **FLOATING
C13840 S.t652 SUB 0.02fF
C13841 S.n12531 SUB 0.89fF $ **FLOATING
C13842 S.t2358 SUB 0.02fF
C13843 S.n12532 SUB 0.89fF $ **FLOATING
C13844 S.t251 SUB 0.02fF
C13845 S.n12533 SUB 0.02fF $ **FLOATING
C13846 S.n12534 SUB 0.37fF $ **FLOATING
C13847 S.t2306 SUB 0.02fF
C13848 S.n12535 SUB 0.89fF $ **FLOATING
C13849 S.t1503 SUB 0.02fF
C13850 S.n12536 SUB 0.89fF $ **FLOATING
C13851 S.t1917 SUB 0.02fF
C13852 S.n12537 SUB 0.02fF $ **FLOATING
C13853 S.n12538 SUB 0.37fF $ **FLOATING
C13854 S.t1450 SUB 0.02fF
C13855 S.n12539 SUB 0.89fF $ **FLOATING
C13856 S.t642 SUB 0.02fF
C13857 S.n12540 SUB 0.89fF $ **FLOATING
C13858 S.t1057 SUB 0.02fF
C13859 S.n12541 SUB 0.02fF $ **FLOATING
C13860 S.n12542 SUB 0.37fF $ **FLOATING
C13861 S.t593 SUB 0.02fF
C13862 S.n12543 SUB 0.89fF $ **FLOATING
C13863 S.t1645 SUB 0.02fF
C13864 S.n12544 SUB 0.44fF $ **FLOATING
C13865 S.t35 SUB 171.33fF
C13866 S.t1110 SUB 0.02fF
C13867 S.n12545 SUB 1.31fF $ **FLOATING
C13868 S.n12546 SUB 0.25fF $ **FLOATING
C13869 S.n12547 SUB 4.43fF $ **FLOATING
C13870 S.n12548 SUB 2.52fF $ **FLOATING
C13871 S.n12549 SUB 6.81fF $ **FLOATING
C13872 S.n12550 SUB 2.92fF $ **FLOATING
C13873 S.n12551 SUB 0.25fF $ **FLOATING
C13874 S.n12552 SUB 0.09fF $ **FLOATING
C13875 S.n12553 SUB 0.20fF $ **FLOATING
C13876 S.n12554 SUB 0.78fF $ **FLOATING
C13877 S.n12555 SUB 1.93fF $ **FLOATING
C13878 S.n12556 SUB 1.88fF $ **FLOATING
C13879 S.n12557 SUB 0.12fF $ **FLOATING
C13880 S.t264 SUB 0.02fF
C13881 S.n12558 SUB 0.14fF $ **FLOATING
C13882 S.t1526 SUB 0.02fF
C13883 S.n12560 SUB 0.24fF $ **FLOATING
C13884 S.n12561 SUB 0.36fF $ **FLOATING
C13885 S.n12562 SUB 0.61fF $ **FLOATING
C13886 S.n12563 SUB 2.67fF $ **FLOATING
C13887 S.n12564 SUB 2.99fF $ **FLOATING
C13888 S.t80 SUB 0.02fF
C13889 S.n12565 SUB 0.24fF $ **FLOATING
C13890 S.n12566 SUB 0.91fF $ **FLOATING
C13891 S.n12567 SUB 0.05fF $ **FLOATING
C13892 S.t1532 SUB 0.02fF
C13893 S.n12568 SUB 0.12fF $ **FLOATING
C13894 S.n12569 SUB 0.14fF $ **FLOATING
C13895 S.n12571 SUB 20.78fF $ **FLOATING
C13896 S.n12572 SUB 1.76fF $ **FLOATING
C13897 S.n12573 SUB 3.05fF $ **FLOATING
C13898 S.t664 SUB 0.02fF
C13899 S.n12574 SUB 0.24fF $ **FLOATING
C13900 S.n12575 SUB 0.36fF $ **FLOATING
C13901 S.n12576 SUB 0.61fF $ **FLOATING
C13902 S.n12577 SUB 0.12fF $ **FLOATING
C13903 S.t130 SUB 0.02fF
C13904 S.n12578 SUB 0.14fF $ **FLOATING
C13905 S.n12580 SUB 0.18fF $ **FLOATING
C13906 S.n12581 SUB 0.20fF $ **FLOATING
C13907 S.n12582 SUB 0.23fF $ **FLOATING
C13908 S.n12583 SUB 0.66fF $ **FLOATING
C13909 S.n12584 SUB 0.91fF $ **FLOATING
C13910 S.n12585 SUB 0.23fF $ **FLOATING
C13911 S.n12586 SUB 0.09fF $ **FLOATING
C13912 S.n12587 SUB 0.21fF $ **FLOATING
C13913 S.n12588 SUB 0.07fF $ **FLOATING
C13914 S.n12589 SUB 0.06fF $ **FLOATING
C13915 S.n12590 SUB 0.07fF $ **FLOATING
C13916 S.n12591 SUB 1.99fF $ **FLOATING
C13917 S.t316 SUB 0.02fF
C13918 S.n12592 SUB 0.12fF $ **FLOATING
C13919 S.n12593 SUB 0.14fF $ **FLOATING
C13920 S.t1978 SUB 0.02fF
C13921 S.n12595 SUB 0.24fF $ **FLOATING
C13922 S.n12596 SUB 0.91fF $ **FLOATING
C13923 S.n12597 SUB 0.05fF $ **FLOATING
C13924 S.n12598 SUB 1.95fF $ **FLOATING
C13925 S.n12599 SUB 0.12fF $ **FLOATING
C13926 S.t232 SUB 0.02fF
C13927 S.n12600 SUB 0.14fF $ **FLOATING
C13928 S.t2236 SUB 0.02fF
C13929 S.n12602 SUB 1.22fF $ **FLOATING
C13930 S.n12603 SUB 1.96fF $ **FLOATING
C13931 S.n12604 SUB 0.06fF $ **FLOATING
C13932 S.n12605 SUB 0.10fF $ **FLOATING
C13933 S.n12606 SUB 0.60fF $ **FLOATING
C13934 S.n12607 SUB 3.03fF $ **FLOATING
C13935 S.n12608 SUB 0.93fF $ **FLOATING
C13936 S.n12609 SUB 0.84fF $ **FLOATING
C13937 S.n12610 SUB 0.02fF $ **FLOATING
C13938 S.n12611 SUB 0.97fF $ **FLOATING
C13939 S.t128 SUB 21.38fF
C13940 S.n12612 SUB 19.94fF $ **FLOATING
C13941 S.n12614 SUB 1.22fF $ **FLOATING
C13942 S.n12615 SUB 1.45fF $ **FLOATING
C13943 S.n12616 SUB 2.90fF $ **FLOATING
C13944 S.n12617 SUB 2.42fF $ **FLOATING
C13945 S.n12618 SUB 3.85fF $ **FLOATING
C13946 S.n12619 SUB 0.25fF $ **FLOATING
C13947 S.n12620 SUB 0.01fF $ **FLOATING
C13948 S.t1108 SUB 0.02fF
C13949 S.n12621 SUB 0.25fF $ **FLOATING
C13950 S.t1472 SUB 0.02fF
C13951 S.n12622 SUB 0.95fF $ **FLOATING
C13952 S.n12623 SUB 0.70fF $ **FLOATING
C13953 S.n12624 SUB 0.04fF $ **FLOATING
C13954 S.n12625 SUB 0.10fF $ **FLOATING
C13955 S.n12626 SUB 0.29fF $ **FLOATING
C13956 S.n12627 SUB 0.25fF $ **FLOATING
C13957 S.n12628 SUB 0.12fF $ **FLOATING
C13958 S.n12629 SUB 0.05fF $ **FLOATING
C13959 S.n12630 SUB 0.18fF $ **FLOATING
C13960 S.n12631 SUB 1.26fF $ **FLOATING
C13961 S.n12632 SUB 2.77fF $ **FLOATING
C13962 S.n12633 SUB 0.12fF $ **FLOATING
C13963 S.t2467 SUB 0.02fF
C13964 S.n12634 SUB 0.14fF $ **FLOATING
C13965 S.t822 SUB 0.02fF
C13966 S.n12636 SUB 0.24fF $ **FLOATING
C13967 S.n12637 SUB 0.36fF $ **FLOATING
C13968 S.n12638 SUB 0.61fF $ **FLOATING
C13969 S.n12639 SUB 2.62fF $ **FLOATING
C13970 S.n12640 SUB 2.05fF $ **FLOATING
C13971 S.t181 SUB 0.02fF
C13972 S.n12641 SUB 0.24fF $ **FLOATING
C13973 S.n12642 SUB 0.91fF $ **FLOATING
C13974 S.n12643 SUB 0.05fF $ **FLOATING
C13975 S.t747 SUB 0.02fF
C13976 S.n12644 SUB 0.12fF $ **FLOATING
C13977 S.n12645 SUB 0.14fF $ **FLOATING
C13978 S.n12647 SUB 0.04fF $ **FLOATING
C13979 S.n12648 SUB 0.10fF $ **FLOATING
C13980 S.n12649 SUB 0.29fF $ **FLOATING
C13981 S.n12650 SUB 0.25fF $ **FLOATING
C13982 S.n12651 SUB 0.12fF $ **FLOATING
C13983 S.n12652 SUB 0.05fF $ **FLOATING
C13984 S.n12653 SUB 0.17fF $ **FLOATING
C13985 S.n12654 SUB 1.15fF $ **FLOATING
C13986 S.n12655 SUB 1.87fF $ **FLOATING
C13987 S.n12656 SUB 0.12fF $ **FLOATING
C13988 S.t2336 SUB 0.02fF
C13989 S.n12657 SUB 0.14fF $ **FLOATING
C13990 S.t818 SUB 0.02fF
C13991 S.n12659 SUB 0.24fF $ **FLOATING
C13992 S.n12660 SUB 0.36fF $ **FLOATING
C13993 S.n12661 SUB 0.61fF $ **FLOATING
C13994 S.n12662 SUB 2.53fF $ **FLOATING
C13995 S.n12663 SUB 1.94fF $ **FLOATING
C13996 S.t1115 SUB 0.02fF
C13997 S.n12664 SUB 0.24fF $ **FLOATING
C13998 S.n12665 SUB 0.91fF $ **FLOATING
C13999 S.n12666 SUB 0.05fF $ **FLOATING
C14000 S.t589 SUB 0.02fF
C14001 S.n12667 SUB 0.12fF $ **FLOATING
C14002 S.n12668 SUB 0.14fF $ **FLOATING
C14003 S.n12670 SUB 20.78fF $ **FLOATING
C14004 S.n12671 SUB 1.95fF $ **FLOATING
C14005 S.n12672 SUB 2.54fF $ **FLOATING
C14006 S.t2149 SUB 0.02fF
C14007 S.n12673 SUB 0.24fF $ **FLOATING
C14008 S.n12674 SUB 0.36fF $ **FLOATING
C14009 S.n12675 SUB 0.61fF $ **FLOATING
C14010 S.n12676 SUB 0.12fF $ **FLOATING
C14011 S.t1038 SUB 0.02fF
C14012 S.n12677 SUB 0.14fF $ **FLOATING
C14013 S.n12679 SUB 2.41fF $ **FLOATING
C14014 S.n12680 SUB 2.30fF $ **FLOATING
C14015 S.t1825 SUB 0.02fF
C14016 S.n12681 SUB 0.12fF $ **FLOATING
C14017 S.n12682 SUB 0.14fF $ **FLOATING
C14018 S.t1406 SUB 0.02fF
C14019 S.n12684 SUB 0.24fF $ **FLOATING
C14020 S.n12685 SUB 0.91fF $ **FLOATING
C14021 S.n12686 SUB 0.05fF $ **FLOATING
C14022 S.n12687 SUB 1.95fF $ **FLOATING
C14023 S.n12688 SUB 2.54fF $ **FLOATING
C14024 S.t1289 SUB 0.02fF
C14025 S.n12689 SUB 0.24fF $ **FLOATING
C14026 S.n12690 SUB 0.36fF $ **FLOATING
C14027 S.n12691 SUB 0.61fF $ **FLOATING
C14028 S.n12692 SUB 0.12fF $ **FLOATING
C14029 S.t141 SUB 0.02fF
C14030 S.n12693 SUB 0.14fF $ **FLOATING
C14031 S.n12695 SUB 2.41fF $ **FLOATING
C14032 S.n12696 SUB 2.30fF $ **FLOATING
C14033 S.t961 SUB 0.02fF
C14034 S.n12697 SUB 0.12fF $ **FLOATING
C14035 S.n12698 SUB 0.14fF $ **FLOATING
C14036 S.t539 SUB 0.02fF
C14037 S.n12700 SUB 0.24fF $ **FLOATING
C14038 S.n12701 SUB 0.91fF $ **FLOATING
C14039 S.n12702 SUB 0.05fF $ **FLOATING
C14040 S.n12703 SUB 1.95fF $ **FLOATING
C14041 S.n12704 SUB 2.54fF $ **FLOATING
C14042 S.t402 SUB 0.02fF
C14043 S.n12705 SUB 0.24fF $ **FLOATING
C14044 S.n12706 SUB 0.36fF $ **FLOATING
C14045 S.n12707 SUB 0.61fF $ **FLOATING
C14046 S.n12708 SUB 0.12fF $ **FLOATING
C14047 S.t1811 SUB 0.02fF
C14048 S.n12709 SUB 0.14fF $ **FLOATING
C14049 S.n12711 SUB 2.41fF $ **FLOATING
C14050 S.n12712 SUB 2.30fF $ **FLOATING
C14051 S.t15 SUB 0.02fF
C14052 S.n12713 SUB 0.12fF $ **FLOATING
C14053 S.n12714 SUB 0.14fF $ **FLOATING
C14054 S.t2181 SUB 0.02fF
C14055 S.n12716 SUB 0.24fF $ **FLOATING
C14056 S.n12717 SUB 0.91fF $ **FLOATING
C14057 S.n12718 SUB 0.05fF $ **FLOATING
C14058 S.n12719 SUB 1.95fF $ **FLOATING
C14059 S.n12720 SUB 2.54fF $ **FLOATING
C14060 S.t2051 SUB 0.02fF
C14061 S.n12721 SUB 0.24fF $ **FLOATING
C14062 S.n12722 SUB 0.36fF $ **FLOATING
C14063 S.n12723 SUB 0.61fF $ **FLOATING
C14064 S.n12724 SUB 0.12fF $ **FLOATING
C14065 S.t944 SUB 0.02fF
C14066 S.n12725 SUB 0.14fF $ **FLOATING
C14067 S.n12727 SUB 2.41fF $ **FLOATING
C14068 S.n12728 SUB 2.30fF $ **FLOATING
C14069 S.t1724 SUB 0.02fF
C14070 S.n12729 SUB 0.12fF $ **FLOATING
C14071 S.n12730 SUB 0.14fF $ **FLOATING
C14072 S.t1320 SUB 0.02fF
C14073 S.n12732 SUB 0.24fF $ **FLOATING
C14074 S.n12733 SUB 0.91fF $ **FLOATING
C14075 S.n12734 SUB 0.05fF $ **FLOATING
C14076 S.n12735 SUB 1.95fF $ **FLOATING
C14077 S.n12736 SUB 2.54fF $ **FLOATING
C14078 S.t1191 SUB 0.02fF
C14079 S.n12737 SUB 0.24fF $ **FLOATING
C14080 S.n12738 SUB 0.36fF $ **FLOATING
C14081 S.n12739 SUB 0.61fF $ **FLOATING
C14082 S.n12740 SUB 0.12fF $ **FLOATING
C14083 S.t193 SUB 0.02fF
C14084 S.n12741 SUB 0.14fF $ **FLOATING
C14085 S.n12743 SUB 2.41fF $ **FLOATING
C14086 S.n12744 SUB 2.30fF $ **FLOATING
C14087 S.t852 SUB 0.02fF
C14088 S.n12745 SUB 0.12fF $ **FLOATING
C14089 S.n12746 SUB 0.14fF $ **FLOATING
C14090 S.t439 SUB 0.02fF
C14091 S.n12748 SUB 0.24fF $ **FLOATING
C14092 S.n12749 SUB 0.91fF $ **FLOATING
C14093 S.n12750 SUB 0.05fF $ **FLOATING
C14094 S.n12751 SUB 1.95fF $ **FLOATING
C14095 S.n12752 SUB 2.54fF $ **FLOATING
C14096 S.t224 SUB 0.02fF
C14097 S.n12753 SUB 0.24fF $ **FLOATING
C14098 S.n12754 SUB 0.36fF $ **FLOATING
C14099 S.n12755 SUB 0.61fF $ **FLOATING
C14100 S.n12756 SUB 0.12fF $ **FLOATING
C14101 S.t1889 SUB 0.02fF
C14102 S.n12757 SUB 0.14fF $ **FLOATING
C14103 S.n12759 SUB 2.41fF $ **FLOATING
C14104 S.n12760 SUB 2.30fF $ **FLOATING
C14105 S.t2492 SUB 0.02fF
C14106 S.n12761 SUB 0.12fF $ **FLOATING
C14107 S.n12762 SUB 0.14fF $ **FLOATING
C14108 S.t2064 SUB 0.02fF
C14109 S.n12764 SUB 0.24fF $ **FLOATING
C14110 S.n12765 SUB 0.91fF $ **FLOATING
C14111 S.n12766 SUB 0.05fF $ **FLOATING
C14112 S.n12767 SUB 1.95fF $ **FLOATING
C14113 S.n12768 SUB 2.54fF $ **FLOATING
C14114 S.t1891 SUB 0.02fF
C14115 S.n12769 SUB 0.24fF $ **FLOATING
C14116 S.n12770 SUB 0.36fF $ **FLOATING
C14117 S.n12771 SUB 0.61fF $ **FLOATING
C14118 S.n12772 SUB 0.12fF $ **FLOATING
C14119 S.t1027 SUB 0.02fF
C14120 S.n12773 SUB 0.14fF $ **FLOATING
C14121 S.n12775 SUB 2.41fF $ **FLOATING
C14122 S.n12776 SUB 2.30fF $ **FLOATING
C14123 S.t1655 SUB 0.02fF
C14124 S.n12777 SUB 0.12fF $ **FLOATING
C14125 S.n12778 SUB 0.14fF $ **FLOATING
C14126 S.t1201 SUB 0.02fF
C14127 S.n12780 SUB 0.24fF $ **FLOATING
C14128 S.n12781 SUB 0.91fF $ **FLOATING
C14129 S.n12782 SUB 0.05fF $ **FLOATING
C14130 S.n12783 SUB 1.95fF $ **FLOATING
C14131 S.n12784 SUB 2.54fF $ **FLOATING
C14132 S.t1028 SUB 0.02fF
C14133 S.n12785 SUB 0.24fF $ **FLOATING
C14134 S.n12786 SUB 0.36fF $ **FLOATING
C14135 S.n12787 SUB 0.61fF $ **FLOATING
C14136 S.n12788 SUB 0.12fF $ **FLOATING
C14137 S.t127 SUB 0.02fF
C14138 S.n12789 SUB 0.14fF $ **FLOATING
C14139 S.n12791 SUB 2.41fF $ **FLOATING
C14140 S.n12792 SUB 2.30fF $ **FLOATING
C14141 S.t785 SUB 0.02fF
C14142 S.n12793 SUB 0.12fF $ **FLOATING
C14143 S.n12794 SUB 0.14fF $ **FLOATING
C14144 S.t324 SUB 0.02fF
C14145 S.n12796 SUB 0.24fF $ **FLOATING
C14146 S.n12797 SUB 0.91fF $ **FLOATING
C14147 S.n12798 SUB 0.05fF $ **FLOATING
C14148 S.n12799 SUB 1.95fF $ **FLOATING
C14149 S.n12800 SUB 2.54fF $ **FLOATING
C14150 S.t129 SUB 0.02fF
C14151 S.n12801 SUB 0.24fF $ **FLOATING
C14152 S.n12802 SUB 0.36fF $ **FLOATING
C14153 S.n12803 SUB 0.61fF $ **FLOATING
C14154 S.n12804 SUB 0.12fF $ **FLOATING
C14155 S.t1798 SUB 0.02fF
C14156 S.n12805 SUB 0.14fF $ **FLOATING
C14157 S.n12807 SUB 2.41fF $ **FLOATING
C14158 S.n12808 SUB 2.30fF $ **FLOATING
C14159 S.t2435 SUB 0.02fF
C14160 S.n12809 SUB 0.12fF $ **FLOATING
C14161 S.n12810 SUB 0.14fF $ **FLOATING
C14162 S.t1983 SUB 0.02fF
C14163 S.n12812 SUB 0.24fF $ **FLOATING
C14164 S.n12813 SUB 0.91fF $ **FLOATING
C14165 S.n12814 SUB 0.05fF $ **FLOATING
C14166 S.n12815 SUB 1.95fF $ **FLOATING
C14167 S.n12816 SUB 2.54fF $ **FLOATING
C14168 S.t1799 SUB 0.02fF
C14169 S.n12817 SUB 0.24fF $ **FLOATING
C14170 S.n12818 SUB 0.36fF $ **FLOATING
C14171 S.n12819 SUB 0.61fF $ **FLOATING
C14172 S.n12820 SUB 0.12fF $ **FLOATING
C14173 S.t928 SUB 0.02fF
C14174 S.n12821 SUB 0.14fF $ **FLOATING
C14175 S.n12823 SUB 2.41fF $ **FLOATING
C14176 S.n12824 SUB 2.30fF $ **FLOATING
C14177 S.t1571 SUB 0.02fF
C14178 S.n12825 SUB 0.12fF $ **FLOATING
C14179 S.n12826 SUB 0.14fF $ **FLOATING
C14180 S.t1135 SUB 0.02fF
C14181 S.n12828 SUB 0.24fF $ **FLOATING
C14182 S.n12829 SUB 0.91fF $ **FLOATING
C14183 S.n12830 SUB 0.05fF $ **FLOATING
C14184 S.n12831 SUB 1.95fF $ **FLOATING
C14185 S.n12832 SUB 2.54fF $ **FLOATING
C14186 S.t929 SUB 0.02fF
C14187 S.n12833 SUB 0.24fF $ **FLOATING
C14188 S.n12834 SUB 0.36fF $ **FLOATING
C14189 S.n12835 SUB 0.61fF $ **FLOATING
C14190 S.n12836 SUB 0.12fF $ **FLOATING
C14191 S.t2569 SUB 0.02fF
C14192 S.n12837 SUB 0.14fF $ **FLOATING
C14193 S.n12839 SUB 2.41fF $ **FLOATING
C14194 S.n12840 SUB 2.30fF $ **FLOATING
C14195 S.t842 SUB 0.02fF
C14196 S.n12841 SUB 0.12fF $ **FLOATING
C14197 S.n12842 SUB 0.14fF $ **FLOATING
C14198 S.t256 SUB 0.02fF
C14199 S.n12844 SUB 0.24fF $ **FLOATING
C14200 S.n12845 SUB 0.91fF $ **FLOATING
C14201 S.n12846 SUB 0.05fF $ **FLOATING
C14202 S.n12847 SUB 1.95fF $ **FLOATING
C14203 S.n12848 SUB 2.54fF $ **FLOATING
C14204 S.t2572 SUB 0.02fF
C14205 S.n12849 SUB 0.24fF $ **FLOATING
C14206 S.n12850 SUB 0.36fF $ **FLOATING
C14207 S.n12851 SUB 0.61fF $ **FLOATING
C14208 S.n12852 SUB 0.12fF $ **FLOATING
C14209 S.t1693 SUB 0.02fF
C14210 S.n12853 SUB 0.14fF $ **FLOATING
C14211 S.n12855 SUB 2.41fF $ **FLOATING
C14212 S.n12856 SUB 2.30fF $ **FLOATING
C14213 S.t2485 SUB 0.02fF
C14214 S.n12857 SUB 0.12fF $ **FLOATING
C14215 S.n12858 SUB 0.14fF $ **FLOATING
C14216 S.t1922 SUB 0.02fF
C14217 S.n12860 SUB 0.24fF $ **FLOATING
C14218 S.n12861 SUB 0.91fF $ **FLOATING
C14219 S.n12862 SUB 0.05fF $ **FLOATING
C14220 S.n12863 SUB 2.41fF $ **FLOATING
C14221 S.n12864 SUB 1.98fF $ **FLOATING
C14222 S.n12865 SUB 0.12fF $ **FLOATING
C14223 S.t823 SUB 0.02fF
C14224 S.n12866 SUB 0.14fF $ **FLOATING
C14225 S.t1697 SUB 0.02fF
C14226 S.n12868 SUB 0.24fF $ **FLOATING
C14227 S.n12869 SUB 0.36fF $ **FLOATING
C14228 S.n12870 SUB 0.61fF $ **FLOATING
C14229 S.n12871 SUB 2.55fF $ **FLOATING
C14230 S.n12872 SUB 2.31fF $ **FLOATING
C14231 S.t1611 SUB 0.02fF
C14232 S.n12873 SUB 0.12fF $ **FLOATING
C14233 S.n12874 SUB 0.14fF $ **FLOATING
C14234 S.t1062 SUB 0.02fF
C14235 S.n12876 SUB 0.24fF $ **FLOATING
C14236 S.n12877 SUB 0.91fF $ **FLOATING
C14237 S.n12878 SUB 0.05fF $ **FLOATING
C14238 S.t14 SUB 48.31fF
C14239 S.t902 SUB 0.02fF
C14240 S.n12879 SUB 0.12fF $ **FLOATING
C14241 S.n12880 SUB 0.14fF $ **FLOATING
C14242 S.t610 SUB 0.02fF
C14243 S.n12882 SUB 0.24fF $ **FLOATING
C14244 S.n12883 SUB 0.91fF $ **FLOATING
C14245 S.n12884 SUB 0.05fF $ **FLOATING
C14246 S.t1376 SUB 0.02fF
C14247 S.n12885 SUB 0.24fF $ **FLOATING
C14248 S.n12886 SUB 0.36fF $ **FLOATING
C14249 S.n12887 SUB 0.61fF $ **FLOATING
C14250 S.n12888 SUB 0.30fF $ **FLOATING
C14251 S.n12889 SUB 1.09fF $ **FLOATING
C14252 S.n12890 SUB 0.15fF $ **FLOATING
C14253 S.n12891 SUB 2.10fF $ **FLOATING
C14254 S.n12892 SUB 2.12fF $ **FLOATING
C14255 S.n12893 SUB 1.79fF $ **FLOATING
C14256 S.n12894 SUB 1.88fF $ **FLOATING
C14257 S.n12895 SUB 0.12fF $ **FLOATING
C14258 S.t1800 SUB 0.02fF
C14259 S.n12896 SUB 0.14fF $ **FLOATING
C14260 S.t2318 SUB 0.02fF
C14261 S.n12898 SUB 0.24fF $ **FLOATING
C14262 S.n12899 SUB 0.36fF $ **FLOATING
C14263 S.n12900 SUB 0.61fF $ **FLOATING
C14264 S.n12901 SUB 0.92fF $ **FLOATING
C14265 S.n12902 SUB 0.32fF $ **FLOATING
C14266 S.n12903 SUB 0.92fF $ **FLOATING
C14267 S.n12904 SUB 1.09fF $ **FLOATING
C14268 S.n12905 SUB 0.15fF $ **FLOATING
C14269 S.n12906 SUB 4.96fF $ **FLOATING
C14270 S.t1981 SUB 0.02fF
C14271 S.n12907 SUB 0.12fF $ **FLOATING
C14272 S.n12908 SUB 0.14fF $ **FLOATING
C14273 S.t1125 SUB 0.02fF
C14274 S.n12910 SUB 0.24fF $ **FLOATING
C14275 S.n12911 SUB 0.91fF $ **FLOATING
C14276 S.n12912 SUB 0.05fF $ **FLOATING
C14277 S.n12913 SUB 1.88fF $ **FLOATING
C14278 S.n12914 SUB 2.67fF $ **FLOATING
C14279 S.t1555 SUB 0.02fF
C14280 S.n12915 SUB 0.24fF $ **FLOATING
C14281 S.n12916 SUB 0.36fF $ **FLOATING
C14282 S.n12917 SUB 0.61fF $ **FLOATING
C14283 S.n12918 SUB 0.12fF $ **FLOATING
C14284 S.t1067 SUB 0.02fF
C14285 S.n12919 SUB 0.14fF $ **FLOATING
C14286 S.n12921 SUB 1.95fF $ **FLOATING
C14287 S.n12922 SUB 2.54fF $ **FLOATING
C14288 S.t503 SUB 0.02fF
C14289 S.n12923 SUB 0.24fF $ **FLOATING
C14290 S.n12924 SUB 0.36fF $ **FLOATING
C14291 S.n12925 SUB 0.61fF $ **FLOATING
C14292 S.t2264 SUB 0.02fF
C14293 S.n12926 SUB 0.24fF $ **FLOATING
C14294 S.n12927 SUB 0.91fF $ **FLOATING
C14295 S.n12928 SUB 0.05fF $ **FLOATING
C14296 S.t2545 SUB 0.02fF
C14297 S.n12929 SUB 0.12fF $ **FLOATING
C14298 S.n12930 SUB 0.14fF $ **FLOATING
C14299 S.n12932 SUB 0.12fF $ **FLOATING
C14300 S.t1898 SUB 0.02fF
C14301 S.n12933 SUB 0.14fF $ **FLOATING
C14302 S.n12935 SUB 2.30fF $ **FLOATING
C14303 S.n12936 SUB 1.77fF $ **FLOATING
C14304 S.n12937 SUB 5.16fF $ **FLOATING
C14305 S.t1131 SUB 0.02fF
C14306 S.n12938 SUB 0.12fF $ **FLOATING
C14307 S.n12939 SUB 0.14fF $ **FLOATING
C14308 S.t357 SUB 0.02fF
C14309 S.n12941 SUB 0.24fF $ **FLOATING
C14310 S.n12942 SUB 0.91fF $ **FLOATING
C14311 S.n12943 SUB 0.05fF $ **FLOATING
C14312 S.n12944 SUB 1.88fF $ **FLOATING
C14313 S.n12945 SUB 2.67fF $ **FLOATING
C14314 S.t693 SUB 0.02fF
C14315 S.n12946 SUB 0.24fF $ **FLOATING
C14316 S.n12947 SUB 0.36fF $ **FLOATING
C14317 S.n12948 SUB 0.61fF $ **FLOATING
C14318 S.n12949 SUB 0.12fF $ **FLOATING
C14319 S.t186 SUB 0.02fF
C14320 S.n12950 SUB 0.14fF $ **FLOATING
C14321 S.n12952 SUB 5.17fF $ **FLOATING
C14322 S.t252 SUB 0.02fF
C14323 S.n12953 SUB 0.12fF $ **FLOATING
C14324 S.n12954 SUB 0.14fF $ **FLOATING
C14325 S.t2011 SUB 0.02fF
C14326 S.n12956 SUB 0.24fF $ **FLOATING
C14327 S.n12957 SUB 0.91fF $ **FLOATING
C14328 S.n12958 SUB 0.05fF $ **FLOATING
C14329 S.n12959 SUB 1.88fF $ **FLOATING
C14330 S.n12960 SUB 2.67fF $ **FLOATING
C14331 S.t2353 SUB 0.02fF
C14332 S.n12961 SUB 0.24fF $ **FLOATING
C14333 S.n12962 SUB 0.36fF $ **FLOATING
C14334 S.n12963 SUB 0.61fF $ **FLOATING
C14335 S.n12964 SUB 0.12fF $ **FLOATING
C14336 S.t1853 SUB 0.02fF
C14337 S.n12965 SUB 0.14fF $ **FLOATING
C14338 S.n12967 SUB 5.17fF $ **FLOATING
C14339 S.t1919 SUB 0.02fF
C14340 S.n12968 SUB 0.12fF $ **FLOATING
C14341 S.n12969 SUB 0.14fF $ **FLOATING
C14342 S.t1159 SUB 0.02fF
C14343 S.n12971 SUB 0.24fF $ **FLOATING
C14344 S.n12972 SUB 0.91fF $ **FLOATING
C14345 S.n12973 SUB 0.05fF $ **FLOATING
C14346 S.n12974 SUB 1.88fF $ **FLOATING
C14347 S.n12975 SUB 2.67fF $ **FLOATING
C14348 S.t1495 SUB 0.02fF
C14349 S.n12976 SUB 0.24fF $ **FLOATING
C14350 S.n12977 SUB 0.36fF $ **FLOATING
C14351 S.n12978 SUB 0.61fF $ **FLOATING
C14352 S.n12979 SUB 0.12fF $ **FLOATING
C14353 S.t989 SUB 0.02fF
C14354 S.n12980 SUB 0.14fF $ **FLOATING
C14355 S.n12982 SUB 5.17fF $ **FLOATING
C14356 S.t1058 SUB 0.02fF
C14357 S.n12983 SUB 0.12fF $ **FLOATING
C14358 S.n12984 SUB 0.14fF $ **FLOATING
C14359 S.t286 SUB 0.02fF
C14360 S.n12986 SUB 0.24fF $ **FLOATING
C14361 S.n12987 SUB 0.91fF $ **FLOATING
C14362 S.n12988 SUB 0.05fF $ **FLOATING
C14363 S.n12989 SUB 1.88fF $ **FLOATING
C14364 S.n12990 SUB 2.67fF $ **FLOATING
C14365 S.t632 SUB 0.02fF
C14366 S.n12991 SUB 0.24fF $ **FLOATING
C14367 S.n12992 SUB 0.36fF $ **FLOATING
C14368 S.n12993 SUB 0.61fF $ **FLOATING
C14369 S.n12994 SUB 0.12fF $ **FLOATING
C14370 S.t73 SUB 0.02fF
C14371 S.n12995 SUB 0.14fF $ **FLOATING
C14372 S.n12997 SUB 5.17fF $ **FLOATING
C14373 S.t171 SUB 0.02fF
C14374 S.n12998 SUB 0.12fF $ **FLOATING
C14375 S.n12999 SUB 0.14fF $ **FLOATING
C14376 S.t1947 SUB 0.02fF
C14377 S.n13001 SUB 0.24fF $ **FLOATING
C14378 S.n13002 SUB 0.91fF $ **FLOATING
C14379 S.n13003 SUB 0.05fF $ **FLOATING
C14380 S.n13004 SUB 1.88fF $ **FLOATING
C14381 S.n13005 SUB 2.67fF $ **FLOATING
C14382 S.t2287 SUB 0.02fF
C14383 S.n13006 SUB 0.24fF $ **FLOATING
C14384 S.n13007 SUB 0.36fF $ **FLOATING
C14385 S.n13008 SUB 0.61fF $ **FLOATING
C14386 S.n13009 SUB 0.12fF $ **FLOATING
C14387 S.t1753 SUB 0.02fF
C14388 S.n13010 SUB 0.14fF $ **FLOATING
C14389 S.n13012 SUB 5.17fF $ **FLOATING
C14390 S.t1951 SUB 0.02fF
C14391 S.n13013 SUB 0.12fF $ **FLOATING
C14392 S.n13014 SUB 0.14fF $ **FLOATING
C14393 S.t1089 SUB 0.02fF
C14394 S.n13016 SUB 0.24fF $ **FLOATING
C14395 S.n13017 SUB 0.91fF $ **FLOATING
C14396 S.n13018 SUB 0.05fF $ **FLOATING
C14397 S.n13019 SUB 1.88fF $ **FLOATING
C14398 S.n13020 SUB 2.67fF $ **FLOATING
C14399 S.t1285 SUB 0.02fF
C14400 S.n13021 SUB 0.24fF $ **FLOATING
C14401 S.n13022 SUB 0.36fF $ **FLOATING
C14402 S.n13023 SUB 0.61fF $ **FLOATING
C14403 S.n13024 SUB 0.12fF $ **FLOATING
C14404 S.t707 SUB 0.02fF
C14405 S.n13025 SUB 0.14fF $ **FLOATING
C14406 S.n13027 SUB 5.17fF $ **FLOATING
C14407 S.t939 SUB 0.02fF
C14408 S.n13028 SUB 0.12fF $ **FLOATING
C14409 S.n13029 SUB 0.14fF $ **FLOATING
C14410 S.t1251 SUB 0.02fF
C14411 S.n13031 SUB 0.24fF $ **FLOATING
C14412 S.n13032 SUB 0.91fF $ **FLOATING
C14413 S.n13033 SUB 0.05fF $ **FLOATING
C14414 S.n13034 SUB 1.88fF $ **FLOATING
C14415 S.n13035 SUB 2.67fF $ **FLOATING
C14416 S.t397 SUB 0.02fF
C14417 S.n13036 SUB 0.24fF $ **FLOATING
C14418 S.n13037 SUB 0.36fF $ **FLOATING
C14419 S.n13038 SUB 0.61fF $ **FLOATING
C14420 S.n13039 SUB 0.12fF $ **FLOATING
C14421 S.t2364 SUB 0.02fF
C14422 S.n13040 SUB 0.14fF $ **FLOATING
C14423 S.n13042 SUB 5.17fF $ **FLOATING
C14424 S.t2578 SUB 0.02fF
C14425 S.n13043 SUB 0.12fF $ **FLOATING
C14426 S.n13044 SUB 0.14fF $ **FLOATING
C14427 S.t369 SUB 0.02fF
C14428 S.n13046 SUB 0.24fF $ **FLOATING
C14429 S.n13047 SUB 0.91fF $ **FLOATING
C14430 S.n13048 SUB 0.05fF $ **FLOATING
C14431 S.n13049 SUB 1.88fF $ **FLOATING
C14432 S.n13050 SUB 2.67fF $ **FLOATING
C14433 S.t2049 SUB 0.02fF
C14434 S.n13051 SUB 0.24fF $ **FLOATING
C14435 S.n13052 SUB 0.36fF $ **FLOATING
C14436 S.n13053 SUB 0.61fF $ **FLOATING
C14437 S.n13054 SUB 0.12fF $ **FLOATING
C14438 S.t1508 SUB 0.02fF
C14439 S.n13055 SUB 0.14fF $ **FLOATING
C14440 S.n13057 SUB 5.17fF $ **FLOATING
C14441 S.t1701 SUB 0.02fF
C14442 S.n13058 SUB 0.12fF $ **FLOATING
C14443 S.n13059 SUB 0.14fF $ **FLOATING
C14444 S.t2022 SUB 0.02fF
C14445 S.n13061 SUB 0.24fF $ **FLOATING
C14446 S.n13062 SUB 0.91fF $ **FLOATING
C14447 S.n13063 SUB 0.05fF $ **FLOATING
C14448 S.n13064 SUB 1.88fF $ **FLOATING
C14449 S.n13065 SUB 2.67fF $ **FLOATING
C14450 S.t1190 SUB 0.02fF
C14451 S.n13066 SUB 0.24fF $ **FLOATING
C14452 S.n13067 SUB 0.36fF $ **FLOATING
C14453 S.n13068 SUB 0.61fF $ **FLOATING
C14454 S.n13069 SUB 0.12fF $ **FLOATING
C14455 S.t648 SUB 0.02fF
C14456 S.n13070 SUB 0.14fF $ **FLOATING
C14457 S.n13072 SUB 5.17fF $ **FLOATING
C14458 S.t828 SUB 0.02fF
C14459 S.n13073 SUB 0.12fF $ **FLOATING
C14460 S.n13074 SUB 0.14fF $ **FLOATING
C14461 S.t1166 SUB 0.02fF
C14462 S.n13076 SUB 0.24fF $ **FLOATING
C14463 S.n13077 SUB 0.91fF $ **FLOATING
C14464 S.n13078 SUB 0.05fF $ **FLOATING
C14465 S.n13079 SUB 1.88fF $ **FLOATING
C14466 S.n13080 SUB 2.67fF $ **FLOATING
C14467 S.t456 SUB 0.02fF
C14468 S.n13081 SUB 0.24fF $ **FLOATING
C14469 S.n13082 SUB 0.36fF $ **FLOATING
C14470 S.n13083 SUB 0.61fF $ **FLOATING
C14471 S.n13084 SUB 0.12fF $ **FLOATING
C14472 S.t2405 SUB 0.02fF
C14473 S.n13085 SUB 0.14fF $ **FLOATING
C14474 S.n13087 SUB 5.17fF $ **FLOATING
C14475 S.t2473 SUB 0.02fF
C14476 S.n13088 SUB 0.12fF $ **FLOATING
C14477 S.n13089 SUB 0.14fF $ **FLOATING
C14478 S.t421 SUB 0.02fF
C14479 S.n13091 SUB 0.24fF $ **FLOATING
C14480 S.n13092 SUB 0.91fF $ **FLOATING
C14481 S.n13093 SUB 0.05fF $ **FLOATING
C14482 S.n13094 SUB 1.88fF $ **FLOATING
C14483 S.n13095 SUB 2.67fF $ **FLOATING
C14484 S.t2101 SUB 0.02fF
C14485 S.n13096 SUB 0.24fF $ **FLOATING
C14486 S.n13097 SUB 0.36fF $ **FLOATING
C14487 S.n13098 SUB 0.61fF $ **FLOATING
C14488 S.n13099 SUB 0.12fF $ **FLOATING
C14489 S.t1543 SUB 0.02fF
C14490 S.n13100 SUB 0.14fF $ **FLOATING
C14491 S.n13102 SUB 5.17fF $ **FLOATING
C14492 S.t1604 SUB 0.02fF
C14493 S.n13103 SUB 0.12fF $ **FLOATING
C14494 S.n13104 SUB 0.14fF $ **FLOATING
C14495 S.t2068 SUB 0.02fF
C14496 S.n13106 SUB 0.24fF $ **FLOATING
C14497 S.n13107 SUB 0.91fF $ **FLOATING
C14498 S.n13108 SUB 0.05fF $ **FLOATING
C14499 S.n13109 SUB 1.88fF $ **FLOATING
C14500 S.n13110 SUB 2.67fF $ **FLOATING
C14501 S.t1236 SUB 0.02fF
C14502 S.n13111 SUB 0.24fF $ **FLOATING
C14503 S.n13112 SUB 0.36fF $ **FLOATING
C14504 S.n13113 SUB 0.61fF $ **FLOATING
C14505 S.n13114 SUB 0.12fF $ **FLOATING
C14506 S.t682 SUB 0.02fF
C14507 S.n13115 SUB 0.14fF $ **FLOATING
C14508 S.n13117 SUB 5.17fF $ **FLOATING
C14509 S.t740 SUB 0.02fF
C14510 S.n13118 SUB 0.12fF $ **FLOATING
C14511 S.n13119 SUB 0.14fF $ **FLOATING
C14512 S.t1207 SUB 0.02fF
C14513 S.n13121 SUB 0.24fF $ **FLOATING
C14514 S.n13122 SUB 0.91fF $ **FLOATING
C14515 S.n13123 SUB 0.05fF $ **FLOATING
C14516 S.n13124 SUB 0.36fF $ **FLOATING
C14517 S.n13125 SUB 0.47fF $ **FLOATING
C14518 S.n13126 SUB 1.14fF $ **FLOATING
C14519 S.n13127 SUB 1.88fF $ **FLOATING
C14520 S.n13128 SUB 0.12fF $ **FLOATING
C14521 S.t2341 SUB 0.02fF
C14522 S.n13129 SUB 0.14fF $ **FLOATING
C14523 S.t356 SUB 0.02fF
C14524 S.n13131 SUB 0.24fF $ **FLOATING
C14525 S.n13132 SUB 0.36fF $ **FLOATING
C14526 S.n13133 SUB 0.61fF $ **FLOATING
C14527 S.n13134 SUB 2.67fF $ **FLOATING
C14528 S.n13135 SUB 3.93fF $ **FLOATING
C14529 S.t2390 SUB 0.02fF
C14530 S.n13136 SUB 0.12fF $ **FLOATING
C14531 S.n13137 SUB 0.14fF $ **FLOATING
C14532 S.t329 SUB 0.02fF
C14533 S.n13139 SUB 0.24fF $ **FLOATING
C14534 S.n13140 SUB 0.91fF $ **FLOATING
C14535 S.n13141 SUB 0.05fF $ **FLOATING
C14536 S.t72 SUB 47.92fF
C14537 S.t2023 SUB 0.02fF
C14538 S.n13142 SUB 0.01fF $ **FLOATING
C14539 S.n13143 SUB 0.26fF $ **FLOATING
C14540 S.t395 SUB 0.02fF
C14541 S.n13145 SUB 1.19fF $ **FLOATING
C14542 S.n13146 SUB 0.05fF $ **FLOATING
C14543 S.t427 SUB 0.02fF
C14544 S.n13147 SUB 0.64fF $ **FLOATING
C14545 S.n13148 SUB 0.61fF $ **FLOATING
C14546 S.n13149 SUB 13.61fF $ **FLOATING
C14547 S.n13150 SUB 13.61fF $ **FLOATING
C14548 S.n13151 SUB 0.60fF $ **FLOATING
C14549 S.n13152 SUB 0.44fF $ **FLOATING
C14550 S.n13153 SUB 0.59fF $ **FLOATING
C14551 S.n13154 SUB 3.43fF $ **FLOATING
C14552 S.n13155 SUB 0.29fF $ **FLOATING
C14553 S.t180 SUB 21.38fF
C14554 S.n13156 SUB 21.67fF $ **FLOATING
C14555 S.n13157 SUB 0.77fF $ **FLOATING
C14556 S.n13158 SUB 0.28fF $ **FLOATING
C14557 S.n13159 SUB 4.50fF $ **FLOATING
C14558 S.n13160 SUB 2.33fF $ **FLOATING
C14559 S.n13161 SUB 5.58fF $ **FLOATING
C14560 S.n13162 SUB 16.08fF $ **FLOATING
C14561 S.n13163 SUB 9.28fF $ **FLOATING
C14562 S.n13164 SUB 9.29fF $ **FLOATING
C14563 S.n13165 SUB 9.29fF $ **FLOATING
C14564 S.n13166 SUB 9.29fF $ **FLOATING
C14565 S.n13167 SUB 9.29fF $ **FLOATING
C14566 S.n13168 SUB 9.29fF $ **FLOATING
C14567 S.n13169 SUB 9.29fF $ **FLOATING
C14568 S.n13170 SUB 9.29fF $ **FLOATING
C14569 S.n13171 SUB 9.29fF $ **FLOATING
C14570 S.n13172 SUB 9.29fF $ **FLOATING
C14571 S.n13173 SUB 9.29fF $ **FLOATING
C14572 S.n13174 SUB 9.29fF $ **FLOATING
C14573 S.n13175 SUB 9.29fF $ **FLOATING
C14574 S.n13176 SUB 9.29fF $ **FLOATING
C14575 S.n13177 SUB 9.39fF $ **FLOATING
C14576 S.n13178 SUB 17.77fF $ **FLOATING
.ends

