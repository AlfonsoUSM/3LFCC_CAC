magic
tech sky130A
timestamp 1679234436
<< checkpaint >>
rect -6555 -6605 7705 7655
<< dnwell >>
rect -3475 -3525 4625 4575
<< nwell >>
rect -5925 2225 7075 7025
rect -5925 -1175 -1125 2225
rect 2275 -1175 7075 2225
rect -5925 -5975 7075 -1175
<< pwell >>
rect -1125 1100 0 2225
rect 1100 1100 2275 2225
rect -1125 -1175 0 0
rect 1100 -1175 2275 0
<< mvnmos >>
rect 1100 1131 1150 1569
rect -469 -50 -31 0
rect 1181 -50 1619 0
rect 1100 -519 1150 -81
<< mvndiff >>
rect 1179 1569 1621 1571
rect -29 1563 0 1569
rect -29 1164 -23 1563
rect -64 1137 -23 1164
rect -6 1137 0 1563
rect -64 1131 0 1137
rect 1097 1131 1100 1569
rect 1150 1563 1621 1569
rect 1150 1137 1156 1563
rect 1173 1515 1621 1563
rect 1173 1185 1235 1515
rect 1565 1185 1621 1515
rect 1173 1137 1621 1185
rect 1150 1131 1621 1137
rect -64 1129 -31 1131
rect -469 1123 -31 1129
rect -469 1106 -463 1123
rect -37 1106 -31 1123
rect -469 1100 -31 1106
rect 1179 1129 1621 1131
rect 1181 1123 1619 1129
rect 1181 1106 1187 1123
rect 1613 1106 1619 1123
rect 1181 1100 1619 1106
rect -469 0 -31 3
rect 1181 0 1619 3
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 1181 -56 1619 -50
rect 1181 -73 1187 -56
rect 1613 -73 1619 -56
rect 1181 -79 1619 -73
rect 1181 -81 1214 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 1097 -519 1100 -81
rect 1150 -87 1214 -81
rect 1150 -513 1156 -87
rect 1173 -114 1214 -87
rect 1173 -513 1179 -114
rect 1150 -519 1179 -513
rect -471 -521 -29 -519
<< mvndiffc >>
rect -23 1137 -6 1563
rect 1156 1137 1173 1563
rect -463 1106 -37 1123
rect 1187 1106 1613 1123
rect -463 -73 -37 -56
rect 1187 -73 1613 -56
rect -23 -513 -6 -87
rect 1156 -513 1173 -87
<< mvpsubdiff >>
rect -1025 2113 0 2125
rect -1025 1117 -1013 2113
rect -19 1837 0 2113
rect -737 1825 0 1837
rect 1100 2113 2175 2125
rect 1100 1825 1887 1837
rect -737 1117 -725 1825
rect -1025 1100 -725 1117
rect 1235 1503 1565 1515
rect 1235 1197 1247 1503
rect 1553 1197 1565 1503
rect 1235 1185 1565 1197
rect 1875 1117 1887 1825
rect 2163 1117 2175 2113
rect 1875 1100 2175 1117
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 1875 -775 1887 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 1100 -787 1887 -775
rect 2163 -1063 2175 0
rect 1100 -1075 2175 -1063
<< mvnsubdiff >>
rect -5525 6613 6675 6625
rect -5525 -5563 -5513 6613
rect -1537 2625 2687 2637
rect -1537 -1575 -1525 2625
rect 2675 -1575 2687 2625
rect -1537 -1587 2687 -1575
rect 6663 -5563 6675 6613
rect -5525 -5575 6675 -5563
<< mvpsubdiffcont >>
rect -1013 1837 -19 2113
rect -1013 1117 -737 1837
rect 1100 1837 2163 2113
rect 1247 1197 1553 1503
rect 1887 1117 2163 1837
rect -1013 -787 -737 0
rect -403 -453 -97 -147
rect -1013 -1063 -17 -787
rect 1887 -787 2163 0
rect 1100 -1063 2163 -787
<< mvnsubdiffcont >>
rect -5513 2637 6663 6613
rect -5513 -1587 -1537 2637
rect 2687 -1587 6663 2637
rect -5513 -5563 6663 -1587
<< poly >>
rect -550 1642 0 1650
rect -550 1608 -542 1642
rect -508 1608 0 1642
rect -550 1600 0 1608
rect 1100 1642 1700 1650
rect 1100 1608 1108 1642
rect 1142 1608 1658 1642
rect 1692 1608 1700 1642
rect 1100 1600 1700 1608
rect -550 1100 -500 1600
rect 1100 1569 1150 1600
rect 1100 1100 1150 1131
rect 1650 1100 1700 1600
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -50 0 0
rect 1100 -8 1181 0
rect 1100 -42 1108 -8
rect 1142 -42 1181 -8
rect 1100 -50 1181 -42
rect 1619 -8 1700 0
rect 1619 -42 1658 -8
rect 1692 -42 1700 -8
rect 1619 -50 1700 -42
rect -550 -550 -500 -50
rect 1100 -81 1150 -50
rect 1100 -550 1150 -519
rect 1650 -550 1700 -50
rect -550 -558 0 -550
rect -550 -592 -542 -558
rect -508 -592 0 -558
rect -550 -600 0 -592
rect 1100 -558 1700 -550
rect 1100 -592 1108 -558
rect 1142 -592 1658 -558
rect 1692 -592 1700 -558
rect 1100 -600 1700 -592
<< polycont >>
rect -542 1608 -508 1642
rect 1108 1608 1142 1642
rect 1658 1608 1692 1642
rect -542 -42 -508 -8
rect 1108 -42 1142 -8
rect 1658 -42 1692 -8
rect -542 -592 -508 -558
rect 1108 -592 1142 -558
rect 1658 -592 1692 -558
<< locali >>
rect -5525 6613 6675 6625
rect -5525 -5563 -5513 6613
rect -1537 2625 2687 2637
rect -1537 -1575 -1525 2625
rect -1025 2113 0 2125
rect -1025 1117 -1013 2113
rect -19 1837 0 2113
rect -737 1825 0 1837
rect 1100 2113 2175 2125
rect 1100 1825 1887 1837
rect -737 1117 -725 1825
rect -550 1642 -500 1650
rect -550 1608 -542 1642
rect -508 1608 -500 1642
rect -550 1600 -500 1608
rect 1100 1642 1150 1650
rect 1100 1608 1108 1642
rect 1142 1608 1150 1642
rect 1100 1600 1150 1608
rect 1650 1642 1700 1650
rect 1650 1608 1658 1642
rect 1692 1608 1700 1642
rect 1650 1600 1700 1608
rect 1173 1571 1627 1577
rect -23 1563 -6 1571
rect -64 1137 -23 1164
rect -64 1129 -6 1137
rect 1156 1563 1627 1571
rect 1173 1515 1627 1563
rect 1173 1185 1235 1515
rect 1565 1185 1627 1515
rect 1173 1137 1627 1185
rect 1156 1129 1627 1137
rect -64 1123 -29 1129
rect 1173 1123 1627 1129
rect -1025 1100 -725 1117
rect -471 1106 -463 1123
rect -37 1106 -29 1123
rect 1179 1106 1187 1123
rect 1613 1106 1621 1123
rect 1875 1117 1887 1825
rect 2163 1117 2175 2113
rect 1875 1100 2175 1117
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 1100 -8 1150 0
rect 1100 -42 1108 -8
rect 1142 -42 1150 -8
rect 1100 -50 1150 -42
rect 1650 -8 1700 0
rect 1650 -42 1658 -8
rect 1692 -42 1700 -8
rect 1650 -50 1700 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 1179 -73 1187 -56
rect 1613 -73 1621 -56
rect -477 -79 -23 -73
rect 1179 -79 1214 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 1156 -87 1214 -79
rect 1173 -114 1214 -87
rect 1156 -521 1173 -513
rect -477 -527 -23 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 1100 -558 1150 -550
rect 1100 -592 1108 -558
rect 1142 -592 1150 -558
rect 1100 -600 1150 -592
rect 1650 -558 1700 -550
rect 1650 -592 1658 -558
rect 1692 -592 1700 -558
rect 1650 -600 1700 -592
rect 1875 -775 1887 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 1100 -787 1887 -775
rect 2163 -1063 2175 0
rect 1100 -1075 2175 -1063
rect 2675 -1575 2687 2625
rect -1537 -1587 2687 -1575
rect 6663 -5563 6675 6613
rect -5525 -5575 6675 -5563
<< viali >>
rect -5513 2637 6663 6613
rect -5513 -1587 -1537 2637
rect -1013 1837 -19 2113
rect -1013 1119 -737 1837
rect 1100 1837 2163 2113
rect -542 1608 -508 1642
rect 1108 1608 1142 1642
rect 1658 1608 1692 1642
rect -23 1137 -6 1563
rect 1156 1137 1173 1563
rect 1235 1503 1565 1515
rect 1235 1197 1247 1503
rect 1247 1197 1553 1503
rect 1553 1197 1565 1503
rect 1235 1185 1565 1197
rect -463 1106 -37 1123
rect 1187 1106 1613 1123
rect 1887 1119 2163 1837
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 1108 -42 1142 -8
rect 1658 -42 1692 -8
rect -463 -73 -37 -56
rect 1187 -73 1613 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 1156 -513 1173 -87
rect -542 -592 -508 -558
rect 1108 -592 1142 -558
rect 1658 -592 1692 -558
rect -1013 -1063 -19 -787
rect 1887 -787 2163 0
rect 1100 -1063 2163 -787
rect 2687 -1587 6663 2637
rect -5513 -5563 6663 -1587
<< metal1 >>
rect -5525 6613 6675 6625
rect -5525 -5563 -5513 6613
rect -1537 2625 2687 2637
rect -1537 -1575 -1525 2625
rect -1025 2113 0 2125
rect -1025 1119 -1013 2113
rect -19 1837 0 2113
rect -737 1825 0 1837
rect 1100 2113 2175 2125
rect 1100 1825 1887 1837
rect -737 1119 -725 1825
rect -550 1642 -500 1650
rect -550 1608 -542 1642
rect -508 1608 -500 1642
rect -550 1600 -500 1608
rect 1100 1642 1150 1650
rect 1100 1608 1108 1642
rect 1142 1608 1150 1642
rect 1100 1600 1150 1608
rect 1650 1642 1700 1650
rect 1650 1608 1658 1642
rect 1692 1608 1700 1642
rect 1650 1600 1700 1608
rect -474 1569 -26 1574
rect 1176 1569 1624 1574
rect -474 1563 -3 1569
rect -474 1515 -23 1563
rect -474 1185 -415 1515
rect -85 1185 -23 1515
rect -474 1137 -23 1185
rect -6 1137 -3 1563
rect -474 1131 -3 1137
rect 1153 1563 1624 1569
rect 1153 1137 1156 1563
rect 1173 1515 1624 1563
rect 1173 1185 1235 1515
rect 1565 1185 1624 1515
rect 1173 1137 1624 1185
rect 1153 1131 1624 1137
rect -474 1126 -26 1131
rect 1176 1126 1624 1131
rect -1025 1100 -725 1119
rect -469 1123 -31 1126
rect -469 1106 -463 1123
rect -37 1106 -31 1123
rect -469 1103 -31 1106
rect 1181 1123 1619 1126
rect 1181 1106 1187 1123
rect 1613 1106 1619 1123
rect 1181 1103 1619 1106
rect 1875 1119 1887 1825
rect 2163 1119 2175 2113
rect 1875 1100 2175 1119
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 1100 -8 1150 0
rect 1100 -42 1108 -8
rect 1142 -42 1150 -8
rect 1100 -50 1150 -42
rect 1650 -8 1700 0
rect 1650 -42 1658 -8
rect 1692 -42 1700 -8
rect 1650 -50 1700 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 1181 -56 1619 -53
rect 1181 -73 1187 -56
rect 1613 -73 1619 -56
rect 1181 -76 1619 -73
rect -474 -81 -26 -76
rect 1176 -81 1624 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 1153 -87 1624 -81
rect 1153 -513 1156 -87
rect 1173 -135 1624 -87
rect 1173 -465 1235 -135
rect 1565 -465 1624 -135
rect 1173 -513 1624 -465
rect 1153 -519 1624 -513
rect -474 -524 -26 -519
rect 1176 -524 1624 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 1100 -558 1150 -550
rect 1100 -592 1108 -558
rect 1142 -592 1150 -558
rect 1100 -600 1150 -592
rect 1650 -558 1700 -550
rect 1650 -592 1658 -558
rect 1692 -592 1700 -558
rect 1650 -600 1700 -592
rect 1875 -775 1887 0
rect -737 -787 0 -775
rect -19 -1063 0 -787
rect -1025 -1075 0 -1063
rect 1100 -787 1887 -775
rect 2163 -1063 2175 0
rect 1100 -1075 2175 -1063
rect 2675 -1575 2687 2625
rect -1537 -1587 2687 -1575
rect 6663 -5563 6675 6613
rect -5525 -5575 6675 -5563
<< via1 >>
rect -5513 2637 6663 6613
rect -5513 1117 -1537 2625
rect 1188 1925 1288 2025
rect -542 1608 -508 1642
rect 1108 1608 1142 1642
rect 1658 1608 1692 1642
rect -415 1185 -85 1515
rect 1235 1185 1565 1515
rect 1975 1138 2075 1238
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 1108 -42 1142 -8
rect 1658 -42 1692 -8
rect -415 -465 -85 -135
rect 1235 -465 1565 -135
rect -542 -592 -508 -558
rect 1108 -592 1142 -558
rect 1658 -592 1692 -558
rect -138 -975 -38 -875
rect 2687 -1587 6663 2637
rect -495 -5563 6663 -1587
<< metal2 >>
rect -5525 6613 6675 6625
rect -5525 2637 -5513 6613
rect -5525 2625 2687 2637
rect -5525 1117 -5513 2625
rect -1537 1117 -1525 2625
rect 1178 2025 1298 2035
rect 1178 1925 1188 2025
rect 1288 1925 1298 2025
rect 1178 1915 1298 1925
rect -725 1642 0 1825
rect -725 1608 -542 1642
rect -508 1608 0 1642
rect -725 1600 0 1608
rect 1100 1642 1875 1825
rect 1100 1608 1108 1642
rect 1142 1608 1658 1642
rect 1692 1608 1875 1642
rect 1100 1600 1875 1608
rect -725 1100 -500 1600
rect -425 1515 -75 1525
rect -425 1185 -415 1515
rect -85 1185 -75 1515
rect -425 1175 -75 1185
rect 1100 1100 1150 1600
rect 1225 1515 1575 1525
rect 1225 1185 1235 1515
rect 1565 1185 1575 1515
rect 1225 1175 1575 1185
rect 1650 1100 1875 1600
rect 1965 1238 2085 1248
rect 1965 1138 1975 1238
rect 2075 1138 2085 1238
rect 1965 1128 2085 1138
rect -725 -8 0 0
rect -725 -42 -542 -8
rect -508 -42 0 -8
rect -725 -50 0 -42
rect 1100 -8 1875 0
rect 1100 -42 1108 -8
rect 1142 -42 1658 -8
rect 1692 -42 1875 -8
rect 1100 -50 1875 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 1100 -550 1150 -50
rect 1225 -135 1575 -125
rect 1225 -465 1235 -135
rect 1565 -465 1575 -135
rect 1225 -475 1575 -465
rect 1650 -550 1875 -50
rect -725 -558 0 -550
rect -725 -592 -542 -558
rect -508 -592 0 -558
rect -725 -775 0 -592
rect 1100 -558 1875 -550
rect 1100 -592 1108 -558
rect 1142 -592 1658 -558
rect 1692 -592 1875 -558
rect 1100 -775 1875 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
rect 2675 -1575 2687 2625
rect -507 -1587 2687 -1575
rect -507 -5563 -495 -1587
rect 6663 -5563 6675 6613
rect -507 -5575 6675 -5563
<< via2 >>
rect 1188 1925 1288 2025
rect -310 1290 -190 1410
rect 1340 1290 1460 1410
rect 1975 1138 2075 1238
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 1340 -360 1460 -240
rect -138 -975 -38 -875
<< metal3 >>
rect -2525 2625 1675 3625
rect -2525 1738 -1525 2625
rect -638 1738 -186 2625
rect -2525 1414 -186 1738
rect -88 1512 0 2125
tri -186 1414 -88 1512 sw
tri -88 1424 0 1512 ne
rect 1100 2025 1464 2125
rect 1100 1925 1188 2025
rect 1288 1925 1464 2025
rect 1100 1424 1464 1925
rect -2525 1410 -88 1414
rect -2525 1290 -310 1410
rect -190 1326 -88 1410
tri -88 1326 0 1414 sw
rect -190 1290 0 1326
rect -2525 1286 0 1290
rect -2525 -575 -1525 1286
tri -412 1188 -314 1286 ne
rect -314 1188 0 1286
rect -1025 1100 -412 1188
tri -412 1100 -324 1188 sw
tri -314 1100 -226 1188 ne
rect -226 1100 0 1188
tri 1100 1326 1198 1424 ne
rect 1198 1414 1464 1424
tri 1464 1414 1562 1512 sw
rect 2675 1414 3675 1625
rect 1198 1410 3675 1414
rect 1198 1326 1340 1410
tri 1100 1238 1188 1326 sw
tri 1198 1238 1286 1326 ne
rect 1286 1290 1340 1326
rect 1460 1290 3675 1410
rect 1286 1238 3675 1290
rect 1100 1158 1188 1238
tri 1188 1158 1268 1238 sw
tri 1286 1158 1366 1238 ne
rect 1366 1158 1975 1238
rect 1100 1100 1268 1158
tri 1268 1100 1326 1158 sw
tri 1366 1100 1424 1158 ne
rect 1424 1138 1975 1158
rect 2075 1138 3675 1238
rect 1424 1100 3675 1138
rect 2675 0 3675 1100
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 1100 -40 1326 0
tri 1326 -40 1366 0 sw
tri 1424 -40 1464 0 ne
rect 1464 -40 3675 0
rect 1100 -138 1366 -40
tri 1366 -138 1464 -40 sw
tri 1464 -138 1562 -40 ne
rect 1562 -138 3675 -40
rect 1100 -226 1464 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 1100 -324 1198 -226 ne
rect 1198 -236 1464 -226
tri 1464 -236 1562 -138 sw
rect 1198 -240 2175 -236
rect 1198 -324 1340 -240
tri 1100 -364 1140 -324 sw
tri 1198 -364 1238 -324 ne
rect 1238 -360 1340 -324
rect 1460 -360 2175 -240
rect 1238 -364 2175 -360
rect 1100 -462 1140 -364
tri 1140 -462 1238 -364 sw
tri 1238 -462 1336 -364 ne
rect 1100 -1575 1238 -462
rect 1336 -688 2175 -364
rect 1336 -1075 1788 -688
rect 2675 -1575 3675 -138
rect -525 -2575 3675 -1575
<< via3 >>
rect 1188 1925 1288 2025
rect -310 1290 -190 1410
rect 1340 1290 1460 1410
rect 1975 1138 2075 1238
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect -138 -975 -38 -875
rect 1340 -360 1460 -240
<< metal4 >>
rect -2525 2625 1675 3625
rect -2525 1738 -1525 2625
rect -638 1738 -186 2625
rect -2525 1414 -186 1738
rect -88 1512 0 2125
tri -186 1414 -88 1512 sw
tri -88 1424 0 1512 ne
rect 1100 2025 1464 2125
rect 1100 1925 1188 2025
rect 1288 1925 1464 2025
rect 1100 1424 1464 1925
rect -2525 1410 -88 1414
rect -2525 1290 -310 1410
rect -190 1326 -88 1410
tri -88 1326 0 1414 sw
rect -190 1290 0 1326
rect -2525 1286 0 1290
rect -2525 -575 -1525 1286
tri -412 1188 -314 1286 ne
rect -314 1188 0 1286
rect -1025 1100 -412 1188
tri -412 1100 -324 1188 sw
tri -314 1100 -226 1188 ne
rect -226 1100 0 1188
tri 1100 1326 1198 1424 ne
rect 1198 1414 1464 1424
tri 1464 1414 1562 1512 sw
rect 2675 1414 3675 1625
rect 1198 1410 3675 1414
rect 1198 1326 1340 1410
tri 1100 1238 1188 1326 sw
tri 1198 1238 1286 1326 ne
rect 1286 1290 1340 1326
rect 1460 1290 3675 1410
rect 1286 1238 3675 1290
rect 1100 1158 1188 1238
tri 1188 1158 1268 1238 sw
tri 1286 1158 1366 1238 ne
rect 1366 1158 1975 1238
rect 1100 1100 1268 1158
tri 1268 1100 1326 1158 sw
tri 1366 1100 1424 1158 ne
rect 1424 1138 1975 1158
rect 2075 1138 3675 1238
rect 1424 1100 3675 1138
rect 2675 0 3675 1100
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 1100 -40 1326 0
tri 1326 -40 1366 0 sw
tri 1424 -40 1464 0 ne
rect 1464 -40 3675 0
rect 1100 -138 1366 -40
tri 1366 -138 1464 -40 sw
tri 1464 -138 1562 -40 ne
rect 1562 -138 3675 -40
rect 1100 -226 1464 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 1100 -324 1198 -226 ne
rect 1198 -236 1464 -226
tri 1464 -236 1562 -138 sw
rect 1198 -240 2175 -236
rect 1198 -324 1340 -240
tri 1100 -364 1140 -324 sw
tri 1198 -364 1238 -324 ne
rect 1238 -360 1340 -324
rect 1460 -360 2175 -240
rect 1238 -364 2175 -360
rect 1100 -462 1140 -364
tri 1140 -462 1238 -364 sw
tri 1238 -462 1336 -364 ne
rect 1100 -1575 1238 -462
rect 1336 -688 2175 -364
rect 1336 -1075 1788 -688
rect 2675 -1575 3675 -138
rect -525 -2575 3675 -1575
<< via4 >>
rect -310 1290 -190 1410
rect 1340 1290 1460 1410
rect -310 -360 -190 -240
rect 1340 -360 1460 -240
<< metal5 >>
rect -2525 2625 1675 3625
rect -2525 1703 -1525 2625
rect -603 1703 -292 2625
rect -2525 1410 -292 1703
tri -292 1410 -154 1548 sw
rect -53 1547 0 2125
tri -53 1494 0 1547 ne
rect 1100 1494 1358 2125
rect -2525 1392 -310 1410
rect -2525 -575 -1525 1392
tri -448 1290 -346 1392 ne
rect -346 1290 -310 1392
rect -190 1290 -154 1410
rect -1025 1100 -447 1153
tri -447 1100 -394 1153 sw
tri -346 1100 -156 1290 ne
rect -156 1256 -154 1290
tri -154 1256 0 1410 sw
rect -156 1100 0 1256
tri 1100 1256 1338 1494 ne
rect 1338 1410 1358 1494
tri 1358 1410 1496 1548 sw
rect 1338 1290 1340 1410
rect 1460 1308 1496 1410
tri 1496 1308 1598 1410 sw
rect 2675 1308 3675 1625
rect 1460 1290 3675 1308
rect 1338 1256 3675 1290
tri 1100 1100 1256 1256 sw
tri 1338 1100 1494 1256 ne
rect 1494 1100 3675 1256
rect 2675 0 3675 1100
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 0 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -156 0 -103 ne
rect 1100 -103 1256 0
tri 1256 -103 1359 0 sw
tri 1494 -103 1597 0 ne
rect 1597 -103 3675 0
rect 1100 -156 1359 -103
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
rect -208 -1575 0 -394
tri 1100 -394 1338 -156 ne
rect 1338 -240 1359 -156
tri 1359 -240 1496 -103 sw
rect 1338 -360 1340 -240
rect 1460 -342 1496 -240
tri 1496 -342 1598 -240 sw
rect 1460 -360 2175 -342
rect 1338 -394 2175 -360
tri 1100 -497 1203 -394 sw
rect 1100 -1575 1203 -497
tri 1338 -498 1442 -394 ne
rect 1442 -653 2175 -394
rect 1442 -1075 1753 -653
rect 2675 -1575 3675 -103
rect -525 -2575 3675 -1575
use nmos_drain_frame_lt  nmos_drain_frame_lt_0 waffle_cells
timestamp 1675431365
transform 1 0 -550 0 1 0
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_1
timestamp 1675431365
transform 0 -1 1100 -1 0 1650
box -975 -113 663 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_0 waffle_cells
timestamp 1675431051
transform 0 -1 550 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_1
timestamp 1675431051
transform 1 0 1100 0 1 550
box -113 -113 1575 663
use nmos_drain_in  nmos_drain_in_0 waffle_cells
timestamp 1675431861
transform 1 0 0 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_1
timestamp 1675431861
transform 1 0 550 0 1 0
box -113 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_0 waffle_cells
timestamp 1675431308
transform 0 -1 550 -1 0 1650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_1
timestamp 1675431308
transform 1 0 -550 0 1 550
box -975 -113 663 663
use nmos_source_frame_rb  nmos_source_frame_rb_0 waffle_cells
timestamp 1675430904
transform 1 0 1100 0 1 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_1
timestamp 1675430904
transform 0 -1 1100 -1 0 0
box -113 -113 1575 663
use nmos_source_in  nmos_source_in_0 waffle_cells
timestamp 1675431769
transform 1 0 0 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_1
timestamp 1675431769
transform 1 0 550 0 1 550
box -113 -113 663 663
<< properties >>
string MASKHINTS_HVI -140 2200 0 2340 -140 -140 0 0 2200 -140 2340 0 2200 2200 2340 2340
string MASKHINTS_HVNTM -1007 -1107 -21 -1079 -1007 -1079 -979 -121 2321 3179 3307 3207 3279 2221 3307 3179 -170 2230 -30 2370
<< end >>
