* NGSPICE file created from mag_files/POSTLAYOUT/nmos_flat_8x8.ext - technology: sky130A

.subckt nmos_flat_8x8 G S D DNW VSUBS
X0 S.t126 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X1 S.t125 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2 D G S.t124 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3 D G S.t123 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4 D G S.t122 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5 D G S.t121 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6 S.t120 G D S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7 D G S.t119 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8 S.t118 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9 S.t117 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10 S.t116 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11 S.t115 G D S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12 D G S.t114 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13 S.t113 G D S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X14 S.t112 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X15 D G S.t111 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X16 D G S.t110 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X17 D G S.t109 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X18 S.t108 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X19 S.t107 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X20 S.t106 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X21 D G S.t105 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X22 S.t104 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X23 D G S.t103 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X24 D G S.t102 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X25 D G S.t101 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X26 D G S.t100 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X27 D G S.t99 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X28 D G S.t98 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X29 D G S.t97 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X30 S.t96 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X31 D G S.t95 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X32 S.t94 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X33 S.t93 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X34 S.t92 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X35 S.t91 G D S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X36 S.t90 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X37 S.t89 G D S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X38 S.t88 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X39 D G S.t87 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X40 D G S.t86 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X41 D G S.t85 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X42 D G S.t84 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X43 D G S.t83 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X44 D G S.t82 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X45 S.t81 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X46 D G S.t80 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X47 S.t79 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X48 D G S.t78 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X49 D G S.t77 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X50 S.t76 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X51 S.t75 G D S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X52 D G S.t74 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X53 S.t73 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X54 S.t72 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X55 S.t71 G D S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X56 D G S.t70 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X57 S.t69 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X58 D G S.t68 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X59 D G S.t67 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X60 D G S.t66 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X61 D G S.t65 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X62 D G S.t64 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X63 D G S.t63 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X64 S.t62 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X65 D G S.t61 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X66 D G S.t60 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X67 S.t59 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X68 S.t58 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X69 S.t57 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X70 S.t56 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X71 S.t55 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X72 D G S.t54 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X73 S.t53 G D S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X74 D G S.t52 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X75 D G S.t51 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X76 D G S.t50 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X77 S.t49 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X78 D G S.t48 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X79 S.t46 G D S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X80 S.t45 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X81 S.t44 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X82 D G S.t43 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X83 S.t41 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X84 D G S.t39 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X85 D G S.t38 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X86 S.t37 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X87 D G S.t36 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X88 D G S.t35 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X89 S.t33 G D S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X90 S.t31 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X91 D G S.t30 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X92 S.t28 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X93 S.t27 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X94 S.t26 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X95 D G S.t25 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X96 S.t24 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X97 D G S.t23 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X98 D G S.t22 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X99 D G S.t21 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X100 D G S.t20 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X101 S.t18 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X102 D G S.t16 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X103 S.t14 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X104 S.t12 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X105 D G S.t11 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X106 S.t9 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X107 S.t7 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X108 S.t6 G D S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X109 S.t4 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X110 D G S.t3 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X111 S.t1 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
R0 S.t47 S.t8 216.071
R1 S.n162 S.t15 188.571
R2 S.n60 S.t13 188.571
R3 S.n483 S.t19 188.571
R4 S.n557 S.t2 188.571
R5 S.n413 S.t10 188.571
R6 S.n256 S.t29 188.571
R7 S.t40 S.n150 182.285
R8 S.t0 S.n91 182.285
R9 S.t42 S.n513 182.285
R10 S.t5 S.n604 182.285
R11 S.t17 S.n382 182.285
R12 S.t34 S.n288 182.285
R13 S.t32 S.n424 182.285
R14 S.n160 S.n158 169.353
R15 S.n481 S.n480 169.353
R16 S.n411 S.n410 169.353
R17 S.n160 S.n159 169.353
R18 S.n409 S.n408 137.98
R19 S.n479 S.n478 137.98
R20 S.n157 S.n156 137.98
R21 S.n58 S.n57 135.611
R22 S.n555 S.n554 135.611
R23 S.n254 S.n253 135.611
R24 S.n264 S.n263 91.65
R25 S.n70 S.n69 91.65
R26 S.n567 S.n566 91.65
R27 S.n404 S.n403 91.389
R28 S.n637 S.n636 91.389
R29 S.n175 S.n174 91.389
R30 S.n231 S.n230 87.222
R31 S.n212 S.n211 87.222
R32 S.n16 S.n15 87.222
R33 S.n465 S.n464 86.961
R34 S.n450 S.n449 86.961
R35 S.n439 S.n438 86.961
R36 S.n423 S.t85 3.904
R37 S.n422 S.t64 3.904
R38 S.n404 S.t102 3.904
R39 S.n352 S.t25 3.904
R40 S.n465 S.t60 3.904
R41 S.n463 S.t36 3.904
R42 S.n299 S.n298 3.904
R43 S.n307 S.t38 3.904
R44 S.n310 S.t11 3.904
R45 S.n302 S.n301 3.904
R46 S.n390 S.n389 3.904
R47 S.n398 S.t80 3.904
R48 S.n401 S.t3 3.904
R49 S.n393 S.n392 3.904
R50 S.n591 S.n590 3.904
R51 S.n602 S.t100 3.904
R52 S.n599 S.t54 3.904
R53 S.n594 S.n593 3.904
R54 S.n637 S.t124 3.904
R55 S.n639 S.t70 3.904
R56 S.n232 S.t109 3.904
R57 S.n135 S.n134 3.904
R58 S.n148 S.t83 3.904
R59 S.n145 S.t21 3.904
R60 S.n132 S.n131 3.904
R61 S.n360 S.n359 3.904
R62 S.n380 S.t39 3.904
R63 S.n377 S.t68 3.904
R64 S.n357 S.n356 3.904
R65 S.n576 S.n575 3.904
R66 S.n585 S.t123 3.904
R67 S.n582 S.t20 3.904
R68 S.n573 S.n572 3.904
R69 S.n496 S.n495 3.904
R70 S.n511 S.t84 3.904
R71 S.n508 S.t67 3.904
R72 S.n493 S.n492 3.904
R73 S.n122 S.n121 3.904
R74 S.n119 S.t121 3.904
R75 S.n116 S.t16 3.904
R76 S.n50 S.n49 3.904
R77 S.n210 S.t87 3.904
R78 S.n24 S.n23 3.904
R79 S.n180 S.t51 3.904
R80 S.n183 S.t23 3.904
R81 S.n186 S.n185 3.904
R82 S.n71 S.t99 3.904
R83 S.n81 S.n80 3.904
R84 S.n89 S.t52 3.904
R85 S.n86 S.t65 3.904
R86 S.n78 S.n77 3.904
R87 S.n525 S.n524 3.904
R88 S.n533 S.t122 3.904
R89 S.n536 S.t103 3.904
R90 S.n528 S.n527 3.904
R91 S.n568 S.t66 3.904
R92 S.n14 S.t48 3.904
R93 S.n29 S.n28 3.904
R94 S.n45 S.t119 3.904
R95 S.n42 S.t101 3.904
R96 S.n32 S.n31 3.904
R97 S.n175 S.t74 3.904
R98 S.n177 S.t105 3.904
R99 S.n100 S.n99 3.904
R100 S.n110 S.t50 3.904
R101 S.n113 S.t111 3.904
R102 S.n103 S.n102 3.904
R103 S.n623 S.n622 3.904
R104 S.n631 S.t43 3.904
R105 S.n634 S.t77 3.904
R106 S.n626 S.n625 3.904
R107 S.n544 S.n543 3.904
R108 S.n606 S.t86 3.904
R109 S.n609 S.t98 3.904
R110 S.n612 S.n611 3.904
R111 S.n334 S.n333 3.904
R112 S.n350 S.t114 3.904
R113 S.n347 S.t22 3.904
R114 S.n337 S.n336 3.904
R115 S.n245 S.n244 3.904
R116 S.n314 S.t82 3.904
R117 S.n317 S.t61 3.904
R118 S.n320 S.n319 3.904
R119 S.n450 S.t95 3.904
R120 S.n445 S.t78 3.904
R121 S.n439 S.t30 3.904
R122 S.n437 S.t110 3.904
R123 S.n275 S.n274 3.904
R124 S.n286 S.t35 3.904
R125 S.n283 S.t63 3.904
R126 S.n278 S.n277 3.904
R127 S.n247 S.t97 3.904
R128 S.n264 S.t89 3.643
R129 S.n242 S.t26 3.643
R130 S.n462 S.t33 3.643
R131 S.n299 S.t120 3.643
R132 S.n307 S.n306 3.643
R133 S.n310 S.n309 3.643
R134 S.n302 S.t49 3.643
R135 S.n390 S.t18 3.643
R136 S.n398 S.n397 3.643
R137 S.n401 S.n400 3.643
R138 S.n393 S.t79 3.643
R139 S.n591 S.t71 3.643
R140 S.n602 S.n601 3.643
R141 S.n599 S.n598 3.643
R142 S.n594 S.t117 3.643
R143 S.n641 S.t108 3.643
R144 S.n229 S.t92 3.643
R145 S.n214 S.t62 3.643
R146 S.n231 S.t12 3.643
R147 S.n233 S.t76 3.643
R148 S.n135 S.t107 3.643
R149 S.n148 S.n147 3.643
R150 S.n145 S.n144 3.643
R151 S.n132 S.t55 3.643
R152 S.n360 S.t37 3.643
R153 S.n380 S.n379 3.643
R154 S.n377 S.n376 3.643
R155 S.n357 S.t69 3.643
R156 S.n576 S.t91 3.643
R157 S.n585 S.n584 3.643
R158 S.n582 S.n581 3.643
R159 S.n573 S.t59 3.643
R160 S.n496 S.t81 3.643
R161 S.n511 S.n510 3.643
R162 S.n508 S.n507 3.643
R163 S.n493 S.t106 3.643
R164 S.n122 S.t90 3.643
R165 S.n119 S.n118 3.643
R166 S.n116 S.n115 3.643
R167 S.n50 S.t58 3.643
R168 S.n212 S.t9 3.643
R169 S.n213 S.t56 3.643
R170 S.n24 S.t41 3.643
R171 S.n180 S.n179 3.643
R172 S.n183 S.n182 3.643
R173 S.n186 S.t72 3.643
R174 S.n70 S.t57 3.643
R175 S.n52 S.t14 3.643
R176 S.n81 S.t1 3.643
R177 S.n89 S.n88 3.643
R178 S.n86 S.n85 3.643
R179 S.n78 S.t94 3.643
R180 S.n525 S.t118 3.643
R181 S.n533 S.n532 3.643
R182 S.n536 S.n535 3.643
R183 S.n528 S.t28 3.643
R184 S.n567 S.t6 3.643
R185 S.n546 S.t96 3.643
R186 S.n16 S.t93 3.643
R187 S.n17 S.t125 3.643
R188 S.n29 S.t116 3.643
R189 S.n45 S.n44 3.643
R190 S.n42 S.n41 3.643
R191 S.n32 S.t27 3.643
R192 S.n167 S.t31 3.643
R193 S.n100 S.t4 3.643
R194 S.n110 S.n109 3.643
R195 S.n113 S.n112 3.643
R196 S.n103 S.t73 3.643
R197 S.n623 S.t44 3.643
R198 S.n631 S.n630 3.643
R199 S.n634 S.n633 3.643
R200 S.n626 S.t104 3.643
R201 S.n544 S.t53 3.643
R202 S.n606 S.n605 3.643
R203 S.n609 S.n608 3.643
R204 S.n612 S.t7 3.643
R205 S.n334 S.t112 3.643
R206 S.n350 S.n349 3.643
R207 S.n347 S.n346 3.643
R208 S.n337 S.t24 3.643
R209 S.n245 S.t46 3.643
R210 S.n314 S.n313 3.643
R211 S.n317 S.n316 3.643
R212 S.n320 S.t88 3.643
R213 S.n444 S.t75 3.643
R214 S.n440 S.t115 3.643
R215 S.n275 S.t113 3.643
R216 S.n286 S.n285 3.643
R217 S.n283 S.n282 3.643
R218 S.n278 S.t45 3.643
R219 S.n312 S.t126 3.643
R220 S.n60 S.n58 2.799
R221 S.n557 S.n555 2.799
R222 S.n256 S.n254 2.799
R223 S.n222 S.n221 2.645
R224 S.n54 S.n53 2.645
R225 S.n551 S.n550 2.645
R226 S.n474 S.n471 0.178
R227 S.n164 S.n163 0.172
R228 S.n224 S.n220 0.164
R229 S.n477 S.n476 0.143
R230 S.n241 S.n238 0.123
R231 S.n443 S.n442 0.11
R232 S.n477 S.n419 0.11
R233 S.n75 S.n74 0.109
R234 S.n107 S.n106 0.109
R235 S.n650 S.n649 0.104
R236 S.n250 S.n249 0.093
R237 S.n549 S.n548 0.093
R238 S.n266 S.n265 0.092
R239 S.n290 S.n289 0.092
R240 S S.n651 0.09
R241 S.n436 S.n435 0.087
R242 S.n226 S.n224 0.084
R243 S.n165 S.n162 0.082
R244 S.n486 S.n483 0.082
R245 S.n417 S.n413 0.082
R246 S.n421 S.n420 0.08
R247 S.n65 S.n64 0.076
R248 S.n562 S.n561 0.074
R249 S.n261 S.n260 0.074
R250 S.t32 S.n448 0.068
R251 S.n236 S.n235 0.067
R252 S.n206 S.n204 0.067
R253 S.n10 S.n8 0.067
R254 S.n10 S.n9 0.067
R255 S.n206 S.n205 0.067
R256 S.n165 S.n155 0.067
R257 S.n165 S.n153 0.067
R258 S.n417 S.n407 0.067
R259 S.n417 S.n416 0.067
R260 S.n236 S.n234 0.067
R261 S.n195 S.n194 0.066
R262 S.n166 S.n151 0.065
R263 S.n217 S.n215 0.065
R264 S.n130 S.n129 0.064
R265 S.n5 S.n4 0.063
R266 S.n487 S.n486 0.063
R267 S.n40 S.n27 0.063
R268 S.n143 S.n142 0.063
R269 S.n128 S.n127 0.063
R270 S.n506 S.n505 0.063
R271 S.n237 S.n236 0.062
R272 S.n13 S.n10 0.062
R273 S.n207 S.n206 0.061
R274 S.n226 S.n225 0.06
R275 S.n371 S.n370 0.059
R276 S.n515 S.n514 0.059
R277 S.n418 S.n417 0.058
R278 S.n166 S.n165 0.058
R279 S.n228 S.n214 0.055
R280 S.n640 S.n639 0.055
R281 S.n178 S.n177 0.055
R282 S.n405 S.n242 0.054
R283 S.n68 S.n52 0.054
R284 S.n565 S.n546 0.054
R285 S.n475 S.n474 0.054
R286 S.n206 S.n203 0.054
R287 S.n311 S.n310 0.054
R288 S.n402 S.n401 0.054
R289 S.n600 S.n599 0.054
R290 S.n146 S.n145 0.054
R291 S.n378 S.n377 0.054
R292 S.n583 S.n582 0.054
R293 S.n509 S.n508 0.054
R294 S.n117 S.n116 0.054
R295 S.n184 S.n183 0.054
R296 S.n87 S.n86 0.054
R297 S.n537 S.n536 0.054
R298 S.n43 S.n42 0.054
R299 S.n114 S.n113 0.054
R300 S.n635 S.n634 0.054
R301 S.n610 S.n609 0.054
R302 S.n348 S.n347 0.054
R303 S.n318 S.n317 0.054
R304 S.n284 S.n283 0.054
R305 S.n466 S.n422 0.053
R306 S.t34 S.n247 0.052
R307 S.n63 S.n62 0.052
R308 S.n560 S.n559 0.052
R309 S.n259 S.n258 0.052
R310 S.t34 S.n312 0.051
R311 S.n428 S.n427 0.051
R312 S.n457 S.n456 0.051
R313 S.n459 S.n458 0.051
R314 S.n155 S.n154 0.051
R315 S.n153 S.n152 0.051
R316 S.n531 S.n518 0.05
R317 S.n375 S.n374 0.05
R318 S.n139 S.n138 0.05
R319 S.n305 S.n303 0.047
R320 S.n396 S.n394 0.047
R321 S.n597 S.n595 0.047
R322 S.n647 S.n642 0.047
R323 S.n143 S.n133 0.047
R324 S.n375 S.n358 0.047
R325 S.n580 S.n574 0.047
R326 S.n506 S.n494 0.047
R327 S.n128 S.n51 0.047
R328 S.n195 S.n187 0.047
R329 S.n84 S.n79 0.047
R330 S.n531 S.n529 0.047
R331 S.n40 S.n33 0.047
R332 S.n173 S.n168 0.047
R333 S.n108 S.n104 0.047
R334 S.n629 S.n627 0.047
R335 S.n616 S.n613 0.047
R336 S.n345 S.n338 0.047
R337 S.n325 S.n321 0.047
R338 S.n281 S.n279 0.047
R339 S.n13 S.n12 0.046
R340 S.n209 S.n208 0.046
R341 S.n629 S.n616 0.046
R342 S.n453 S.n452 0.045
R343 S.n426 S.n425 0.045
R344 S.n345 S.n327 0.044
R345 S.n443 S.n441 0.044
R346 S.n518 S.n517 0.043
R347 S.n374 S.n373 0.043
R348 S.n191 S.n190 0.043
R349 S.n7 S.n6 0.043
R350 S.n502 S.n499 0.042
R351 S.n197 S.n196 0.042
R352 S.n252 S.n251 0.042
R353 S.n4 S.n3 0.041
R354 S.n170 S.n169 0.041
R355 S.n63 S.n54 0.04
R356 S.n560 S.n551 0.04
R357 S.n223 S.n222 0.039
R358 S.n430 S.n429 0.039
R359 S.n62 S.n55 0.039
R360 S.n559 S.n552 0.039
R361 S.n61 S.n56 0.038
R362 S.n558 S.n553 0.038
R363 S.n470 S.n467 0.038
R364 S.n549 S.n547 0.038
R365 S.n250 S.n248 0.038
R366 S.n207 S.n198 0.038
R367 S.n331 S.n328 0.037
R368 S.n620 S.n617 0.037
R369 S.n173 S.n170 0.036
R370 S.n387 S.n386 0.035
R371 S.n353 S.n352 0.035
R372 S.n72 S.n71 0.035
R373 S.n569 S.n568 0.035
R374 S.n22 S.n20 0.035
R375 S.t32 S.n463 0.035
R376 S.t47 S.n232 0.035
R377 S.t47 S.n210 0.035
R378 S.t47 S.n14 0.035
R379 S.t32 S.n445 0.035
R380 S.t32 S.n437 0.035
R381 S.n447 S.n446 0.035
R382 S.n325 S.n322 0.034
R383 S.n345 S.n340 0.034
R384 S.t32 S.n462 0.034
R385 S.t47 S.n233 0.034
R386 S.t47 S.n213 0.034
R387 S.t47 S.n17 0.034
R388 S.t32 S.n444 0.034
R389 S.t32 S.n440 0.034
R390 S.n227 S.n218 0.033
R391 S.n562 S.n549 0.032
R392 S.n261 S.n250 0.032
R393 S.t17 S.n353 0.031
R394 S.t0 S.n72 0.031
R395 S.t5 S.n569 0.031
R396 S.n240 S.n239 0.031
R397 S.n241 S.n240 0.031
R398 S.n172 S.n171 0.031
R399 S.n651 S.n650 0.031
R400 S.n650 S.n477 0.031
R401 S.n343 S.n342 0.031
R402 S.n502 S.n501 0.029
R403 S.n368 S.n367 0.028
R404 S.n162 S.n157 0.028
R405 S.n483 S.n479 0.028
R406 S.n413 S.n409 0.028
R407 S.n620 S.n619 0.027
R408 S.n331 S.n330 0.027
R409 S.n327 S.n326 0.027
R410 S.n36 S.n35 0.027
R411 S.n195 S.n192 0.027
R412 S.n647 S.n646 0.027
R413 S.n342 S.n341 0.027
R414 S.n340 S.n339 0.027
R415 S.n531 S.n522 0.026
R416 S.n597 S.n588 0.026
R417 S.n128 S.n125 0.026
R418 S.n506 S.n503 0.026
R419 S.n580 S.n579 0.026
R420 S.n375 S.n369 0.026
R421 S.n272 S.n271 0.026
R422 S.n296 S.n295 0.026
R423 S.n485 S.n484 0.024
R424 S.n415 S.n414 0.024
R425 S.n473 S.n472 0.024
R426 S.n646 S.n645 0.024
R427 S.n644 S.n643 0.023
R428 S.n461 S.n453 0.023
R429 S.n37 S.n36 0.023
R430 S.n192 S.n188 0.023
R431 S.n434 S.n426 0.023
R432 S.n517 S.n516 0.022
R433 S.n373 S.n372 0.022
R434 S.n521 S.n520 0.022
R435 S.n368 S.n363 0.021
R436 S.n138 S.n137 0.021
R437 S.n501 S.n500 0.021
R438 S.n499 S.n498 0.021
R439 S.n367 S.n366 0.021
R440 S.n142 S.n141 0.021
R441 S.n190 S.n189 0.021
R442 S.n433 S.n430 0.02
R443 S.n460 S.n454 0.02
R444 S.n3 S.n2 0.02
R445 S.n386 S.n385 0.02
R446 S.n518 S.n515 0.02
R447 S.n374 S.n371 0.02
R448 S.n162 S.n161 0.02
R449 S.n483 S.n482 0.02
R450 S.n413 S.n412 0.02
R451 S.n12 S.n11 0.02
R452 S.n195 S.n22 0.019
R453 S.n541 S.n540 0.019
R454 S S.n241 0.018
R455 S.n97 S.n96 0.018
R456 S.n94 S.n93 0.017
R457 S.n217 S.n216 0.017
R458 S.n269 S.n268 0.017
R459 S.n293 S.n292 0.017
R460 S.n619 S.n618 0.015
R461 S.n330 S.n329 0.015
R462 S.n363 S.n362 0.015
R463 S.n520 S.n519 0.015
R464 S.n39 S.n38 0.015
R465 S.n96 S.n95 0.015
R466 S.n539 S.n538 0.015
R467 S.t32 S.n447 0.015
R468 S.n649 S.n648 0.014
R469 S.n489 S.n488 0.014
R470 S.n629 S.n620 0.014
R471 S.n345 S.n331 0.014
R472 S.n429 S.n428 0.012
R473 S.n458 S.n457 0.012
R474 S.n143 S.n140 0.012
R475 S.n305 S.n296 0.011
R476 S.n281 S.n272 0.011
R477 S.n108 S.n94 0.01
R478 S.n84 S.n76 0.01
R479 S.n227 S.n217 0.01
R480 S.n108 S.n105 0.01
R481 S.n281 S.n269 0.01
R482 S.n305 S.n293 0.01
R483 S.n647 S.n644 0.01
R484 S.n20 S.n18 0.01
R485 S.n20 S.n19 0.01
R486 S.n419 S.n406 0.009
R487 S.n647 S.n487 0.009
R488 S.n268 S.n267 0.008
R489 S.n292 S.n291 0.008
R490 S.n433 S.n432 0.008
R491 S.n460 S.n459 0.008
R492 S.n84 S.n75 0.008
R493 S.n27 S.n26 0.008
R494 S.n38 S.n34 0.008
R495 S.n38 S.n37 0.008
R496 S.n108 S.n107 0.008
R497 S.n173 S.n172 0.008
R498 S.n384 S.n383 0.008
R499 S.n127 S.n126 0.008
R500 S.n505 S.n504 0.008
R501 S.n365 S.n364 0.008
R502 S.n194 S.n193 0.008
R503 S.n648 S.n647 0.007
R504 S.n93 S.n92 0.007
R505 S.n385 S.n384 0.006
R506 S.n366 S.n365 0.006
R507 S.n434 S.n433 0.006
R508 S.n461 S.n460 0.006
R509 S.n432 S.n431 0.005
R510 S.n459 S.n455 0.005
R511 S.n227 S.n226 0.005
R512 S.t47 S.n207 0.005
R513 S.n303 S.n302 0.004
R514 S.n394 S.n393 0.004
R515 S.n595 S.n594 0.004
R516 S.n642 S.n641 0.004
R517 S.n133 S.n132 0.004
R518 S.n358 S.n357 0.004
R519 S.n574 S.n573 0.004
R520 S.n494 S.n493 0.004
R521 S.n51 S.n50 0.004
R522 S.n187 S.n186 0.004
R523 S.n79 S.n78 0.004
R524 S.n529 S.n528 0.004
R525 S.n33 S.n32 0.004
R526 S.n168 S.n167 0.004
R527 S.n104 S.n103 0.004
R528 S.n627 S.n626 0.004
R529 S.n613 S.n612 0.004
R530 S.n338 S.n337 0.004
R531 S.n321 S.n320 0.004
R532 S.n279 S.n278 0.004
R533 S.n143 S.n130 0.004
R534 S.t47 S.n13 0.004
R535 S.n67 S.n66 0.004
R536 S.n84 S.n83 0.004
R537 S.n564 S.n562 0.004
R538 S.t34 S.n261 0.004
R539 S.n22 S.n21 0.004
R540 S.n541 S.n539 0.004
R541 S.t47 S.n229 0.004
R542 S.t47 S.n231 0.004
R543 S.t47 S.n212 0.004
R544 S.t0 S.n70 0.004
R545 S.t5 S.n567 0.004
R546 S.t47 S.n16 0.004
R547 S.t32 S.n465 0.004
R548 S.t32 S.n450 0.004
R549 S.t32 S.n439 0.004
R550 S.t47 S.n0 0.004
R551 S.t32 S.n443 0.004
R552 S.t17 S.n404 0.004
R553 S.t47 S.n237 0.004
R554 S.n564 S.n563 0.004
R555 S.n308 S.n307 0.003
R556 S.n399 S.n398 0.003
R557 S.n603 S.n602 0.003
R558 S.n638 S.n637 0.003
R559 S.n149 S.n148 0.003
R560 S.n381 S.n380 0.003
R561 S.n586 S.n585 0.003
R562 S.n512 S.n511 0.003
R563 S.n120 S.n119 0.003
R564 S.n181 S.n180 0.003
R565 S.n90 S.n89 0.003
R566 S.n534 S.n533 0.003
R567 S.n46 S.n45 0.003
R568 S.n176 S.n175 0.003
R569 S.n111 S.n110 0.003
R570 S.n632 S.n631 0.003
R571 S.n607 S.n606 0.003
R572 S.n351 S.n350 0.003
R573 S.n315 S.n314 0.003
R574 S.n287 S.n286 0.003
R575 S.n305 S.n300 0.003
R576 S.n396 S.n391 0.003
R577 S.n597 S.n592 0.003
R578 S.n143 S.n136 0.003
R579 S.n375 S.n361 0.003
R580 S.n580 S.n577 0.003
R581 S.n506 S.n497 0.003
R582 S.n128 S.n123 0.003
R583 S.n195 S.n25 0.003
R584 S.n84 S.n82 0.003
R585 S.n531 S.n526 0.003
R586 S.n40 S.n30 0.003
R587 S.n108 S.n101 0.003
R588 S.n629 S.n624 0.003
R589 S.n616 S.n545 0.003
R590 S.n345 S.n335 0.003
R591 S.n325 S.n246 0.003
R592 S.n281 S.n276 0.003
R593 S.n173 S.n166 0.003
R594 S.n476 S.n475 0.003
R595 S.n476 S.n421 0.003
R596 S.n67 S.n65 0.003
R597 S.n616 S.n541 0.003
R598 S.n419 S.n418 0.003
R599 S.t34 S.n264 0.003
R600 S.t32 S.n423 0.003
R601 S.t34 S.n262 0.003
R602 S.t32 S.n451 0.003
R603 S.n522 S.n521 0.003
R604 S.n396 S.n387 0.003
R605 S.t32 S.n436 0.003
R606 S.n140 S.n139 0.003
R607 S.n84 S.n73 0.002
R608 S.n325 S.n243 0.002
R609 S.n345 S.n332 0.002
R610 S.n616 S.n542 0.002
R611 S.n629 S.n621 0.002
R612 S.n597 S.n589 0.002
R613 S.n396 S.n388 0.002
R614 S.n305 S.n297 0.002
R615 S.n196 S.n195 0.002
R616 S.n531 S.n523 0.002
R617 S.n267 S.n266 0.002
R618 S.n291 S.n290 0.002
R619 S.t47 S.n209 0.002
R620 S.t47 S.n5 0.002
R621 S.n629 S.n628 0.002
R622 S.n369 S.n368 0.002
R623 S.n597 S.n596 0.002
R624 S.n396 S.n395 0.002
R625 S.n305 S.n304 0.002
R626 S.n580 S.n571 0.002
R627 S.n506 S.n491 0.002
R628 S.n129 S.n128 0.002
R629 S.n281 S.n280 0.002
R630 S.n40 S.n39 0.002
R631 S.n108 S.n97 0.002
R632 S.n647 S.n489 0.002
R633 S.n202 S.n200 0.002
R634 S.t32 S.n434 0.002
R635 S.t32 S.n461 0.002
R636 S.n375 S.n355 0.002
R637 S.n531 S.n530 0.002
R638 S.n327 S.n325 0.002
R639 S.n375 S.n354 0.002
R640 S.n580 S.n570 0.002
R641 S.n506 S.n490 0.002
R642 S.n128 S.n48 0.002
R643 S.n143 S.n47 0.002
R644 S.n281 S.n273 0.002
R645 S.n476 S.n466 0.002
R646 S.n4 S.n1 0.002
R647 S.n469 S.n468 0.001
R648 S.n228 S.n227 0.001
R649 S.t47 S.n228 0.001
R650 S.n466 S.t32 0.001
R651 S.n125 S.n124 0.001
R652 S.n503 S.n502 0.001
R653 S.n579 S.n578 0.001
R654 S.n108 S.n98 0.001
R655 S.t47 S.n197 0.001
R656 S.t47 S.n7 0.001
R657 S.n202 S.n201 0.001
R658 S.n238 S.t47 0.001
R659 S.n62 S.n61 0.001
R660 S.n559 S.n558 0.001
R661 S.n471 S.n470 0.001
R662 S.n68 S.n67 0.001
R663 S.n565 S.n564 0.001
R664 S.n419 S.n405 0.001
R665 S.n202 S.n199 0.001
R666 S.n325 S.n324 0.001
R667 S.n345 S.n344 0.001
R668 S.n616 S.n615 0.001
R669 S.n271 S.n270 0.001
R670 S.n295 S.n294 0.001
R671 S.n60 S.n59 0.001
R672 S.n557 S.n556 0.001
R673 S.n256 S.n255 0.001
R674 S.n405 S.t17 0.001
R675 S.t0 S.n68 0.001
R676 S.t5 S.n565 0.001
R677 S.n470 S.n469 0.001
R678 S.n61 S.n60 0.001
R679 S.n558 S.n557 0.001
R680 S.n258 S.n252 0.001
R681 S.n588 S.n587 0.001
R682 S.n161 S.n160 0.001
R683 S.n482 S.n481 0.001
R684 S.n412 S.n411 0.001
R685 S.n192 S.n191 0.001
R686 S.n203 S.n202 0.001
R687 S.n300 S.n299 0.001
R688 S.n391 S.n390 0.001
R689 S.n592 S.n591 0.001
R690 S.n136 S.n135 0.001
R691 S.n361 S.n360 0.001
R692 S.n577 S.n576 0.001
R693 S.n497 S.n496 0.001
R694 S.n123 S.n122 0.001
R695 S.n25 S.n24 0.001
R696 S.n82 S.n81 0.001
R697 S.n526 S.n525 0.001
R698 S.n30 S.n29 0.001
R699 S.n101 S.n100 0.001
R700 S.n624 S.n623 0.001
R701 S.n545 S.n544 0.001
R702 S.n335 S.n334 0.001
R703 S.n246 S.n245 0.001
R704 S.n276 S.n275 0.001
R705 S.n260 S.n259 0.001
R706 S.n561 S.n560 0.001
R707 S.n64 S.n63 0.001
R708 S.t34 S.n308 0.001
R709 S.t34 S.n311 0.001
R710 S.t17 S.n399 0.001
R711 S.t17 S.n402 0.001
R712 S.t5 S.n603 0.001
R713 S.t5 S.n600 0.001
R714 S.n600 S.n597 0.001
R715 S.n638 S.t42 0.001
R716 S.n647 S.n640 0.001
R717 S.t40 S.n149 0.001
R718 S.t40 S.n146 0.001
R719 S.n146 S.n143 0.001
R720 S.t17 S.n381 0.001
R721 S.t17 S.n378 0.001
R722 S.n378 S.n375 0.001
R723 S.t5 S.n586 0.001
R724 S.t5 S.n583 0.001
R725 S.n583 S.n580 0.001
R726 S.t42 S.n512 0.001
R727 S.t42 S.n509 0.001
R728 S.n509 S.n506 0.001
R729 S.n117 S.t0 0.001
R730 S.n128 S.n117 0.001
R731 S.n181 S.t40 0.001
R732 S.n195 S.n184 0.001
R733 S.t0 S.n90 0.001
R734 S.t0 S.n87 0.001
R735 S.n87 S.n84 0.001
R736 S.t42 S.n534 0.001
R737 S.t42 S.n537 0.001
R738 S.t40 S.n46 0.001
R739 S.t40 S.n43 0.001
R740 S.n43 S.n40 0.001
R741 S.t40 S.n176 0.001
R742 S.t40 S.n178 0.001
R743 S.t0 S.n111 0.001
R744 S.t0 S.n114 0.001
R745 S.t42 S.n632 0.001
R746 S.t42 S.n635 0.001
R747 S.n607 S.t5 0.001
R748 S.n616 S.n610 0.001
R749 S.t17 S.n351 0.001
R750 S.t17 S.n348 0.001
R751 S.n348 S.n345 0.001
R752 S.n315 S.t34 0.001
R753 S.n325 S.n318 0.001
R754 S.n324 S.n323 0.001
R755 S.n344 S.n343 0.001
R756 S.n615 S.n614 0.001
R757 S.n220 S.n219 0.001
R758 S.n224 S.n223 0.001
R759 S.n417 S.n415 0.001
R760 S.n486 S.n485 0.001
R761 S.n165 S.n164 0.001
R762 S.n474 S.n473 0.001
R763 S.n257 S.n256 0.001
R764 S.n308 S.n305 0.001
R765 S.n399 S.n396 0.001
R766 S.n647 S.n638 0.001
R767 S.n128 S.n120 0.001
R768 S.n534 S.n531 0.001
R769 S.n195 S.n181 0.001
R770 S.n176 S.n173 0.001
R771 S.n325 S.n315 0.001
R772 S.n616 S.n607 0.001
R773 S.n632 S.n629 0.001
R774 S.n111 S.n108 0.001
R775 S.n258 S.n257 0.001
R776 S.t34 S.n287 0.001
R777 S.t34 S.n284 0.001
R778 S.n284 S.n281 0.001
C0 DNW D 142.40fF
C1 G S 735.54fF
C2 D S 181.34fF
C3 DNW S 544.96fF
C4 G D 212.13fF
C5 G DNW 3.95fF
C6 D SUB 14.16fF
C7 G SUB -88.18fF
C8 S SUB -276.62fF
C9 DNW SUB 2658.03fF $ **FLOATING
C10 S.n0 SUB 2.07fF
C11 S.t8 SUB 8.16fF
C12 S.n1 SUB 0.56fF
C13 S.n2 SUB 1.00fF
C14 S.n3 SUB 0.27fF
C15 S.n4 SUB 2.21fF
C16 S.n5 SUB 1.93fF
C17 S.n6 SUB 1.91fF
C18 S.n7 SUB 3.35fF
C19 S.n8 SUB 11.43fF
C20 S.n9 SUB 11.43fF
C21 S.n10 SUB 7.09fF
C22 S.n11 SUB 0.18fF
C23 S.n12 SUB 2.22fF
C24 S.n13 SUB 2.06fF
C25 S.t48 SUB 0.03fF
C26 S.n14 SUB 1.14fF
C27 S.n15 SUB 0.02fF
C28 S.t93 SUB 0.03fF
C29 S.n16 SUB 0.47fF
C30 S.t125 SUB 0.03fF
C31 S.n17 SUB 1.13fF
C32 S.n18 SUB 0.21fF
C33 S.n19 SUB 1.98fF
C34 S.n20 SUB 0.10fF
C35 S.n21 SUB 0.96fF
C36 S.n22 SUB 0.03fF
C37 S.n23 SUB 0.15fF
C38 S.t41 SUB 0.03fF
C39 S.n24 SUB 0.18fF
C40 S.n26 SUB 0.32fF
C41 S.n27 SUB 0.11fF
C42 S.n28 SUB 0.15fF
C43 S.t116 SUB 0.03fF
C44 S.n29 SUB 0.18fF
C45 S.t27 SUB 0.03fF
C46 S.n31 SUB 0.31fF
C47 S.n32 SUB 0.45fF
C48 S.n33 SUB 0.77fF
C49 S.n34 SUB 0.81fF
C50 S.n35 SUB 0.47fF
C51 S.n36 SUB 0.32fF
C52 S.n37 SUB 0.28fF
C53 S.n38 SUB 0.77fF
C54 S.n39 SUB 0.35fF
C55 S.n40 SUB 2.47fF
C56 S.t101 SUB 0.03fF
C57 S.n41 SUB 0.30fF
C58 S.n42 SUB 1.16fF
C59 S.n43 SUB 0.06fF
C60 S.t119 SUB 0.03fF
C61 S.n44 SUB 0.15fF
C62 S.n45 SUB 0.18fF
C63 S.n47 SUB 2.35fF
C64 S.n48 SUB 2.40fF
C65 S.t58 SUB 0.03fF
C66 S.n49 SUB 0.31fF
C67 S.n50 SUB 0.45fF
C68 S.n51 SUB 0.77fF
C69 S.t14 SUB 0.03fF
C70 S.n52 SUB 1.55fF
C71 S.n53 SUB 0.45fF
C72 S.n54 SUB 0.80fF
C73 S.n55 SUB 1.47fF
C74 S.n56 SUB 1.39fF
C75 S.n57 SUB 0.75fF
C76 S.n58 SUB 0.02fF
C77 S.n59 SUB 1.23fF
C78 S.t13 SUB 7.26fF
C79 S.n60 SUB 8.79fF
C80 S.n62 SUB 0.48fF
C81 S.n63 SUB 0.30fF
C82 S.n64 SUB 3.71fF
C83 S.n65 SUB 2.39fF
C84 S.n66 SUB 2.92fF
C85 S.n67 SUB 5.58fF
C86 S.n68 SUB 0.32fF
C87 S.n69 SUB 0.02fF
C88 S.t57 SUB 0.03fF
C89 S.n70 SUB 0.32fF
C90 S.t99 SUB 0.03fF
C91 S.n71 SUB 1.22fF
C92 S.n72 SUB 0.90fF
C93 S.n73 SUB 2.39fF
C94 S.n74 SUB 0.91fF
C95 S.n75 SUB 0.45fF
C96 S.n76 SUB 1.58fF
C97 S.t94 SUB 0.03fF
C98 S.n77 SUB 0.31fF
C99 S.n78 SUB 0.45fF
C100 S.n79 SUB 0.77fF
C101 S.n80 SUB 0.15fF
C102 S.t1 SUB 0.03fF
C103 S.n81 SUB 0.18fF
C104 S.n83 SUB 2.88fF
C105 S.n84 SUB 2.58fF
C106 S.t65 SUB 0.03fF
C107 S.n85 SUB 0.30fF
C108 S.n86 SUB 1.16fF
C109 S.n87 SUB 0.06fF
C110 S.t52 SUB 0.03fF
C111 S.n88 SUB 0.15fF
C112 S.n89 SUB 0.18fF
C113 S.n91 SUB 7.06fF
C114 S.n92 SUB 0.04fF
C115 S.n93 SUB 0.18fF
C116 S.n94 SUB 0.74fF
C117 S.n95 SUB 0.15fF
C118 S.n96 SUB 0.68fF
C119 S.n97 SUB 0.52fF
C120 S.n98 SUB 2.49fF
C121 S.n99 SUB 0.15fF
C122 S.t4 SUB 0.03fF
C123 S.n100 SUB 0.18fF
C124 S.t73 SUB 0.03fF
C125 S.n102 SUB 0.31fF
C126 S.n103 SUB 0.45fF
C127 S.n104 SUB 0.77fF
C128 S.n105 SUB 1.99fF
C129 S.n106 SUB 0.90fF
C130 S.n107 SUB 0.36fF
C131 S.n108 SUB 2.51fF
C132 S.t50 SUB 0.03fF
C133 S.n109 SUB 0.15fF
C134 S.n110 SUB 0.18fF
C135 S.t111 SUB 0.03fF
C136 S.n112 SUB 0.30fF
C137 S.n113 SUB 1.16fF
C138 S.n114 SUB 0.06fF
C139 S.t0 SUB 15.18fF
C140 S.t16 SUB 0.03fF
C141 S.n115 SUB 0.30fF
C142 S.n116 SUB 1.16fF
C143 S.n117 SUB 0.06fF
C144 S.t121 SUB 0.03fF
C145 S.n118 SUB 0.15fF
C146 S.n119 SUB 0.18fF
C147 S.n121 SUB 0.15fF
C148 S.t90 SUB 0.03fF
C149 S.n122 SUB 0.18fF
C150 S.n124 SUB 1.47fF
C151 S.n125 SUB 0.28fF
C152 S.n126 SUB 0.32fF
C153 S.n127 SUB 0.11fF
C154 S.n128 SUB 2.40fF
C155 S.n129 SUB 3.50fF
C156 S.n130 SUB 3.17fF
C157 S.t55 SUB 0.03fF
C158 S.n131 SUB 0.31fF
C159 S.n132 SUB 0.45fF
C160 S.n133 SUB 0.77fF
C161 S.n134 SUB 0.15fF
C162 S.t107 SUB 0.03fF
C163 S.n135 SUB 0.18fF
C164 S.n137 SUB 0.87fF
C165 S.n138 SUB 0.35fF
C166 S.n139 SUB 2.21fF
C167 S.n140 SUB 0.27fF
C168 S.n141 SUB 0.24fF
C169 S.n142 SUB 0.12fF
C170 S.n143 SUB 2.37fF
C171 S.t21 SUB 0.03fF
C172 S.n144 SUB 0.30fF
C173 S.n145 SUB 1.16fF
C174 S.n146 SUB 0.06fF
C175 S.t83 SUB 0.03fF
C176 S.n147 SUB 0.15fF
C177 S.n148 SUB 0.18fF
C178 S.n150 SUB 7.06fF
C179 S.n151 SUB 1.45fF
C180 S.n152 SUB 11.43fF
C181 S.n153 SUB 25.94fF
C182 S.n154 SUB 11.43fF
C183 S.n155 SUB 25.94fF
C184 S.n156 SUB 0.76fF
C185 S.n157 SUB 0.28fF
C186 S.n158 SUB 1.12fF
C187 S.n159 SUB 1.12fF
C188 S.n160 SUB 1.90fF
C189 S.n161 SUB 0.37fF
C190 S.t15 SUB 7.26fF
C191 S.n162 SUB 10.59fF
C192 S.n163 SUB 0.27fF
C193 S.n164 SUB 1.80fF
C194 S.n165 SUB 5.41fF
C195 S.n166 SUB 2.29fF
C196 S.t31 SUB 0.03fF
C197 S.n167 SUB 0.81fF
C198 S.n168 SUB 0.77fF
C199 S.n169 SUB 1.54fF
C200 S.n170 SUB 0.47fF
C201 S.n171 SUB 1.44fF
C202 S.n172 SUB 0.49fF
C203 S.n173 SUB 5.39fF
C204 S.t74 SUB 0.03fF
C205 S.n174 SUB 0.02fF
C206 S.n175 SUB 0.33fF
C207 S.t105 SUB 0.03fF
C208 S.n177 SUB 1.52fF
C209 S.n178 SUB 0.06fF
C210 S.t40 SUB 14.69fF
C211 S.t51 SUB 0.03fF
C212 S.n179 SUB 0.15fF
C213 S.n180 SUB 0.18fF
C214 S.t23 SUB 0.03fF
C215 S.n182 SUB 0.30fF
C216 S.n183 SUB 1.16fF
C217 S.n184 SUB 0.06fF
C218 S.t72 SUB 0.03fF
C219 S.n185 SUB 0.31fF
C220 S.n186 SUB 0.45fF
C221 S.n187 SUB 0.77fF
C222 S.n188 SUB 0.80fF
C223 S.n189 SUB 1.00fF
C224 S.n190 SUB 0.25fF
C225 S.n191 SUB 0.39fF
C226 S.n192 SUB 0.33fF
C227 S.n193 SUB 0.32fF
C228 S.n194 SUB 0.11fF
C229 S.n195 SUB 2.27fF
C230 S.n196 SUB 2.55fF
C231 S.n197 SUB 3.35fF
C232 S.n198 SUB 1.83fF
C233 S.n199 SUB 5.45fF
C234 S.n200 SUB 5.98fF
C235 S.n201 SUB 2.79fF
C236 S.n202 SUB 37.12fF
C237 S.n203 SUB 5.42fF
C238 S.n204 SUB 17.33fF
C239 S.n205 SUB 17.33fF
C240 S.n206 SUB 7.21fF
C241 S.n207 SUB 2.02fF
C242 S.n208 SUB 1.01fF
C243 S.n209 SUB 2.36fF
C244 S.t87 SUB 0.03fF
C245 S.n210 SUB 1.14fF
C246 S.n211 SUB 0.02fF
C247 S.t9 SUB 0.03fF
C248 S.n212 SUB 0.47fF
C249 S.t56 SUB 0.03fF
C250 S.n213 SUB 1.13fF
C251 S.t62 SUB 0.03fF
C252 S.n214 SUB 1.66fF
C253 S.n215 SUB 1.14fF
C254 S.n216 SUB 1.74fF
C255 S.n217 SUB 0.83fF
C256 S.n218 SUB 0.20fF
C257 S.n219 SUB 24.77fF
C258 S.n220 SUB 2.83fF
C259 S.n221 SUB 0.45fF
C260 S.n222 SUB 0.80fF
C261 S.n223 SUB 0.67fF
C262 S.n224 SUB 3.83fF
C263 S.n225 SUB 15.84fF
C264 S.n226 SUB 2.66fF
C265 S.n227 SUB 9.20fF
C266 S.n228 SUB 0.32fF
C267 S.t92 SUB 0.03fF
C268 S.n229 SUB 0.56fF
C269 S.n230 SUB 0.02fF
C270 S.t12 SUB 0.03fF
C271 S.n231 SUB 0.47fF
C272 S.t109 SUB 0.03fF
C273 S.n232 SUB 1.14fF
C274 S.t76 SUB 0.03fF
C275 S.n233 SUB 1.13fF
C276 S.n234 SUB 26.49fF
C277 S.n235 SUB 26.49fF
C278 S.n236 SUB 7.37fF
C279 S.n237 SUB 2.50fF
C280 S.t47 SUB 36.17fF
C281 S.n238 SUB 4.16fF
C282 S.n239 SUB 20.98fF
C283 S.n240 SUB 12.02fF
C284 S.n241 SUB 9.85fF
C285 S.t26 SUB 0.03fF
C286 S.n242 SUB 1.55fF
C287 S.n243 SUB 2.48fF
C288 S.n244 SUB 0.15fF
C289 S.t46 SUB 0.03fF
C290 S.n245 SUB 0.18fF
C291 S.t97 SUB 0.03fF
C292 S.n247 SUB 1.53fF
C293 S.n248 SUB 0.08fF
C294 S.n249 SUB 0.12fF
C295 S.n250 SUB 0.77fF
C296 S.n251 SUB 1.39fF
C297 S.n252 SUB 1.18fF
C298 S.n253 SUB 1.07fF
C299 S.n254 SUB 0.02fF
C300 S.n255 SUB 1.23fF
C301 S.t29 SUB 7.26fF
C302 S.n256 SUB 8.40fF
C303 S.n258 SUB 1.56fF
C304 S.n259 SUB 1.84fF
C305 S.n260 SUB 3.69fF
C306 S.n261 SUB 3.08fF
C307 S.n262 SUB 2.50fF
C308 S.n263 SUB 0.02fF
C309 S.t89 SUB 0.03fF
C310 S.n264 SUB 0.32fF
C311 S.n265 SUB 0.05fF
C312 S.n266 SUB 0.12fF
C313 S.n267 SUB 0.37fF
C314 S.n268 SUB 0.32fF
C315 S.n269 SUB 0.15fF
C316 S.n270 SUB 0.07fF
C317 S.n271 SUB 0.22fF
C318 S.n272 SUB 1.46fF
C319 S.n273 SUB 2.39fF
C320 S.n274 SUB 0.15fF
C321 S.t113 SUB 0.03fF
C322 S.n275 SUB 0.18fF
C323 S.t45 SUB 0.03fF
C324 S.n277 SUB 0.31fF
C325 S.n278 SUB 0.45fF
C326 S.n279 SUB 0.77fF
C327 S.n280 SUB 3.25fF
C328 S.n281 SUB 2.47fF
C329 S.t63 SUB 0.03fF
C330 S.n282 SUB 0.30fF
C331 S.n283 SUB 1.16fF
C332 S.n284 SUB 0.06fF
C333 S.t35 SUB 0.03fF
C334 S.n285 SUB 0.15fF
C335 S.n286 SUB 0.18fF
C336 S.n288 SUB 7.06fF
C337 S.n289 SUB 0.05fF
C338 S.n290 SUB 0.12fF
C339 S.n291 SUB 0.37fF
C340 S.n292 SUB 0.32fF
C341 S.n293 SUB 0.15fF
C342 S.n294 SUB 0.07fF
C343 S.n295 SUB 0.22fF
C344 S.n296 SUB 1.60fF
C345 S.n297 SUB 3.53fF
C346 S.n298 SUB 0.15fF
C347 S.t120 SUB 0.03fF
C348 S.n299 SUB 0.18fF
C349 S.t49 SUB 0.03fF
C350 S.n301 SUB 0.31fF
C351 S.n302 SUB 0.45fF
C352 S.n303 SUB 0.77fF
C353 S.n304 SUB 3.32fF
C354 S.n305 SUB 2.61fF
C355 S.t38 SUB 0.03fF
C356 S.n306 SUB 0.15fF
C357 S.n307 SUB 0.18fF
C358 S.t11 SUB 0.03fF
C359 S.n309 SUB 0.30fF
C360 S.n310 SUB 1.16fF
C361 S.n311 SUB 0.06fF
C362 S.t126 SUB 0.03fF
C363 S.n312 SUB 1.52fF
C364 S.t34 SUB 21.04fF
C365 S.t82 SUB 0.03fF
C366 S.n313 SUB 0.15fF
C367 S.n314 SUB 0.18fF
C368 S.t61 SUB 0.03fF
C369 S.n316 SUB 0.30fF
C370 S.n317 SUB 1.16fF
C371 S.n318 SUB 0.06fF
C372 S.t88 SUB 0.03fF
C373 S.n319 SUB 0.31fF
C374 S.n320 SUB 0.45fF
C375 S.n321 SUB 0.77fF
C376 S.n322 SUB 0.38fF
C377 S.n323 SUB 1.39fF
C378 S.n324 SUB 0.20fF
C379 S.n325 SUB 2.68fF
C380 S.n326 SUB 2.70fF
C381 S.n327 SUB 2.27fF
C382 S.n328 SUB 0.59fF
C383 S.n329 SUB 0.13fF
C384 S.n330 SUB 0.45fF
C385 S.n331 SUB 1.45fF
C386 S.n332 SUB 2.39fF
C387 S.n333 SUB 0.15fF
C388 S.t112 SUB 0.03fF
C389 S.n334 SUB 0.18fF
C390 S.t24 SUB 0.03fF
C391 S.n336 SUB 0.31fF
C392 S.n337 SUB 0.45fF
C393 S.n338 SUB 0.77fF
C394 S.n339 SUB 1.18fF
C395 S.n340 SUB 0.41fF
C396 S.n341 SUB 0.41fF
C397 S.n342 SUB 1.18fF
C398 S.n343 SUB 1.39fF
C399 S.n344 SUB 0.20fF
C400 S.n345 SUB 4.71fF
C401 S.t22 SUB 0.03fF
C402 S.n346 SUB 0.30fF
C403 S.n347 SUB 1.16fF
C404 S.n348 SUB 0.06fF
C405 S.t114 SUB 0.03fF
C406 S.n349 SUB 0.15fF
C407 S.n350 SUB 0.18fF
C408 S.t25 SUB 0.03fF
C409 S.n352 SUB 1.22fF
C410 S.n353 SUB 0.90fF
C411 S.n354 SUB 2.21fF
C412 S.n355 SUB 3.88fF
C413 S.t69 SUB 0.03fF
C414 S.n356 SUB 0.31fF
C415 S.n357 SUB 0.45fF
C416 S.n358 SUB 0.77fF
C417 S.n359 SUB 0.15fF
C418 S.t37 SUB 0.03fF
C419 S.n360 SUB 0.18fF
C420 S.n362 SUB 0.23fF
C421 S.n363 SUB 0.26fF
C422 S.n364 SUB 0.32fF
C423 S.n365 SUB 0.11fF
C424 S.n366 SUB 0.29fF
C425 S.n367 SUB 0.84fF
C426 S.n368 SUB 1.15fF
C427 S.n369 SUB 0.29fF
C428 S.n370 SUB 0.12fF
C429 S.n371 SUB 0.26fF
C430 S.n372 SUB 0.09fF
C431 S.n373 SUB 0.07fF
C432 S.n374 SUB 0.09fF
C433 S.n375 SUB 2.53fF
C434 S.t68 SUB 0.03fF
C435 S.n376 SUB 0.30fF
C436 S.n377 SUB 1.16fF
C437 S.n378 SUB 0.06fF
C438 S.t39 SUB 0.03fF
C439 S.n379 SUB 0.15fF
C440 S.n380 SUB 0.18fF
C441 S.n382 SUB 7.06fF
C442 S.n383 SUB 0.32fF
C443 S.n384 SUB 0.11fF
C444 S.n385 SUB 0.26fF
C445 S.n386 SUB 0.99fF
C446 S.n387 SUB 2.46fF
C447 S.n388 SUB 2.39fF
C448 S.n389 SUB 0.15fF
C449 S.t18 SUB 0.03fF
C450 S.n390 SUB 0.18fF
C451 S.t79 SUB 0.03fF
C452 S.n392 SUB 0.31fF
C453 S.n393 SUB 0.45fF
C454 S.n394 SUB 0.77fF
C455 S.n395 SUB 3.40fF
C456 S.n396 SUB 3.81fF
C457 S.t80 SUB 0.03fF
C458 S.n397 SUB 0.15fF
C459 S.n398 SUB 0.18fF
C460 S.t3 SUB 0.03fF
C461 S.n400 SUB 0.30fF
C462 S.n401 SUB 1.16fF
C463 S.n402 SUB 0.06fF
C464 S.t102 SUB 0.03fF
C465 S.n403 SUB 0.02fF
C466 S.n404 SUB 0.33fF
C467 S.t17 SUB 15.17fF
C468 S.n405 SUB 0.32fF
C469 S.n406 SUB 3.72fF
C470 S.n407 SUB 17.33fF
C471 S.n408 SUB 0.76fF
C472 S.n409 SUB 0.56fF
C473 S.n410 SUB 0.75fF
C474 S.n411 SUB 1.90fF
C475 S.n412 SUB 0.37fF
C476 S.t10 SUB 7.26fF
C477 S.n413 SUB 10.59fF
C478 S.n414 SUB 0.98fF
C479 S.n415 SUB 0.35fF
C480 S.n416 SUB 17.33fF
C481 S.n417 SUB 5.73fF
C482 S.n418 SUB 2.97fF
C483 S.n419 SUB 5.82fF
C484 S.n420 SUB 5.64fF
C485 S.n421 SUB 3.21fF
C486 S.t64 SUB 0.03fF
C487 S.n422 SUB 1.63fF
C488 S.t85 SUB 0.03fF
C489 S.n423 SUB 0.56fF
C490 S.n424 SUB 7.06fF
C491 S.n425 SUB 0.03fF
C492 S.n426 SUB 0.03fF
C493 S.n427 SUB 0.04fF
C494 S.n428 SUB 0.04fF
C495 S.n429 SUB 0.03fF
C496 S.n430 SUB 0.02fF
C497 S.n431 SUB 0.79fF
C498 S.n432 SUB 0.31fF
C499 S.n433 SUB 0.19fF
C500 S.n434 SUB 0.23fF
C501 S.n435 SUB 60.94fF
C502 S.n436 SUB 5.97fF
C503 S.t110 SUB 0.03fF
C504 S.n437 SUB 1.14fF
C505 S.t30 SUB 0.03fF
C506 S.n438 SUB 0.02fF
C507 S.n439 SUB 0.47fF
C508 S.t115 SUB 0.03fF
C509 S.n440 SUB 1.13fF
C510 S.n441 SUB 1.18fF
C511 S.n442 SUB 5.20fF
C512 S.n443 SUB 2.35fF
C513 S.t75 SUB 0.03fF
C514 S.n444 SUB 1.13fF
C515 S.t78 SUB 0.03fF
C516 S.n445 SUB 1.14fF
C517 S.n446 SUB 1.52fF
C518 S.n447 SUB 0.42fF
C519 S.n448 SUB 0.40fF
C520 S.t95 SUB 0.03fF
C521 S.n449 SUB 0.02fF
C522 S.n450 SUB 0.47fF
C523 S.n451 SUB 5.80fF
C524 S.n452 SUB 0.03fF
C525 S.n453 SUB 0.03fF
C526 S.n454 SUB 0.02fF
C527 S.n455 SUB 0.79fF
C528 S.n456 SUB 0.04fF
C529 S.n457 SUB 0.04fF
C530 S.n458 SUB 0.03fF
C531 S.n459 SUB 0.31fF
C532 S.n460 SUB 0.19fF
C533 S.n461 SUB 0.23fF
C534 S.t33 SUB 0.03fF
C535 S.n462 SUB 1.13fF
C536 S.t36 SUB 0.03fF
C537 S.n463 SUB 1.14fF
C538 S.t60 SUB 0.03fF
C539 S.n464 SUB 0.02fF
C540 S.n465 SUB 0.47fF
C541 S.t32 SUB 46.43fF
C542 S.n466 SUB 0.60fF
C543 S.n467 SUB 8.10fF
C544 S.n468 SUB 2.20fF
C545 S.n469 SUB 14.66fF
C546 S.n471 SUB 3.04fF
C547 S.n472 SUB 0.98fF
C548 S.n473 SUB 0.67fF
C549 S.n474 SUB 14.81fF
C550 S.n475 SUB 3.21fF
C551 S.n476 SUB 8.82fF
C552 S.n477 SUB 20.55fF
C553 S.n478 SUB 0.76fF
C554 S.n479 SUB 0.28fF
C555 S.n480 SUB 0.75fF
C556 S.n481 SUB 1.90fF
C557 S.n482 SUB 0.37fF
C558 S.t19 SUB 7.26fF
C559 S.n483 SUB 10.59fF
C560 S.n484 SUB 0.98fF
C561 S.n485 SUB 0.35fF
C562 S.n486 SUB 5.43fF
C563 S.n487 SUB 3.57fF
C564 S.n488 SUB 0.88fF
C565 S.n489 SUB 0.53fF
C566 S.n490 SUB 2.40fF
C567 S.n491 SUB 3.40fF
C568 S.t106 SUB 0.03fF
C569 S.n492 SUB 0.31fF
C570 S.n493 SUB 0.45fF
C571 S.n494 SUB 0.77fF
C572 S.n495 SUB 0.15fF
C573 S.t81 SUB 0.03fF
C574 S.n496 SUB 0.18fF
C575 S.n498 SUB 0.89fF
C576 S.n499 SUB 0.29fF
C577 S.n500 SUB 0.29fF
C578 S.n501 SUB 0.89fF
C579 S.n502 SUB 1.47fF
C580 S.n503 SUB 0.28fF
C581 S.n504 SUB 0.32fF
C582 S.n505 SUB 0.11fF
C583 S.n506 SUB 2.40fF
C584 S.t67 SUB 0.03fF
C585 S.n507 SUB 0.30fF
C586 S.n508 SUB 1.16fF
C587 S.n509 SUB 0.06fF
C588 S.t84 SUB 0.03fF
C589 S.n510 SUB 0.15fF
C590 S.n511 SUB 0.18fF
C591 S.n513 SUB 7.06fF
C592 S.n514 SUB 0.12fF
C593 S.n515 SUB 0.26fF
C594 S.n516 SUB 0.09fF
C595 S.n517 SUB 0.07fF
C596 S.n518 SUB 0.09fF
C597 S.n519 SUB 0.23fF
C598 S.n520 SUB 0.25fF
C599 S.n521 SUB 1.32fF
C600 S.n522 SUB 0.69fF
C601 S.n523 SUB 2.97fF
C602 S.n524 SUB 0.15fF
C603 S.t118 SUB 0.03fF
C604 S.n525 SUB 0.18fF
C605 S.t28 SUB 0.03fF
C606 S.n527 SUB 0.31fF
C607 S.n528 SUB 0.45fF
C608 S.n529 SUB 0.77fF
C609 S.n530 SUB 2.20fF
C610 S.n531 SUB 3.11fF
C611 S.t122 SUB 0.03fF
C612 S.n532 SUB 0.15fF
C613 S.n533 SUB 0.18fF
C614 S.t103 SUB 0.03fF
C615 S.n535 SUB 0.30fF
C616 S.n536 SUB 1.16fF
C617 S.n537 SUB 0.06fF
C618 S.n538 SUB 0.15fF
C619 S.n539 SUB 0.12fF
C620 S.n540 SUB 0.15fF
C621 S.n541 SUB 0.23fF
C622 S.n542 SUB 2.39fF
C623 S.n543 SUB 0.15fF
C624 S.t53 SUB 0.03fF
C625 S.n544 SUB 0.18fF
C626 S.t96 SUB 0.03fF
C627 S.n546 SUB 1.55fF
C628 S.n547 SUB 0.08fF
C629 S.n548 SUB 0.12fF
C630 S.n549 SUB 0.77fF
C631 S.n550 SUB 0.45fF
C632 S.n551 SUB 0.80fF
C633 S.n552 SUB 1.47fF
C634 S.n553 SUB 1.39fF
C635 S.n554 SUB 0.75fF
C636 S.n555 SUB 0.02fF
C637 S.n556 SUB 1.23fF
C638 S.t2 SUB 7.26fF
C639 S.n557 SUB 8.79fF
C640 S.n559 SUB 0.48fF
C641 S.n560 SUB 0.30fF
C642 S.n561 SUB 3.69fF
C643 S.n562 SUB 3.08fF
C644 S.n563 SUB 3.15fF
C645 S.n564 SUB 5.46fF
C646 S.n565 SUB 0.32fF
C647 S.n566 SUB 0.02fF
C648 S.t6 SUB 0.03fF
C649 S.n567 SUB 0.32fF
C650 S.t66 SUB 0.03fF
C651 S.n568 SUB 1.22fF
C652 S.n569 SUB 0.90fF
C653 S.n570 SUB 2.40fF
C654 S.n571 SUB 3.40fF
C655 S.t59 SUB 0.03fF
C656 S.n572 SUB 0.31fF
C657 S.n573 SUB 0.45fF
C658 S.n574 SUB 0.77fF
C659 S.n575 SUB 0.15fF
C660 S.t91 SUB 0.03fF
C661 S.n576 SUB 0.18fF
C662 S.n578 SUB 1.47fF
C663 S.n579 SUB 0.28fF
C664 S.n580 SUB 2.40fF
C665 S.t20 SUB 0.03fF
C666 S.n581 SUB 0.30fF
C667 S.n582 SUB 1.16fF
C668 S.n583 SUB 0.06fF
C669 S.t123 SUB 0.03fF
C670 S.n584 SUB 0.15fF
C671 S.n585 SUB 0.18fF
C672 S.n587 SUB 0.98fF
C673 S.n588 SUB 0.56fF
C674 S.n589 SUB 1.89fF
C675 S.n590 SUB 0.15fF
C676 S.t71 SUB 0.03fF
C677 S.n591 SUB 0.18fF
C678 S.t117 SUB 0.03fF
C679 S.n593 SUB 0.31fF
C680 S.n594 SUB 0.45fF
C681 S.n595 SUB 0.77fF
C682 S.n596 SUB 3.00fF
C683 S.n597 SUB 2.54fF
C684 S.t54 SUB 0.03fF
C685 S.n598 SUB 0.30fF
C686 S.n599 SUB 1.16fF
C687 S.n600 SUB 0.06fF
C688 S.t100 SUB 0.03fF
C689 S.n601 SUB 0.15fF
C690 S.n602 SUB 0.18fF
C691 S.n604 SUB 7.06fF
C692 S.t5 SUB 15.18fF
C693 S.t86 SUB 0.03fF
C694 S.n605 SUB 0.15fF
C695 S.n606 SUB 0.18fF
C696 S.t98 SUB 0.03fF
C697 S.n608 SUB 0.30fF
C698 S.n609 SUB 1.16fF
C699 S.n610 SUB 0.06fF
C700 S.t7 SUB 0.03fF
C701 S.n611 SUB 0.31fF
C702 S.n612 SUB 0.45fF
C703 S.n613 SUB 0.77fF
C704 S.n614 SUB 1.97fF
C705 S.n615 SUB 0.20fF
C706 S.n616 SUB 3.94fF
C707 S.n617 SUB 0.59fF
C708 S.n618 SUB 0.13fF
C709 S.n619 SUB 0.45fF
C710 S.n620 SUB 1.45fF
C711 S.n621 SUB 2.39fF
C712 S.n622 SUB 0.15fF
C713 S.t44 SUB 0.03fF
C714 S.n623 SUB 0.18fF
C715 S.t104 SUB 0.03fF
C716 S.n625 SUB 0.31fF
C717 S.n626 SUB 0.45fF
C718 S.n627 SUB 0.77fF
C719 S.n628 SUB 1.62fF
C720 S.n629 SUB 6.00fF
C721 S.t43 SUB 0.03fF
C722 S.n630 SUB 0.15fF
C723 S.n631 SUB 0.18fF
C724 S.t77 SUB 0.03fF
C725 S.n633 SUB 0.30fF
C726 S.n634 SUB 1.16fF
C727 S.n635 SUB 0.06fF
C728 S.t42 SUB 14.69fF
C729 S.t124 SUB 0.03fF
C730 S.n636 SUB 0.02fF
C731 S.n637 SUB 0.33fF
C732 S.t70 SUB 0.03fF
C733 S.n639 SUB 1.52fF
C734 S.n640 SUB 0.06fF
C735 S.t108 SUB 0.03fF
C736 S.n641 SUB 0.81fF
C737 S.n642 SUB 0.77fF
C738 S.n643 SUB 1.91fF
C739 S.n644 SUB 0.45fF
C740 S.n645 SUB 1.65fF
C741 S.n646 SUB 0.20fF
C742 S.n647 SUB 2.41fF
C743 S.n648 SUB 0.10fF
C744 S.n649 SUB 2.18fF
C745 S.n650 SUB 11.69fF
C746 S.n651 SUB 22.64fF
.ends

