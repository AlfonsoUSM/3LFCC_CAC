magic
tech sky130A
timestamp 1679664366
<< checkpaint >>
rect -630 26170 14730 56430
rect -630 -630 13630 26170
<< metal2 >>
rect 3000 50060 5200 50600
rect 3000 49870 4960 50060
rect 3000 49000 5200 49870
rect 3000 31760 5740 32000
rect 5930 31760 6800 32000
rect 3000 30400 6800 31760
rect 3000 21440 6800 22800
rect 3000 21200 5740 21440
rect 5930 21200 6800 21440
rect 3000 5749 4962 6000
rect 3000 5200 5300 5749
<< metal3 >>
rect 6000 51600 12900 54600
rect 1000 45700 4000 48600
rect 9900 47700 12900 51600
rect 1000 36700 7900 45700
rect 1000 32800 4000 36700
rect 9900 30800 12900 34700
rect 3900 27800 12900 30800
rect 6000 22800 12400 27800
rect 1000 17400 4000 20800
rect 9400 19400 12400 22800
rect 1000 9400 7400 17400
rect 1000 7000 4000 9400
rect 9400 4000 12400 7400
rect 6000 1000 12400 4000
<< metal4 >>
rect 6000 51600 12900 54600
rect 1000 45700 4000 48600
rect 9900 47700 12900 51600
rect 1000 36700 7900 45700
rect 1000 32800 4000 36700
rect 9900 30800 12900 34700
rect 3900 27800 12900 30800
rect 6000 22800 12400 27800
rect 1000 17400 4000 20800
rect 9400 19400 12400 22800
rect 1000 9400 7400 17400
rect 1000 7000 4000 9400
rect 9400 4000 12400 7400
rect 6000 1000 12400 4000
<< metal5 >>
rect 6000 51600 12900 54600
rect 1000 45700 4000 48600
rect 9900 47700 12900 51600
rect 1000 36700 7900 45700
rect 1000 32800 4000 36700
rect 9900 30800 12900 34700
rect 3900 27800 12900 30800
rect 6000 22800 12400 27800
rect 1000 17400 4000 20800
rect 9400 19400 12400 22800
rect 1000 9400 7400 17400
rect 1000 7000 4000 9400
rect 9400 4000 12400 7400
rect 6000 1000 12400 4000
use nmos_waffle_4x4  nmos_waffle_4x4_0
timestamp 1679664275
transform 1 0 5925 0 1 5975
box -5925 -5975 7075 7025
use nmos_waffle_4x4  nmos_waffle_4x4_1
timestamp 1679664275
transform 0 1 5975 -1 0 20475
box -5925 -5975 7075 7025
use pmos_waffle_6x6  pmos_waffle_6x6_0
timestamp 1679664290
transform 0 1 5975 1 0 32725
box -5925 -5975 8175 8125
use pmos_waffle_6x6  pmos_waffle_6x6_1
timestamp 1679664290
transform 1 0 5925 0 -1 49825
box -5925 -5975 8175 8125
<< labels >>
rlabel metal5 6000 52600 7000 53600 7 VP
rlabel metal2 3000 49600 4000 50600 7 s1
rlabel metal5 1000 40700 2000 41700 7 fc1
rlabel metal2 3000 30800 4000 31800 7 s2
rlabel metal5 6000 25800 7000 26800 7 out
rlabel metal2 3000 21800 4000 22800 7 s3
rlabel metal5 1000 12900 2000 13900 7 fc2
rlabel metal2 3000 5500 4000 6000 7 s4
rlabel metal5 6000 2000 7000 3000 7 VN
<< end >>
