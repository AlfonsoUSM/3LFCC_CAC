**.subckt NMOS_RONcalc
XM1 VDS VGS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='mul' m='mul'
VGS VGS GND {VGS}
.save i(vgs)
VSS VSS GND 0
VDS VDS VSS 1
.save i(vss)
**** begin user architecture code


.param VGS = 5
.param mul = 364
.option temp=70
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.control
compose voltage values (2.5) 5
foreach volt $&voltage
alterparam VGS=$volt
reset
save i(VDS)
dc VDS 0 3 0.0001
wrdata input_files/SPICE_files/NMOS/PRELAYOUT/NMOS_R_on_calc_PRELAYOUT.txt i(VDS)
set appendwrite
end

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
.control
quit
.endc