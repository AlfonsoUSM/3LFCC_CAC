* NGSPICE file created from mag_files/POSTLAYOUT/pmos_flat_12x12.ext - technology: sky130A

.subckt pmos_flat_12x12 G S D PW
X0 S.t286 G D S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1 S.t285 G D S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2 S.t284 G D S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3 D G S.t283 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4 D G S.t282 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5 D G S.t281 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6 S.t280 G D S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7 S.t279 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8 D G S.t278 S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9 D G S.t277 S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10 S.t276 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11 S.t275 G D S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12 S.t274 G D S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13 D G S.t273 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14 S.t272 G D S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X15 D G S.t271 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X16 D G S.t270 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X17 D G S.t269 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X18 D G S.t268 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X19 D G S.t267 S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X20 D G S.t266 S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X21 D G S.t265 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X22 D G S.t264 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X23 S.t263 G D S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X24 D G S.t262 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X25 D G S.t261 S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X26 S.t260 G D S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X27 D G S.t259 S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X28 S.t258 G D S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X29 S.t257 G D S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X30 D G S.t256 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X31 D G S.t255 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X32 S.t254 G D S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X33 S.t253 G D S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X34 S.t252 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X35 D G S.t251 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X36 S.t250 G D S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X37 D G S.t249 S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X38 S.t248 G D S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X39 D G S.t247 S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X40 S.t246 G D S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X41 S.t245 G D S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X42 S.t244 G D S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X43 D G S.t243 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X44 D G S.t242 S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X45 S.t241 G D S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X46 D G S.t240 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X47 S.t239 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X48 S.t238 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X49 D G S.t237 S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X50 S.t236 G D S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X51 S.t235 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X52 S.t234 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X53 S.t233 G D S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X54 S.t232 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X55 S.t231 G D S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X56 S.t230 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X57 D G S.t229 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X58 S.t228 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X59 D G S.t227 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X60 D G S.t226 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X61 D G S.t225 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X62 D G S.t224 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X63 D G S.t223 S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X64 D G S.t222 S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X65 S.t221 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X66 D G S.t220 S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X67 D G S.t219 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X68 D G S.t218 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X69 D G S.t217 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X70 D G S.t216 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X71 D G S.t215 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X72 D G S.t214 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X73 S.t213 G D S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X74 S.t212 G D S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X75 D G S.t211 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X76 D G S.t210 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X77 S.t209 G D S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X78 D G S.t208 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X79 D G S.t207 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X80 S.t206 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X81 S.t205 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X82 S.t204 G D S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X83 S.t203 G D S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X84 S.t202 G D S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X85 S.t201 G D S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X86 S.t200 G D S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X87 S.t199 G D S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X88 S.t198 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X89 S.t197 G D S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X90 D G S.t196 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X91 S.t195 G D S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X92 D G S.t194 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X93 S.t193 G D S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X94 S.t192 G D S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X95 D G S.t191 S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X96 D G S.t190 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X97 D G S.t189 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X98 S.t188 G D S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X99 D G S.t187 S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X100 D G S.t186 S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X101 S.t185 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X102 S.t184 G D S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X103 S.t183 G D S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X104 D G S.t182 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X105 D G S.t181 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X106 S.t180 G D S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X107 D G S.t179 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X108 D G S.t178 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X109 D G S.t177 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X110 S.t176 G D S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X111 D G S.t175 S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X112 D G S.t174 S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X113 S.t173 G D S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X114 D G S.t172 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X115 D G S.t171 S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X116 S.t170 G D S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X117 D G S.t169 S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X118 S.t168 G D S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X119 S.t167 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X120 S.t166 G D S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X121 S.t165 G D S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X122 D G S.t164 S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X123 S.t163 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X124 D G S.t162 S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X125 S.t161 G D S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X126 D G S.t160 S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X127 S.t159 G D S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X128 D G S.t158 S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X129 S.t157 G D S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X130 S.t156 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X131 S.t155 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X132 S.t154 G D S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X133 S.t153 G D S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X134 S.t152 G D S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X135 S.t151 G D S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X136 D G S.t150 S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X137 D G S.t149 S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X138 D G S.t148 S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X139 D G S.t147 S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X140 S.t146 G D S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X141 D G S.t145 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X142 S.t144 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X143 D G S.t143 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X144 D G S.t142 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X145 D G S.t141 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X146 D G S.t140 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X147 D G S.t139 S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X148 D G S.t138 S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X149 D G S.t137 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X150 D G S.t136 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X151 D G S.t135 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X152 D G S.t134 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X153 D G S.t133 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X154 D G S.t132 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X155 S.t131 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X156 S.t130 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X157 S.t129 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X158 D G S.t128 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X159 D G S.t127 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X160 D G S.t126 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X161 S.t125 G D S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X162 S.t124 G D S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X163 D G S.t123 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X164 S.t122 G D S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X165 D G S.t121 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X166 D G S.t120 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X167 S.t119 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X168 S.t118 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X169 S.t117 G D S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X170 S.t116 G D S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X171 S.t115 G D S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X172 S.t114 G D S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X173 S.t113 G D S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X174 S.t112 G D S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X175 S.t111 G D S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X176 D G S.t110 S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X177 S.t109 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X178 S.t108 G D S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X179 S.t107 G D S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X180 S.t106 G D S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X181 D G S.t105 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X182 D G S.t104 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X183 D G S.t103 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X184 D G S.t102 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X185 D G S.t101 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X186 S.t100 G D S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X187 S.t99 G D S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X188 S.t98 G D S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X189 D G S.t96 S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X190 D G S.t95 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X191 D G S.t94 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X192 D G S.t93 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X193 D G S.t92 S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X194 D G S.t91 S.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X195 S.t89 G D S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X196 S.t88 G D S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X197 S.t87 G D S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X198 D G S.t86 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X199 S.t85 G D S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X200 S.t84 G D S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X201 D G S.t83 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X202 D G S.t82 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X203 S.t81 G D S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X204 D G S.t80 S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X205 S.t79 G D S.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X206 S.t77 G D S.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X207 D G S.t75 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X208 D G S.t74 S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X209 S.t73 G D S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X210 S.t72 G D S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X211 D G S.t71 S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X212 S.t70 G D S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X213 S.t69 G D S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X214 D G S.t68 S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X215 S.t67 G D S.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X216 D G S.t65 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X217 S.t63 G D S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X218 S.t62 G D S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X219 D G S.t61 S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X220 S.t60 G D S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X221 S.t59 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X222 S.t58 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X223 D G S.t57 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X224 S.t56 G D S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X225 S.t55 G D S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X226 S.t53 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X227 S.t52 G D S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X228 D G S.t51 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X229 D G S.t50 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X230 S.t49 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X231 D G S.t48 S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X232 D G S.t47 S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X233 D G S.t46 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X234 D G S.t45 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X235 D G S.t44 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X236 D G S.t43 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X237 D G S.t42 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X238 S.t41 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X239 D G S.t40 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X240 D G S.t39 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X241 D G S.t38 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X242 D G S.t37 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X243 S.t35 G D S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X244 D G S.t33 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X245 D G S.t32 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X246 D G S.t30 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X247 S.t28 G D S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X248 S.t27 G D S.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X249 D G S.t25 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X250 D G S.t23 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X251 D G S.t22 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X252 D G S.t20 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X253 S.t18 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X254 S.t17 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X255 S.t16 G D S.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X256 S.t14 G D S.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X257 S.t12 G D S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X258 S.t11 G D S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X259 S.t9 G D S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X260 D G S.t7 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X261 S.t5 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X262 S.t3 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X263 S.t1 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
R0 S.n963 S.n962 153.554
R1 S.n523 S.n522 153.554
R2 S.n743 S.n742 153.554
R3 S.n1347 S.n1346 153.554
R4 S.n108 S.n107 153.554
R5 S.n1105 S.n1104 153.118
R6 S.n1458 S.n1457 153.118
R7 S.n259 S.n258 153.118
R8 S.n610 S.n609 153.118
R9 S.n875 S.n874 153.118
R10 S.n344 S.n343 146.135
R11 S.n314 S.n313 146.135
R12 S.n335 S.n334 146.135
R13 S.n317 S.n316 146.135
R14 S.n358 S.n357 146.135
R15 S.n1196 S.n1195 145.699
R16 S.n1162 S.n1161 145.699
R17 S.n1172 S.n1171 145.699
R18 S.n1180 S.n1179 145.699
R19 S.n1150 S.n1149 145.699
R20 S.n242 S.n241 101.08
R21 S.n384 S.n383 101.08
R22 S.n636 S.n635 101.08
R23 S.n1217 S.n1216 101.08
R24 S.n1112 S.n1111 101.08
R25 S.n246 S.n245 98.123
R26 S.n1201 S.n1200 88.439
R27 S.n1110 S.n1109 68.586
R28 S.n1215 S.n1214 68.586
R29 S.n634 S.n633 68.586
R30 S.n382 S.n381 68.586
R31 S.n240 S.n239 68.586
R32 S.n96 S.n95 65.312
R33 S.n511 S.n510 65.312
R34 S.n731 S.n730 65.312
R35 S.n1335 S.n1334 65.312
R36 S.n973 S.n972 65.312
R37 S.t10 S.t13 33.493
R38 S.n244 S.t29 29.23
R39 S.n98 S.t2 29.23
R40 S.n386 S.t36 29.23
R41 S.n513 S.t8 29.23
R42 S.n638 S.t24 29.23
R43 S.n733 S.t15 29.23
R44 S.n1219 S.t31 29.23
R45 S.n1337 S.t0 29.23
R46 S.n1114 S.t6 29.23
R47 S.n975 S.t21 29.23
R48 S.t54 S.n206 28.256
R49 S.t34 S.n169 28.256
R50 S.t19 S.n462 28.256
R51 S.t90 S.n562 28.256
R52 S.t78 S.n700 28.256
R53 S.t4 S.n785 28.256
R54 S.t76 S.n1256 28.256
R55 S.t97 S.n1393 28.256
R56 S.t26 S.n1083 28.256
R57 S.t64 S.n936 28.256
R58 S.t66 S.n1125 28.256
R59 S.n1202 S.n1201 10.138
R60 S.n503 S.t110 6.541
R61 S.n580 S.n579 6.541
R62 S.n1124 S.t174 6.541
R63 S.n1123 S.t128 6.541
R64 S.n1105 S.t220 6.541
R65 S.n1055 S.t45 6.541
R66 S.n1196 S.t120 6.541
R67 S.n1194 S.t68 6.541
R68 S.n947 S.n946 6.541
R69 S.n955 S.t75 6.541
R70 S.n958 S.t7 6.541
R71 S.n950 S.n949 6.541
R72 S.n1091 S.n1090 6.541
R73 S.n1099 S.t164 6.541
R74 S.n1102 S.t283 6.541
R75 S.n1094 S.n1093 6.541
R76 S.n1373 S.n1372 6.541
R77 S.n1391 S.t215 6.541
R78 S.n1388 S.t101 6.541
R79 S.n1376 S.n1375 6.541
R80 S.n1458 S.t267 6.541
R81 S.n1460 S.t147 6.541
R82 S.n341 S.t251 6.541
R83 S.n76 S.n75 6.541
R84 S.n204 S.t256 6.541
R85 S.n201 S.t61 6.541
R86 S.n79 S.n78 6.541
R87 S.n445 S.n444 6.541
R88 S.n460 S.t83 6.541
R89 S.n457 S.t38 6.541
R90 S.n442 S.n441 6.541
R91 S.n960 S.t133 6.541
R92 S.n1063 S.n1062 6.541
R93 S.n1081 S.t261 6.541
R94 S.n1078 S.t51 6.541
R95 S.n1060 S.n1059 6.541
R96 S.n1356 S.n1355 6.541
R97 S.n1367 S.t194 6.541
R98 S.n1364 S.t219 6.541
R99 S.n1353 S.n1352 6.541
R100 S.n1239 S.n1238 6.541
R101 S.n1254 S.t96 6.541
R102 S.n1251 S.t48 6.541
R103 S.n1236 S.n1235 6.541
R104 S.n772 S.n771 6.541
R105 S.n783 S.t190 6.541
R106 S.n780 S.t216 6.541
R107 S.n769 S.n768 6.541
R108 S.n681 S.n680 6.541
R109 S.n698 S.t92 6.541
R110 S.n695 S.t42 6.541
R111 S.n678 S.n677 6.541
R112 S.n551 S.n550 6.541
R113 S.n560 S.t186 6.541
R114 S.n557 S.t214 6.541
R115 S.n548 S.n547 6.541
R116 S.n87 S.n86 6.541
R117 S.n188 S.t178 6.541
R118 S.n191 S.t211 6.541
R119 S.n194 S.n193 6.541
R120 S.n306 S.t189 6.541
R121 S.n17 S.n16 6.541
R122 S.n45 S.t270 6.541
R123 S.n42 S.t47 6.541
R124 S.n20 S.n19 6.541
R125 S.n472 S.n471 6.541
R126 S.n484 S.t105 6.541
R127 S.n487 S.t50 6.541
R128 S.n469 S.n468 6.541
R129 S.n524 S.t224 6.541
R130 S.n114 S.n113 6.541
R131 S.n129 S.t196 6.541
R132 S.n126 S.t218 6.541
R133 S.n117 S.n116 6.541
R134 S.n141 S.n140 6.541
R135 S.n149 S.t102 6.541
R136 S.n146 S.t135 6.541
R137 S.n138 S.n137 6.541
R138 S.n399 S.n398 6.541
R139 S.n417 S.t271 6.541
R140 S.n414 S.t226 6.541
R141 S.n396 S.n395 6.541
R142 S.n702 S.n701 6.541
R143 S.n716 S.t278 6.541
R144 S.n719 S.t229 6.541
R145 S.n705 S.n704 6.541
R146 S.n744 S.t143 6.541
R147 S.n270 S.n269 6.541
R148 S.n267 S.t181 6.541
R149 S.n264 S.t222 6.541
R150 S.n8 S.n7 6.541
R151 S.n159 S.n158 6.541
R152 S.n167 S.t268 6.541
R153 S.n164 S.t30 6.541
R154 S.n156 S.n155 6.541
R155 S.n426 S.n425 6.541
R156 S.n437 S.t182 6.541
R157 S.n434 S.t141 6.541
R158 S.n429 S.n428 6.541
R159 S.n530 S.n529 6.541
R160 S.n543 S.t277 6.541
R161 S.n540 S.t37 6.541
R162 S.n533 S.n532 6.541
R163 S.n652 S.n651 6.541
R164 S.n664 S.t187 6.541
R165 S.n661 S.t145 6.541
R166 S.n655 S.n654 6.541
R167 S.n750 S.n749 6.541
R168 S.n764 S.t282 6.541
R169 S.n761 S.t40 6.541
R170 S.n753 S.n752 6.541
R171 S.n1268 S.n1267 6.541
R172 S.n1276 S.t191 6.541
R173 S.n1279 S.t150 6.541
R174 S.n1271 S.n1270 6.541
R175 S.n1348 S.t44 6.541
R176 S.n323 S.t265 6.541
R177 S.n50 S.n49 6.541
R178 S.n66 S.t82 6.541
R179 S.n63 S.t139 6.541
R180 S.n53 S.n52 6.541
R181 S.n318 S.t94 6.541
R182 S.n356 S.t281 6.541
R183 S.n216 S.n215 6.541
R184 S.n229 S.t104 6.541
R185 S.n232 S.t149 6.541
R186 S.n219 S.n218 6.541
R187 S.n109 S.t43 6.541
R188 S.n259 S.t240 6.541
R189 S.n261 S.t148 6.541
R190 S.n172 S.n171 6.541
R191 S.n182 S.t123 6.541
R192 S.n185 S.t273 6.541
R193 S.n175 S.n174 6.541
R194 S.n596 S.n595 6.541
R195 S.n604 S.t255 6.541
R196 S.n607 S.t179 6.541
R197 S.n599 S.n598 6.541
R198 S.n491 S.n490 6.541
R199 S.n582 S.t91 6.541
R200 S.n585 S.t126 6.541
R201 S.n588 S.n587 6.541
R202 S.n840 S.n839 6.541
R203 S.n852 S.t259 6.541
R204 S.n855 S.t217 6.541
R205 S.n843 S.n842 6.541
R206 S.n723 S.n722 6.541
R207 S.n825 S.t95 6.541
R208 S.n828 S.t134 6.541
R209 S.n831 S.n830 6.541
R210 S.n1284 S.n1283 6.541
R211 S.n1296 S.t266 6.541
R212 S.n1299 S.t223 6.541
R213 S.n1287 S.n1286 6.541
R214 S.n1396 S.n1395 6.541
R215 S.n1406 S.t103 6.541
R216 S.n1409 S.t136 6.541
R217 S.n1399 S.n1398 6.541
R218 S.n1038 S.n1037 6.541
R219 S.n1053 S.t171 6.541
R220 S.n1050 S.t227 6.541
R221 S.n1041 S.n1040 6.541
R222 S.n934 S.n933 6.541
R223 S.n1023 S.t93 6.541
R224 S.n1026 S.t23 6.541
R225 S.n1029 S.n1028 6.541
R226 S.n1162 S.t132 6.541
R227 S.n1156 S.t71 6.541
R228 S.n610 S.t20 6.541
R229 S.n612 S.t46 6.541
R230 S.n566 S.n565 6.541
R231 S.n574 S.t237 6.541
R232 S.n577 S.t137 6.541
R233 S.n569 S.n568 6.541
R234 S.n863 S.n862 6.541
R235 S.n867 S.t169 6.541
R236 S.n870 S.t33 6.541
R237 S.n860 S.n859 6.541
R238 S.n1172 S.t22 6.541
R239 S.n1167 S.t247 6.541
R240 S.n921 S.n920 6.541
R241 S.n918 S.t262 6.541
R242 S.n915 S.t208 6.541
R243 S.n912 S.n911 6.541
R244 S.n907 S.n906 6.541
R245 S.n930 S.t74 6.541
R246 S.n927 S.t142 6.541
R247 S.n904 S.n903 6.541
R248 S.n1417 S.n1416 6.541
R249 S.n1421 S.t269 6.541
R250 S.n1424 S.t32 6.541
R251 S.n1414 S.n1413 6.541
R252 S.n1307 S.n1306 6.541
R253 S.n1312 S.t175 6.541
R254 S.n1315 S.t138 6.541
R255 S.n1304 S.n1303 6.541
R256 S.n792 S.n791 6.541
R257 S.n796 S.t264 6.541
R258 S.n799 S.t25 6.541
R259 S.n789 S.n788 6.541
R260 S.n875 S.t158 6.541
R261 S.n872 S.t225 6.541
R262 S.n802 S.n801 6.541
R263 S.n819 S.t86 6.541
R264 S.n822 S.t243 6.541
R265 S.n805 S.n804 6.541
R266 S.n1443 S.n1442 6.541
R267 S.n1452 S.t80 6.541
R268 S.n1455 S.t160 6.541
R269 S.n1446 S.n1445 6.541
R270 S.n1180 S.t207 6.541
R271 S.n1177 S.t162 6.541
R272 S.n986 S.n985 6.541
R273 S.n994 S.t172 6.541
R274 S.n997 S.t121 6.541
R275 S.n989 S.n988 6.541
R276 S.n888 S.n887 6.541
R277 S.n899 S.t249 6.541
R278 S.n896 S.t39 6.541
R279 S.n891 S.n890 6.541
R280 S.n1324 S.n1323 6.541
R281 S.n1427 S.t177 6.541
R282 S.n1430 S.t210 6.541
R283 S.n1433 S.n1432 6.541
R284 S.n1150 S.t57 6.541
R285 S.n1148 S.t242 6.541
R286 S.n1009 S.n1008 6.541
R287 S.n1017 S.t65 6.541
R288 S.n1020 S.t127 6.541
R289 S.n1012 S.n1011 6.541
R290 S.n496 S.t140 6.541
R291 S.n494 S.n493 6.541
R292 S.n503 S.n502 6.105
R293 S.n580 S.t209 6.105
R294 S.n882 S.t49 6.105
R295 S.n1193 S.t67 6.105
R296 S.n947 S.t258 6.105
R297 S.n955 S.n954 6.105
R298 S.n958 S.n957 6.105
R299 S.n950 S.t85 6.105
R300 S.n1091 S.t27 6.105
R301 S.n1099 S.n1098 6.105
R302 S.n1102 S.n1101 6.105
R303 S.n1094 S.t163 6.105
R304 S.n1373 S.t146 6.105
R305 S.n1391 S.n1390 6.105
R306 S.n1388 S.n1387 6.105
R307 S.n1376 S.t252 6.105
R308 S.n1462 S.t234 6.105
R309 S.n300 S.t11 6.105
R310 S.n283 S.t212 6.105
R311 S.n344 S.t56 6.105
R312 S.n340 S.t180 6.105
R313 S.n76 S.t55 6.105
R314 S.n204 S.n203 6.105
R315 S.n201 S.n200 6.105
R316 S.n79 S.t131 6.105
R317 S.n445 S.t73 6.105
R318 S.n460 S.n459 6.105
R319 S.n457 S.n456 6.105
R320 S.n442 S.t151 6.105
R321 S.n963 S.t108 6.105
R322 S.n964 S.t197 6.105
R323 S.n1063 S.t253 6.105
R324 S.n1081 S.n1080 6.105
R325 S.n1078 S.n1077 6.105
R326 S.n1060 S.t53 6.105
R327 S.n1356 S.t113 6.105
R328 S.n1367 S.n1366 6.105
R329 S.n1364 S.n1363 6.105
R330 S.n1353 S.t18 6.105
R331 S.n1239 S.t81 6.105
R332 S.n1254 S.n1253 6.105
R333 S.n1251 S.n1250 6.105
R334 S.n1236 S.t156 6.105
R335 S.n772 S.t109 6.105
R336 S.n783 S.n782 6.105
R337 S.n780 S.n779 6.105
R338 S.n769 S.t16 6.105
R339 S.n681 S.t79 6.105
R340 S.n698 S.n697 6.105
R341 S.n695 S.n694 6.105
R342 S.n678 S.t153 6.105
R343 S.n551 S.t106 6.105
R344 S.n560 S.n559 6.105
R345 S.n557 S.n556 6.105
R346 S.n548 S.t9 6.105
R347 S.n87 S.t99 6.105
R348 S.n188 S.n187 6.105
R349 S.n191 S.n190 6.105
R350 S.n194 S.t3 6.105
R351 S.n314 S.t14 6.105
R352 S.n305 S.t111 6.105
R353 S.n17 S.t257 6.105
R354 S.n45 S.n44 6.105
R355 S.n42 S.n41 6.105
R356 S.n20 S.t155 6.105
R357 S.n472 S.t89 6.105
R358 S.n484 S.n483 6.105
R359 S.n487 S.n486 6.105
R360 S.n469 S.t157 6.105
R361 S.n523 S.t117 6.105
R362 S.n504 S.t28 6.105
R363 S.n114 S.t112 6.105
R364 S.n129 S.n128 6.105
R365 S.n126 S.n125 6.105
R366 S.n117 S.t17 6.105
R367 S.n141 S.t284 6.105
R368 S.n149 S.n148 6.105
R369 S.n146 S.n145 6.105
R370 S.n138 S.t205 6.105
R371 S.n399 S.t260 6.105
R372 S.n417 S.n416 6.105
R373 S.n414 S.n413 6.105
R374 S.n396 S.t60 6.105
R375 S.n702 S.t263 6.105
R376 S.n716 S.n715 6.105
R377 S.n719 S.n718 6.105
R378 S.n705 S.t63 6.105
R379 S.n743 S.t5 6.105
R380 S.n725 S.t213 6.105
R381 S.n270 S.t168 6.105
R382 S.n267 S.n266 6.105
R383 S.n264 S.n263 6.105
R384 S.n8 S.t58 6.105
R385 S.n159 S.t192 6.105
R386 S.n167 S.n166 6.105
R387 S.n164 S.n163 6.105
R388 S.n156 S.t118 6.105
R389 S.n426 S.t170 6.105
R390 S.n437 S.n436 6.105
R391 S.n434 S.n433 6.105
R392 S.n429 S.t233 6.105
R393 S.n530 S.t195 6.105
R394 S.n543 S.n542 6.105
R395 S.n540 S.n539 6.105
R396 S.n533 S.t122 6.105
R397 S.n652 S.t173 6.105
R398 S.n664 S.n663 6.105
R399 S.n661 S.n660 6.105
R400 S.n655 S.t236 6.105
R401 S.n750 S.t198 6.105
R402 S.n764 S.n763 6.105
R403 S.n761 S.n760 6.105
R404 S.n753 S.t125 6.105
R405 S.n1268 S.t176 6.105
R406 S.n1276 S.n1275 6.105
R407 S.n1279 S.n1278 6.105
R408 S.n1271 S.t239 6.105
R409 S.n1347 S.t202 6.105
R410 S.n1326 S.t130 6.105
R411 S.n335 S.t115 6.105
R412 S.n322 S.t188 6.105
R413 S.n50 S.t72 6.105
R414 S.n66 S.n65 6.105
R415 S.n63 S.n62 6.105
R416 S.n53 S.t230 6.105
R417 S.n317 S.t203 6.105
R418 S.n315 S.t280 6.105
R419 S.n358 S.t124 6.105
R420 S.n359 S.t200 6.105
R421 S.n216 S.t84 6.105
R422 S.n229 S.n228 6.105
R423 S.n232 S.n231 6.105
R424 S.n219 S.t238 6.105
R425 S.n108 S.t201 6.105
R426 S.n89 S.t129 6.105
R427 S.n250 S.t235 6.105
R428 S.n172 S.t35 6.105
R429 S.n182 S.n181 6.105
R430 S.n185 S.n184 6.105
R431 S.n175 S.t167 6.105
R432 S.n596 S.t116 6.105
R433 S.n604 S.n603 6.105
R434 S.n607 S.n606 6.105
R435 S.n599 S.t241 6.105
R436 S.n491 S.t272 6.105
R437 S.n582 S.n581 6.105
R438 S.n585 S.n584 6.105
R439 S.n588 S.t199 6.105
R440 S.n840 S.t250 6.105
R441 S.n852 S.n851 6.105
R442 S.n855 S.n854 6.105
R443 S.n843 S.t52 6.105
R444 S.n723 S.t276 6.105
R445 S.n825 S.n824 6.105
R446 S.n828 S.n827 6.105
R447 S.n831 S.t204 6.105
R448 S.n1284 S.t254 6.105
R449 S.n1296 S.n1295 6.105
R450 S.n1299 S.n1298 6.105
R451 S.n1287 S.t59 6.105
R452 S.n1396 S.t285 6.105
R453 S.n1406 S.n1405 6.105
R454 S.n1409 S.n1408 6.105
R455 S.n1399 S.t206 6.105
R456 S.n1038 S.t165 6.105
R457 S.n1053 S.n1052 6.105
R458 S.n1050 S.n1049 6.105
R459 S.n1041 S.t228 6.105
R460 S.n934 S.t275 6.105
R461 S.n1023 S.n1022 6.105
R462 S.n1026 S.n1025 6.105
R463 S.n1029 S.t107 6.105
R464 S.n1155 S.t69 6.105
R465 S.n614 S.t154 6.105
R466 S.n566 S.t161 6.105
R467 S.n574 S.n573 6.105
R468 S.n577 S.n576 6.105
R469 S.n569 S.t12 6.105
R470 S.n863 S.t231 6.105
R471 S.n867 S.n866 6.105
R472 S.n870 S.n869 6.105
R473 S.n860 S.t100 6.105
R474 S.n1168 S.t244 6.105
R475 S.n921 S.t184 6.105
R476 S.n918 S.n917 6.105
R477 S.n915 S.n914 6.105
R478 S.n912 S.t274 6.105
R479 S.n907 S.t70 6.105
R480 S.n930 S.n929 6.105
R481 S.n927 S.n926 6.105
R482 S.n904 S.t144 6.105
R483 S.n1417 S.t193 6.105
R484 S.n1421 S.n1420 6.105
R485 S.n1424 S.n1423 6.105
R486 S.n1414 S.t119 6.105
R487 S.n1307 S.t166 6.105
R488 S.n1312 S.n1311 6.105
R489 S.n1315 S.n1314 6.105
R490 S.n1304 S.t232 6.105
R491 S.n792 S.t185 6.105
R492 S.n796 S.n795 6.105
R493 S.n799 S.n798 6.105
R494 S.n789 S.t114 6.105
R495 S.n643 S.t62 6.105
R496 S.n802 S.t279 6.105
R497 S.n819 S.n818 6.105
R498 S.n822 S.n821 6.105
R499 S.n805 S.t152 6.105
R500 S.n1443 S.t77 6.105
R501 S.n1452 S.n1451 6.105
R502 S.n1455 S.n1454 6.105
R503 S.n1446 S.t221 6.105
R504 S.n1176 S.t159 6.105
R505 S.n986 S.t88 6.105
R506 S.n994 S.n993 6.105
R507 S.n997 S.n996 6.105
R508 S.n989 S.t183 6.105
R509 S.n888 S.t246 6.105
R510 S.n899 S.n898 6.105
R511 S.n896 S.n895 6.105
R512 S.n891 S.t41 6.105
R513 S.n1324 S.t98 6.105
R514 S.n1427 S.n1426 6.105
R515 S.n1430 S.n1429 6.105
R516 S.n1433 S.t1 6.105
R517 S.n1151 S.t248 6.105
R518 S.n1009 S.t245 6.105
R519 S.n1017 S.n1016 6.105
R520 S.n1020 S.n1019 6.105
R521 S.n1012 S.t87 6.105
R522 S.n496 S.n495 6.105
R523 S.n494 S.t286 6.105
R524 S.n98 S.n96 4.263
R525 S.n513 S.n511 4.263
R526 S.n733 S.n731 4.263
R527 S.n1337 S.n1335 4.263
R528 S.n975 S.n973 4.263
R529 S.n287 S.n286 2.645
R530 S.n92 S.n91 2.645
R531 S.n507 S.n506 2.645
R532 S.n727 S.n726 2.645
R533 S.n1331 S.n1330 2.645
R534 S.n624 S.n623 0.21
R535 S.n1208 S.n1205 0.178
R536 S.n289 S.n285 0.164
R537 S.n1211 S.n1210 0.141
R538 S.n247 S.n246 0.136
R539 S.n713 S.n712 0.133
R540 S.n658 S.n657 0.133
R541 S.n379 S.n374 0.123
R542 S.n1482 S.n621 0.116
R543 S.n1481 S.n881 0.111
R544 S.n1154 S.n1153 0.11
R545 S.n1480 S.n1479 0.11
R546 S.n1211 S.n1120 0.11
R547 S.n133 S.n132 0.109
R548 S.n758 S.n756 0.109
R549 S.n153 S.n152 0.109
R550 S.n179 S.n178 0.109
R551 S.n1384 S.n1379 0.106
R552 S.n36 S.n31 0.104
R553 S.n35 S.n32 0.097
R554 S.n1472 S.n1471 0.095
R555 S.n1166 S.n1165 0.093
R556 S.n968 S.n967 0.093
R557 S.n1329 S.n1328 0.093
R558 S.n1000 S.n999 0.092
R559 S.n938 S.n937 0.092
R560 S S.n1483 0.09
R561 S.n1147 S.n1146 0.087
R562 S.n1164 S.n1163 0.085
R563 S.n248 S.n244 0.082
R564 S.n389 S.n386 0.082
R565 S.n641 S.n638 0.082
R566 S.n1222 S.n1219 0.082
R567 S.n1118 S.n1114 0.082
R568 S.n1122 S.n1121 0.08
R569 S.n738 S.n737 0.076
R570 S.n980 S.n979 0.074
R571 S.n518 S.n517 0.074
R572 S.n1342 S.n1341 0.074
R573 S.n103 S.n102 0.074
R574 S.n1170 S.n1169 0.073
R575 S.n1175 S.n1174 0.073
R576 S.n257 S.n256 0.071
R577 S.n1382 S.n1381 0.07
R578 S.t66 S.n1160 0.068
R579 S.n338 S.n336 0.067
R580 S.n338 S.n337 0.067
R581 S.n303 S.n301 0.067
R582 S.n332 S.n330 0.067
R583 S.n332 S.n331 0.067
R584 S.n362 S.n361 0.067
R585 S.n303 S.n302 0.067
R586 S.n354 S.n352 0.067
R587 S.n354 S.n353 0.067
R588 S.n248 S.n238 0.067
R589 S.n248 S.n236 0.067
R590 S.n641 S.n632 0.067
R591 S.n641 S.n631 0.067
R592 S.n1118 S.n1108 0.067
R593 S.n1222 S.n1213 0.067
R594 S.n1222 S.n1212 0.067
R595 S.n1118 S.n1117 0.067
R596 S.n362 S.n360 0.067
R597 S.n296 S.n295 0.066
R598 S.n275 S.n3 0.066
R599 S.n249 S.n234 0.065
R600 S.n198 S.n197 0.064
R601 S.n333 S.n329 0.063
R602 S.n1223 S.n1222 0.063
R603 S.n333 S.n332 0.063
R604 S.n455 S.n454 0.063
R605 S.n693 S.n692 0.063
R606 S.n778 S.n777 0.063
R607 S.n1249 S.n1248 0.063
R608 S.n1362 S.n1361 0.063
R609 S.n199 S.n69 0.063
R610 S.n196 S.n83 0.063
R611 S.n432 S.n420 0.063
R612 S.n659 S.n646 0.063
R613 S.n61 S.n48 0.063
R614 S.n227 S.n226 0.063
R615 S.n120 S.n119 0.062
R616 S.n339 S.n338 0.062
R617 S.n304 S.n303 0.062
R618 S.n373 S.n362 0.061
R619 S.n355 S.n354 0.06
R620 S.n1072 S.n1071 0.059
R621 S.n1258 S.n1257 0.059
R622 S.n1119 S.n1118 0.058
R623 S.n249 S.n248 0.058
R624 S.n347 S.n346 0.056
R625 S.n299 S.n283 0.055
R626 S.n1461 S.n1460 0.055
R627 S.n262 S.n261 0.055
R628 S.n613 S.n612 0.055
R629 S.n873 S.n872 0.055
R630 S.n1106 S.n882 0.054
R631 S.n982 S.n964 0.054
R632 S.n521 S.n504 0.054
R633 S.n741 S.n725 0.054
R634 S.n1345 S.n1326 0.054
R635 S.n106 S.n89 0.054
R636 S.n1209 S.n1208 0.054
R637 S.n959 S.n958 0.054
R638 S.n1103 S.n1102 0.054
R639 S.n1389 S.n1388 0.054
R640 S.n202 S.n201 0.054
R641 S.n458 S.n457 0.054
R642 S.n1079 S.n1078 0.054
R643 S.n1365 S.n1364 0.054
R644 S.n1252 S.n1251 0.054
R645 S.n781 S.n780 0.054
R646 S.n696 S.n695 0.054
R647 S.n558 S.n557 0.054
R648 S.n192 S.n191 0.054
R649 S.n43 S.n42 0.054
R650 S.n488 S.n487 0.054
R651 S.n127 S.n126 0.054
R652 S.n147 S.n146 0.054
R653 S.n415 S.n414 0.054
R654 S.n720 S.n719 0.054
R655 S.n265 S.n264 0.054
R656 S.n165 S.n164 0.054
R657 S.n435 S.n434 0.054
R658 S.n541 S.n540 0.054
R659 S.n662 S.n661 0.054
R660 S.n762 S.n761 0.054
R661 S.n1280 S.n1279 0.054
R662 S.n64 S.n63 0.054
R663 S.n233 S.n232 0.054
R664 S.n186 S.n185 0.054
R665 S.n608 S.n607 0.054
R666 S.n586 S.n585 0.054
R667 S.n856 S.n855 0.054
R668 S.n829 S.n828 0.054
R669 S.n1300 S.n1299 0.054
R670 S.n1410 S.n1409 0.054
R671 S.n1051 S.n1050 0.054
R672 S.n1027 S.n1026 0.054
R673 S.n578 S.n577 0.054
R674 S.n871 S.n870 0.054
R675 S.n916 S.n915 0.054
R676 S.n928 S.n927 0.054
R677 S.n1425 S.n1424 0.054
R678 S.n1316 S.n1315 0.054
R679 S.n800 S.n799 0.054
R680 S.n823 S.n822 0.054
R681 S.n1456 S.n1455 0.054
R682 S.n998 S.n997 0.054
R683 S.n897 S.n896 0.054
R684 S.n1431 S.n1430 0.054
R685 S.n1021 S.n1020 0.054
R686 S.n1197 S.n1123 0.053
R687 S.t90 S.n496 0.052
R688 S.n101 S.n100 0.052
R689 S.n516 S.n515 0.052
R690 S.n736 S.n735 0.052
R691 S.n1340 S.n1339 0.052
R692 S.n978 S.n977 0.052
R693 S.n392 S.n391 0.052
R694 S.n879 S.n878 0.052
R695 S.n1477 S.n1476 0.052
R696 S.n1381 S.n1380 0.052
R697 S.t90 S.n580 0.051
R698 S.n480 S.n478 0.051
R699 S.n210 S.n208 0.051
R700 S.n1131 S.n1130 0.051
R701 S.n1133 S.n1132 0.051
R702 S.n1186 S.n1185 0.051
R703 S.n238 S.n237 0.051
R704 S.n236 S.n235 0.051
R705 S.n1076 S.n1075 0.05
R706 S.n482 S.n481 0.05
R707 S.n1274 S.n1261 0.05
R708 S.n227 S.n211 0.05
R709 S.n72 S.n71 0.05
R710 S.n136 S.n135 0.049
R711 S.n624 S.n622 0.049
R712 S.n816 S.n815 0.048
R713 S.n390 S.n389 0.048
R714 S.n642 S.n641 0.048
R715 S.n309 S.n308 0.047
R716 S.n953 S.n951 0.047
R717 S.n1097 S.n1095 0.047
R718 S.n1386 S.n1377 0.047
R719 S.n1479 S.n1463 0.047
R720 S.n199 S.n80 0.047
R721 S.n455 S.n443 0.047
R722 S.n1076 S.n1061 0.047
R723 S.n1362 S.n1354 0.047
R724 S.n1249 S.n1237 0.047
R725 S.n778 S.n770 0.047
R726 S.n693 S.n679 0.047
R727 S.n555 S.n549 0.047
R728 S.n196 S.n195 0.047
R729 S.n40 S.n21 0.047
R730 S.n482 S.n470 0.047
R731 S.n124 S.n118 0.047
R732 S.n144 S.n139 0.047
R733 S.n412 S.n397 0.047
R734 S.n714 S.n706 0.047
R735 S.n275 S.n9 0.047
R736 S.n162 S.n157 0.047
R737 S.n432 S.n430 0.047
R738 S.n538 S.n534 0.047
R739 S.n659 S.n656 0.047
R740 S.n759 S.n754 0.047
R741 S.n1274 S.n1272 0.047
R742 S.n61 S.n54 0.047
R743 S.n227 S.n220 0.047
R744 S.n257 S.n251 0.047
R745 S.n180 S.n176 0.047
R746 S.n602 S.n600 0.047
R747 S.n593 S.n589 0.047
R748 S.n850 S.n844 0.047
R749 S.n836 S.n832 0.047
R750 S.n1294 S.n1288 0.047
R751 S.n1404 S.n1400 0.047
R752 S.n1048 S.n1042 0.047
R753 S.n1034 S.n1030 0.047
R754 S.n620 S.n615 0.047
R755 S.n572 S.n570 0.047
R756 S.n865 S.n861 0.047
R757 S.n923 S.n913 0.047
R758 S.n925 S.n905 0.047
R759 S.n1419 S.n1415 0.047
R760 S.n1310 S.n1305 0.047
R761 S.n794 S.n790 0.047
R762 S.n881 S.n644 0.047
R763 S.n817 S.n806 0.047
R764 S.n1450 S.n1447 0.047
R765 S.n992 S.n990 0.047
R766 S.n894 S.n892 0.047
R767 S.n1436 S.n1434 0.047
R768 S.n1015 S.n1013 0.047
R769 S.n321 S.n320 0.046
R770 S.n602 S.n593 0.046
R771 S.n1449 S.n1448 0.045
R772 S.n1182 S.n1181 0.045
R773 S.n409 S.n401 0.045
R774 S.n273 S.n272 0.045
R775 S.n1184 S.n1183 0.045
R776 S.n121 S.n120 0.045
R777 S.n1127 S.n1126 0.045
R778 S.n1450 S.n1436 0.044
R779 S.n850 S.n837 0.044
R780 S.n1294 S.n1281 0.044
R781 S.n1048 S.n1035 0.044
R782 S.n1310 S.n1309 0.044
R783 S.n925 S.n924 0.044
R784 S.n1154 S.n1152 0.044
R785 S.n312 S.n310 0.044
R786 S.n373 S.n372 0.043
R787 S.n1075 S.n1074 0.043
R788 S.n1261 S.n1260 0.043
R789 S.n244 S.n240 0.043
R790 S.n386 S.n382 0.043
R791 S.n638 S.n634 0.043
R792 S.n1219 S.n1215 0.043
R793 S.n1114 S.n1110 0.043
R794 S.n351 S.n350 0.043
R795 S.n325 S.n324 0.043
R796 S.n223 S.n222 0.042
R797 S.n1245 S.n1242 0.042
R798 S.n689 S.n684 0.042
R799 S.n451 S.n448 0.042
R800 S.n277 S.n276 0.042
R801 S.n648 S.n647 0.042
R802 S.n422 S.n421 0.042
R803 S.n971 S.n970 0.042
R804 S.n329 S.n328 0.041
R805 S.n467 S.n466 0.041
R806 S.n349 S.n348 0.041
R807 S.n253 S.n252 0.041
R808 S.n297 S.n289 0.04
R809 S.n101 S.n92 0.04
R810 S.n516 S.n507 0.04
R811 S.n736 S.n727 0.04
R812 S.n1340 S.n1331 0.04
R813 S.n978 S.n969 0.04
R814 S.n1139 S.n1138 0.04
R815 S.n1137 S.n1136 0.04
R816 S.n1174 S.n1173 0.039
R817 S.n288 S.n287 0.039
R818 S.n1468 S.n1467 0.039
R819 S.n1188 S.n1187 0.039
R820 S.n100 S.n93 0.039
R821 S.n515 S.n508 0.039
R822 S.n735 S.n728 0.039
R823 S.n1339 S.n1332 0.039
R824 S.n968 S.n966 0.038
R825 S.n1329 S.n1327 0.038
R826 S.n1233 S.n1232 0.038
R827 S.n675 S.n674 0.038
R828 S.n711 S.n710 0.037
R829 S.n1468 S.n1465 0.037
R830 S.n1467 S.n1466 0.037
R831 S.n885 S.n884 0.037
R832 S.n1440 S.n1439 0.037
R833 S.n257 S.n253 0.036
R834 S.n527 S.n526 0.036
R835 S.n747 S.n746 0.036
R836 S.n1088 S.n1087 0.035
R837 S.n1056 S.n1055 0.035
R838 S.n961 S.n960 0.035
R839 S.n525 S.n524 0.035
R840 S.n745 S.n744 0.035
R841 S.n1349 S.n1348 0.035
R842 S.n110 S.n109 0.035
R843 S.n1469 S.n1468 0.035
R844 S.n1233 S.n1228 0.035
R845 S.n675 S.n670 0.035
R846 S.n482 S.n467 0.035
R847 S.n34 S.n33 0.035
R848 S.t66 S.n1194 0.035
R849 S.t10 S.n341 0.035
R850 S.t10 S.n306 0.035
R851 S.t10 S.n323 0.035
R852 S.t10 S.n318 0.035
R853 S.t10 S.n356 0.035
R854 S.t66 S.n1156 0.035
R855 S.t66 S.n1167 0.035
R856 S.t66 S.n1177 0.035
R857 S.t66 S.n1148 0.035
R858 S.n1159 S.n1158 0.035
R859 S.n629 S.n628 0.034
R860 S.n1034 S.n1031 0.034
R861 S.n1048 S.n1044 0.034
R862 S.n1404 S.n1401 0.034
R863 S.n1294 S.n1290 0.034
R864 S.n836 S.n833 0.034
R865 S.n850 S.n846 0.034
R866 S.n593 S.n590 0.034
R867 S.n620 S.n380 0.034
R868 S.n881 S.n880 0.034
R869 S.n1479 S.n1478 0.034
R870 S.n518 S.n505 0.034
R871 S.n103 S.n90 0.034
R872 S.t66 S.n1193 0.034
R873 S.t10 S.n340 0.034
R874 S.t10 S.n305 0.034
R875 S.t10 S.n322 0.034
R876 S.t10 S.n315 0.034
R877 S.t10 S.n359 0.034
R878 S.t66 S.n1155 0.034
R879 S.t66 S.n1168 0.034
R880 S.t66 S.n1176 0.034
R881 S.t66 S.n1151 0.034
R882 S.n297 S.n296 0.033
R883 S.n980 S.n968 0.032
R884 S.n1342 S.n1329 0.032
R885 S.n475 S.n474 0.031
R886 S.t26 S.n1056 0.031
R887 S.t64 S.n961 0.031
R888 S.t90 S.n525 0.031
R889 S.t4 S.n745 0.031
R890 S.t97 S.n1349 0.031
R891 S.t34 S.n110 0.031
R892 S.n1228 S.n1227 0.031
R893 S.n670 S.n669 0.031
R894 S.n376 S.n375 0.031
R895 S.n377 S.n376 0.031
R896 S.n378 S.n377 0.031
R897 S.n379 S.n378 0.031
R898 S.n255 S.n254 0.031
R899 S.n1483 S.n1482 0.031
R900 S.n1482 S.n1481 0.031
R901 S.n1481 S.n1480 0.031
R902 S.n1480 S.n1211 0.031
R903 S.n1046 S.n1045 0.031
R904 S.n1292 S.n1291 0.031
R905 S.n848 S.n847 0.031
R906 S.n404 S.n403 0.03
R907 S.n365 S.n364 0.03
R908 S.n99 S.n94 0.03
R909 S.n514 S.n509 0.03
R910 S.n734 S.n729 0.03
R911 S.n1338 S.n1333 0.03
R912 S.n451 S.n450 0.029
R913 S.n689 S.n688 0.029
R914 S.n1245 S.n1244 0.029
R915 S.n403 S.n402 0.029
R916 S.n364 S.n363 0.029
R917 S.n1228 S.n1225 0.028
R918 S.n670 S.n667 0.028
R919 S.n1069 S.n1068 0.028
R920 S.n885 S.n883 0.027
R921 S.n1440 S.n1438 0.027
R922 S.n1205 S.n1204 0.027
R923 S.n312 S.n311 0.027
R924 S.n57 S.n56 0.027
R925 S.n275 S.n6 0.027
R926 S.n620 S.n619 0.027
R927 S.n846 S.n845 0.027
R928 S.n1290 S.n1289 0.027
R929 S.n1044 S.n1043 0.027
R930 S.n455 S.n452 0.026
R931 S.n555 S.n554 0.026
R932 S.n693 S.n690 0.026
R933 S.n778 S.n775 0.026
R934 S.n1249 S.n1246 0.026
R935 S.n1362 S.n1359 0.026
R936 S.n1076 S.n1070 0.026
R937 S.n196 S.n85 0.026
R938 S.n482 S.n476 0.026
R939 S.n501 S.n500 0.026
R940 S.n758 S.n757 0.026
R941 S.n537 S.n536 0.026
R942 S.n432 S.n423 0.026
R943 S.n659 S.n649 0.026
R944 S.n1274 S.n1265 0.026
R945 S.n227 S.n214 0.026
R946 S.n227 S.n224 0.026
R947 S.n1386 S.n1370 0.026
R948 S.n1006 S.n1005 0.026
R949 S.n213 S.n212 0.026
R950 S.n944 S.n943 0.026
R951 S.n24 S.n23 0.026
R952 S.t10 S.n349 0.025
R953 S.n13 S.n12 0.025
R954 S.n282 S.n281 0.024
R955 S.n388 S.n387 0.024
R956 S.n640 S.n639 0.024
R957 S.n1221 S.n1220 0.024
R958 S.n1116 S.n1115 0.024
R959 S.n1207 S.n1206 0.024
R960 S.n619 S.n618 0.024
R961 S.n281 S.n280 0.024
R962 S.n1379 S.n1378 0.023
R963 S.n1477 S.n1464 0.023
R964 S.n1192 S.n1184 0.023
R965 S.n122 S.n121 0.023
R966 S.n14 S.n11 0.023
R967 S.n58 S.n57 0.023
R968 S.n6 S.n4 0.023
R969 S.t10 S.n282 0.023
R970 S.n136 S.n134 0.023
R971 S.n1159 S.n1157 0.023
R972 S.n392 S.n390 0.023
R973 S.n617 S.n616 0.023
R974 S.n879 S.n877 0.023
R975 S.n1135 S.n1127 0.023
R976 S.n1074 S.n1073 0.022
R977 S.n1260 S.n1259 0.022
R978 S.n36 S.n35 0.022
R979 S.n368 S.n367 0.022
R980 S.n407 S.n406 0.022
R981 S.n480 S.n479 0.022
R982 S.n210 S.n209 0.022
R983 S.n1264 S.n1263 0.022
R984 S.n1069 S.n1066 0.021
R985 S.n450 S.n449 0.021
R986 S.n448 S.n447 0.021
R987 S.n688 S.n687 0.021
R988 S.n684 S.n683 0.021
R989 S.n1244 S.n1243 0.021
R990 S.n1242 S.n1241 0.021
R991 S.n1068 S.n1067 0.021
R992 S.n71 S.n70 0.021
R993 S.n1227 S.n1226 0.021
R994 S.n669 S.n668 0.021
R995 S.n69 S.n68 0.021
R996 S.n481 S.n480 0.021
R997 S.n711 S.n708 0.021
R998 S.n211 S.n210 0.021
R999 S.n1166 S.n1164 0.021
R1000 S.n37 S.n30 0.021
R1001 S.n625 S.n624 0.021
R1002 S.n26 S.n25 0.02
R1003 S.n1134 S.n1128 0.02
R1004 S.n1191 S.n1188 0.02
R1005 S.n328 S.n327 0.02
R1006 S.n222 S.n221 0.02
R1007 S.n1087 S.n1086 0.02
R1008 S.n1075 S.n1072 0.02
R1009 S.n481 S.n477 0.02
R1010 S.n1261 S.n1258 0.02
R1011 S.n211 S.n207 0.02
R1012 S.n320 S.n319 0.02
R1013 S.t10 S.n312 0.019
R1014 S.n274 S.n273 0.019
R1015 S.n1321 S.n1320 0.019
R1016 S.n411 S.n410 0.019
R1017 S.n1 S.n0 0.018
R1018 S.n11 S.n10 0.018
R1019 S S.n379 0.018
R1020 S.n813 S.n812 0.018
R1021 S.n279 S.n278 0.018
R1022 S.n810 S.n809 0.017
R1023 S.n39 S.n38 0.017
R1024 S.n1003 S.n1002 0.017
R1025 S.n941 S.n940 0.017
R1026 S.n817 S.n814 0.017
R1027 S.n1474 S.n1473 0.017
R1028 S.n244 S.n243 0.017
R1029 S.n386 S.n385 0.017
R1030 S.n638 S.n637 0.017
R1031 S.n1219 S.n1218 0.017
R1032 S.n1114 S.n1113 0.017
R1033 S.n1473 S.n1472 0.017
R1034 S.n1438 S.n1437 0.015
R1035 S.n1066 S.n1065 0.015
R1036 S.n1263 S.n1262 0.015
R1037 S.n60 S.n59 0.015
R1038 S.t66 S.n1159 0.015
R1039 S.n1319 S.n1318 0.015
R1040 S.n1318 S.n1317 0.015
R1041 S.n812 S.n811 0.015
R1042 S.n881 S.n642 0.015
R1043 S.n369 S.n368 0.015
R1044 S.n368 S.n365 0.015
R1045 S.n409 S.n408 0.015
R1046 S.n408 S.n407 0.015
R1047 S.n407 S.n404 0.015
R1048 S.n1230 S.n1229 0.015
R1049 S.n672 S.n671 0.015
R1050 S.n372 S.n371 0.014
R1051 S.n628 S.n626 0.014
R1052 S.n894 S.n885 0.014
R1053 S.n1450 S.n1440 0.014
R1054 S.n1385 S.n1384 0.014
R1055 S.n1234 S.n1233 0.013
R1056 S.n676 S.n675 0.013
R1057 S.n710 S.n709 0.013
R1058 S.n30 S.n29 0.013
R1059 S.n1384 S.n1383 0.013
R1060 S.t10 S.n345 0.012
R1061 S.n642 S.n630 0.012
R1062 S.n1470 S.n1469 0.012
R1063 S.n1231 S.n1230 0.012
R1064 S.n673 S.n672 0.012
R1065 S.n199 S.n73 0.012
R1066 S.n35 S.n34 0.012
R1067 S.n1132 S.n1131 0.012
R1068 S.n1187 S.n1186 0.012
R1069 S.n1383 S.n1382 0.012
R1070 S.n40 S.n24 0.011
R1071 S.n953 S.n944 0.011
R1072 S.n1015 S.n1006 0.011
R1073 S.n817 S.n810 0.01
R1074 S.n465 S.n464 0.01
R1075 S.n14 S.n13 0.01
R1076 S.t90 S.n499 0.01
R1077 S.n759 S.n755 0.01
R1078 S.n538 S.n535 0.01
R1079 S.n162 S.n154 0.01
R1080 S.n144 S.n136 0.01
R1081 S.n40 S.n39 0.01
R1082 S.n180 S.n177 0.01
R1083 S.n620 S.n617 0.01
R1084 S.n620 S.n392 0.01
R1085 S.n881 S.n879 0.01
R1086 S.n1015 S.n1003 0.01
R1087 S.n953 S.n941 0.01
R1088 S.n1479 S.n1477 0.01
R1089 S.n1472 S.n1470 0.01
R1090 S.n1120 S.n1107 0.009
R1091 S.n1475 S.n1474 0.009
R1092 S.n714 S.n711 0.009
R1093 S.t66 S.n1166 0.009
R1094 S.n1479 S.n1223 0.009
R1095 S.n38 S.n37 0.008
R1096 S.n1002 S.n1001 0.008
R1097 S.n940 S.n939 0.008
R1098 S.n1134 S.n1133 0.008
R1099 S.n1191 S.n1190 0.008
R1100 S.n1232 S.n1231 0.008
R1101 S.n674 S.n673 0.008
R1102 S.n454 S.n453 0.008
R1103 S.n686 S.n685 0.008
R1104 S.n692 S.n691 0.008
R1105 S.n777 S.n776 0.008
R1106 S.n1248 S.n1247 0.008
R1107 S.n1361 S.n1360 0.008
R1108 S.n83 S.n82 0.008
R1109 S.t90 S.n501 0.008
R1110 S.n759 S.n758 0.008
R1111 S.n538 S.n537 0.008
R1112 S.n162 S.n153 0.008
R1113 S.n420 S.n419 0.008
R1114 S.n646 S.n645 0.008
R1115 S.n48 S.n47 0.008
R1116 S.n59 S.n55 0.008
R1117 S.n59 S.n58 0.008
R1118 S.n144 S.n133 0.008
R1119 S.n226 S.n225 0.008
R1120 S.n180 S.n179 0.008
R1121 S.n257 S.n255 0.008
R1122 S.n817 S.n816 0.008
R1123 S.n1085 S.n1084 0.008
R1124 S.n3 S.n2 0.008
R1125 S.n3 S.n1 0.007
R1126 S.n123 S.n122 0.007
R1127 S.n371 S.n370 0.007
R1128 S.n809 S.n808 0.007
R1129 S.n214 S.n213 0.007
R1130 S.t66 S.n1178 0.006
R1131 S.n687 S.n686 0.006
R1132 S.n1086 S.n1085 0.006
R1133 S.n124 S.n123 0.006
R1134 S.n1135 S.n1134 0.006
R1135 S.n1192 S.n1191 0.006
R1136 S.n27 S.n26 0.006
R1137 S.n40 S.n14 0.006
R1138 S.t10 S.n309 0.005
R1139 S.n1133 S.n1129 0.005
R1140 S.n1190 S.n1189 0.005
R1141 S.t10 S.n373 0.005
R1142 S.n951 S.n950 0.004
R1143 S.n1095 S.n1094 0.004
R1144 S.n1377 S.n1376 0.004
R1145 S.n1463 S.n1462 0.004
R1146 S.n80 S.n79 0.004
R1147 S.n443 S.n442 0.004
R1148 S.n1061 S.n1060 0.004
R1149 S.n1354 S.n1353 0.004
R1150 S.n1237 S.n1236 0.004
R1151 S.n770 S.n769 0.004
R1152 S.n679 S.n678 0.004
R1153 S.n549 S.n548 0.004
R1154 S.n195 S.n194 0.004
R1155 S.n21 S.n20 0.004
R1156 S.n470 S.n469 0.004
R1157 S.n118 S.n117 0.004
R1158 S.n139 S.n138 0.004
R1159 S.n397 S.n396 0.004
R1160 S.n706 S.n705 0.004
R1161 S.n9 S.n8 0.004
R1162 S.n157 S.n156 0.004
R1163 S.n430 S.n429 0.004
R1164 S.n534 S.n533 0.004
R1165 S.n656 S.n655 0.004
R1166 S.n754 S.n753 0.004
R1167 S.n1272 S.n1271 0.004
R1168 S.n54 S.n53 0.004
R1169 S.n220 S.n219 0.004
R1170 S.n251 S.n250 0.004
R1171 S.n176 S.n175 0.004
R1172 S.n600 S.n599 0.004
R1173 S.n589 S.n588 0.004
R1174 S.n844 S.n843 0.004
R1175 S.n832 S.n831 0.004
R1176 S.n1288 S.n1287 0.004
R1177 S.n1400 S.n1399 0.004
R1178 S.n1042 S.n1041 0.004
R1179 S.n1030 S.n1029 0.004
R1180 S.n615 S.n614 0.004
R1181 S.n570 S.n569 0.004
R1182 S.n861 S.n860 0.004
R1183 S.n913 S.n912 0.004
R1184 S.n905 S.n904 0.004
R1185 S.n1415 S.n1414 0.004
R1186 S.n1305 S.n1304 0.004
R1187 S.n790 S.n789 0.004
R1188 S.n644 S.n643 0.004
R1189 S.n806 S.n805 0.004
R1190 S.n1447 S.n1446 0.004
R1191 S.n990 S.n989 0.004
R1192 S.n892 S.n891 0.004
R1193 S.n1434 S.n1433 0.004
R1194 S.n1013 S.n1012 0.004
R1195 S.t10 S.n279 0.004
R1196 S.n199 S.n198 0.004
R1197 S.t10 S.n321 0.004
R1198 S.n520 S.n519 0.004
R1199 S.n105 S.n104 0.004
R1200 S.n367 S.n366 0.004
R1201 S.n406 S.n405 0.004
R1202 S.n981 S.n980 0.004
R1203 S.n520 S.n518 0.004
R1204 S.n162 S.n161 0.004
R1205 S.n538 S.n527 0.004
R1206 S.n759 S.n747 0.004
R1207 S.n1344 S.n1342 0.004
R1208 S.n105 S.n103 0.004
R1209 S.n29 S.n28 0.004
R1210 S.n1321 S.n1319 0.004
R1211 S.n630 S.n629 0.004
R1212 S.n881 S.n625 0.004
R1213 S.n411 S.n409 0.004
R1214 S.t66 S.n1170 0.004
R1215 S.t66 S.n1175 0.004
R1216 S.t10 S.n300 0.004
R1217 S.t10 S.n344 0.004
R1218 S.t64 S.n963 0.004
R1219 S.t10 S.n314 0.004
R1220 S.t90 S.n523 0.004
R1221 S.t4 S.n743 0.004
R1222 S.t97 S.n1347 0.004
R1223 S.t10 S.n335 0.004
R1224 S.t10 S.n317 0.004
R1225 S.t10 S.n358 0.004
R1226 S.t34 S.n108 0.004
R1227 S.t66 S.n1196 0.004
R1228 S.t66 S.n1162 0.004
R1229 S.t66 S.n1172 0.004
R1230 S.t66 S.n1180 0.004
R1231 S.t66 S.n1150 0.004
R1232 S.t10 S.n342 0.004
R1233 S.t66 S.n1154 0.004
R1234 S.t90 S.n494 0.004
R1235 S.t26 S.n1105 0.004
R1236 S.t10 S.n355 0.004
R1237 S.t10 S.n339 0.004
R1238 S.t10 S.n304 0.004
R1239 S.n740 S.n739 0.004
R1240 S.n1344 S.n1343 0.004
R1241 S.n956 S.n955 0.003
R1242 S.n1100 S.n1099 0.003
R1243 S.n1392 S.n1391 0.003
R1244 S.n1459 S.n1458 0.003
R1245 S.n205 S.n204 0.003
R1246 S.n461 S.n460 0.003
R1247 S.n1082 S.n1081 0.003
R1248 S.n1368 S.n1367 0.003
R1249 S.n1255 S.n1254 0.003
R1250 S.n784 S.n783 0.003
R1251 S.n699 S.n698 0.003
R1252 S.n561 S.n560 0.003
R1253 S.n189 S.n188 0.003
R1254 S.n46 S.n45 0.003
R1255 S.n485 S.n484 0.003
R1256 S.n130 S.n129 0.003
R1257 S.n150 S.n149 0.003
R1258 S.n418 S.n417 0.003
R1259 S.n717 S.n716 0.003
R1260 S.n268 S.n267 0.003
R1261 S.n168 S.n167 0.003
R1262 S.n438 S.n437 0.003
R1263 S.n544 S.n543 0.003
R1264 S.n665 S.n664 0.003
R1265 S.n765 S.n764 0.003
R1266 S.n1277 S.n1276 0.003
R1267 S.n67 S.n66 0.003
R1268 S.n230 S.n229 0.003
R1269 S.n260 S.n259 0.003
R1270 S.n183 S.n182 0.003
R1271 S.n605 S.n604 0.003
R1272 S.n583 S.n582 0.003
R1273 S.n853 S.n852 0.003
R1274 S.n826 S.n825 0.003
R1275 S.n1297 S.n1296 0.003
R1276 S.n1407 S.n1406 0.003
R1277 S.n1054 S.n1053 0.003
R1278 S.n1024 S.n1023 0.003
R1279 S.n611 S.n610 0.003
R1280 S.n575 S.n574 0.003
R1281 S.n868 S.n867 0.003
R1282 S.n919 S.n918 0.003
R1283 S.n931 S.n930 0.003
R1284 S.n1422 S.n1421 0.003
R1285 S.n1313 S.n1312 0.003
R1286 S.n797 S.n796 0.003
R1287 S.n876 S.n875 0.003
R1288 S.n820 S.n819 0.003
R1289 S.n1453 S.n1452 0.003
R1290 S.n995 S.n994 0.003
R1291 S.n900 S.n899 0.003
R1292 S.n1428 S.n1427 0.003
R1293 S.n1018 S.n1017 0.003
R1294 S.n953 S.n948 0.003
R1295 S.n1097 S.n1092 0.003
R1296 S.n1386 S.n1374 0.003
R1297 S.n199 S.n77 0.003
R1298 S.n455 S.n446 0.003
R1299 S.n1076 S.n1064 0.003
R1300 S.n1362 S.n1357 0.003
R1301 S.n1249 S.n1240 0.003
R1302 S.n778 S.n773 0.003
R1303 S.n693 S.n682 0.003
R1304 S.n555 S.n552 0.003
R1305 S.n196 S.n88 0.003
R1306 S.n40 S.n18 0.003
R1307 S.n482 S.n473 0.003
R1308 S.n124 S.n115 0.003
R1309 S.n144 S.n142 0.003
R1310 S.n412 S.n400 0.003
R1311 S.n714 S.n703 0.003
R1312 S.n275 S.n271 0.003
R1313 S.n162 S.n160 0.003
R1314 S.n432 S.n427 0.003
R1315 S.n538 S.n531 0.003
R1316 S.n659 S.n653 0.003
R1317 S.n759 S.n751 0.003
R1318 S.n1274 S.n1269 0.003
R1319 S.n61 S.n51 0.003
R1320 S.n227 S.n217 0.003
R1321 S.n180 S.n173 0.003
R1322 S.n602 S.n597 0.003
R1323 S.n593 S.n492 0.003
R1324 S.n850 S.n841 0.003
R1325 S.n836 S.n724 0.003
R1326 S.n1294 S.n1285 0.003
R1327 S.n1404 S.n1397 0.003
R1328 S.n1048 S.n1039 0.003
R1329 S.n1034 S.n935 0.003
R1330 S.n572 S.n567 0.003
R1331 S.n865 S.n864 0.003
R1332 S.n923 S.n922 0.003
R1333 S.n925 S.n908 0.003
R1334 S.n1419 S.n1418 0.003
R1335 S.n1310 S.n1308 0.003
R1336 S.n794 S.n793 0.003
R1337 S.n817 S.n803 0.003
R1338 S.n1450 S.n1444 0.003
R1339 S.n992 S.n987 0.003
R1340 S.n894 S.n889 0.003
R1341 S.n1436 S.n1325 0.003
R1342 S.n1015 S.n1010 0.003
R1343 S.n257 S.n249 0.003
R1344 S.n349 S.n347 0.003
R1345 S.n1210 S.n1209 0.003
R1346 S.n1210 S.n1122 0.003
R1347 S.n740 S.n738 0.003
R1348 S.n28 S.n27 0.003
R1349 S.n1436 S.n1321 0.003
R1350 S.n412 S.n411 0.003
R1351 S.n1120 S.n1119 0.003
R1352 S.t90 S.n503 0.003
R1353 S.t66 S.n1124 0.003
R1354 S.n981 S.n965 0.003
R1355 S.n1265 S.n1264 0.003
R1356 S.n1097 S.n1088 0.003
R1357 S.t66 S.n1147 0.003
R1358 S.t66 S.n1182 0.003
R1359 S.n476 S.n475 0.003
R1360 S.n73 S.n72 0.003
R1361 S.n370 S.n369 0.003
R1362 S.n276 S.n275 0.002
R1363 S.n144 S.n131 0.002
R1364 S.n412 S.n393 0.002
R1365 S.t90 S.n498 0.002
R1366 S.n759 S.n748 0.002
R1367 S.n659 S.n650 0.002
R1368 S.n538 S.n528 0.002
R1369 S.n432 S.n424 0.002
R1370 S.n162 S.n151 0.002
R1371 S.n1034 S.n932 0.002
R1372 S.n1048 S.n1036 0.002
R1373 S.n1404 S.n1394 0.002
R1374 S.n1294 S.n1282 0.002
R1375 S.n836 S.n721 0.002
R1376 S.n850 S.n838 0.002
R1377 S.n593 S.n489 0.002
R1378 S.n602 S.n594 0.002
R1379 S.n923 S.n909 0.002
R1380 S.n925 S.n901 0.002
R1381 S.n1419 S.n1411 0.002
R1382 S.n1310 S.n1301 0.002
R1383 S.n794 S.n786 0.002
R1384 S.n865 S.n857 0.002
R1385 S.n572 S.n564 0.002
R1386 S.n1436 S.n1322 0.002
R1387 S.n894 S.n886 0.002
R1388 S.n992 S.n984 0.002
R1389 S.n817 S.n807 0.002
R1390 S.n1450 S.n1441 0.002
R1391 S.n1386 S.n1371 0.002
R1392 S.n1097 S.n1089 0.002
R1393 S.n953 S.n945 0.002
R1394 S.n714 S.n707 0.002
R1395 S.n1274 S.n1266 0.002
R1396 S.n37 S.n36 0.002
R1397 S.n1001 S.n1000 0.002
R1398 S.n939 S.n938 0.002
R1399 S.n1141 S.n1140 0.002
R1400 S.n1144 S.n1143 0.002
R1401 S.t10 S.n333 0.002
R1402 S.n602 S.n601 0.002
R1403 S.n1070 S.n1069 0.002
R1404 S.n455 S.n440 0.002
R1405 S.n865 S.n858 0.002
R1406 S.n1436 S.n1435 0.002
R1407 S.n894 S.n893 0.002
R1408 S.n992 S.n991 0.002
R1409 S.n1386 S.n1385 0.002
R1410 S.n1097 S.n1096 0.002
R1411 S.n953 S.n952 0.002
R1412 S.n1362 S.n1351 0.002
R1413 S.n1249 S.n1234 0.002
R1414 S.n778 S.n767 0.002
R1415 S.n693 S.n676 0.002
R1416 S.n555 S.n546 0.002
R1417 S.n197 S.n196 0.002
R1418 S.n923 S.n910 0.002
R1419 S.n925 S.n902 0.002
R1420 S.n1419 S.n1412 0.002
R1421 S.n1310 S.n1302 0.002
R1422 S.n794 S.n787 0.002
R1423 S.n572 S.n571 0.002
R1424 S.n1450 S.n1449 0.002
R1425 S.n1015 S.n1014 0.002
R1426 S.n61 S.n60 0.002
R1427 S.n817 S.n813 0.002
R1428 S.n275 S.n274 0.002
R1429 S.n294 S.n291 0.002
R1430 S.t66 S.n1135 0.002
R1431 S.t66 S.n1192 0.002
R1432 S.n621 S.n620 0.002
R1433 S.n1076 S.n1058 0.002
R1434 S.n298 S.n297 0.002
R1435 S.n714 S.n713 0.002
R1436 S.n412 S.n394 0.002
R1437 S.n1274 S.n1273 0.002
R1438 S.n659 S.n658 0.002
R1439 S.n432 S.n431 0.002
R1440 S.n992 S.n983 0.002
R1441 S.n180 S.n170 0.002
R1442 S.n837 S.n836 0.002
R1443 S.n1035 S.n1034 0.002
R1444 S.n572 S.n563 0.002
R1445 S.n924 S.n923 0.002
R1446 S.n144 S.n143 0.002
R1447 S.t90 S.n497 0.002
R1448 S.n1199 S.n1198 0.002
R1449 S.n1076 S.n1057 0.002
R1450 S.n1362 S.n1350 0.002
R1451 S.n1249 S.n1224 0.002
R1452 S.n778 S.n766 0.002
R1453 S.n693 S.n666 0.002
R1454 S.n555 S.n545 0.002
R1455 S.n455 S.n439 0.002
R1456 S.n196 S.n81 0.002
R1457 S.n199 S.n74 0.002
R1458 S.n482 S.n463 0.002
R1459 S.n124 S.n111 0.002
R1460 S.n40 S.n15 0.002
R1461 S.n1015 S.n1007 0.002
R1462 S.n1210 S.n1197 0.002
R1463 S.n329 S.n326 0.002
R1464 S.n299 S.n298 0.001
R1465 S.n1146 S.n1142 0.001
R1466 S.n1146 S.n1145 0.001
R1467 S.t10 S.n299 0.001
R1468 S.n649 S.n648 0.001
R1469 S.n423 S.n422 0.001
R1470 S.n1197 S.t66 0.001
R1471 S.n628 S.n627 0.001
R1472 S.n1205 S.n1199 0.001
R1473 S.n1476 S.n1475 0.001
R1474 S.n224 S.n223 0.001
R1475 S.n452 S.n451 0.001
R1476 S.n554 S.n553 0.001
R1477 S.n690 S.n689 0.001
R1478 S.n775 S.n774 0.001
R1479 S.n1246 S.n1245 0.001
R1480 S.n1359 S.n1358 0.001
R1481 S.n85 S.n84 0.001
R1482 S.n100 S.n99 0.001
R1483 S.n515 S.n514 0.001
R1484 S.n735 S.n734 0.001
R1485 S.n1339 S.n1338 0.001
R1486 S.t10 S.n277 0.001
R1487 S.n374 S.t10 0.001
R1488 S.t10 S.n307 0.001
R1489 S.t10 S.n325 0.001
R1490 S.t10 S.n351 0.001
R1491 S.n295 S.n294 0.001
R1492 S.n982 S.n981 0.001
R1493 S.n521 S.n520 0.001
R1494 S.n741 S.n740 0.001
R1495 S.n1345 S.n1344 0.001
R1496 S.n106 S.n105 0.001
R1497 S.n1120 S.n1106 0.001
R1498 S.n294 S.n293 0.001
R1499 S.n482 S.n465 0.001
R1500 S.n23 S.n22 0.001
R1501 S.n1034 S.n1033 0.001
R1502 S.n1048 S.n1047 0.001
R1503 S.n1404 S.n1403 0.001
R1504 S.n1294 S.n1293 0.001
R1505 S.n836 S.n835 0.001
R1506 S.n850 S.n849 0.001
R1507 S.n593 S.n592 0.001
R1508 S.n1005 S.n1004 0.001
R1509 S.n943 S.n942 0.001
R1510 S.n98 S.n97 0.001
R1511 S.n513 S.n512 0.001
R1512 S.n733 S.n732 0.001
R1513 S.n1337 S.n1336 0.001
R1514 S.n975 S.n974 0.001
R1515 S.n1106 S.t26 0.001
R1516 S.t64 S.n982 0.001
R1517 S.t90 S.n521 0.001
R1518 S.t4 S.n741 0.001
R1519 S.t97 S.n1345 0.001
R1520 S.t34 S.n106 0.001
R1521 S.n977 S.n971 0.001
R1522 S.n1146 S.n1139 0.001
R1523 S.n99 S.n98 0.001
R1524 S.n514 S.n513 0.001
R1525 S.n734 S.n733 0.001
R1526 S.n1338 S.n1337 0.001
R1527 S.n1370 S.n1369 0.001
R1528 S.n124 S.n112 0.001
R1529 S.n6 S.n5 0.001
R1530 S.n243 S.n242 0.001
R1531 S.n385 S.n384 0.001
R1532 S.n637 S.n636 0.001
R1533 S.n1218 S.n1217 0.001
R1534 S.n1113 S.n1112 0.001
R1535 S.n294 S.n290 0.001
R1536 S.n948 S.n947 0.001
R1537 S.n1092 S.n1091 0.001
R1538 S.n1374 S.n1373 0.001
R1539 S.n77 S.n76 0.001
R1540 S.n446 S.n445 0.001
R1541 S.n1064 S.n1063 0.001
R1542 S.n1357 S.n1356 0.001
R1543 S.n1240 S.n1239 0.001
R1544 S.n773 S.n772 0.001
R1545 S.n682 S.n681 0.001
R1546 S.n552 S.n551 0.001
R1547 S.n88 S.n87 0.001
R1548 S.n18 S.n17 0.001
R1549 S.n473 S.n472 0.001
R1550 S.n115 S.n114 0.001
R1551 S.n142 S.n141 0.001
R1552 S.n400 S.n399 0.001
R1553 S.n703 S.n702 0.001
R1554 S.n271 S.n270 0.001
R1555 S.n160 S.n159 0.001
R1556 S.n427 S.n426 0.001
R1557 S.n531 S.n530 0.001
R1558 S.n653 S.n652 0.001
R1559 S.n751 S.n750 0.001
R1560 S.n1269 S.n1268 0.001
R1561 S.n51 S.n50 0.001
R1562 S.n217 S.n216 0.001
R1563 S.n173 S.n172 0.001
R1564 S.n597 S.n596 0.001
R1565 S.n492 S.n491 0.001
R1566 S.n841 S.n840 0.001
R1567 S.n724 S.n723 0.001
R1568 S.n1285 S.n1284 0.001
R1569 S.n1397 S.n1396 0.001
R1570 S.n1039 S.n1038 0.001
R1571 S.n935 S.n934 0.001
R1572 S.n567 S.n566 0.001
R1573 S.n864 S.n863 0.001
R1574 S.n922 S.n921 0.001
R1575 S.n908 S.n907 0.001
R1576 S.n1418 S.n1417 0.001
R1577 S.n1308 S.n1307 0.001
R1578 S.n793 S.n792 0.001
R1579 S.n803 S.n802 0.001
R1580 S.n1444 S.n1443 0.001
R1581 S.n987 S.n986 0.001
R1582 S.n889 S.n888 0.001
R1583 S.n1325 S.n1324 0.001
R1584 S.n1010 S.n1009 0.001
R1585 S.n1142 S.n1141 0.001
R1586 S.n1145 S.n1144 0.001
R1587 S.n979 S.n978 0.001
R1588 S.n1341 S.n1340 0.001
R1589 S.n737 S.n736 0.001
R1590 S.n517 S.n516 0.001
R1591 S.n102 S.n101 0.001
R1592 S.n294 S.n292 0.001
R1593 S.t64 S.n956 0.001
R1594 S.t64 S.n959 0.001
R1595 S.t26 S.n1100 0.001
R1596 S.t26 S.n1103 0.001
R1597 S.t97 S.n1392 0.001
R1598 S.t97 S.n1389 0.001
R1599 S.n1389 S.n1386 0.001
R1600 S.n1459 S.t76 0.001
R1601 S.n1479 S.n1461 0.001
R1602 S.t54 S.n205 0.001
R1603 S.t54 S.n202 0.001
R1604 S.n202 S.n199 0.001
R1605 S.t19 S.n461 0.001
R1606 S.t19 S.n458 0.001
R1607 S.n458 S.n455 0.001
R1608 S.t26 S.n1082 0.001
R1609 S.t26 S.n1079 0.001
R1610 S.n1079 S.n1076 0.001
R1611 S.t97 S.n1368 0.001
R1612 S.t97 S.n1365 0.001
R1613 S.n1365 S.n1362 0.001
R1614 S.t76 S.n1255 0.001
R1615 S.t76 S.n1252 0.001
R1616 S.n1252 S.n1249 0.001
R1617 S.t4 S.n784 0.001
R1618 S.t4 S.n781 0.001
R1619 S.n781 S.n778 0.001
R1620 S.t78 S.n699 0.001
R1621 S.t78 S.n696 0.001
R1622 S.n696 S.n693 0.001
R1623 S.t90 S.n561 0.001
R1624 S.t90 S.n558 0.001
R1625 S.n558 S.n555 0.001
R1626 S.n189 S.t34 0.001
R1627 S.n196 S.n192 0.001
R1628 S.t54 S.n46 0.001
R1629 S.t54 S.n43 0.001
R1630 S.n43 S.n40 0.001
R1631 S.t19 S.n485 0.001
R1632 S.t19 S.n488 0.001
R1633 S.t34 S.n130 0.001
R1634 S.t34 S.n127 0.001
R1635 S.n127 S.n124 0.001
R1636 S.t34 S.n150 0.001
R1637 S.t34 S.n147 0.001
R1638 S.n147 S.n144 0.001
R1639 S.t19 S.n418 0.001
R1640 S.t19 S.n415 0.001
R1641 S.n415 S.n412 0.001
R1642 S.t78 S.n717 0.001
R1643 S.t78 S.n720 0.001
R1644 S.n265 S.t54 0.001
R1645 S.n275 S.n265 0.001
R1646 S.t34 S.n168 0.001
R1647 S.t34 S.n165 0.001
R1648 S.n165 S.n162 0.001
R1649 S.t19 S.n438 0.001
R1650 S.t19 S.n435 0.001
R1651 S.n435 S.n432 0.001
R1652 S.t90 S.n544 0.001
R1653 S.t90 S.n541 0.001
R1654 S.n541 S.n538 0.001
R1655 S.t78 S.n665 0.001
R1656 S.t78 S.n662 0.001
R1657 S.n662 S.n659 0.001
R1658 S.t4 S.n765 0.001
R1659 S.t4 S.n762 0.001
R1660 S.n762 S.n759 0.001
R1661 S.t76 S.n1277 0.001
R1662 S.t76 S.n1280 0.001
R1663 S.t54 S.n67 0.001
R1664 S.t54 S.n64 0.001
R1665 S.n64 S.n61 0.001
R1666 S.t54 S.n230 0.001
R1667 S.t54 S.n233 0.001
R1668 S.t54 S.n260 0.001
R1669 S.t54 S.n262 0.001
R1670 S.t34 S.n183 0.001
R1671 S.t34 S.n186 0.001
R1672 S.t19 S.n605 0.001
R1673 S.t19 S.n608 0.001
R1674 S.n583 S.t90 0.001
R1675 S.n593 S.n586 0.001
R1676 S.t78 S.n853 0.001
R1677 S.t78 S.n856 0.001
R1678 S.n826 S.t4 0.001
R1679 S.n836 S.n829 0.001
R1680 S.t76 S.n1297 0.001
R1681 S.t76 S.n1300 0.001
R1682 S.t97 S.n1407 0.001
R1683 S.t97 S.n1410 0.001
R1684 S.t26 S.n1054 0.001
R1685 S.t26 S.n1051 0.001
R1686 S.n1051 S.n1048 0.001
R1687 S.n1024 S.t64 0.001
R1688 S.n1034 S.n1027 0.001
R1689 S.n1033 S.n1032 0.001
R1690 S.n1047 S.n1046 0.001
R1691 S.n1403 S.n1402 0.001
R1692 S.n1293 S.n1292 0.001
R1693 S.n835 S.n834 0.001
R1694 S.n849 S.n848 0.001
R1695 S.n592 S.n591 0.001
R1696 S.n611 S.t19 0.001
R1697 S.n620 S.n613 0.001
R1698 S.t90 S.n575 0.001
R1699 S.t90 S.n578 0.001
R1700 S.t78 S.n868 0.001
R1701 S.t78 S.n871 0.001
R1702 S.n923 S.n916 0.001
R1703 S.t26 S.n931 0.001
R1704 S.t26 S.n928 0.001
R1705 S.n928 S.n925 0.001
R1706 S.t97 S.n1422 0.001
R1707 S.t97 S.n1425 0.001
R1708 S.t76 S.n1313 0.001
R1709 S.t76 S.n1316 0.001
R1710 S.t4 S.n797 0.001
R1711 S.t4 S.n800 0.001
R1712 S.n873 S.t78 0.001
R1713 S.n881 S.n873 0.001
R1714 S.t4 S.n820 0.001
R1715 S.t4 S.n823 0.001
R1716 S.t76 S.n1453 0.001
R1717 S.t76 S.n1456 0.001
R1718 S.t64 S.n995 0.001
R1719 S.t64 S.n998 0.001
R1720 S.t26 S.n900 0.001
R1721 S.t26 S.n897 0.001
R1722 S.n897 S.n894 0.001
R1723 S.n1428 S.t97 0.001
R1724 S.n1436 S.n1431 0.001
R1725 S.n285 S.n284 0.001
R1726 S.n289 S.n288 0.001
R1727 S.n1118 S.n1116 0.001
R1728 S.n1222 S.n1221 0.001
R1729 S.n248 S.n247 0.001
R1730 S.n389 S.n388 0.001
R1731 S.n641 S.n640 0.001
R1732 S.n1208 S.n1207 0.001
R1733 S.n1146 S.n1137 0.001
R1734 S.n976 S.n975 0.001
R1735 S.n1204 S.n1203 0.001
R1736 S.n956 S.n953 0.001
R1737 S.n1100 S.n1097 0.001
R1738 S.n1479 S.n1459 0.001
R1739 S.n196 S.n189 0.001
R1740 S.n1277 S.n1274 0.001
R1741 S.n717 S.n714 0.001
R1742 S.n275 S.n268 0.001
R1743 S.n485 S.n482 0.001
R1744 S.n230 S.n227 0.001
R1745 S.n260 S.n257 0.001
R1746 S.n1034 S.n1024 0.001
R1747 S.n1407 S.n1404 0.001
R1748 S.n1297 S.n1294 0.001
R1749 S.n836 S.n826 0.001
R1750 S.n853 S.n850 0.001
R1751 S.n593 S.n583 0.001
R1752 S.n605 S.n602 0.001
R1753 S.n183 S.n180 0.001
R1754 S.n620 S.n611 0.001
R1755 S.n923 S.n919 0.001
R1756 S.n1422 S.n1419 0.001
R1757 S.n1313 S.n1310 0.001
R1758 S.n797 S.n794 0.001
R1759 S.n868 S.n865 0.001
R1760 S.n575 S.n572 0.001
R1761 S.n881 S.n876 0.001
R1762 S.n820 S.n817 0.001
R1763 S.n1453 S.n1450 0.001
R1764 S.n1436 S.n1428 0.001
R1765 S.n995 S.n992 0.001
R1766 S.n977 S.n976 0.001
R1767 S.n1204 S.n1202 0.001
R1768 S.t64 S.n1018 0.001
R1769 S.t64 S.n1021 0.001
R1770 S.n1018 S.n1015 0.001
C0 S G 1532.33fF
C1 D S 372.66fF
C2 D G 464.98fF
C3 D PW 250.67fF
C4 G PW -177.02fF
C5 S PW 296.86fF
C6 S.n0 PW 0.39fF
C7 S.n1 PW 0.18fF
C8 S.n2 PW 0.26fF
C9 S.n3 PW 0.09fF
C10 S.n4 PW 0.65fF
C11 S.n5 PW 0.36fF
C12 S.n6 PW 0.27fF
C13 S.t58 PW 0.02fF
C14 S.n7 PW 0.25fF
C15 S.n8 PW 0.37fF
C16 S.n9 PW 0.63fF
C17 S.n10 PW 0.67fF
C18 S.n11 PW 0.45fF
C19 S.n12 PW 1.74fF
C20 S.n13 PW 0.49fF
C21 S.n14 PW 0.47fF
C22 S.n15 PW 1.90fF
C23 S.n16 PW 0.12fF
C24 S.t257 PW 0.02fF
C25 S.n17 PW 0.14fF
C26 S.t155 PW 0.02fF
C27 S.n19 PW 0.25fF
C28 S.n20 PW 0.37fF
C29 S.n21 PW 0.63fF
C30 S.n22 PW 0.05fF
C31 S.n23 PW 0.18fF
C32 S.n24 PW 1.63fF
C33 S.n25 PW 0.02fF
C34 S.n26 PW 0.12fF
C35 S.n27 PW 0.19fF
C36 S.n28 PW 0.12fF
C37 S.n29 PW 0.26fF
C38 S.n30 PW 0.82fF
C39 S.n31 PW 0.03fF
C40 S.n32 PW 0.02fF
C41 S.n33 PW 0.01fF
C42 S.n34 PW 0.02fF
C43 S.n35 PW 0.03fF
C44 S.n36 PW 0.10fF
C45 S.n37 PW 0.07fF
C46 S.n38 PW 0.26fF
C47 S.n39 PW 0.12fF
C48 S.n40 PW 2.00fF
C49 S.t47 PW 0.02fF
C50 S.n41 PW 0.25fF
C51 S.n42 PW 0.94fF
C52 S.n43 PW 0.05fF
C53 S.t270 PW 0.02fF
C54 S.n44 PW 0.12fF
C55 S.n45 PW 0.15fF
C56 S.n47 PW 0.26fF
C57 S.n48 PW 0.09fF
C58 S.n49 PW 0.12fF
C59 S.t72 PW 0.02fF
C60 S.n50 PW 0.14fF
C61 S.t230 PW 0.02fF
C62 S.n52 PW 0.25fF
C63 S.n53 PW 0.37fF
C64 S.n54 PW 0.63fF
C65 S.n55 PW 0.66fF
C66 S.n56 PW 0.38fF
C67 S.n57 PW 0.26fF
C68 S.n58 PW 0.23fF
C69 S.n59 PW 0.62fF
C70 S.n60 PW 0.28fF
C71 S.n61 PW 2.00fF
C72 S.t139 PW 0.02fF
C73 S.n62 PW 0.25fF
C74 S.n63 PW 0.94fF
C75 S.n64 PW 0.05fF
C76 S.t82 PW 0.02fF
C77 S.n65 PW 0.12fF
C78 S.n66 PW 0.15fF
C79 S.n68 PW 0.19fF
C80 S.n69 PW 0.10fF
C81 S.n70 PW 0.70fF
C82 S.n71 PW 0.29fF
C83 S.n72 PW 1.79fF
C84 S.n73 PW 0.22fF
C85 S.n74 PW 1.90fF
C86 S.n75 PW 0.12fF
C87 S.t55 PW 0.02fF
C88 S.n76 PW 0.14fF
C89 S.t131 PW 0.02fF
C90 S.n78 PW 0.25fF
C91 S.n79 PW 0.37fF
C92 S.n80 PW 0.63fF
C93 S.n81 PW 1.95fF
C94 S.n82 PW 0.26fF
C95 S.n83 PW 0.09fF
C96 S.n84 PW 1.19fF
C97 S.n85 PW 0.23fF
C98 S.n86 PW 0.12fF
C99 S.t99 PW 0.02fF
C100 S.n87 PW 0.14fF
C101 S.t129 PW 0.02fF
C102 S.n89 PW 1.25fF
C103 S.n90 PW 0.62fF
C104 S.n91 PW 0.37fF
C105 S.n92 PW 0.65fF
C106 S.n93 PW 1.16fF
C107 S.n94 PW 1.42fF
C108 S.n95 PW 0.61fF
C109 S.n96 PW 0.02fF
C110 S.n97 PW 1.00fF
C111 S.t2 PW 8.19fF
C112 S.n98 PW 9.08fF
C113 S.n100 PW 0.39fF
C114 S.n101 PW 0.24fF
C115 S.n102 PW 2.98fF
C116 S.n103 PW 2.53fF
C117 S.n104 PW 2.37fF
C118 S.n105 PW 4.42fF
C119 S.n106 PW 0.26fF
C120 S.n107 PW 0.01fF
C121 S.t201 PW 0.02fF
C122 S.n108 PW 0.26fF
C123 S.t43 PW 0.02fF
C124 S.n109 PW 0.98fF
C125 S.n110 PW 0.73fF
C126 S.n111 PW 1.95fF
C127 S.n112 PW 2.02fF
C128 S.n113 PW 0.12fF
C129 S.t112 PW 0.02fF
C130 S.n114 PW 0.14fF
C131 S.t17 PW 0.02fF
C132 S.n116 PW 0.25fF
C133 S.n117 PW 0.37fF
C134 S.n118 PW 0.63fF
C135 S.n119 PW 0.01fF
C136 S.n120 PW 0.03fF
C137 S.n121 PW 0.02fF
C138 S.n122 PW 0.64fF
C139 S.n123 PW 0.88fF
C140 S.n124 PW 2.70fF
C141 S.t218 PW 0.02fF
C142 S.n125 PW 0.25fF
C143 S.n126 PW 0.94fF
C144 S.n127 PW 0.05fF
C145 S.t196 PW 0.02fF
C146 S.n128 PW 0.12fF
C147 S.n129 PW 0.15fF
C148 S.n131 PW 1.94fF
C149 S.n132 PW 0.42fF
C150 S.n133 PW 0.36fF
C151 S.n134 PW 0.93fF
C152 S.n135 PW 0.81fF
C153 S.n136 PW 1.00fF
C154 S.t205 PW 0.02fF
C155 S.n137 PW 0.25fF
C156 S.n138 PW 0.37fF
C157 S.n139 PW 0.63fF
C158 S.n140 PW 0.12fF
C159 S.t284 PW 0.02fF
C160 S.n141 PW 0.14fF
C161 S.n143 PW 2.69fF
C162 S.n144 PW 2.23fF
C163 S.t135 PW 0.02fF
C164 S.n145 PW 0.25fF
C165 S.n146 PW 0.94fF
C166 S.n147 PW 0.05fF
C167 S.t102 PW 0.02fF
C168 S.n148 PW 0.12fF
C169 S.n149 PW 0.15fF
C170 S.n151 PW 1.94fF
C171 S.n152 PW 0.73fF
C172 S.n153 PW 0.36fF
C173 S.n154 PW 1.28fF
C174 S.t118 PW 0.02fF
C175 S.n155 PW 0.25fF
C176 S.n156 PW 0.37fF
C177 S.n157 PW 0.63fF
C178 S.n158 PW 0.12fF
C179 S.t192 PW 0.02fF
C180 S.n159 PW 0.14fF
C181 S.n161 PW 2.37fF
C182 S.n162 PW 2.09fF
C183 S.t30 PW 0.02fF
C184 S.n163 PW 0.25fF
C185 S.n164 PW 0.94fF
C186 S.n165 PW 0.05fF
C187 S.t268 PW 0.02fF
C188 S.n166 PW 0.12fF
C189 S.n167 PW 0.15fF
C190 S.n169 PW 7.96fF
C191 S.n170 PW 2.81fF
C192 S.n171 PW 0.12fF
C193 S.t35 PW 0.02fF
C194 S.n172 PW 0.14fF
C195 S.t167 PW 0.02fF
C196 S.n174 PW 0.25fF
C197 S.n175 PW 0.37fF
C198 S.n176 PW 0.63fF
C199 S.n177 PW 1.61fF
C200 S.n178 PW 0.73fF
C201 S.n179 PW 0.29fF
C202 S.n180 PW 2.17fF
C203 S.t123 PW 0.02fF
C204 S.n181 PW 0.12fF
C205 S.n182 PW 0.15fF
C206 S.t273 PW 0.02fF
C207 S.n184 PW 0.25fF
C208 S.n185 PW 0.94fF
C209 S.n186 PW 0.05fF
C210 S.t34 PW 17.65fF
C211 S.t178 PW 0.02fF
C212 S.n187 PW 0.12fF
C213 S.n188 PW 0.15fF
C214 S.t211 PW 0.02fF
C215 S.n190 PW 0.25fF
C216 S.n191 PW 0.94fF
C217 S.n192 PW 0.05fF
C218 S.t3 PW 0.02fF
C219 S.n193 PW 0.25fF
C220 S.n194 PW 0.37fF
C221 S.n195 PW 0.63fF
C222 S.n196 PW 1.94fF
C223 S.n197 PW 2.82fF
C224 S.n198 PW 2.57fF
C225 S.n199 PW 1.92fF
C226 S.t61 PW 0.02fF
C227 S.n200 PW 0.25fF
C228 S.n201 PW 0.94fF
C229 S.n202 PW 0.05fF
C230 S.t256 PW 0.02fF
C231 S.n203 PW 0.12fF
C232 S.n204 PW 0.15fF
C233 S.n206 PW 7.96fF
C234 S.n207 PW 0.21fF
C235 S.n208 PW 0.21fF
C236 S.n209 PW 0.07fF
C237 S.n210 PW 0.09fF
C238 S.n211 PW 0.10fF
C239 S.n212 PW 0.26fF
C240 S.n213 PW 0.21fF
C241 S.n214 PW 0.46fF
C242 S.n215 PW 0.12fF
C243 S.t84 PW 0.02fF
C244 S.n216 PW 0.14fF
C245 S.t238 PW 0.02fF
C246 S.n218 PW 0.25fF
C247 S.n219 PW 0.37fF
C248 S.n220 PW 0.63fF
C249 S.n221 PW 0.81fF
C250 S.n222 PW 0.21fF
C251 S.n223 PW 1.27fF
C252 S.n224 PW 0.46fF
C253 S.n225 PW 0.26fF
C254 S.n226 PW 0.09fF
C255 S.n227 PW 1.87fF
C256 S.t104 PW 0.02fF
C257 S.n228 PW 0.12fF
C258 S.n229 PW 0.15fF
C259 S.t149 PW 0.02fF
C260 S.n231 PW 0.25fF
C261 S.n232 PW 0.94fF
C262 S.n233 PW 0.05fF
C263 S.n234 PW 1.17fF
C264 S.n235 PW 9.26fF
C265 S.n236 PW 21.01fF
C266 S.n237 PW 9.26fF
C267 S.n238 PW 21.01fF
C268 S.n239 PW 0.62fF
C269 S.n240 PW 0.24fF
C270 S.n241 PW 0.91fF
C271 S.n242 PW 1.83fF
C272 S.n243 PW 0.30fF
C273 S.t29 PW 8.19fF
C274 S.n244 PW 10.54fF
C275 S.n245 PW 0.91fF
C276 S.n246 PW 0.27fF
C277 S.n247 PW 1.40fF
C278 S.n248 PW 4.38fF
C279 S.n249 PW 1.86fF
C280 S.t235 PW 0.02fF
C281 S.n250 PW 0.66fF
C282 S.n251 PW 0.63fF
C283 S.n252 PW 1.24fF
C284 S.n253 PW 0.38fF
C285 S.n254 PW 1.22fF
C286 S.n255 PW 0.40fF
C287 S.n256 PW 2.01fF
C288 S.n257 PW 4.35fF
C289 S.t240 PW 0.02fF
C290 S.n258 PW 0.01fF
C291 S.n259 PW 0.26fF
C292 S.t148 PW 0.02fF
C293 S.n261 PW 1.23fF
C294 S.n262 PW 0.05fF
C295 S.t54 PW 17.26fF
C296 S.t222 PW 0.02fF
C297 S.n263 PW 0.25fF
C298 S.n264 PW 0.94fF
C299 S.n265 PW 0.05fF
C300 S.t181 PW 0.02fF
C301 S.n266 PW 0.12fF
C302 S.n267 PW 0.15fF
C303 S.n269 PW 0.12fF
C304 S.t168 PW 0.02fF
C305 S.n270 PW 0.14fF
C306 S.n272 PW 0.04fF
C307 S.n273 PW 0.50fF
C308 S.n274 PW 0.39fF
C309 S.n275 PW 2.02fF
C310 S.n276 PW 1.54fF
C311 S.n277 PW 2.71fF
C312 S.n278 PW 0.38fF
C313 S.n279 PW 0.85fF
C314 S.n280 PW 1.17fF
C315 S.n282 PW 0.41fF
C316 S.t212 PW 0.02fF
C317 S.n283 PW 1.35fF
C318 S.n284 PW 25.16fF
C319 S.n285 PW 2.30fF
C320 S.n286 PW 0.37fF
C321 S.n287 PW 0.64fF
C322 S.n288 PW 0.54fF
C323 S.n289 PW 3.78fF
C324 S.n290 PW 4.38fF
C325 S.n291 PW 4.84fF
C326 S.n292 PW 4.44fF
C327 S.n293 PW 4.41fF
C328 S.n294 PW 44.75fF
C329 S.n295 PW 2.26fF
C330 S.n296 PW 13.34fF
C331 S.n297 PW 1.96fF
C332 S.n298 PW 9.70fF
C333 S.n299 PW 0.26fF
C334 S.t11 PW 0.02fF
C335 S.n300 PW 0.45fF
C336 S.n301 PW 9.26fF
C337 S.n302 PW 9.26fF
C338 S.n303 PW 5.48fF
C339 S.n304 PW 1.90fF
C340 S.t111 PW 0.02fF
C341 S.n305 PW 0.92fF
C342 S.t189 PW 0.02fF
C343 S.n306 PW 0.92fF
C344 S.n307 PW 3.37fF
C345 S.n308 PW 0.26fF
C346 S.n309 PW 0.26fF
C347 S.n310 PW 1.09fF
C348 S.n311 PW 0.36fF
C349 S.n312 PW 0.47fF
C350 S.n313 PW 0.02fF
C351 S.t14 PW 0.02fF
C352 S.n314 PW 0.38fF
C353 S.t280 PW 0.02fF
C354 S.n315 PW 0.92fF
C355 S.n316 PW 0.02fF
C356 S.t203 PW 0.02fF
C357 S.n317 PW 0.38fF
C358 S.t94 PW 0.02fF
C359 S.n318 PW 0.92fF
C360 S.n319 PW 0.14fF
C361 S.n320 PW 1.80fF
C362 S.n321 PW 1.67fF
C363 S.t188 PW 0.02fF
C364 S.n322 PW 0.92fF
C365 S.t265 PW 0.02fF
C366 S.n323 PW 0.92fF
C367 S.n324 PW 1.55fF
C368 S.n325 PW 2.71fF
C369 S.n326 PW 0.46fF
C370 S.n327 PW 0.81fF
C371 S.n328 PW 0.22fF
C372 S.n329 PW 1.79fF
C373 S.n330 PW 9.26fF
C374 S.n331 PW 9.26fF
C375 S.n332 PW 5.73fF
C376 S.n333 PW 1.56fF
C377 S.n334 PW 0.02fF
C378 S.t115 PW 0.02fF
C379 S.n335 PW 0.38fF
C380 S.n336 PW 21.45fF
C381 S.n337 PW 21.45fF
C382 S.n338 PW 6.01fF
C383 S.n339 PW 2.02fF
C384 S.t180 PW 0.02fF
C385 S.n340 PW 0.92fF
C386 S.t251 PW 0.02fF
C387 S.n341 PW 0.92fF
C388 S.n342 PW 1.67fF
C389 S.n343 PW 0.02fF
C390 S.t56 PW 0.02fF
C391 S.n344 PW 0.38fF
C392 S.t13 PW 9.21fF
C393 S.n345 PW 0.99fF
C394 S.n346 PW 0.96fF
C395 S.n347 PW 0.35fF
C396 S.n348 PW 0.44fF
C397 S.n349 PW 0.31fF
C398 S.n350 PW 2.02fF
C399 S.n351 PW 2.71fF
C400 S.n352 PW 14.04fF
C401 S.n353 PW 14.04fF
C402 S.n354 PW 5.53fF
C403 S.n355 PW 2.12fF
C404 S.t281 PW 0.02fF
C405 S.n356 PW 0.92fF
C406 S.n357 PW 0.02fF
C407 S.t124 PW 0.02fF
C408 S.n358 PW 0.38fF
C409 S.t200 PW 0.02fF
C410 S.n359 PW 0.92fF
C411 S.n360 PW 9.26fF
C412 S.n361 PW 9.26fF
C413 S.n362 PW 5.95fF
C414 S.n363 PW 0.11fF
C415 S.n364 PW 0.37fF
C416 S.n365 PW 0.39fF
C417 S.n366 PW 0.03fF
C418 S.n367 PW 0.03fF
C419 S.n368 PW 0.11fF
C420 S.n369 PW 0.12fF
C421 S.n370 PW 0.03fF
C422 S.n371 PW 0.07fF
C423 S.n372 PW 1.46fF
C424 S.n373 PW 1.82fF
C425 S.t10 PW 43.34fF
C426 S.n374 PW 3.37fF
C427 S.n375 PW 16.99fF
C428 S.n376 PW 9.74fF
C429 S.n377 PW 9.73fF
C430 S.n378 PW 9.74fF
C431 S.n379 PW 7.98fF
C432 S.n380 PW 0.25fF
C433 S.n381 PW 0.62fF
C434 S.n382 PW 0.24fF
C435 S.n383 PW 0.61fF
C436 S.n384 PW 1.83fF
C437 S.n385 PW 0.30fF
C438 S.t36 PW 8.19fF
C439 S.n386 PW 10.54fF
C440 S.n387 PW 0.79fF
C441 S.n388 PW 0.28fF
C442 S.n389 PW 4.13fF
C443 S.n390 PW 1.55fF
C444 S.n391 PW 1.35fF
C445 S.n392 PW 0.28fF
C446 S.n393 PW 1.94fF
C447 S.n394 PW 1.63fF
C448 S.t60 PW 0.02fF
C449 S.n395 PW 0.25fF
C450 S.n396 PW 0.37fF
C451 S.n397 PW 0.63fF
C452 S.n398 PW 0.12fF
C453 S.t260 PW 0.02fF
C454 S.n399 PW 0.14fF
C455 S.n401 PW 0.04fF
C456 S.n402 PW 0.11fF
C457 S.n403 PW 0.37fF
C458 S.n404 PW 0.39fF
C459 S.n405 PW 0.03fF
C460 S.n406 PW 0.03fF
C461 S.n407 PW 0.11fF
C462 S.n408 PW 0.12fF
C463 S.n409 PW 0.07fF
C464 S.n410 PW 0.12fF
C465 S.n411 PW 0.19fF
C466 S.n412 PW 4.16fF
C467 S.t226 PW 0.02fF
C468 S.n413 PW 0.25fF
C469 S.n414 PW 0.94fF
C470 S.n415 PW 0.05fF
C471 S.t271 PW 0.02fF
C472 S.n416 PW 0.12fF
C473 S.n417 PW 0.15fF
C474 S.n419 PW 0.26fF
C475 S.n420 PW 0.09fF
C476 S.n421 PW 0.21fF
C477 S.n422 PW 1.32fF
C478 S.n423 PW 0.55fF
C479 S.n424 PW 1.94fF
C480 S.n425 PW 0.12fF
C481 S.t170 PW 0.02fF
C482 S.n426 PW 0.14fF
C483 S.t233 PW 0.02fF
C484 S.n428 PW 0.25fF
C485 S.n429 PW 0.37fF
C486 S.n430 PW 0.63fF
C487 S.n431 PW 1.63fF
C488 S.n432 PW 2.53fF
C489 S.t141 PW 0.02fF
C490 S.n433 PW 0.25fF
C491 S.n434 PW 0.94fF
C492 S.n435 PW 0.05fF
C493 S.t182 PW 0.02fF
C494 S.n436 PW 0.12fF
C495 S.n437 PW 0.15fF
C496 S.n439 PW 1.95fF
C497 S.n440 PW 2.76fF
C498 S.t151 PW 0.02fF
C499 S.n441 PW 0.25fF
C500 S.n442 PW 0.37fF
C501 S.n443 PW 0.63fF
C502 S.n444 PW 0.12fF
C503 S.t73 PW 0.02fF
C504 S.n445 PW 0.14fF
C505 S.n447 PW 0.72fF
C506 S.n448 PW 0.23fF
C507 S.n449 PW 0.23fF
C508 S.n450 PW 0.72fF
C509 S.n451 PW 1.19fF
C510 S.n452 PW 0.23fF
C511 S.n453 PW 0.26fF
C512 S.n454 PW 0.09fF
C513 S.n455 PW 1.95fF
C514 S.t38 PW 0.02fF
C515 S.n456 PW 0.25fF
C516 S.n457 PW 0.94fF
C517 S.n458 PW 0.05fF
C518 S.t83 PW 0.02fF
C519 S.n459 PW 0.12fF
C520 S.n460 PW 0.15fF
C521 S.n462 PW 7.96fF
C522 S.n463 PW 1.77fF
C523 S.n464 PW 0.67fF
C524 S.n465 PW 0.71fF
C525 S.n466 PW 0.75fF
C526 S.n467 PW 0.38fF
C527 S.t157 PW 0.02fF
C528 S.n468 PW 0.25fF
C529 S.n469 PW 0.37fF
C530 S.n470 PW 0.63fF
C531 S.n471 PW 0.12fF
C532 S.t89 PW 0.02fF
C533 S.n472 PW 0.14fF
C534 S.n474 PW 0.29fF
C535 S.n475 PW 0.77fF
C536 S.n476 PW 0.62fF
C537 S.n477 PW 0.21fF
C538 S.n478 PW 0.21fF
C539 S.n479 PW 0.07fF
C540 S.n480 PW 0.09fF
C541 S.n481 PW 0.10fF
C542 S.n482 PW 1.73fF
C543 S.t105 PW 0.02fF
C544 S.n483 PW 0.12fF
C545 S.n484 PW 0.15fF
C546 S.t50 PW 0.02fF
C547 S.n486 PW 0.25fF
C548 S.n487 PW 0.94fF
C549 S.n488 PW 0.05fF
C550 S.n489 PW 1.94fF
C551 S.n490 PW 0.12fF
C552 S.t272 PW 0.02fF
C553 S.n491 PW 0.14fF
C554 S.n493 PW 0.12fF
C555 S.t286 PW 0.02fF
C556 S.n494 PW 0.14fF
C557 S.t140 PW 0.02fF
C558 S.n495 PW 0.25fF
C559 S.n496 PW 0.95fF
C560 S.n497 PW 1.49fF
C561 S.n498 PW 1.94fF
C562 S.n499 PW 1.43fF
C563 S.n500 PW 1.18fF
C564 S.n501 PW 0.36fF
C565 S.t110 PW 0.02fF
C566 S.n502 PW 0.12fF
C567 S.n503 PW 0.15fF
C568 S.t28 PW 0.02fF
C569 S.n504 PW 1.25fF
C570 S.n505 PW 0.62fF
C571 S.n506 PW 0.37fF
C572 S.n507 PW 0.65fF
C573 S.n508 PW 1.16fF
C574 S.n509 PW 1.42fF
C575 S.n510 PW 0.61fF
C576 S.n511 PW 0.02fF
C577 S.n512 PW 1.00fF
C578 S.t8 PW 8.19fF
C579 S.n513 PW 9.08fF
C580 S.n515 PW 0.39fF
C581 S.n516 PW 0.24fF
C582 S.n517 PW 2.98fF
C583 S.n518 PW 2.53fF
C584 S.n519 PW 2.61fF
C585 S.n520 PW 4.06fF
C586 S.n521 PW 0.26fF
C587 S.n522 PW 0.01fF
C588 S.t117 PW 0.02fF
C589 S.n523 PW 0.26fF
C590 S.t224 PW 0.02fF
C591 S.n524 PW 0.98fF
C592 S.n525 PW 0.73fF
C593 S.n526 PW 0.81fF
C594 S.n527 PW 2.37fF
C595 S.n528 PW 1.94fF
C596 S.n529 PW 0.12fF
C597 S.t195 PW 0.02fF
C598 S.n530 PW 0.14fF
C599 S.t122 PW 0.02fF
C600 S.n532 PW 0.25fF
C601 S.n533 PW 0.37fF
C602 S.n534 PW 0.63fF
C603 S.n535 PW 1.43fF
C604 S.n536 PW 1.18fF
C605 S.n537 PW 0.36fF
C606 S.n538 PW 2.09fF
C607 S.t37 PW 0.02fF
C608 S.n539 PW 0.25fF
C609 S.n540 PW 0.94fF
C610 S.n541 PW 0.05fF
C611 S.t277 PW 0.02fF
C612 S.n542 PW 0.12fF
C613 S.n543 PW 0.15fF
C614 S.n545 PW 1.95fF
C615 S.n546 PW 2.76fF
C616 S.t9 PW 0.02fF
C617 S.n547 PW 0.25fF
C618 S.n548 PW 0.37fF
C619 S.n549 PW 0.63fF
C620 S.n550 PW 0.12fF
C621 S.t106 PW 0.02fF
C622 S.n551 PW 0.14fF
C623 S.n553 PW 1.19fF
C624 S.n554 PW 0.23fF
C625 S.n555 PW 1.94fF
C626 S.t214 PW 0.02fF
C627 S.n556 PW 0.25fF
C628 S.n557 PW 0.94fF
C629 S.n558 PW 0.05fF
C630 S.t186 PW 0.02fF
C631 S.n559 PW 0.12fF
C632 S.n560 PW 0.15fF
C633 S.n562 PW 7.96fF
C634 S.n563 PW 2.81fF
C635 S.n564 PW 1.87fF
C636 S.n565 PW 0.12fF
C637 S.t161 PW 0.02fF
C638 S.n566 PW 0.14fF
C639 S.t12 PW 0.02fF
C640 S.n568 PW 0.25fF
C641 S.n569 PW 0.37fF
C642 S.n570 PW 0.63fF
C643 S.n571 PW 2.44fF
C644 S.n572 PW 2.37fF
C645 S.t237 PW 0.02fF
C646 S.n573 PW 0.12fF
C647 S.n574 PW 0.15fF
C648 S.t137 PW 0.02fF
C649 S.n576 PW 0.25fF
C650 S.n577 PW 0.94fF
C651 S.n578 PW 0.05fF
C652 S.t209 PW 0.02fF
C653 S.n579 PW 0.25fF
C654 S.n580 PW 0.94fF
C655 S.t90 PW 19.97fF
C656 S.t91 PW 0.02fF
C657 S.n581 PW 0.12fF
C658 S.n582 PW 0.15fF
C659 S.t126 PW 0.02fF
C660 S.n584 PW 0.25fF
C661 S.n585 PW 0.94fF
C662 S.n586 PW 0.05fF
C663 S.t199 PW 0.02fF
C664 S.n587 PW 0.25fF
C665 S.n588 PW 0.37fF
C666 S.n589 PW 0.63fF
C667 S.n590 PW 0.33fF
C668 S.n591 PW 1.59fF
C669 S.n592 PW 0.16fF
C670 S.n593 PW 5.13fF
C671 S.n594 PW 1.94fF
C672 S.n595 PW 0.12fF
C673 S.t116 PW 0.02fF
C674 S.n596 PW 0.14fF
C675 S.t241 PW 0.02fF
C676 S.n598 PW 0.25fF
C677 S.n599 PW 0.37fF
C678 S.n600 PW 0.63fF
C679 S.n601 PW 1.31fF
C680 S.n602 PW 6.16fF
C681 S.t255 PW 0.02fF
C682 S.n603 PW 0.12fF
C683 S.n604 PW 0.15fF
C684 S.t179 PW 0.02fF
C685 S.n606 PW 0.25fF
C686 S.n607 PW 0.94fF
C687 S.n608 PW 0.05fF
C688 S.t19 PW 17.26fF
C689 S.t20 PW 0.02fF
C690 S.n609 PW 0.01fF
C691 S.n610 PW 0.26fF
C692 S.t46 PW 0.02fF
C693 S.n612 PW 1.23fF
C694 S.n613 PW 0.05fF
C695 S.t154 PW 0.02fF
C696 S.n614 PW 0.66fF
C697 S.n615 PW 0.63fF
C698 S.n616 PW 1.55fF
C699 S.n617 PW 0.36fF
C700 S.n618 PW 1.34fF
C701 S.n619 PW 0.16fF
C702 S.n620 PW 1.81fF
C703 S.n621 PW 2.36fF
C704 S.n622 PW 0.02fF
C705 S.n623 PW 0.03fF
C706 S.n624 PW 0.25fF
C707 S.n625 PW 0.13fF
C708 S.n626 PW 0.58fF
C709 S.n627 PW 0.03fF
C710 S.n628 PW 0.89fF
C711 S.n629 PW 0.23fF
C712 S.n630 PW 0.15fF
C713 S.n631 PW 9.26fF
C714 S.n632 PW 9.26fF
C715 S.n633 PW 0.62fF
C716 S.n634 PW 0.24fF
C717 S.n635 PW 0.61fF
C718 S.n636 PW 1.83fF
C719 S.n637 PW 0.30fF
C720 S.t24 PW 8.19fF
C721 S.n638 PW 10.54fF
C722 S.n639 PW 0.79fF
C723 S.n640 PW 0.28fF
C724 S.n641 PW 4.13fF
C725 S.n642 PW 1.17fF
C726 S.t62 PW 0.02fF
C727 S.n643 PW 0.66fF
C728 S.n644 PW 0.63fF
C729 S.n645 PW 0.26fF
C730 S.n646 PW 0.09fF
C731 S.n647 PW 0.21fF
C732 S.n648 PW 1.32fF
C733 S.n649 PW 0.55fF
C734 S.n650 PW 1.94fF
C735 S.n651 PW 0.12fF
C736 S.t173 PW 0.02fF
C737 S.n652 PW 0.14fF
C738 S.t236 PW 0.02fF
C739 S.n654 PW 0.25fF
C740 S.n655 PW 0.37fF
C741 S.n656 PW 0.63fF
C742 S.n657 PW 0.73fF
C743 S.n658 PW 1.63fF
C744 S.n659 PW 2.53fF
C745 S.t145 PW 0.02fF
C746 S.n660 PW 0.25fF
C747 S.n661 PW 0.94fF
C748 S.n662 PW 0.05fF
C749 S.t187 PW 0.02fF
C750 S.n663 PW 0.12fF
C751 S.n664 PW 0.15fF
C752 S.n666 PW 1.95fF
C753 S.n667 PW 0.06fF
C754 S.n668 PW 0.03fF
C755 S.n669 PW 0.04fF
C756 S.n670 PW 1.02fF
C757 S.n671 PW 0.02fF
C758 S.n672 PW 0.01fF
C759 S.n673 PW 0.02fF
C760 S.n674 PW 0.09fF
C761 S.n675 PW 0.37fF
C762 S.n676 PW 1.91fF
C763 S.t153 PW 0.02fF
C764 S.n677 PW 0.25fF
C765 S.n678 PW 0.37fF
C766 S.n679 PW 0.63fF
C767 S.n680 PW 0.12fF
C768 S.t79 PW 0.02fF
C769 S.n681 PW 0.14fF
C770 S.n683 PW 0.72fF
C771 S.n684 PW 0.23fF
C772 S.n685 PW 0.26fF
C773 S.n686 PW 0.09fF
C774 S.n687 PW 0.23fF
C775 S.n688 PW 0.72fF
C776 S.n689 PW 1.19fF
C777 S.n690 PW 0.23fF
C778 S.n691 PW 0.26fF
C779 S.n692 PW 0.09fF
C780 S.n693 PW 1.94fF
C781 S.t42 PW 0.02fF
C782 S.n694 PW 0.25fF
C783 S.n695 PW 0.94fF
C784 S.n696 PW 0.05fF
C785 S.t92 PW 0.02fF
C786 S.n697 PW 0.12fF
C787 S.n698 PW 0.15fF
C788 S.n700 PW 7.96fF
C789 S.n701 PW 0.12fF
C790 S.t263 PW 0.02fF
C791 S.n702 PW 0.14fF
C792 S.t63 PW 0.02fF
C793 S.n704 PW 0.25fF
C794 S.n705 PW 0.37fF
C795 S.n706 PW 0.63fF
C796 S.n707 PW 2.46fF
C797 S.n708 PW 2.28fF
C798 S.n709 PW 0.20fF
C799 S.n710 PW 1.62fF
C800 S.n711 PW 0.33fF
C801 S.n712 PW 0.73fF
C802 S.n713 PW 1.78fF
C803 S.n714 PW 2.49fF
C804 S.t278 PW 0.02fF
C805 S.n715 PW 0.12fF
C806 S.n716 PW 0.15fF
C807 S.t229 PW 0.02fF
C808 S.n718 PW 0.25fF
C809 S.n719 PW 0.94fF
C810 S.n720 PW 0.05fF
C811 S.n721 PW 1.94fF
C812 S.n722 PW 0.12fF
C813 S.t276 PW 0.02fF
C814 S.n723 PW 0.14fF
C815 S.t213 PW 0.02fF
C816 S.n725 PW 1.25fF
C817 S.n726 PW 0.37fF
C818 S.n727 PW 0.65fF
C819 S.n728 PW 1.16fF
C820 S.n729 PW 1.42fF
C821 S.n730 PW 0.61fF
C822 S.n731 PW 0.02fF
C823 S.n732 PW 1.00fF
C824 S.t15 PW 8.19fF
C825 S.n733 PW 9.08fF
C826 S.n735 PW 0.39fF
C827 S.n736 PW 0.24fF
C828 S.n737 PW 3.01fF
C829 S.n738 PW 2.06fF
C830 S.n739 PW 2.55fF
C831 S.n740 PW 4.51fF
C832 S.n741 PW 0.26fF
C833 S.n742 PW 0.01fF
C834 S.t5 PW 0.02fF
C835 S.n743 PW 0.26fF
C836 S.t143 PW 0.02fF
C837 S.n744 PW 0.98fF
C838 S.n745 PW 0.73fF
C839 S.n746 PW 0.81fF
C840 S.n747 PW 2.33fF
C841 S.n748 PW 1.94fF
C842 S.n749 PW 0.12fF
C843 S.t198 PW 0.02fF
C844 S.n750 PW 0.14fF
C845 S.t125 PW 0.02fF
C846 S.n752 PW 0.25fF
C847 S.n753 PW 0.37fF
C848 S.n754 PW 0.63fF
C849 S.n755 PW 1.43fF
C850 S.n756 PW 0.73fF
C851 S.n757 PW 1.18fF
C852 S.n758 PW 0.36fF
C853 S.n759 PW 2.09fF
C854 S.t40 PW 0.02fF
C855 S.n760 PW 0.25fF
C856 S.n761 PW 0.94fF
C857 S.n762 PW 0.05fF
C858 S.t282 PW 0.02fF
C859 S.n763 PW 0.12fF
C860 S.n764 PW 0.15fF
C861 S.n766 PW 1.95fF
C862 S.n767 PW 1.94fF
C863 S.t16 PW 0.02fF
C864 S.n768 PW 0.25fF
C865 S.n769 PW 0.37fF
C866 S.n770 PW 0.63fF
C867 S.n771 PW 0.12fF
C868 S.t109 PW 0.02fF
C869 S.n772 PW 0.14fF
C870 S.n774 PW 1.19fF
C871 S.n775 PW 0.23fF
C872 S.n776 PW 0.26fF
C873 S.n777 PW 0.09fF
C874 S.n778 PW 1.94fF
C875 S.t216 PW 0.02fF
C876 S.n779 PW 0.25fF
C877 S.n780 PW 0.94fF
C878 S.n781 PW 0.05fF
C879 S.t190 PW 0.02fF
C880 S.n782 PW 0.12fF
C881 S.n783 PW 0.15fF
C882 S.n785 PW 7.96fF
C883 S.n786 PW 1.94fF
C884 S.n787 PW 2.76fF
C885 S.t114 PW 0.02fF
C886 S.n788 PW 0.25fF
C887 S.n789 PW 0.37fF
C888 S.n790 PW 0.63fF
C889 S.n791 PW 0.12fF
C890 S.t185 PW 0.02fF
C891 S.n792 PW 0.14fF
C892 S.n794 PW 5.34fF
C893 S.t264 PW 0.02fF
C894 S.n795 PW 0.12fF
C895 S.n796 PW 0.15fF
C896 S.t25 PW 0.02fF
C897 S.n798 PW 0.25fF
C898 S.n799 PW 0.94fF
C899 S.n800 PW 0.05fF
C900 S.n801 PW 0.12fF
C901 S.t279 PW 0.02fF
C902 S.n802 PW 0.14fF
C903 S.t152 PW 0.02fF
C904 S.n804 PW 0.25fF
C905 S.n805 PW 0.37fF
C906 S.n806 PW 0.63fF
C907 S.n807 PW 1.65fF
C908 S.n808 PW 0.03fF
C909 S.n809 PW 0.14fF
C910 S.n810 PW 0.60fF
C911 S.n811 PW 0.12fF
C912 S.n812 PW 0.55fF
C913 S.n813 PW 0.42fF
C914 S.n814 PW 0.25fF
C915 S.n815 PW 0.25fF
C916 S.n816 PW 0.70fF
C917 S.n817 PW 2.04fF
C918 S.t86 PW 0.02fF
C919 S.n818 PW 0.12fF
C920 S.n819 PW 0.15fF
C921 S.t243 PW 0.02fF
C922 S.n821 PW 0.25fF
C923 S.n822 PW 0.94fF
C924 S.n823 PW 0.05fF
C925 S.t4 PW 17.65fF
C926 S.t95 PW 0.02fF
C927 S.n824 PW 0.12fF
C928 S.n825 PW 0.15fF
C929 S.t134 PW 0.02fF
C930 S.n827 PW 0.25fF
C931 S.n828 PW 0.94fF
C932 S.n829 PW 0.05fF
C933 S.t204 PW 0.02fF
C934 S.n830 PW 0.25fF
C935 S.n831 PW 0.37fF
C936 S.n832 PW 0.63fF
C937 S.n833 PW 0.33fF
C938 S.n834 PW 1.12fF
C939 S.n835 PW 0.16fF
C940 S.n836 PW 2.17fF
C941 S.n837 PW 3.03fF
C942 S.n838 PW 1.94fF
C943 S.n839 PW 0.12fF
C944 S.t250 PW 0.02fF
C945 S.n840 PW 0.14fF
C946 S.t52 PW 0.02fF
C947 S.n842 PW 0.25fF
C948 S.n843 PW 0.37fF
C949 S.n844 PW 0.63fF
C950 S.n845 PW 0.95fF
C951 S.n846 PW 0.33fF
C952 S.n847 PW 0.95fF
C953 S.n848 PW 1.12fF
C954 S.n849 PW 0.16fF
C955 S.n850 PW 4.83fF
C956 S.t259 PW 0.02fF
C957 S.n851 PW 0.12fF
C958 S.n852 PW 0.15fF
C959 S.t217 PW 0.02fF
C960 S.n854 PW 0.25fF
C961 S.n855 PW 0.94fF
C962 S.n856 PW 0.05fF
C963 S.n857 PW 1.94fF
C964 S.n858 PW 2.76fF
C965 S.t100 PW 0.02fF
C966 S.n859 PW 0.25fF
C967 S.n860 PW 0.37fF
C968 S.n861 PW 0.63fF
C969 S.n862 PW 0.12fF
C970 S.t231 PW 0.02fF
C971 S.n863 PW 0.14fF
C972 S.n865 PW 5.63fF
C973 S.t169 PW 0.02fF
C974 S.n866 PW 0.12fF
C975 S.n867 PW 0.15fF
C976 S.t33 PW 0.02fF
C977 S.n869 PW 0.25fF
C978 S.n870 PW 0.94fF
C979 S.n871 PW 0.05fF
C980 S.t78 PW 17.26fF
C981 S.t225 PW 0.02fF
C982 S.n872 PW 1.23fF
C983 S.n873 PW 0.05fF
C984 S.t158 PW 0.02fF
C985 S.n874 PW 0.01fF
C986 S.n875 PW 0.26fF
C987 S.n877 PW 1.55fF
C988 S.n878 PW 1.29fF
C989 S.n879 PW 0.28fF
C990 S.n880 PW 0.25fF
C991 S.n881 PW 4.52fF
C992 S.t49 PW 0.02fF
C993 S.n882 PW 1.25fF
C994 S.n883 PW 0.37fF
C995 S.n884 PW 0.48fF
C996 S.n885 PW 1.17fF
C997 S.n886 PW 1.94fF
C998 S.n887 PW 0.12fF
C999 S.t246 PW 0.02fF
C1000 S.n888 PW 0.14fF
C1001 S.t41 PW 0.02fF
C1002 S.n890 PW 0.25fF
C1003 S.n891 PW 0.37fF
C1004 S.n892 PW 0.63fF
C1005 S.n893 PW 2.75fF
C1006 S.n894 PW 4.05fF
C1007 S.t39 PW 0.02fF
C1008 S.n895 PW 0.25fF
C1009 S.n896 PW 0.94fF
C1010 S.n897 PW 0.05fF
C1011 S.t249 PW 0.02fF
C1012 S.n898 PW 0.12fF
C1013 S.n899 PW 0.15fF
C1014 S.n901 PW 1.94fF
C1015 S.n902 PW 2.75fF
C1016 S.t144 PW 0.02fF
C1017 S.n903 PW 0.25fF
C1018 S.n904 PW 0.37fF
C1019 S.n905 PW 0.63fF
C1020 S.n906 PW 0.12fF
C1021 S.t70 PW 0.02fF
C1022 S.n907 PW 0.14fF
C1023 S.n909 PW 2.01fF
C1024 S.n910 PW 2.62fF
C1025 S.t274 PW 0.02fF
C1026 S.n911 PW 0.25fF
C1027 S.n912 PW 0.37fF
C1028 S.n913 PW 0.63fF
C1029 S.t208 PW 0.02fF
C1030 S.n914 PW 0.25fF
C1031 S.n915 PW 0.94fF
C1032 S.n916 PW 0.05fF
C1033 S.t262 PW 0.02fF
C1034 S.n917 PW 0.12fF
C1035 S.n918 PW 0.15fF
C1036 S.n920 PW 0.12fF
C1037 S.t184 PW 0.02fF
C1038 S.n921 PW 0.14fF
C1039 S.n923 PW 2.37fF
C1040 S.n924 PW 1.83fF
C1041 S.n925 PW 5.32fF
C1042 S.t142 PW 0.02fF
C1043 S.n926 PW 0.25fF
C1044 S.n927 PW 0.94fF
C1045 S.n928 PW 0.05fF
C1046 S.t74 PW 0.02fF
C1047 S.n929 PW 0.12fF
C1048 S.n930 PW 0.15fF
C1049 S.n932 PW 2.01fF
C1050 S.n933 PW 0.12fF
C1051 S.t275 PW 0.02fF
C1052 S.n934 PW 0.14fF
C1053 S.n936 PW 7.96fF
C1054 S.n937 PW 0.04fF
C1055 S.n938 PW 0.10fF
C1056 S.n939 PW 0.30fF
C1057 S.n940 PW 0.26fF
C1058 S.n941 PW 0.12fF
C1059 S.n942 PW 0.05fF
C1060 S.n943 PW 0.18fF
C1061 S.n944 PW 1.30fF
C1062 S.n945 PW 2.86fF
C1063 S.n946 PW 0.12fF
C1064 S.t258 PW 0.02fF
C1065 S.n947 PW 0.14fF
C1066 S.t85 PW 0.02fF
C1067 S.n949 PW 0.25fF
C1068 S.n950 PW 0.37fF
C1069 S.n951 PW 0.63fF
C1070 S.n952 PW 2.70fF
C1071 S.n953 PW 2.12fF
C1072 S.t75 PW 0.02fF
C1073 S.n954 PW 0.12fF
C1074 S.n955 PW 0.15fF
C1075 S.t7 PW 0.02fF
C1076 S.n957 PW 0.25fF
C1077 S.n958 PW 0.94fF
C1078 S.n959 PW 0.05fF
C1079 S.t133 PW 0.02fF
C1080 S.n960 PW 0.98fF
C1081 S.n961 PW 0.73fF
C1082 S.n962 PW 0.01fF
C1083 S.t108 PW 0.02fF
C1084 S.n963 PW 0.26fF
C1085 S.t197 PW 0.02fF
C1086 S.n964 PW 1.25fF
C1087 S.n965 PW 2.02fF
C1088 S.n966 PW 0.06fF
C1089 S.n967 PW 0.10fF
C1090 S.n968 PW 0.62fF
C1091 S.n969 PW 1.40fF
C1092 S.n970 PW 1.42fF
C1093 S.n971 PW 0.92fF
C1094 S.n972 PW 0.87fF
C1095 S.n973 PW 0.02fF
C1096 S.n974 PW 1.00fF
C1097 S.t21 PW 8.19fF
C1098 S.n975 PW 8.77fF
C1099 S.n977 PW 0.70fF
C1100 S.n978 PW 0.24fF
C1101 S.n979 PW 2.99fF
C1102 S.n980 PW 2.50fF
C1103 S.n981 PW 3.97fF
C1104 S.n982 PW 0.26fF
C1105 S.n983 PW 2.48fF
C1106 S.n984 PW 2.04fF
C1107 S.n985 PW 0.12fF
C1108 S.t88 PW 0.02fF
C1109 S.n986 PW 0.14fF
C1110 S.t183 PW 0.02fF
C1111 S.n988 PW 0.25fF
C1112 S.n989 PW 0.37fF
C1113 S.n990 PW 0.63fF
C1114 S.n991 PW 2.63fF
C1115 S.n992 PW 2.38fF
C1116 S.t172 PW 0.02fF
C1117 S.n993 PW 0.12fF
C1118 S.n994 PW 0.15fF
C1119 S.t121 PW 0.02fF
C1120 S.n996 PW 0.25fF
C1121 S.n997 PW 0.94fF
C1122 S.n998 PW 0.05fF
C1123 S.n999 PW 0.04fF
C1124 S.n1000 PW 0.10fF
C1125 S.n1001 PW 0.30fF
C1126 S.n1002 PW 0.26fF
C1127 S.n1003 PW 0.12fF
C1128 S.n1004 PW 0.05fF
C1129 S.n1005 PW 0.18fF
C1130 S.n1006 PW 1.18fF
C1131 S.n1007 PW 1.93fF
C1132 S.n1008 PW 0.12fF
C1133 S.t245 PW 0.02fF
C1134 S.n1009 PW 0.14fF
C1135 S.t87 PW 0.02fF
C1136 S.n1011 PW 0.25fF
C1137 S.n1012 PW 0.37fF
C1138 S.n1013 PW 0.63fF
C1139 S.n1014 PW 2.63fF
C1140 S.n1015 PW 2.00fF
C1141 S.t65 PW 0.02fF
C1142 S.n1016 PW 0.12fF
C1143 S.n1017 PW 0.15fF
C1144 S.t127 PW 0.02fF
C1145 S.n1019 PW 0.25fF
C1146 S.n1020 PW 0.94fF
C1147 S.n1021 PW 0.05fF
C1148 S.t64 PW 17.65fF
C1149 S.t93 PW 0.02fF
C1150 S.n1022 PW 0.12fF
C1151 S.n1023 PW 0.15fF
C1152 S.t23 PW 0.02fF
C1153 S.n1025 PW 0.25fF
C1154 S.n1026 PW 0.94fF
C1155 S.n1027 PW 0.05fF
C1156 S.t107 PW 0.02fF
C1157 S.n1028 PW 0.25fF
C1158 S.n1029 PW 0.37fF
C1159 S.n1030 PW 0.63fF
C1160 S.n1031 PW 0.31fF
C1161 S.n1032 PW 1.12fF
C1162 S.n1033 PW 0.16fF
C1163 S.n1034 PW 2.17fF
C1164 S.n1035 PW 1.84fF
C1165 S.n1036 PW 1.94fF
C1166 S.n1037 PW 0.12fF
C1167 S.t165 PW 0.02fF
C1168 S.n1038 PW 0.14fF
C1169 S.t228 PW 0.02fF
C1170 S.n1040 PW 0.25fF
C1171 S.n1041 PW 0.37fF
C1172 S.n1042 PW 0.63fF
C1173 S.n1043 PW 0.95fF
C1174 S.n1044 PW 0.33fF
C1175 S.n1045 PW 0.95fF
C1176 S.n1046 PW 1.12fF
C1177 S.n1047 PW 0.16fF
C1178 S.n1048 PW 5.12fF
C1179 S.t227 PW 0.02fF
C1180 S.n1049 PW 0.25fF
C1181 S.n1050 PW 0.94fF
C1182 S.n1051 PW 0.05fF
C1183 S.t171 PW 0.02fF
C1184 S.n1052 PW 0.12fF
C1185 S.n1053 PW 0.15fF
C1186 S.t45 PW 0.02fF
C1187 S.n1055 PW 0.98fF
C1188 S.n1056 PW 0.73fF
C1189 S.n1057 PW 1.82fF
C1190 S.n1058 PW 3.14fF
C1191 S.t53 PW 0.02fF
C1192 S.n1059 PW 0.25fF
C1193 S.n1060 PW 0.37fF
C1194 S.n1061 PW 0.63fF
C1195 S.n1062 PW 0.12fF
C1196 S.t253 PW 0.02fF
C1197 S.n1063 PW 0.14fF
C1198 S.n1065 PW 0.19fF
C1199 S.n1066 PW 0.21fF
C1200 S.n1067 PW 0.23fF
C1201 S.n1068 PW 0.68fF
C1202 S.n1069 PW 0.93fF
C1203 S.n1070 PW 0.23fF
C1204 S.n1071 PW 0.10fF
C1205 S.n1072 PW 0.21fF
C1206 S.n1073 PW 0.07fF
C1207 S.n1074 PW 0.06fF
C1208 S.n1075 PW 0.07fF
C1209 S.n1076 PW 2.05fF
C1210 S.t51 PW 0.02fF
C1211 S.n1077 PW 0.25fF
C1212 S.n1078 PW 0.94fF
C1213 S.n1079 PW 0.05fF
C1214 S.t261 PW 0.02fF
C1215 S.n1080 PW 0.12fF
C1216 S.n1081 PW 0.15fF
C1217 S.n1083 PW 7.96fF
C1218 S.n1084 PW 0.26fF
C1219 S.n1085 PW 0.09fF
C1220 S.n1086 PW 0.21fF
C1221 S.n1087 PW 0.80fF
C1222 S.n1088 PW 2.00fF
C1223 S.n1089 PW 1.94fF
C1224 S.n1090 PW 0.12fF
C1225 S.t27 PW 0.02fF
C1226 S.n1091 PW 0.14fF
C1227 S.t163 PW 0.02fF
C1228 S.n1093 PW 0.25fF
C1229 S.n1094 PW 0.37fF
C1230 S.n1095 PW 0.63fF
C1231 S.n1096 PW 2.75fF
C1232 S.n1097 PW 3.09fF
C1233 S.t164 PW 0.02fF
C1234 S.n1098 PW 0.12fF
C1235 S.n1099 PW 0.15fF
C1236 S.t283 PW 0.02fF
C1237 S.n1101 PW 0.25fF
C1238 S.n1102 PW 0.94fF
C1239 S.n1103 PW 0.05fF
C1240 S.t220 PW 0.02fF
C1241 S.n1104 PW 0.01fF
C1242 S.n1105 PW 0.26fF
C1243 S.t26 PW 17.65fF
C1244 S.n1106 PW 0.26fF
C1245 S.n1107 PW 3.01fF
C1246 S.n1108 PW 14.04fF
C1247 S.n1109 PW 0.62fF
C1248 S.n1110 PW 0.49fF
C1249 S.n1111 PW 0.61fF
C1250 S.n1112 PW 1.83fF
C1251 S.n1113 PW 0.30fF
C1252 S.t6 PW 8.19fF
C1253 S.n1114 PW 10.54fF
C1254 S.n1115 PW 0.79fF
C1255 S.n1116 PW 0.28fF
C1256 S.n1117 PW 14.04fF
C1257 S.n1118 PW 4.64fF
C1258 S.n1119 PW 2.40fF
C1259 S.n1120 PW 4.71fF
C1260 S.n1121 PW 4.60fF
C1261 S.n1122 PW 2.60fF
C1262 S.t128 PW 0.02fF
C1263 S.n1123 PW 1.32fF
C1264 S.t174 PW 0.02fF
C1265 S.n1124 PW 0.45fF
C1266 S.n1125 PW 7.96fF
C1267 S.n1126 PW 0.03fF
C1268 S.n1127 PW 0.02fF
C1269 S.n1128 PW 0.02fF
C1270 S.n1129 PW 0.64fF
C1271 S.n1130 PW 0.03fF
C1272 S.n1131 PW 0.03fF
C1273 S.n1132 PW 0.02fF
C1274 S.n1133 PW 0.25fF
C1275 S.n1134 PW 0.15fF
C1276 S.n1135 PW 0.18fF
C1277 S.n1136 PW 1.29fF
C1278 S.n1137 PW 0.24fF
C1279 S.n1138 PW 1.29fF
C1280 S.n1139 PW 0.24fF
C1281 S.n1141 PW 1.51fF
C1282 S.n1142 PW 0.41fF
C1283 S.n1144 PW 1.74fF
C1284 S.n1145 PW 0.41fF
C1285 S.n1146 PW 58.92fF
C1286 S.n1147 PW 4.84fF
C1287 S.t242 PW 0.02fF
C1288 S.n1148 PW 0.92fF
C1289 S.t57 PW 0.02fF
C1290 S.n1149 PW 0.02fF
C1291 S.n1150 PW 0.38fF
C1292 S.t248 PW 0.02fF
C1293 S.n1151 PW 0.92fF
C1294 S.n1152 PW 0.95fF
C1295 S.n1153 PW 4.24fF
C1296 S.n1154 PW 1.91fF
C1297 S.t69 PW 0.02fF
C1298 S.n1155 PW 0.92fF
C1299 S.t71 PW 0.02fF
C1300 S.n1156 PW 0.92fF
C1301 S.n1157 PW 2.19fF
C1302 S.n1158 PW 1.23fF
C1303 S.n1159 PW 0.34fF
C1304 S.n1160 PW 0.32fF
C1305 S.t132 PW 0.02fF
C1306 S.n1161 PW 0.02fF
C1307 S.n1162 PW 0.38fF
C1308 S.n1163 PW 0.21fF
C1309 S.n1164 PW 2.26fF
C1310 S.n1165 PW 1.31fF
C1311 S.n1166 PW 0.32fF
C1312 S.t247 PW 0.02fF
C1313 S.n1167 PW 0.92fF
C1314 S.t244 PW 0.02fF
C1315 S.n1168 PW 0.92fF
C1316 S.n1169 PW 3.99fF
C1317 S.n1170 PW 2.88fF
C1318 S.t22 PW 0.02fF
C1319 S.n1171 PW 0.02fF
C1320 S.n1172 PW 0.38fF
C1321 S.n1173 PW 1.02fF
C1322 S.n1174 PW 3.72fF
C1323 S.n1175 PW 2.89fF
C1324 S.t159 PW 0.02fF
C1325 S.n1176 PW 0.92fF
C1326 S.t162 PW 0.02fF
C1327 S.n1177 PW 0.92fF
C1328 S.n1178 PW 2.50fF
C1329 S.t207 PW 0.02fF
C1330 S.n1179 PW 0.02fF
C1331 S.n1180 PW 0.38fF
C1332 S.n1181 PW 4.10fF
C1333 S.n1182 PW 2.87fF
C1334 S.n1183 PW 0.03fF
C1335 S.n1184 PW 0.02fF
C1336 S.n1185 PW 0.03fF
C1337 S.n1186 PW 0.03fF
C1338 S.n1187 PW 0.02fF
C1339 S.n1188 PW 0.02fF
C1340 S.n1189 PW 0.64fF
C1341 S.n1190 PW 0.25fF
C1342 S.n1191 PW 0.15fF
C1343 S.n1192 PW 0.18fF
C1344 S.t67 PW 0.02fF
C1345 S.n1193 PW 0.92fF
C1346 S.t68 PW 0.02fF
C1347 S.n1194 PW 0.92fF
C1348 S.t120 PW 0.02fF
C1349 S.n1195 PW 0.02fF
C1350 S.n1196 PW 0.38fF
C1351 S.t66 PW 56.97fF
C1352 S.n1197 PW 0.48fF
C1353 S.n1198 PW 2.53fF
C1354 S.n1200 PW 0.87fF
C1355 S.n1201 PW 0.13fF
C1356 S.n1202 PW 1.11fF
C1357 S.n1203 PW 8.73fF
C1358 S.n1205 PW 14.84fF
C1359 S.n1206 PW 0.79fF
C1360 S.n1207 PW 0.54fF
C1361 S.n1208 PW 12.00fF
C1362 S.n1209 PW 2.60fF
C1363 S.n1210 PW 7.20fF
C1364 S.n1211 PW 16.58fF
C1365 S.n1212 PW 9.26fF
C1366 S.n1213 PW 9.26fF
C1367 S.n1214 PW 0.62fF
C1368 S.n1215 PW 0.24fF
C1369 S.n1216 PW 0.61fF
C1370 S.n1217 PW 1.83fF
C1371 S.n1218 PW 0.30fF
C1372 S.t31 PW 8.19fF
C1373 S.n1219 PW 10.54fF
C1374 S.n1220 PW 0.79fF
C1375 S.n1221 PW 0.28fF
C1376 S.n1222 PW 4.40fF
C1377 S.n1223 PW 2.89fF
C1378 S.n1224 PW 1.95fF
C1379 S.n1225 PW 0.06fF
C1380 S.n1226 PW 0.03fF
C1381 S.n1227 PW 0.04fF
C1382 S.n1228 PW 1.02fF
C1383 S.n1229 PW 0.02fF
C1384 S.n1230 PW 0.01fF
C1385 S.n1231 PW 0.02fF
C1386 S.n1232 PW 0.09fF
C1387 S.n1233 PW 0.37fF
C1388 S.n1234 PW 1.91fF
C1389 S.t156 PW 0.02fF
C1390 S.n1235 PW 0.25fF
C1391 S.n1236 PW 0.37fF
C1392 S.n1237 PW 0.63fF
C1393 S.n1238 PW 0.12fF
C1394 S.t81 PW 0.02fF
C1395 S.n1239 PW 0.14fF
C1396 S.n1241 PW 0.72fF
C1397 S.n1242 PW 0.23fF
C1398 S.n1243 PW 0.23fF
C1399 S.n1244 PW 0.72fF
C1400 S.n1245 PW 1.19fF
C1401 S.n1246 PW 0.23fF
C1402 S.n1247 PW 0.26fF
C1403 S.n1248 PW 0.09fF
C1404 S.n1249 PW 1.94fF
C1405 S.t48 PW 0.02fF
C1406 S.n1250 PW 0.25fF
C1407 S.n1251 PW 0.94fF
C1408 S.n1252 PW 0.05fF
C1409 S.t96 PW 0.02fF
C1410 S.n1253 PW 0.12fF
C1411 S.n1254 PW 0.15fF
C1412 S.n1256 PW 7.96fF
C1413 S.n1257 PW 0.10fF
C1414 S.n1258 PW 0.21fF
C1415 S.n1259 PW 0.07fF
C1416 S.n1260 PW 0.06fF
C1417 S.n1261 PW 0.07fF
C1418 S.n1262 PW 0.19fF
C1419 S.n1263 PW 0.20fF
C1420 S.n1264 PW 1.07fF
C1421 S.n1265 PW 0.55fF
C1422 S.n1266 PW 2.41fF
C1423 S.n1267 PW 0.12fF
C1424 S.t176 PW 0.02fF
C1425 S.n1268 PW 0.14fF
C1426 S.t239 PW 0.02fF
C1427 S.n1270 PW 0.25fF
C1428 S.n1271 PW 0.37fF
C1429 S.n1272 PW 0.63fF
C1430 S.n1273 PW 1.78fF
C1431 S.n1274 PW 2.52fF
C1432 S.t191 PW 0.02fF
C1433 S.n1275 PW 0.12fF
C1434 S.n1276 PW 0.15fF
C1435 S.t150 PW 0.02fF
C1436 S.n1278 PW 0.25fF
C1437 S.n1279 PW 0.94fF
C1438 S.n1280 PW 0.05fF
C1439 S.n1281 PW 3.03fF
C1440 S.n1282 PW 1.94fF
C1441 S.n1283 PW 0.12fF
C1442 S.t254 PW 0.02fF
C1443 S.n1284 PW 0.14fF
C1444 S.t59 PW 0.02fF
C1445 S.n1286 PW 0.25fF
C1446 S.n1287 PW 0.37fF
C1447 S.n1288 PW 0.63fF
C1448 S.n1289 PW 0.95fF
C1449 S.n1290 PW 0.33fF
C1450 S.n1291 PW 0.95fF
C1451 S.n1292 PW 1.12fF
C1452 S.n1293 PW 0.16fF
C1453 S.n1294 PW 5.12fF
C1454 S.t266 PW 0.02fF
C1455 S.n1295 PW 0.12fF
C1456 S.n1296 PW 0.15fF
C1457 S.t223 PW 0.02fF
C1458 S.n1298 PW 0.25fF
C1459 S.n1299 PW 0.94fF
C1460 S.n1300 PW 0.05fF
C1461 S.n1301 PW 1.94fF
C1462 S.n1302 PW 2.75fF
C1463 S.t232 PW 0.02fF
C1464 S.n1303 PW 0.25fF
C1465 S.n1304 PW 0.37fF
C1466 S.n1305 PW 0.63fF
C1467 S.n1306 PW 0.12fF
C1468 S.t166 PW 0.02fF
C1469 S.n1307 PW 0.14fF
C1470 S.n1309 PW 3.03fF
C1471 S.n1310 PW 5.04fF
C1472 S.t175 PW 0.02fF
C1473 S.n1311 PW 0.12fF
C1474 S.n1312 PW 0.15fF
C1475 S.t138 PW 0.02fF
C1476 S.n1314 PW 0.25fF
C1477 S.n1315 PW 0.94fF
C1478 S.n1316 PW 0.05fF
C1479 S.n1317 PW 0.11fF
C1480 S.n1318 PW 0.12fF
C1481 S.n1319 PW 0.10fF
C1482 S.n1320 PW 0.12fF
C1483 S.n1321 PW 0.19fF
C1484 S.n1322 PW 1.94fF
C1485 S.n1323 PW 0.12fF
C1486 S.t98 PW 0.02fF
C1487 S.n1324 PW 0.14fF
C1488 S.t130 PW 0.02fF
C1489 S.n1326 PW 1.25fF
C1490 S.n1327 PW 0.06fF
C1491 S.n1328 PW 0.10fF
C1492 S.n1329 PW 0.62fF
C1493 S.n1330 PW 0.37fF
C1494 S.n1331 PW 0.65fF
C1495 S.n1332 PW 1.16fF
C1496 S.n1333 PW 1.42fF
C1497 S.n1334 PW 0.61fF
C1498 S.n1335 PW 0.02fF
C1499 S.n1336 PW 1.00fF
C1500 S.t0 PW 8.19fF
C1501 S.n1337 PW 9.08fF
C1502 S.n1339 PW 0.39fF
C1503 S.n1340 PW 0.24fF
C1504 S.n1341 PW 2.99fF
C1505 S.n1342 PW 2.50fF
C1506 S.n1343 PW 2.55fF
C1507 S.n1344 PW 4.42fF
C1508 S.n1345 PW 0.26fF
C1509 S.n1346 PW 0.01fF
C1510 S.t202 PW 0.02fF
C1511 S.n1347 PW 0.26fF
C1512 S.t44 PW 0.02fF
C1513 S.n1348 PW 0.98fF
C1514 S.n1349 PW 0.73fF
C1515 S.n1350 PW 1.95fF
C1516 S.n1351 PW 1.94fF
C1517 S.t18 PW 0.02fF
C1518 S.n1352 PW 0.25fF
C1519 S.n1353 PW 0.37fF
C1520 S.n1354 PW 0.63fF
C1521 S.n1355 PW 0.12fF
C1522 S.t113 PW 0.02fF
C1523 S.n1356 PW 0.14fF
C1524 S.n1358 PW 1.19fF
C1525 S.n1359 PW 0.23fF
C1526 S.n1360 PW 0.26fF
C1527 S.n1361 PW 0.09fF
C1528 S.n1362 PW 1.94fF
C1529 S.t219 PW 0.02fF
C1530 S.n1363 PW 0.25fF
C1531 S.n1364 PW 0.94fF
C1532 S.n1365 PW 0.05fF
C1533 S.t194 PW 0.02fF
C1534 S.n1366 PW 0.12fF
C1535 S.n1367 PW 0.15fF
C1536 S.n1369 PW 0.80fF
C1537 S.n1370 PW 0.46fF
C1538 S.n1371 PW 1.63fF
C1539 S.n1372 PW 0.12fF
C1540 S.t146 PW 0.02fF
C1541 S.n1373 PW 0.14fF
C1542 S.t252 PW 0.02fF
C1543 S.n1375 PW 0.25fF
C1544 S.n1376 PW 0.37fF
C1545 S.n1377 PW 0.63fF
C1546 S.n1378 PW 0.01fF
C1547 S.n1379 PW 0.07fF
C1548 S.n1380 PW 0.01fF
C1549 S.n1381 PW 0.02fF
C1550 S.n1382 PW 0.02fF
C1551 S.n1383 PW 0.25fF
C1552 S.n1384 PW 1.19fF
C1553 S.n1385 PW 1.38fF
C1554 S.n1386 PW 2.05fF
C1555 S.t101 PW 0.02fF
C1556 S.n1387 PW 0.25fF
C1557 S.n1388 PW 0.94fF
C1558 S.n1389 PW 0.05fF
C1559 S.t215 PW 0.02fF
C1560 S.n1390 PW 0.12fF
C1561 S.n1391 PW 0.15fF
C1562 S.n1393 PW 7.96fF
C1563 S.n1394 PW 1.94fF
C1564 S.n1395 PW 0.12fF
C1565 S.t285 PW 0.02fF
C1566 S.n1396 PW 0.14fF
C1567 S.t206 PW 0.02fF
C1568 S.n1398 PW 0.25fF
C1569 S.n1399 PW 0.37fF
C1570 S.n1400 PW 0.63fF
C1571 S.n1401 PW 0.33fF
C1572 S.n1402 PW 1.12fF
C1573 S.n1403 PW 0.16fF
C1574 S.n1404 PW 2.17fF
C1575 S.t103 PW 0.02fF
C1576 S.n1405 PW 0.12fF
C1577 S.n1406 PW 0.15fF
C1578 S.t136 PW 0.02fF
C1579 S.n1408 PW 0.25fF
C1580 S.n1409 PW 0.94fF
C1581 S.n1410 PW 0.05fF
C1582 S.n1411 PW 1.94fF
C1583 S.n1412 PW 2.75fF
C1584 S.t119 PW 0.02fF
C1585 S.n1413 PW 0.25fF
C1586 S.n1414 PW 0.37fF
C1587 S.n1415 PW 0.63fF
C1588 S.n1416 PW 0.12fF
C1589 S.t193 PW 0.02fF
C1590 S.n1417 PW 0.14fF
C1591 S.n1419 PW 2.37fF
C1592 S.t269 PW 0.02fF
C1593 S.n1420 PW 0.12fF
C1594 S.n1421 PW 0.15fF
C1595 S.t32 PW 0.02fF
C1596 S.n1423 PW 0.25fF
C1597 S.n1424 PW 0.94fF
C1598 S.n1425 PW 0.05fF
C1599 S.t97 PW 17.65fF
C1600 S.t177 PW 0.02fF
C1601 S.n1426 PW 0.12fF
C1602 S.n1427 PW 0.15fF
C1603 S.t210 PW 0.02fF
C1604 S.n1429 PW 0.25fF
C1605 S.n1430 PW 0.94fF
C1606 S.n1431 PW 0.05fF
C1607 S.t1 PW 0.02fF
C1608 S.n1432 PW 0.25fF
C1609 S.n1433 PW 0.37fF
C1610 S.n1434 PW 0.63fF
C1611 S.n1435 PW 2.74fF
C1612 S.n1436 PW 3.38fF
C1613 S.n1437 PW 0.11fF
C1614 S.n1438 PW 0.37fF
C1615 S.n1439 PW 0.48fF
C1616 S.n1440 PW 1.17fF
C1617 S.n1441 PW 1.93fF
C1618 S.n1442 PW 0.12fF
C1619 S.t77 PW 0.02fF
C1620 S.n1443 PW 0.14fF
C1621 S.t221 PW 0.02fF
C1622 S.n1445 PW 0.25fF
C1623 S.n1446 PW 0.37fF
C1624 S.n1447 PW 0.63fF
C1625 S.n1448 PW 1.31fF
C1626 S.n1449 PW 2.46fF
C1627 S.n1450 PW 4.33fF
C1628 S.t80 PW 0.02fF
C1629 S.n1451 PW 0.12fF
C1630 S.n1452 PW 0.15fF
C1631 S.t160 PW 0.02fF
C1632 S.n1454 PW 0.25fF
C1633 S.n1455 PW 0.94fF
C1634 S.n1456 PW 0.05fF
C1635 S.t76 PW 17.26fF
C1636 S.t267 PW 0.02fF
C1637 S.n1457 PW 0.01fF
C1638 S.n1458 PW 0.26fF
C1639 S.t147 PW 0.02fF
C1640 S.n1460 PW 1.23fF
C1641 S.n1461 PW 0.05fF
C1642 S.t234 PW 0.02fF
C1643 S.n1462 PW 0.66fF
C1644 S.n1463 PW 0.63fF
C1645 S.n1464 PW 1.55fF
C1646 S.n1465 PW 0.02fF
C1647 S.n1466 PW 0.01fF
C1648 S.n1467 PW 0.01fF
C1649 S.n1468 PW 0.01fF
C1650 S.n1469 PW 0.02fF
C1651 S.n1470 PW 0.02fF
C1652 S.n1471 PW 0.03fF
C1653 S.n1472 PW 0.04fF
C1654 S.n1473 PW 0.17fF
C1655 S.n1474 PW 0.10fF
C1656 S.n1475 PW 0.17fF
C1657 S.n1476 PW 0.15fF
C1658 S.n1477 PW 0.28fF
C1659 S.n1478 PW 0.25fF
C1660 S.n1479 PW 4.84fF
C1661 S.n1480 PW 9.58fF
C1662 S.n1481 PW 9.58fF
C1663 S.n1482 PW 9.68fF
C1664 S.n1483 PW 18.33fF
.ends

