* NGSPICE file created from mag_files/POSTLAYOUT/power_stage_flat.ext - technology: sky130A

.subckt mag_files/POSTLAYOUT/power_stage_flat s1 s2 s3 s4 fc1 fc2 out VP VN
X0 fc1 s1 VP.t1350 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1 fc2.t390 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3 VP.t1349 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4 fc1 s1 VP.t1348 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7 VN.t390 s4 fc2.t504 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9 VP.t1347 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10 fc1 s1 VP.t1346 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11 VP.t1345 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12 fc2.t389 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14 out s3 fc2.t388 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X15 fc1 s1 VP.t1344 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X16 fc1 s1 VP.t1343 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X17 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X18 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X19 fc1 s1 VP.t1342 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X20 fc1 s1 VP.t1341 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X21 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X22 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X23 fc1 s1 VP.t1340 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X24 VP.t1339 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X25 fc2.t387 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X26 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X27 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X28 fc1 s1 VP.t1338 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X29 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X30 fc1 s1 VP.t1337 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X31 VP.t1336 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X32 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X33 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X34 VP.t1335 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X35 fc1 s1 VP.t1334 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X36 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X37 fc2.t386 s3 out fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X38 fc1 s1 VP.t1333 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X39 VN.t389 s4 fc2.t656 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X40 out s3 fc2.t385 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X41 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X42 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X43 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X44 fc1 s1 VP.t1332 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X45 VN.t388 s4 fc2.t468 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X46 VN.t387 s4 fc2.t537 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X47 VP.t1331 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X48 VP.t1330 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X49 VP.t1329 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X50 VP.t1328 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X51 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X52 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X53 fc1 s1 VP.t1327 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X54 VP.t1326 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X55 VP.t1325 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X56 out s3 fc2.t384 fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X57 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X58 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X59 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X60 fc2.t383 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X61 VN.t386 s4 fc2.t568 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X62 VP.t1324 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X63 fc1 s1 VP.t1323 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X64 VP.t1322 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X65 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X66 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X67 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X68 VP.t1321 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X69 fc2.t382 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X70 VP.t1320 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X71 fc1 s1 VP.t1319 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X72 fc2.t538 s4 VN.t385 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X73 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X74 VP.t1318 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X75 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X76 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X77 fc1 s1 VP.t1317 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X78 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X79 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X80 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X81 fc2.t613 s4 VN.t384 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X82 fc1 s1 VP.t1316 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X83 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X84 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X85 VP.t1315 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X86 VP.t1314 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X87 VP.t1313 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X88 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X89 VP.t1312 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X90 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X91 fc2.t381 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X92 VP.t1311 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X93 fc1 s1 VP.t1310 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X94 fc1 s1 VP.t1309 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X95 fc1 s1 VP.t1308 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X96 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X97 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X98 VP.t1307 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X99 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X101 fc1 s1 VP.t1306 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X102 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X103 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X104 fc1 s1 VP.t1305 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X105 fc2.t380 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X106 VP.t1304 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X107 fc1 s1 VP.t1303 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X108 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X109 fc1 s1 VP.t1302 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X110 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X111 out s3 fc2.t379 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X112 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X113 fc1 s1 VP.t1301 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X114 out s3 fc2.t378 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X116 VN.t383 s4 fc2.t634 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X117 VP.t1300 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X118 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X119 fc2.t734 s4 VN.t382 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X120 out s3 fc2.t377 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X121 VP.t1299 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X122 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X123 fc1 s1 VP.t1298 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X124 VP.t1297 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X125 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X126 fc1 s1 VP.t1296 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X127 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X128 fc1 s1 VP.t1295 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X129 VP.t1294 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X130 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X131 VN.t381 s4 fc2.t526 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X132 fc2.t609 s4 VN.t380 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X133 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X134 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X136 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X137 fc1 s1 VP.t1293 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X138 VP.t1292 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X139 VP.t1291 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X140 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X141 fc2.t376 s3 out fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X142 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X143 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X144 fc1 s1 VP.t1290 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X145 fc2.t375 s3 out fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X146 fc2.t374 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X147 VP.t1289 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X148 fc2.t529 s4 VN.t379 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X149 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X150 VP.t1288 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X151 fc1 s1 VP.t1287 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X152 fc2.t559 s4 VN.t378 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X153 VP.t1286 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X154 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X156 VP.t1285 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X157 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X158 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X159 fc2.t745 s4 VN.t377 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X160 out s3 fc2.t373 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X161 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X162 VP.t1284 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X163 VN.t376 s4 fc2.t744 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X164 fc2.t372 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X165 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X166 fc1 s1 VP.t1283 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X167 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X168 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X169 VN.t375 s4 fc2.t576 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X170 fc2.t371 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X171 fc1 s1 VP.t1282 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X172 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X173 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X174 VP.t1281 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X175 fc1 s1 VP.t1280 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X176 VP.t1279 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X177 fc2.t575 s4 VN.t374 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X178 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X179 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X180 VP.t1278 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X181 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X182 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X183 fc1 s1 VP.t1277 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X184 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X185 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X186 fc2.t619 s4 VN.t373 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X187 VP.t1276 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X188 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X189 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X190 out s3 fc2.t370 fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X191 VP.t1275 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X192 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X193 fc2.t663 s4 VN.t372 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X194 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X195 VP.t1274 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X196 fc2.t687 s4 VN.t371 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X197 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X198 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X199 fc1 s1 VP.t1273 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X200 fc1 s1 VP.t1272 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X201 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X202 VN.t370 s4 fc2.t494 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X203 out s3 fc2.t369 fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X204 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X205 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X206 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X207 fc1 s1 VP.t1271 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X208 fc1 s1 VP.t1270 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X209 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X210 VP.t1269 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X211 VN.t369 s4 fc2.t527 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X212 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X213 fc2.t626 s4 VN.t368 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X214 fc1 s1 VP.t1268 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X215 fc1 s1 VP.t1267 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X216 fc1 s1 VP.t1266 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X217 VP.t1265 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X218 VP.t1264 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X219 fc1 s1 VP.t1263 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X220 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X221 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X222 VN.t367 s4 fc2.t691 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X223 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X224 out s3 fc2.t368 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X225 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X226 fc1 s1 VP.t1262 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X227 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X228 fc1 s1 VP.t1261 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X229 VP.t1260 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X230 VP.t1259 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X231 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X232 VP.t1258 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X233 VP.t1257 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X234 VN.t366 s4 fc2.t533 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X235 out s3 fc2.t367 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X236 fc2.t366 s3 out fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X237 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X238 fc1 s1 VP.t1256 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X239 fc2.t365 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X240 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X241 fc1 s1 VP.t1255 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X242 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X243 VP.t1254 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X244 VP.t1253 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X246 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X247 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X248 VP.t1252 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X249 fc2.t364 s3 out fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X250 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X251 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X252 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X253 VP.t1251 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X254 VP.t1250 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X255 fc2.t363 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X256 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X257 VP.t1249 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X258 out s3 fc2.t362 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X260 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X261 out s3 fc2.t361 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X262 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X263 fc1 s1 VP.t1248 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X264 VP.t1247 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X265 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X266 VP.t1246 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X267 VP.t1245 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X268 fc2.t360 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X269 out s3 fc2.t359 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X270 VN.t365 s4 fc2.t535 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X271 fc2.t358 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X272 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X273 fc1 s1 VP.t1244 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X274 VN.t364 s4 fc2.t555 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X275 VN.t363 s4 fc2.t653 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X276 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X277 VP.t1243 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X278 fc1 s1 VP.t1242 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X279 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X280 fc1 s1 VP.t1241 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X281 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X282 VP.t1240 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X283 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X284 out s3 fc2.t357 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X285 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X286 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X287 fc1 s1 VP.t1239 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X288 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X289 VP.t1238 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X290 fc1 s1 VP.t1237 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X291 VP.t1236 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X292 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X293 VN.t362 s4 fc2.t554 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X294 out s3 fc2.t356 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X295 fc2.t355 s3 out fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X296 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X297 fc1 s1 VP.t1235 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X298 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X299 out s3 fc2.t354 fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X300 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X301 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X302 fc1 s1 VP.t1234 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X303 VP.t1233 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X304 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X305 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X306 VP.t1232 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X307 fc1 s1 VP.t1231 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X308 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X309 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X310 fc1 s1 VP.t1230 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X311 VN.t361 s4 fc2.t730 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X312 fc2.t353 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X313 fc1 s1 VP.t1229 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X314 fc2.t598 s4 VN.t360 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X315 VP.t1228 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X316 VN.t359 s4 fc2.t405 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X317 out s3 fc2.t352 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X318 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X319 fc1 s1 VP.t1227 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X320 fc1 s1 VP.t1226 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X321 VP.t1225 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X322 fc1 s1 VP.t1224 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X323 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X324 VP.t1223 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X325 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X326 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X327 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X328 fc2.t720 s4 VN.t358 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X329 fc1 s1 VP.t1222 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X330 VN.t357 s4 fc2.t471 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X331 VP.t1221 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X332 fc1 s1 VP.t1220 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X333 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X334 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X335 fc1 s1 VP.t1219 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X336 out s3 fc2.t351 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X337 VP.t1218 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X338 fc2.t532 s4 VN.t356 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X339 VP.t1217 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X340 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X341 fc1 s1 VP.t1216 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X342 fc2.t391 s4 VN.t355 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X343 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X344 VP.t1215 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X345 VP.t1214 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X346 fc1 s1 VP.t1213 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X347 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X348 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X349 VP.t1212 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X350 VP.t1211 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X351 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X352 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X353 fc1 s1 VP.t1210 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X354 out s3 fc2.t350 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X355 VP.t1209 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X356 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X357 VP.t1208 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X358 VP.t1207 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X359 fc2.t645 s4 VN.t354 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X360 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X361 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X362 out s3 fc2.t349 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X363 VP.t1206 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X364 fc1 s1 VP.t1205 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X365 fc2.t348 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X366 fc2.t557 s4 VN.t353 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X367 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X368 VN.t352 s4 fc2.t675 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X369 fc1 s1 VP.t1204 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X370 fc1 s1 VP.t1203 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X371 fc2.t347 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X372 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X373 fc1 s1 VP.t1202 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X374 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X375 fc1 s1 VP.t1201 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X377 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X378 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X379 VP.t1200 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X380 fc1 s1 VP.t1199 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X381 fc2.t412 s4 VN.t351 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X382 fc2.t346 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X383 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X384 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X385 fc1 s1 VP.t1198 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X386 fc1 s1 VP.t1197 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X387 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X388 out s3 fc2.t345 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X389 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X390 fc1 s1 VP.t1196 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X391 fc1 s1 VP.t1195 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X392 fc1 s1 VP.t1194 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X393 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X394 VN.t350 s4 fc2.t719 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X395 fc1 s1 VP.t1193 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X396 VP.t1192 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X397 out s3 fc2.t344 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X398 VP.t1191 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X399 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X400 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X401 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X402 VP.t1190 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X403 fc1 s1 VP.t1189 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X404 VN.t349 s4 fc2.t416 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X405 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X406 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X407 VP.t1188 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X408 fc1 s1 VP.t1187 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X409 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X410 fc1 s1 VP.t1186 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X411 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X412 fc1 s1 VP.t1185 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X413 fc2.t343 s3 out fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X414 fc1 s1 VP.t1184 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X415 fc2.t743 s4 VN.t348 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X416 out s3 fc2.t342 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X417 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X418 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X419 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X420 fc1 s1 VP.t1183 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X421 fc2.t702 s4 VN.t347 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X422 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X423 VN.t346 s4 fc2.t624 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X424 fc1 s1 VP.t1182 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X425 fc2.t560 s4 VN.t345 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X426 VP.t1181 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X427 VP.t1180 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X428 fc1 s1 VP.t1179 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X429 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X430 fc1 s1 VP.t1178 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X431 VP.t1177 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X432 fc1 s1 VP.t1176 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X433 VP.t1175 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X435 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X436 fc2.t563 s4 VN.t344 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X437 fc1 s1 VP.t1174 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X438 VP.t1173 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X439 VP.t1172 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X440 VP.t1171 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X441 VP.t1170 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X442 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X443 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X444 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X445 fc1 s1 VP.t1169 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X446 VP.t1168 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X447 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X448 VP.t1167 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X449 fc2.t341 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X450 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X451 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X452 fc1 s1 VP.t1166 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X453 VP.t1165 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X454 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X455 fc1 s1 VP.t1164 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X456 VP.t1163 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X457 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X458 fc2.t340 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X459 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X460 VP.t1162 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X461 fc2.t424 s4 VN.t343 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X462 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X463 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X464 fc1 s1 VP.t1161 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X465 fc1 s1 VP.t1160 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X466 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X467 VP.t1159 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X468 fc2.t392 s4 VN.t342 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X469 fc2.t339 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X470 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X471 VP.t1158 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X472 VP.t1157 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X473 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X474 fc2.t406 s4 VN.t341 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X475 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X476 VP.t1156 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X477 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X478 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X479 fc1 s1 VP.t1155 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X480 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X481 fc1 s1 VP.t1154 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X482 fc1 s1 VP.t1153 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X483 VP.t1152 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X484 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X485 out s3 fc2.t338 fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X486 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X487 fc2.t620 s4 VN.t340 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X488 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X489 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X490 fc1 s1 VP.t1151 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X491 fc2.t337 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X492 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X493 fc1 s1 VP.t1150 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X494 VP.t1149 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X495 fc1 s1 VP.t1148 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X496 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X497 VP.t1147 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X498 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X499 fc1 s1 VP.t1146 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X500 out s3 fc2.t336 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X502 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X503 fc2.t658 s4 VN.t339 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X504 out s3 fc2.t335 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X505 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X506 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X507 VP.t1145 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X508 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X509 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X510 fc1 s1 VP.t1144 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X511 VP.t1143 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X512 VP.t1142 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X513 fc1 s1 VP.t1141 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X514 fc2.t334 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X515 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X516 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X517 fc1 s1 VP.t1140 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X518 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X519 out s3 fc2.t333 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X520 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X521 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X522 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X523 fc1 s1 VP.t1139 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X524 VP.t1138 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X525 VP.t1137 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X526 fc2.t332 s3 out fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X527 fc1 s1 VP.t1136 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X528 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X529 fc1 s1 VP.t1135 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X530 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X531 VN.t338 s4 fc2.t671 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X532 fc2.t331 s3 out fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X533 fc2.t330 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X534 fc2.t475 s4 VN.t337 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X535 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X536 VP.t1134 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X537 fc1 s1 VP.t1133 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X538 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X539 fc2.t668 s4 VN.t336 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X540 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X541 VP.t1132 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X542 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X543 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X544 VP.t1131 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X545 fc2.t329 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X546 fc1 s1 VP.t1130 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X547 VP.t1129 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X548 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X549 fc1 s1 VP.t1128 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X550 fc1 s1 VP.t1127 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X551 VP.t1126 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X552 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X553 out s3 fc2.t328 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X554 VP.t1125 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X555 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X556 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X557 fc2.t580 s4 VN.t335 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X558 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X559 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X560 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X561 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X562 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X563 fc2.t327 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X564 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X565 fc1 s1 VP.t1124 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X566 VP.t1123 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X567 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X568 VP.t1122 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X569 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X570 fc1 s1 VP.t1121 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X571 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X572 out s3 fc2.t326 fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X573 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X574 VP.t1120 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X575 VP.t1119 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X576 VN.t334 s4 fc2.t452 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X577 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X578 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X579 VN.t333 s4 fc2.t413 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X580 fc2.t553 s4 VN.t332 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X581 VP.t1118 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X582 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X583 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X584 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X585 fc1 s1 VP.t1117 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X586 fc1 s1 VP.t1116 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X587 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X588 out s3 fc2.t325 fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X590 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X591 fc1 s1 VP.t1115 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X592 fc1 s1 VP.t1114 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X593 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X594 fc1 s1 VP.t1113 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X595 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X596 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X597 fc1 s1 VP.t1112 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X598 fc1 s1 VP.t1111 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X599 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X600 fc1 s1 VP.t1110 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X601 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X602 VP.t1109 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X603 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X604 VN.t331 s4 fc2.t466 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X605 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X606 fc1 s1 VP.t1108 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X607 VN.t330 s4 fc2.t551 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X608 out s3 fc2.t324 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X609 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X610 VN.t329 s4 fc2.t401 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X611 fc1 s1 VP.t1107 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X612 VP.t1106 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X613 VP.t1105 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X614 VP.t1104 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X615 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X616 VP.t1103 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X617 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X618 VN.t328 s4 fc2.t709 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X619 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X620 out s3 fc2.t323 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X621 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X622 fc1 s1 VP.t1102 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X623 fc2.t322 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X624 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X625 fc1 s1 VP.t1101 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X626 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X627 VP.t1100 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X628 VP.t1099 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X629 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X630 VN.t327 s4 fc2.t593 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X631 fc2.t321 s3 out fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X632 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X633 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X634 VP.t1098 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X635 fc1 s1 VP.t1097 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X636 fc2.t320 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X637 VP.t1096 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X638 fc1 s1 VP.t1095 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X639 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X640 VN.t326 s4 fc2.t421 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X641 VN.t325 s4 fc2.t681 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X642 out s3 fc2.t319 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X643 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X644 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X645 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X646 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X647 VN.t324 s4 fc2.t408 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X648 VP.t1094 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X649 VN.t323 s4 fc2.t591 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X650 out s3 fc2.t318 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X651 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X652 fc2.t317 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X653 fc1 s1 VP.t1093 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X654 VP.t1092 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X655 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X656 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X657 VP.t1091 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X658 fc1 s1 VP.t1090 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X659 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X660 fc1 s1 VP.t1089 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X661 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X663 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X664 VP.t1088 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X665 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X666 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X667 fc1 s1 VP.t1087 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X668 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X669 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X670 VP.t1086 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X671 fc1 s1 VP.t1085 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X672 VP.t1084 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X673 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X674 VN.t322 s4 fc2.t725 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X675 out s3 fc2.t316 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X676 fc2.t315 s3 out fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X677 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X678 fc1 s1 VP.t1083 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X679 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X680 out s3 fc2.t314 fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X681 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X682 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X683 VN.t321 s4 fc2.t728 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X684 VN.t320 s4 fc2.t726 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X685 VP.t1082 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X686 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X687 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X688 VP.t1081 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X689 fc1 s1 VP.t1080 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X690 VN.t319 s4 fc2.t705 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X691 fc1 s1 VP.t1079 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X692 fc1 s1 VP.t1078 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X693 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X694 fc1 s1 VP.t1077 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X695 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X696 fc1 s1 VP.t1076 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X697 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X698 fc1 s1 VP.t1075 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X699 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X700 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X701 VP.t1074 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X702 out s3 fc2.t313 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X703 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X704 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X705 fc2.t639 s4 VN.t318 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X706 VN.t317 s4 fc2.t628 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X707 fc1 s1 VP.t1073 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X708 VP.t1072 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X709 VP.t1071 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X710 fc2.t417 s4 VN.t316 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X711 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X712 fc1 s1 VP.t1070 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X713 fc1 s1 VP.t1069 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X714 out s3 fc2.t312 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X715 fc2.t703 s4 VN.t315 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X716 VP.t1068 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X717 fc2.t594 s4 VN.t314 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X718 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X719 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X720 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X721 VP.t1067 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X722 VP.t1066 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X723 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X724 fc2.t311 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X725 VP.t1065 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X726 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X727 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X728 fc1 s1 VP.t1064 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X729 VP.t1063 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X730 out s3 fc2.t310 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X731 VP.t1062 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X732 VP.t1061 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X733 VN.t313 s4 fc2.t590 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X734 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X735 fc1 s1 VP.t1060 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X736 fc2.t309 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X737 out s3 fc2.t308 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X739 fc2.t514 s4 VN.t312 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X740 fc1 s1 VP.t1059 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X741 fc1 s1 VP.t1058 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X742 fc2.t420 s4 VN.t311 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X743 fc1 s1 VP.t1057 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X744 VP.t1056 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X745 fc1 s1 VP.t1055 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X746 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X747 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X748 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X749 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X750 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X751 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X752 VP.t1054 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X753 fc1 s1 VP.t1053 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X754 VP.t1052 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X755 out s3 fc2.t307 fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X756 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X757 fc2.t306 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X758 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X760 fc1 s1 VP.t1051 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X761 fc2.t399 s4 VN.t310 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X762 VP.t1050 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X763 fc1 s1 VP.t1049 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X764 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X765 out s3 fc2.t305 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X766 fc2.t304 s3 out fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X767 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X768 fc1 s1 VP.t1048 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X769 fc1 s1 VP.t1047 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X770 fc1 s1 VP.t1046 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X771 VP.t1045 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X772 VN.t309 s4 fc2.t418 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X773 out s3 fc2.t303 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X774 fc2.t302 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X775 VP.t1044 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X776 VP.t1043 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X777 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X778 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X779 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X780 fc1 s1 VP.t1042 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X781 VP.t1041 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X782 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X783 fc2.t636 s4 VN.t308 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X784 fc2.t448 s4 VN.t307 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X785 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X786 VP.t1040 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X787 fc1 s1 VP.t1039 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X788 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X789 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X790 fc1 s1 VP.t1038 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X791 fc1 s1 VP.t1037 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X792 fc1 s1 VP.t1036 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X793 out s3 fc2.t301 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X794 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X795 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X796 fc1 s1 VP.t1035 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X797 VN.t306 s4 fc2.t500 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X798 fc1 s1 VP.t1034 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X799 VP.t1033 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X800 VP.t1032 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X801 VP.t1031 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X802 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X803 fc1 s1 VP.t1030 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X804 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X805 fc2.t300 s3 out fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X806 fc1 s1 VP.t1029 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X807 VP.t1028 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X808 fc1 s1 VP.t1027 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X809 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X810 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X811 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X812 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X813 fc2.t589 s4 VN.t305 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X814 fc1 s1 VP.t1026 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X815 VP.t1025 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X816 VP.t1024 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X817 VP.t1023 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X818 VP.t1022 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X819 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X820 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X821 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X822 fc1 s1 VP.t1021 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X823 VP.t1020 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X824 VP.t1019 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X825 fc2.t461 s4 VN.t304 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X826 VP.t1018 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X827 fc2.t592 s4 VN.t303 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X828 fc2.t299 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X829 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X830 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X831 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X832 fc1 s1 VP.t1017 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X833 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X834 fc1 s1 VP.t1016 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X835 VP.t1015 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X836 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X837 fc2.t746 s4 VN.t302 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X838 fc2.t510 s4 VN.t301 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X839 fc2.t298 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X840 VP.t1014 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X841 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X842 fc1 s1 VP.t1013 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X843 fc2.t297 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X844 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X845 VP.t1012 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X846 VP.t1011 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X847 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X848 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X849 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X850 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X851 fc1 s1 VP.t1010 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X852 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X853 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X854 fc1 s1 VP.t1009 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X855 fc1 s1 VP.t1008 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X856 VP.t1007 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X857 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X858 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X859 fc2.t704 s4 VN.t300 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X860 fc2.t643 s4 VN.t299 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X861 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X862 fc2.t296 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X863 fc1 s1 VP.t1006 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X864 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X865 fc2.t489 s4 VN.t298 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X866 fc1 s1 VP.t1005 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X867 fc1 s1 VP.t1004 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X868 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X869 VP.t1003 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X870 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X871 fc2.t395 s4 VN.t297 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X872 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X873 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X874 fc1 s1 VP.t1002 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X875 out s3 fc2.t295 fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X876 out s3 fc2.t294 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X877 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X878 fc1 s1 VP.t1001 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X879 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X880 VP.t1000 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X881 fc1 s1 VP.t999 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X882 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X883 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X884 VN.t296 s4 fc2.t419 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X885 VP.t998 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X886 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X887 fc1 s1 VP.t997 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X888 fc1 s1 VP.t996 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X889 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X890 out s3 fc2.t293 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X891 VN.t295 s4 fc2.t682 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X892 out s3 fc2.t292 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X894 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X895 VP.t995 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X896 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X897 fc2.t483 s4 VN.t294 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X898 fc2.t400 s4 VN.t293 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X899 fc1 s1 VP.t994 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X900 fc2.t637 s4 VN.t292 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X901 fc2.t291 s3 out fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X902 fc1 s1 VP.t993 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X904 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X905 VN.t291 s4 fc2.t635 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X906 fc2.t665 s4 VN.t290 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X907 fc2.t290 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X908 VP.t992 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X909 fc1 s1 VP.t991 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X910 VP.t990 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X911 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X912 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X913 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X914 VP.t989 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X915 VP.t988 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X916 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X917 VN.t289 s4 fc2.t683 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X918 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X919 fc2.t289 s3 out fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X920 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X921 VP.t987 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X922 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X923 VN.t288 s4 fc2.t446 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X924 VP.t986 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X925 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X926 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X927 fc1 s1 VP.t985 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X928 VP.t984 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X929 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X930 VP.t983 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X931 VP.t982 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X932 out s3 fc2.t288 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X933 fc1 s1 VP.t981 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X934 VP.t980 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X935 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X936 fc2.t727 s4 VN.t287 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X937 fc2.t661 s4 VN.t286 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X938 fc2.t287 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X939 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X940 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X941 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X942 fc2.t450 s4 VN.t285 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X943 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X944 fc2.t286 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X945 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X946 VP.t979 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X947 fc1 s1 VP.t978 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X948 VP.t977 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X949 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X950 fc2.t660 s4 VN.t284 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X951 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X952 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X953 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X954 VP.t976 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X955 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X956 VP.t975 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X957 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X958 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X959 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X960 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X961 fc1 s1 VP.t974 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X962 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X963 out s3 fc2.t285 fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X964 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X965 fc1 s1 VP.t973 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X966 fc2.t284 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X967 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X968 fc1 s1 VP.t972 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X969 VN.t283 s4 fc2.t438 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X970 fc1 s1 VP.t971 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X971 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X972 VP.t970 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X973 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X974 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X975 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X976 fc1 s1 VP.t969 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X977 fc1 s1 VP.t968 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X978 fc2.t486 s4 VN.t282 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X980 fc1 s1 VP.t967 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X981 VN.t281 s4 fc2.t644 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X982 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X983 fc1 s1 VP.t966 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X984 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X985 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X986 VN.t280 s4 fc2.t670 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X987 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X988 fc1 s1 VP.t965 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X989 VN.t279 s4 fc2.t433 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X990 fc2.t283 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X991 out s3 fc2.t282 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X992 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X993 VP.t964 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X994 fc2.t281 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X995 VP.t963 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X996 fc1 s1 VP.t962 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X997 VP.t961 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X998 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X999 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1000 fc1 s1 VP.t960 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1001 out s3 fc2.t280 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1002 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1003 fc1 s1 VP.t959 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1004 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1005 VP.t958 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1007 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1008 VP.t957 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1009 fc2.t716 s4 VN.t278 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1010 fc2.t279 s3 out fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1011 out s3 fc2.t278 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X1012 fc2.t277 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1013 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1014 fc1 s1 VP.t956 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1015 fc1 s1 VP.t955 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1016 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1017 VP.t954 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1018 VN.t277 s4 fc2.t638 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1019 fc1 s1 VP.t953 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1020 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1021 fc1 s1 VP.t952 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1022 VP.t951 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1023 out s3 fc2.t276 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1024 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1025 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1026 VP.t950 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1027 VP.t949 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1028 fc2.t275 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1029 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1030 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1031 VP.t948 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1032 VP.t947 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1033 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1034 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1035 fc1 s1 VP.t946 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1036 VP.t945 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1037 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1038 out s3 fc2.t274 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1039 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1040 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1041 VP.t944 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1042 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1043 out s3 fc2.t273 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1044 VP.t943 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1045 fc2.t272 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1047 fc2.t271 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1048 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1049 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1050 fc1 s1 VP.t942 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1051 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1052 VN.t276 s4 fc2.t564 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1053 VN.t275 s4 fc2.t396 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1054 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1055 VP.t941 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1056 fc1 s1 VP.t940 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1057 VP.t939 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1058 fc2.t270 s3 out fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1059 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1060 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1061 VN.t274 s4 fc2.t686 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1062 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1063 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1064 fc1 s1 VP.t938 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1065 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1066 VP.t937 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1068 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1069 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1070 fc1 s1 VP.t936 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1071 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1072 VN.t273 s4 fc2.t459 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1073 out s3 fc2.t269 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1074 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1075 fc1 s1 VP.t935 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1076 VP.t934 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1077 fc1 s1 VP.t933 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1078 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1079 fc1 s1 VP.t932 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1080 VP.t931 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1081 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1082 fc1 s1 VP.t930 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1083 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1084 VN.t272 s4 fc2.t454 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1085 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1086 fc1 s1 VP.t929 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1088 VN.t271 s4 fc2.t659 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1089 fc2.t268 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1090 VP.t928 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1091 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1092 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1093 out s3 fc2.t267 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1094 fc1 s1 VP.t927 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1095 VP.t926 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1096 fc1 s1 VP.t925 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1097 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1098 out s3 fc2.t266 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1099 VN.t270 s4 fc2.t455 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1100 fc1 s1 VP.t924 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1101 VP.t923 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1102 fc1 s1 VP.t922 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1103 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1104 VP.t921 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1105 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1106 VN.t269 s4 fc2.t398 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1107 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1108 fc1 s1 VP.t920 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1109 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1110 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1111 VP.t919 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1112 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1113 VP.t918 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1114 VP.t917 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1116 VP.t916 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1117 VP.t915 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1118 VP.t914 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1119 fc2.t265 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1120 out s3 fc2.t264 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1121 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1122 VP.t913 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1123 fc1 s1 VP.t912 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1124 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1125 fc1 s1 VP.t911 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1126 fc1 s1 VP.t910 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1127 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1128 fc1 s1 VP.t909 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1129 VP.t908 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1130 VP.t907 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1131 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1132 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1133 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1134 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1136 fc2.t263 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1137 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1138 VP.t906 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1139 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1140 fc1 s1 VP.t905 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1141 fc1 s1 VP.t904 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1142 VP.t903 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1143 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1144 fc1 s1 VP.t902 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1145 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1146 fc2.t262 s3 out fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1147 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1148 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1149 VN.t268 s4 fc2.t465 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1150 out s3 fc2.t261 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1151 fc1 s1 VP.t901 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1152 VP.t900 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1153 fc1 s1 VP.t899 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1154 VN.t267 s4 fc2.t512 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1155 VP.t898 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1156 VP.t897 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1157 out s3 fc2.t260 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1158 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1159 fc1 s1 VP.t896 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1160 VP.t895 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1161 fc1 s1 VP.t894 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1162 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1163 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1164 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1165 fc1 s1 VP.t893 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1166 fc1 s1 VP.t892 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1167 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1168 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1169 fc1 s1 VP.t891 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1170 VP.t890 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1171 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1172 fc1 s1 VP.t889 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1173 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1174 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1175 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1176 fc1 s1 VP.t888 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1177 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1178 fc1 s1 VP.t887 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1179 VP.t886 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1180 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1181 VP.t885 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1182 fc1 s1 VP.t884 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1183 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1184 fc2.t259 s3 out fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1185 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1186 VP.t883 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1187 fc1 s1 VP.t882 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1188 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1189 out s3 fc2.t258 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1190 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1191 fc2.t583 s4 VN.t266 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1192 VN.t265 s4 fc2.t462 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1193 fc1 s1 VP.t881 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1194 fc2.t497 s4 VN.t264 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1195 VP.t880 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1196 VP.t879 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1197 VP.t878 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1198 VP.t877 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1199 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1200 VP.t876 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1201 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1202 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1203 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1204 VP.t875 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1205 VP.t874 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1206 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1208 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1209 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1210 fc2.t257 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1211 VP.t873 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1212 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1213 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1214 fc1 s1 VP.t872 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1215 VP.t871 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1216 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1217 VP.t870 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1218 fc2.t256 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1219 fc1 s1 VP.t869 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1220 fc2.t685 s4 VN.t263 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1221 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1222 fc1 s1 VP.t868 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1223 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1224 fc1 s1 VP.t867 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1225 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1226 fc2.t443 s4 VN.t262 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1227 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1228 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1229 VP.t866 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1230 fc1 s1 VP.t865 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1231 VP.t864 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1232 out s3 fc2.t255 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X1233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1234 fc2.t579 s4 VN.t261 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1235 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1236 fc2.t254 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1237 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1238 VP.t863 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1239 fc1 s1 VP.t862 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1240 fc1 s1 VP.t861 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1241 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1242 out s3 fc2.t253 fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1243 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1244 VP.t860 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1245 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1246 fc1 s1 VP.t859 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1247 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1248 fc1 s1 VP.t858 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1249 VP.t857 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1250 fc1 s1 VP.t856 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1251 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1252 VN.t260 s4 fc2.t457 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1253 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1254 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1255 fc2.t252 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1256 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1257 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1258 fc1 s1 VP.t855 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1259 out s3 fc2.t251 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1260 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1261 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1262 fc2.t442 s4 VN.t259 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1263 VP.t854 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1264 out s3 fc2.t250 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1265 VP.t853 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1266 VP.t852 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1267 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1268 fc1 s1 VP.t851 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1269 VN.t258 s4 fc2.t449 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1270 fc2.t249 s3 out fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1271 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1272 fc1 s1 VP.t850 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1273 fc1 s1 VP.t849 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1274 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1275 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1276 VN.t257 s4 fc2.t440 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1278 fc1 s1 VP.t848 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1279 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1280 VP.t847 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1281 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1282 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1283 fc2.t248 s3 out fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1284 VP.t846 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1285 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1286 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1287 fc2.t715 s4 VN.t256 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1288 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1289 VP.t845 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1290 fc2.t247 s3 out fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1291 fc2.t246 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1292 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1293 VP.t844 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1295 fc2.t458 s4 VN.t255 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1296 fc1 s1 VP.t843 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1297 VP.t842 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1298 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1299 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1300 VP.t841 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1301 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1302 fc1 s1 VP.t840 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1303 fc2.t487 s4 VN.t254 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1304 out s3 fc2.t245 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1305 VP.t839 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1306 VN.t253 s4 fc2.t511 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1307 fc2.t244 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1308 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1309 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1310 fc2.t496 s4 VN.t252 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1311 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1312 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1313 fc2.t243 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1314 VN.t251 s4 fc2.t451 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1315 VP.t838 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1316 fc1 s1 VP.t837 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1317 VP.t836 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1318 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1319 fc2.t447 s4 VN.t250 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1320 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1321 VP.t835 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1322 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1323 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1324 VP.t834 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1325 VP.t833 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X1326 fc1 s1 VP.t832 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1327 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1328 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1329 VP.t831 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1330 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1331 out s3 fc2.t242 fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1332 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1333 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1334 fc1 s1 VP.t830 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1335 fc2.t473 s4 VN.t249 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1336 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1337 VP.t829 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1338 fc1 s1 VP.t828 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1339 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1340 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1341 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1342 fc1 s1 VP.t827 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1343 fc1 s1 VP.t826 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1344 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1345 VN.t248 s4 fc2.t435 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1346 out s3 fc2.t241 fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1347 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1348 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1349 fc1 s1 VP.t825 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1350 fc1 s1 VP.t824 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1351 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1352 fc1 s1 VP.t823 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1353 fc2.t750 s4 VN.t247 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1354 fc2.t240 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1355 fc1 s1 VP.t822 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1356 VP.t821 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1357 fc2.t239 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1358 VP.t820 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1359 fc1 s1 VP.t819 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1360 VP.t818 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X1361 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1362 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1363 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1364 out s3 fc2.t238 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1365 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1366 fc1 s1 VP.t817 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1367 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X1368 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1369 fc1 s1 VP.t816 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1370 VP.t815 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1371 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1372 VP.t814 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1373 VP.t813 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1374 out s3 fc2.t237 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1375 VN.t246 s4 fc2.t460 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1376 fc2.t236 s3 out fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1377 fc2.t235 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1378 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1379 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1380 fc1 s1 VP.t812 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1381 fc1 s1 VP.t811 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1382 VP.t810 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1383 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1384 VN.t245 s4 fc2.t587 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1385 fc1 s1 VP.t809 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1386 VP.t808 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1387 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1388 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1389 VP.t807 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1390 fc2.t234 s3 out fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1391 out s3 fc2.t233 fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1392 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1393 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1394 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1395 VP.t806 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1396 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1397 fc2.t232 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1398 VP.t805 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1399 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1400 VP.t804 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1401 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1402 fc2.t669 s4 VN.t244 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1403 fc1 s1 VP.t803 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1404 VP.t802 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1405 out s3 fc2.t231 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1406 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1407 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1408 VP.t801 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1409 fc1 s1 VP.t800 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1410 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1411 fc2.t508 s4 VN.t243 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1412 VP.t799 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1413 fc2.t230 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1414 fc2.t229 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1415 VN.t242 s4 fc2.t464 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1416 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1417 fc1 s1 VP.t798 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1418 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1419 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1420 fc1 s1 VP.t797 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1421 fc2.t453 s4 VN.t241 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1422 VN.t240 s4 fc2.t422 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1423 VP.t796 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1424 fc1 s1 VP.t795 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1425 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1426 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1427 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1428 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1429 VN.t239 s4 fc2.t444 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1430 fc1 s1 VP.t794 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1431 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1432 fc1 s1 VP.t793 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1433 VP.t792 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1434 VP.t791 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1435 fc2.t228 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1436 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1437 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1438 VN.t238 s4 fc2.t436 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1439 out s3 fc2.t227 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1440 fc1 s1 VP.t790 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1441 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1442 VP.t789 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1443 VN.t237 s4 fc2.t581 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1444 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1445 fc1 s1 VP.t788 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1446 VP.t787 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1447 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1448 fc1 s1 VP.t786 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1449 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1450 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1451 fc2.t414 s4 VN.t236 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1452 fc1 s1 VP.t785 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1453 fc1 s1 VP.t784 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1454 VP.t783 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1455 fc2.t226 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1456 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1457 out s3 fc2.t225 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1458 fc1 s1 VP.t782 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1459 fc1 s1 VP.t781 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1460 VP.t780 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1461 fc1 s1 VP.t779 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1462 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1463 out s3 fc2.t224 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1464 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1465 VP.t778 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1466 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1467 VP.t777 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1468 fc1 s1 VP.t776 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1469 VN.t235 s4 fc2.t432 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1470 fc1 s1 VP.t775 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1471 VP.t774 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1472 fc1 s1 VP.t773 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1473 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1474 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1475 out s3 fc2.t223 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1476 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1477 fc2.t222 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1478 VP.t772 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1479 VP.t771 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1480 fc1 s1 VP.t770 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1481 fc2.t582 s4 VN.t234 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1482 out s3 fc2.t221 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1483 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1484 VP.t769 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1485 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1486 fc2.t220 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1487 VP.t768 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1488 VP.t767 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1489 VP.t766 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1490 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1491 fc2.t415 s4 VN.t233 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1492 VP.t765 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1493 VP.t764 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1494 out s3 fc2.t219 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1495 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1496 fc1 s1 VP.t763 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1497 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1498 VP.t762 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1499 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1500 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1501 fc1 s1 VP.t761 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1502 fc1 s1 VP.t760 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1503 VP.t759 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1504 VP.t758 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1505 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1506 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1507 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1508 fc2.t751 s4 VN.t232 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1509 out s3 fc2.t218 fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1510 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1511 fc2.t217 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1512 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1513 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1514 VP.t757 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1515 fc2.t445 s4 VN.t231 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1516 VN.t230 s4 fc2.t474 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1517 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1518 fc1 s1 VP.t756 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1519 fc1 s1 VP.t755 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1520 VP.t754 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1521 fc1 s1 VP.t753 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1522 fc1 s1 VP.t752 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1523 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1524 fc2.t216 s3 out fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1525 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1526 fc2.t397 s4 VN.t229 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1527 out s3 fc2.t215 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1528 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1529 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1530 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1531 VP.t751 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1532 fc1 s1 VP.t750 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1533 fc2.t684 s4 VN.t228 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1534 VN.t227 s4 fc2.t492 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1535 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1536 VP.t749 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1537 VP.t748 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1538 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1539 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1540 fc1 s1 VP.t747 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1541 VP.t746 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1542 fc1 s1 VP.t745 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1543 VP.t744 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1544 out s3 fc2.t214 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1545 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1546 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1547 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1548 fc1 s1 VP.t743 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1549 fc1 s1 VP.t742 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1550 fc1 s1 VP.t741 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1551 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1552 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1553 VN.t226 s4 fc2.t467 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1554 VP.t740 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1555 VP.t739 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1556 fc1 s1 VP.t738 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1557 out s3 fc2.t213 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1558 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1559 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1560 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1561 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1562 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1563 fc1 s1 VP.t737 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1564 VP.t736 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1565 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1566 VP.t735 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1567 fc1 s1 VP.t734 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1568 fc1 s1 VP.t733 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1569 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1570 fc1 s1 VP.t732 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1571 fc2.t212 s3 out fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1572 fc1 s1 VP.t731 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1573 fc2.t434 s4 VN.t225 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1574 out s3 fc2.t211 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1575 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1576 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1577 fc2.t641 s4 VN.t224 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1578 fc1 s1 VP.t730 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1579 VN.t223 s4 fc2.t552 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1580 VP.t729 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1581 fc2.t586 s4 VN.t222 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1582 VP.t728 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1583 fc1 s1 VP.t727 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1584 VP.t726 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1585 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1586 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1587 VP.t725 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1588 VP.t724 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1590 fc1 s1 VP.t723 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1591 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1592 VP.t722 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1593 fc1 s1 VP.t721 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1594 VP.t720 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1595 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1596 VP.t719 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1597 VP.t718 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1598 fc1 s1 VP.t717 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1599 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1600 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1601 VP.t716 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1602 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1603 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1604 fc2.t210 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1605 fc1 s1 VP.t715 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1606 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1607 fc1 s1 VP.t714 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1608 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1609 fc2.t209 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1610 VP.t713 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1611 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1612 fc1 s1 VP.t712 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1613 fc1 s1 VP.t711 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1614 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1615 VP.t710 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1616 fc1 s1 VP.t709 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1618 fc2.t566 s4 VN.t221 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1619 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1620 VP.t708 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1622 fc2.t394 s4 VN.t220 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1623 out s3 fc2.t208 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1624 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1625 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1626 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1627 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1628 fc1 s1 VP.t707 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1629 fc1 s1 VP.t706 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1630 fc1 s1 VP.t705 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1631 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1632 out s3 fc2.t207 fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1633 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1634 VP.t704 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1635 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1636 fc2.t717 s4 VN.t219 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1637 out s3 fc2.t206 fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1638 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1639 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1640 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1641 fc1 s1 VP.t703 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1642 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1643 VP.t702 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1644 fc1 s1 VP.t701 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1645 fc1 s1 VP.t700 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1646 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1647 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1648 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1649 VN.t218 s4 fc2.t423 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1650 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1651 fc1 s1 VP.t699 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1652 VP.t698 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1653 fc2.t666 s4 VN.t217 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1654 out s3 fc2.t205 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1655 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1656 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1657 VP.t697 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1658 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X1659 VP.t696 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1660 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1661 VP.t695 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1663 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1664 fc1 s1 VP.t694 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1665 VP.t693 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1666 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1667 fc1 s1 VP.t692 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1668 fc2.t204 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1669 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1670 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1671 fc1 s1 VP.t691 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1672 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1673 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1674 fc1 s1 VP.t690 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1675 VP.t689 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1676 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1677 VN.t216 s4 fc2.t748 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1678 VP.t688 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1679 fc2.t203 s3 out fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1680 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1681 fc1 s1 VP.t687 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1682 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1683 fc2.t488 s4 VN.t215 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1684 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1685 VN.t214 s4 fc2.t584 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1686 fc2.t202 s3 out fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1687 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1688 VP.t686 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1689 VN.t213 s4 fc2.t747 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1690 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1691 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1692 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1693 VP.t685 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1694 VN.t212 s4 fc2.t753 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1695 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1696 VP.t684 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1697 VN.t211 s4 fc2.t696 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1698 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1699 VP.t683 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1700 fc2.t201 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1701 fc2.t498 s4 VN.t210 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1702 VP.t682 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1703 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1704 fc1 s1 VP.t681 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1705 VP.t680 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1706 fc1 s1 VP.t679 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1707 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1708 VP.t678 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1709 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1710 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1711 fc2.t499 s4 VN.t209 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1712 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1713 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1714 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1715 fc1 s1 VP.t677 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1716 VP.t676 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1717 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1718 fc1 s1 VP.t675 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1719 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1720 VP.t674 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1721 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1722 out s3 fc2.t200 fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1723 out s3 fc2.t199 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1724 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1725 VN.t208 s4 fc2.t697 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1726 fc2.t198 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1727 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1728 VN.t207 s4 fc2.t710 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1729 VP.t673 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1730 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1731 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1732 fc1 s1 VP.t672 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1733 out s3 fc2.t197 fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1734 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1735 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1736 fc1 s1 VP.t671 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1737 fc1 s1 VP.t670 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1739 fc1 s1 VP.t669 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1740 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1741 fc1 s1 VP.t668 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1742 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1743 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1744 VP.t667 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1745 fc1 s1 VP.t666 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1746 fc2.t196 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1747 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1748 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1749 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1750 out s3 fc2.t195 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1751 VN.t206 s4 fc2.t711 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1752 out s3 fc2.t194 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1753 VN.t205 s4 fc2.t749 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1754 VP.t665 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1755 VN.t204 s4 fc2.t484 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1756 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1757 fc1 s1 VP.t664 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1758 VP.t663 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1759 VP.t662 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1760 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1761 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1762 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1763 VP.t661 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1764 VN.t203 s4 fc2.t588 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1765 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1766 out s3 fc2.t193 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1767 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1768 fc1 s1 VP.t660 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1769 fc2.t192 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1770 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1771 fc1 s1 VP.t659 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1772 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1773 VP.t658 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1774 fc2.t437 s4 VN.t202 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1775 VP.t657 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1776 VN.t201 s4 fc2.t490 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1777 fc2.t191 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1778 fc2.t190 s3 out fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1779 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1780 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1781 VP.t656 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1782 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1783 VP.t655 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1784 fc1 s1 VP.t654 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1785 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1786 VN.t200 s4 fc2.t595 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1787 fc1 s1 VP.t653 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1788 VN.t199 s4 fc2.t513 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1789 out s3 fc2.t189 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1790 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1791 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1792 fc1 s1 VP.t652 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1793 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1794 VN.t198 s4 fc2.t463 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1795 fc2.t491 s4 VN.t197 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1796 VN.t196 s4 fc2.t652 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1797 VP.t651 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1798 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1799 fc2.t188 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1800 fc1 s1 VP.t650 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1801 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1802 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1803 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1804 VP.t649 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1805 fc1 s1 VP.t648 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1806 VP.t647 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1807 fc1 s1 VP.t646 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1808 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1809 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1810 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1811 VN.t195 s4 fc2.t605 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1812 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1813 VP.t645 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1814 fc1 s1 VP.t644 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1815 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1816 VP.t643 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1817 fc1 s1 VP.t642 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1818 VP.t641 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1819 fc2.t187 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1820 VN.t194 s4 fc2.t543 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1821 out s3 fc2.t186 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1822 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1823 fc1 s1 VP.t640 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1824 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1825 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1826 fc2.t694 s4 VN.t193 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1827 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1828 VP.t639 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1829 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1830 fc1 s1 VP.t638 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1831 fc1 s1 VP.t637 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1832 fc1 s1 VP.t636 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1833 fc2.t185 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1834 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1835 fc1 s1 VP.t635 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1836 fc1 s1 VP.t634 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1837 fc1 s1 VP.t633 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1838 fc1 s1 VP.t632 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1839 VP.t631 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X1840 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1841 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1842 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1843 out s3 fc2.t184 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1844 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1845 VP.t630 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1846 VP.t629 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1847 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1848 fc1 s1 VP.t628 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1849 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1850 VN.t192 s4 fc2.t528 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1851 VP.t627 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1852 VP.t626 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1853 fc1 s1 VP.t625 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1854 fc2.t574 s4 VN.t191 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1855 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1856 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1857 fc1 s1 VP.t624 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1858 out s3 fc2.t183 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1859 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1860 fc2.t182 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1861 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1862 fc2.t456 s4 VN.t190 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1863 VP.t623 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1864 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1865 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1866 out s3 fc2.t181 fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1867 VP.t622 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1868 fc2.t441 s4 VN.t189 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1869 fc2.t180 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1870 VP.t621 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1871 VP.t620 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1872 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1873 VP.t619 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1874 fc2.t599 s4 VN.t188 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1875 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1876 fc1 s1 VP.t618 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1877 VP.t617 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1878 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1879 fc1 s1 VP.t616 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1880 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1881 fc1 s1 VP.t615 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1882 VP.t614 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1883 VP.t613 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1884 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1885 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1886 VN.t187 s4 fc2.t742 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1887 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1888 fc2.t741 s4 VN.t186 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1889 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1890 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1891 fc2.t179 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1892 fc2.t664 s4 VN.t185 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1894 fc1 s1 VP.t612 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1895 fc1 s1 VP.t611 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1896 fc1 s1 VP.t610 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1897 fc2.t544 s4 VN.t184 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1898 VP.t609 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1899 VP.t608 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1900 fc1 s1 VP.t607 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1901 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1902 fc1 s1 VP.t606 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1903 out s3 fc2.t178 fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1904 fc2.t177 s3 out fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1905 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1906 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1907 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1908 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1909 VP.t605 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1910 fc1 s1 VP.t604 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1911 VN.t183 s4 fc2.t708 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1912 VP.t603 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1913 VP.t602 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1914 fc1 s1 VP.t601 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1915 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1916 fc1 s1 VP.t600 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1917 VP.t599 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1918 out s3 fc2.t176 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1919 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1920 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1921 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1922 fc1 s1 VP.t598 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1923 fc1 s1 VP.t597 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1924 fc1 s1 VP.t596 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1925 fc1 s1 VP.t595 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1926 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1927 VN.t182 s4 fc2.t724 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1928 VP.t594 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1929 out s3 fc2.t175 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1930 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1931 VP.t593 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1932 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1933 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1934 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1935 VP.t592 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1936 fc1 s1 VP.t591 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1937 fc2.t480 s4 VN.t181 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1938 fc2.t549 s4 VN.t180 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1939 VP.t590 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1940 fc2.t550 s4 VN.t179 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1941 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1942 fc1 s1 VP.t589 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1943 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1944 fc1 s1 VP.t588 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1945 fc1 s1 VP.t587 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1946 fc2.t516 s4 VN.t178 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1947 fc2.t517 s4 VN.t177 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1948 out s3 fc2.t174 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1949 VN.t176 s4 fc2.t690 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1950 fc1 s1 VP.t586 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1951 VP.t585 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1952 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1953 VP.t584 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1954 VP.t583 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1955 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1956 fc1 s1 VP.t582 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1957 VP.t581 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1958 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1959 fc2.t173 s3 out fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1960 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1961 VP.t580 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1962 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1963 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1964 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1965 VP.t579 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1966 fc1 s1 VP.t578 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1967 VP.t577 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1968 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1969 VP.t576 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1970 VP.t575 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1971 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1972 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1973 fc1 s1 VP.t574 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1974 VP.t573 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1975 fc2.t548 s4 VN.t175 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1976 fc2.t172 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1977 fc2.t171 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1978 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1980 fc1 s1 VP.t572 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1981 fc2.t674 s4 VN.t174 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1982 fc1 s1 VP.t571 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1983 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1984 fc2.t170 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1985 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1986 VP.t570 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1987 fc1 s1 VP.t569 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1988 fc2.t630 s4 VN.t173 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1989 fc1 s1 VP.t568 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1990 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1991 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1992 VP.t567 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1993 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1994 out s3 fc2.t169 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1995 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1996 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1998 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1999 fc1 s1 VP.t566 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2000 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2001 out s3 fc2.t168 fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2002 fc1 s1 VP.t565 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2003 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2004 VP.t564 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2005 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2006 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2007 fc2.t631 s4 VN.t172 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2008 fc2.t410 s4 VN.t171 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2009 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2010 fc1 s1 VP.t563 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2011 fc2.t425 s4 VN.t170 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2012 fc2.t534 s4 VN.t169 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2013 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2014 fc1 s1 VP.t562 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2015 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2016 fc1 s1 VP.t561 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2017 fc1 s1 VP.t560 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2019 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2020 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2021 VN.t168 s4 fc2.t565 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2022 fc2.t689 s4 VN.t167 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2023 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2024 fc1 s1 VP.t559 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2025 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2026 VP.t558 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2027 out s3 fc2.t167 fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2028 out s3 fc2.t166 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2029 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2030 fc1 s1 VP.t557 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2031 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2032 VP.t556 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2033 VP.t555 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2034 fc1 s1 VP.t554 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2035 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2036 VN.t166 s4 fc2.t541 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2037 VP.t553 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2038 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2039 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2040 VN.t165 s4 fc2.t622 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2041 fc1 s1 VP.t552 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2042 out s3 fc2.t165 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2043 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2044 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2045 fc1 s1 VP.t551 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2047 VN.t164 s4 fc2.t633 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2048 out s3 fc2.t164 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2049 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2050 fc1 s1 VP.t550 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2051 VP.t549 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2052 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2053 fc2.t509 s4 VN.t163 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2054 fc2.t427 s4 VN.t162 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2055 fc2.t163 s3 out fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2056 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2057 fc1 s1 VP.t548 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2058 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2059 fc2.t718 s4 VN.t161 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2060 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2061 VN.t160 s4 fc2.t647 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2062 fc1 s1 VP.t547 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2063 fc1 s1 VP.t546 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X2064 VP.t545 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2065 VP.t544 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2066 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2068 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2069 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2070 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2071 VP.t543 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2072 VP.t542 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2073 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2074 VP.t541 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2075 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2076 VP.t540 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2077 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2078 VP.t539 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2079 VP.t538 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2080 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2081 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2082 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2083 fc1 s1 VP.t537 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2084 VP.t536 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2085 VP.t535 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2086 VP.t534 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2087 VP.t533 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2088 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2089 fc2.t521 s4 VN.t159 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2090 fc2.t162 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2091 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2092 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2093 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2094 fc1 s1 VP.t532 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2095 VN.t158 s4 fc2.t469 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2096 VP.t531 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2097 fc1 s1 VP.t530 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2098 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2099 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2100 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2101 out s3 fc2.t161 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2102 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2103 fc1 s1 VP.t529 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2104 fc1 s1 VP.t528 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2105 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2106 VP.t527 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2107 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2108 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2109 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2110 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2111 fc1 s1 VP.t526 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2112 fc1 s1 VP.t525 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2113 out s3 fc2.t160 fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2114 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2116 fc1 s1 VP.t524 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2117 fc2.t159 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2118 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2119 fc1 s1 VP.t523 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2120 VP.t522 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2121 VP.t521 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2122 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2123 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2124 fc1 s1 VP.t520 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2125 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2126 fc2.t721 s4 VN.t157 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2127 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2128 fc1 s1 VP.t519 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2129 VN.t156 s4 fc2.t470 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2130 fc2.t158 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2131 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2132 fc1 s1 VP.t518 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2133 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2134 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2135 VN.t155 s4 fc2.t407 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2136 out s3 fc2.t157 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2137 fc2.t156 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2138 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2139 fc1 s1 VP.t517 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2140 out s3 fc2.t155 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2141 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2142 VP.t516 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2143 fc1 s1 VP.t515 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2144 fc2.t154 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2145 VP.t514 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2146 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2147 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2148 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2149 fc1 s1 VP.t513 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2150 out s3 fc2.t153 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2151 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2152 fc1 s1 VP.t512 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2153 fc1 s1 VP.t511 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2154 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2155 VP.t510 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2156 VP.t509 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2157 fc2.t570 s4 VN.t154 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2158 out s3 fc2.t152 fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2159 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2160 VN.t153 s4 fc2.t482 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2161 fc2.t151 s3 out fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2162 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2163 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2164 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2165 VN.t152 s4 fc2.t735 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2166 VP.t508 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2167 fc1 s1 VP.t507 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2168 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2169 fc1 s1 VP.t506 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2170 VP.t505 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2171 out s3 fc2.t150 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2172 VP.t504 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2173 VP.t503 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2174 fc1 s1 VP.t502 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2175 fc2.t149 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2176 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2177 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2178 VP.t501 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2179 fc2.t729 s4 VN.t151 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2180 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2181 VP.t500 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2182 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2183 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2184 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2185 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2186 VP.t499 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2187 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2188 fc2.t148 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2189 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2190 VP.t498 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2191 fc1 s1 VP.t497 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2192 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2193 VN.t150 s4 fc2.t640 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2194 VP.t496 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2195 fc1 s1 VP.t495 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2196 VP.t494 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2197 fc2.t147 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2198 VN.t149 s4 fc2.t525 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2199 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2200 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2201 fc1 s1 VP.t493 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2202 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2203 fc1 s1 VP.t492 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2205 VP.t491 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2206 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2207 out s3 fc2.t146 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2208 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2209 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2210 fc1 s1 VP.t490 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2211 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2212 fc1 s1 VP.t489 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2213 VP.t488 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2214 fc2.t145 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2215 fc1 s1 VP.t487 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2216 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2217 fc1 s1 VP.t486 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2218 fc1 s1 VP.t485 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2219 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2220 VN.t148 s4 fc2.t542 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2221 out s3 fc2.t144 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2222 fc1 s1 VP.t484 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2223 VP.t483 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2224 VN.t147 s4 fc2.t740 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X2225 VN.t146 s4 fc2.t699 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2226 out s3 fc2.t143 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2227 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2228 VP.t482 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2229 VP.t481 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2230 VP.t480 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2231 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2232 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2233 fc1 s1 VP.t479 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2234 VP.t478 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2235 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2236 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2237 fc1 s1 VP.t477 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2238 out s3 fc2.t142 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2239 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2240 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2241 fc2.t141 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2242 VN.t145 s4 fc2.t621 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2243 VP.t476 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2244 fc1 s1 VP.t475 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2245 VP.t474 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2246 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2247 out s3 fc2.t140 fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2248 VP.t473 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2249 fc2.t139 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2250 VP.t472 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2251 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2252 fc2.t472 s4 VN.t144 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2253 fc1 s1 VP.t471 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X2254 VN.t143 s4 fc2.t506 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2255 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2256 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2257 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2258 fc1 s1 VP.t470 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2260 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2261 VP.t469 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2262 VP.t468 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2263 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2264 VP.t467 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2265 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X2266 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2267 VP.t466 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2268 VP.t465 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2269 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2270 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2271 VP.t464 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2272 VP.t463 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2273 fc2.t138 s3 out fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2274 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2275 VP.t462 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2276 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2277 fc1 s1 VP.t461 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2278 fc1 s1 VP.t460 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2279 fc1 s1 VP.t459 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2280 VP.t458 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2281 VP.t457 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2282 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2283 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2284 fc1 s1 VP.t456 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2285 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2286 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2287 fc2.t137 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2288 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2289 VP.t455 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2290 VN.t142 s4 fc2.t672 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2291 VP.t454 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2292 fc1 s1 VP.t453 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2293 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2294 fc1 s1 VP.t452 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2295 fc1 s1 VP.t451 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X2296 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2297 fc1 s1 VP.t450 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2298 out s3 fc2.t136 fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2299 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2300 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2301 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2302 fc1 s1 VP.t449 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2303 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2304 fc1 s1 VP.t448 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2305 fc1 s1 VP.t447 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2306 VN.t141 s4 fc2.t507 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2307 VP.t446 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2308 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X2309 fc2.t616 s4 VN.t140 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2310 out s3 fc2.t135 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2311 VP.t445 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2312 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2313 fc1 s1 VP.t444 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2314 VP.t443 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2315 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2316 fc1 s1 VP.t442 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2317 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2318 fc1 s1 VP.t441 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2319 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2320 VP.t440 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2321 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2322 fc1 s1 VP.t439 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2323 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2324 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2325 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2326 fc1 s1 VP.t438 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2327 VP.t437 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2328 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2329 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2330 VP.t436 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2331 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2332 fc1 s1 VP.t435 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2333 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2334 VP.t434 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2335 fc2.t134 s3 out fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2336 VP.t433 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2337 out s3 fc2.t133 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2339 fc1 s1 VP.t432 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2340 fc2.t556 s4 VN.t139 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2341 VP.t431 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2342 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2343 VP.t430 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2344 VP.t429 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2345 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2346 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2347 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2348 VP.t428 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2349 fc2.t132 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2350 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2351 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2352 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2353 fc2.t131 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2354 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2355 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2356 VP.t427 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2357 fc1 s1 VP.t426 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2358 VP.t425 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2359 fc2.t601 s4 VN.t138 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2360 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2361 VP.t424 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2362 fc1 s1 VP.t423 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2363 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2364 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2365 fc1 s1 VP.t422 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2366 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2367 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2368 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2369 fc2.t706 s4 VN.t137 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2370 fc1 s1 VP.t421 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2372 out s3 fc2.t130 fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2373 VP.t420 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2374 VP.t419 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2375 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2376 out s3 fc2.t129 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2377 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2378 fc2.t610 s4 VN.t136 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2379 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2380 fc1 s1 VP.t418 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2381 VP.t417 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2382 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2383 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2384 VN.t135 s4 fc2.t411 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2385 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2386 fc1 s1 VP.t416 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2387 fc1 s1 VP.t415 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2388 fc1 s1 VP.t414 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2389 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2390 out s3 fc2.t128 fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2391 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2392 VN.t134 s4 fc2.t722 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2393 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2394 fc1 s1 VP.t413 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2395 VP.t412 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2396 fc1 s1 VP.t411 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2397 VP.t410 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2398 fc1 s1 VP.t409 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2399 VP.t408 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2400 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2401 VP.t407 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2402 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2403 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2404 VN.t133 s4 fc2.t607 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2405 fc2.t127 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2406 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2407 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2408 fc1 s1 VP.t406 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2409 out s3 fc2.t126 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2410 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2411 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2412 VN.t132 s4 fc2.t430 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2413 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2414 fc2.t731 s4 VN.t131 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2415 fc1 s1 VP.t405 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2416 VP.t404 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2417 out s3 fc2.t125 fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2418 VP.t403 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2419 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2420 fc1 s1 VP.t402 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2421 VP.t401 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2422 VN.t130 s4 fc2.t571 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2423 fc2.t124 s3 out fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2424 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2425 fc1 s1 VP.t400 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2426 fc1 s1 VP.t399 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2427 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2428 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2429 VN.t129 s4 fc2.t495 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2430 fc1 s1 VP.t398 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2431 VP.t397 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2432 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2433 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2435 fc2.t123 s3 out fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2436 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2437 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2438 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2439 VP.t396 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2440 fc2.t693 s4 VN.t128 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2441 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2442 VP.t395 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2443 VP.t394 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2444 fc2.t122 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2445 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2446 VP.t393 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2447 VP.t392 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2448 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2449 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2450 fc1 s1 VP.t391 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2451 VP.t390 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2452 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2453 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2454 VP.t389 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2455 VP.t388 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2456 fc2.t679 s4 VN.t127 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2457 VN.t126 s4 fc2.t585 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2458 fc2.t121 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2459 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2460 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2461 VN.t125 s4 fc2.t650 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2462 VP.t387 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2463 fc1 s1 VP.t386 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2464 fc1 s1 VP.t385 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2465 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2466 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2467 VP.t384 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2468 out s3 fc2.t120 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2469 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2470 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2471 fc1 s1 VP.t383 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2472 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2473 VP.t382 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2474 fc1 s1 VP.t381 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2475 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2476 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2477 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2478 fc1 s1 VP.t380 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2479 VP.t379 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2480 out s3 fc2.t119 fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2481 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2482 fc2.t501 s4 VN.t124 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2483 fc1 s1 VP.t378 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2484 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2485 VP.t377 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2486 VP.t376 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2487 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2488 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2489 fc1 s1 VP.t375 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2490 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2491 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2492 fc1 s1 VP.t374 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2493 VN.t123 s4 fc2.t530 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2494 out s3 fc2.t118 fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2495 fc2.t117 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X2496 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2497 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2498 fc1 s1 VP.t373 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2499 out s3 fc2.t116 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2500 fc2.t115 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2502 fc1 s1 VP.t372 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2503 VN.t122 s4 fc2.t393 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2504 fc2.t680 s4 VN.t121 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2505 fc1 s1 VP.t371 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2506 VP.t370 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2507 fc2.t114 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2508 fc1 s1 VP.t369 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2509 VP.t368 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2510 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2511 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2512 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2513 VN.t120 s4 fc2.t667 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2514 out s3 fc2.t113 fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2515 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2516 fc1 s1 VP.t367 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2517 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2518 VP.t366 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2519 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2520 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2521 fc1 s1 VP.t365 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2522 fc1 s1 VP.t364 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2523 fc2.t439 s4 VN.t119 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2524 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2525 VP.t363 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2526 VP.t362 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2527 fc2.t112 s3 out fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2528 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2529 VN.t118 s4 fc2.t409 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2530 fc2.t520 s4 VN.t117 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2531 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2532 VP.t361 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2533 fc1 s1 VP.t360 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2534 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2535 VP.t359 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2536 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2537 VP.t358 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2538 VP.t357 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2539 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2540 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2541 fc1 s1 VP.t356 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2542 fc2.t111 s3 out fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X2543 VP.t355 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2544 VP.t354 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2545 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2546 fc2.t649 s4 VN.t116 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2547 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2548 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2549 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2550 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2551 VP.t353 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2552 fc1 s1 VP.t352 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2553 VN.t115 s4 fc2.t701 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2554 fc2.t110 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2555 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2556 fc1 s1 VP.t351 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2557 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2558 VP.t350 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2559 fc1 s1 VP.t349 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2560 fc2.t754 s4 VN.t114 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2561 fc2.t109 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2562 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2563 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2564 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2565 fc1 s1 VP.t348 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2566 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2567 fc1 s1 VP.t347 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2568 fc1 s1 VP.t346 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2569 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2570 fc2.t108 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2571 VP.t345 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2572 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2573 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2574 fc1 s1 VP.t344 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2575 out s3 fc2.t107 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2576 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2577 VP.t343 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2578 fc1 s1 VP.t342 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2579 VN.t113 s4 fc2.t503 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2580 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2582 fc1 s1 VP.t341 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2583 fc1 s1 VP.t340 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2584 fc1 s1 VP.t339 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2585 fc1 s1 VP.t338 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2586 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2587 out s3 fc2.t106 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2588 fc2.t105 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2590 fc1 s1 VP.t337 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2591 fc2.t608 s4 VN.t112 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2592 VN.t111 s4 fc2.t642 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2593 fc1 s1 VP.t336 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2594 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2595 out s3 fc2.t104 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2596 VP.t335 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2597 VP.t334 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2598 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2599 fc1 s1 VP.t333 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2600 fc1 s1 VP.t332 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2601 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2602 VP.t331 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2603 fc1 s1 VP.t330 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2604 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2605 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2606 out s3 fc2.t103 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2607 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2608 VP.t329 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2609 VP.t328 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2610 VP.t327 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2611 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2612 fc1 s1 VP.t326 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2613 VP.t325 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2614 VN.t110 s4 fc2.t547 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2615 fc1 s1 VP.t324 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2616 VP.t323 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2618 fc2.t102 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2619 out s3 fc2.t101 fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2620 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2621 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2622 fc1 s1 VP.t322 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2623 fc2.t100 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2624 VP.t321 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2625 fc1 s1 VP.t320 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2626 VP.t319 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2627 fc2.t546 s4 VN.t109 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2628 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2629 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2630 fc1 s1 VP.t318 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2631 fc1 s1 VP.t317 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2632 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2633 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2634 VP.t316 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2635 fc2.t688 s4 VN.t108 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2636 fc2.t99 s3 out fc2.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2637 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2638 VP.t315 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2639 VP.t314 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2640 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2641 VP.t313 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2642 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2643 VP.t312 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2644 fc2.t714 s4 VN.t107 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2645 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2646 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2647 VP.t311 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2648 VP.t310 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2649 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2650 VP.t309 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2651 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2652 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2653 fc1 s1 VP.t308 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2654 fc1 s1 VP.t307 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2655 VP.t306 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2656 VP.t305 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2657 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2658 fc2.t515 s4 VN.t106 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X2659 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2660 out s3 fc2.t97 fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2661 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2663 fc2.t96 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2664 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2665 VP.t304 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2666 VN.t105 s4 fc2.t481 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2667 fc2.t629 s4 VN.t104 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2668 VP.t303 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2669 fc1 s1 VP.t302 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2670 fc1 s1 VP.t301 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2671 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2672 fc1 s1 VP.t300 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2673 VP.t299 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2674 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2675 fc1 s1 VP.t298 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2676 fc1 s1 VP.t297 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2677 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2678 fc2.t539 s4 VN.t103 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2679 out s3 fc2.t95 fc2.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2680 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2681 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2682 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2683 fc1 s1 VP.t296 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2684 fc1 s1 VP.t295 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2685 fc2.t657 s4 VN.t102 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2686 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2687 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2688 VP.t294 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2689 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2690 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2691 fc1 s1 VP.t293 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2692 VP.t292 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2693 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2694 VP.t291 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2695 out s3 fc2.t93 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2696 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2697 fc1 s1 VP.t290 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2698 fc1 s1 VP.t289 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2699 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2700 VN.t101 s4 fc2.t524 VN.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2701 VP.t288 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2702 out s3 fc2.t92 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2703 VP.t287 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2704 fc1 s1 VP.t286 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2705 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2706 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2707 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2708 VP.t285 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2709 fc1 s1 VP.t284 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2710 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2711 VP.t283 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2712 fc1 s1 VP.t282 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2713 fc1 s1 VP.t281 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2714 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2715 VP.t280 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2716 VN.t99 s4 fc2.t572 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2717 fc2.t91 s3 out fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2718 fc2.t90 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2719 fc2.t604 s4 VN.t98 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2720 out s3 fc2.t89 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2721 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2722 fc1 s1 VP.t279 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2723 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2724 VP.t278 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2725 fc2.t614 s4 VN.t97 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2726 fc1 s1 VP.t277 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2727 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2728 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2729 VP.t276 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2730 fc2.t88 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2731 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2732 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2733 fc1 s1 VP.t275 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2734 fc1 s1 VP.t274 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2735 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2736 VP.t273 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2737 VP.t272 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2738 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2739 out s3 fc2.t87 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X2740 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2741 fc1 s1 VP.t271 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2742 VP.t270 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2743 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2744 fc2.t562 s4 VN.t96 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2745 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2746 fc1 s1 VP.t269 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2747 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2748 fc2.t86 s3 out fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2749 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2750 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2751 fc1 s1 VP.t268 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2752 VP.t267 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2753 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2754 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2755 fc1 s1 VP.t266 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2756 fc1 s1 VP.t265 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2757 fc2.t732 s4 VN.t95 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2758 VP.t264 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2760 out s3 fc2.t85 fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2761 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2762 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2763 VP.t263 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2764 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2765 out s3 fc2.t84 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2766 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2767 fc2.t632 s4 VN.t94 VN.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2768 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2769 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2770 fc1 s1 VP.t262 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2771 fc1 s1 VP.t261 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2772 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2773 out s3 fc2.t83 fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2774 fc1 s1 VP.t260 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2775 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2776 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2777 fc2.t700 s4 VN.t92 VN.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2778 out s3 fc2.t82 fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2779 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2780 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2781 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2782 fc1 s1 VP.t259 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2783 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2784 fc1 s1 VP.t258 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2785 fc1 s1 VP.t257 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2786 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2787 VP.t256 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2788 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2789 VP.t255 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2790 VN.t90 s4 fc2.t477 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2791 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2792 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2793 fc1 s1 VP.t254 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2794 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2795 VN.t89 s4 fc2.t627 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2796 out s3 fc2.t81 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2797 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2798 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2799 VN.t88 s4 fc2.t478 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2800 VN.t87 s4 fc2.t545 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2801 fc1 s1 VP.t253 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2802 VP.t252 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2803 VP.t251 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2804 VP.t250 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2805 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2806 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2807 VN.t86 s4 fc2.t625 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2808 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2809 fc1 s1 VP.t249 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2810 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2811 fc1 s1 VP.t248 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2812 fc1 s1 VP.t247 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2813 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2814 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2815 fc1 s1 VP.t246 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2816 VP.t245 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2817 VN.t85 s4 fc2.t577 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2818 fc2.t80 s3 out fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2819 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2820 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2821 VP.t244 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2822 fc2.t79 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2823 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2824 fc1 s1 VP.t243 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2825 fc2.t646 s4 VN.t84 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2826 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2827 VP.t242 s1 fc1 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2828 VP.t241 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2829 VP.t240 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2830 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2831 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2832 VN.t83 s4 fc2.t713 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2833 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2834 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2835 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2836 VN.t82 s4 fc2.t733 VN.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2837 VN.t80 s4 fc2.t561 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2838 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2839 VP.t239 s1 fc1 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2840 fc2.t78 s3 out fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2841 out s3 fc2.t77 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2842 fc1 s1 VP.t238 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2843 VP.t237 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2844 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2845 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2846 VP.t236 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2847 fc1 s1 VP.t235 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2848 fc1 s1 VP.t234 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2849 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2850 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2851 VP.t233 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2852 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2853 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2854 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2855 fc1 s1 VP.t232 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2856 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2857 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2858 VP.t231 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2859 fc1 s1 VP.t230 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2860 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2861 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2862 fc1 s1 VP.t229 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2863 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2864 VP.t228 s1 fc1 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2865 fc2.t76 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2866 out s3 fc2.t75 fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2867 out s3 fc2.t74 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2868 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2869 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2870 VN.t79 s4 fc2.t403 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2871 VN.t78 s4 fc2.t479 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2872 VP.t227 s1 fc1 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2873 VP.t226 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2874 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2875 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2876 fc1 s1 VP.t225 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2877 VN.t77 s4 fc2.t573 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2878 out s3 fc2.t73 fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2879 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2880 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2881 fc1 s1 VP.t224 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2882 fc1 s1 VP.t223 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2883 fc2.t72 s3 out fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2884 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2885 fc1 s1 VP.t222 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2886 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2887 fc1 s1 VP.t221 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2888 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2889 fc2.t71 s3 out fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2890 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2891 fc1 s1 VP.t220 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2892 VP.t219 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2894 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2895 VN.t76 s4 fc2.t698 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2896 out s3 fc2.t70 fc2.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2897 out s3 fc2.t68 fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2898 VN.t75 s4 fc2.t402 VN.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2899 VN.t73 s4 fc2.t692 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2900 VP.t218 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2901 VN.t72 s4 fc2.t597 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2902 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2903 fc1 s1 VP.t217 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2904 VP.t216 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2905 fc1 s1 VP.t215 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2906 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2907 VP.t214 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2908 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2909 fc2.t502 s4 VN.t71 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2910 VN.t70 s4 fc2.t648 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2911 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2912 VP.t213 s1 fc1 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2913 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2914 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2915 VP.t212 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2916 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2917 fc2.t654 s4 VN.t69 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2918 VP.t211 s1 fc1 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2919 fc2.t67 s3 out fc2.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2920 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2921 VP.t210 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2922 fc1 s1 VP.t209 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2923 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2924 fc2.t518 s4 VN.t68 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2925 VP.t208 s1 fc1 VP.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2926 fc1 s1 VP.t206 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2927 VN.t67 s4 fc2.t662 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2929 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2930 fc1 s1 VP.t205 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2931 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2932 fc2.t429 s4 VN.t66 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2933 VP.t204 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2934 fc1 s1 VP.t203 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2935 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2936 fc1 s1 VP.t202 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2937 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2938 VP.t201 s1 fc1 VP.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2939 VP.t199 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2940 fc2.t65 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2941 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2942 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2943 fc1 s1 VP.t198 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2944 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2945 VP.t197 s1 fc1 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2946 fc1 s1 VP.t196 VP.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2947 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2948 fc1 s1 VP.t194 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2949 VP.t193 s1 fc1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2950 fc1 s1 VP.t192 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2951 VP.t191 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2952 fc2.t64 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2953 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2954 out s3 fc2.t63 fc2.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2955 out s3 fc2.t61 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2956 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2957 fc1 s1 VP.t190 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2958 fc2.t567 s4 VN.t65 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2959 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2960 fc1 s1 VP.t189 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2961 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2962 fc1 s1 VP.t188 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2963 fc1 s1 VP.t187 VP.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2964 VP.t185 s1 fc1 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2965 fc2.t60 s3 out fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2966 out s3 fc2.t59 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2967 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2968 fc1 s1 VP.t184 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2969 VN.t64 s4 fc2.t476 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2970 fc1 s1 VP.t183 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2971 VP.t182 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2972 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2973 fc1 s1 VP.t181 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2974 VP.t180 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2975 VP.t179 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2976 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2977 fc2.t655 s4 VN.t63 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2978 fc2.t58 s3 out fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2979 fc1 s1 VP.t178 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2980 fc1 s1 VP.t177 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2981 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2982 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2983 fc1 s1 VP.t176 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2984 fc2.t493 s4 VN.t62 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X2985 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2986 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2987 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2988 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2989 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2990 VP.t175 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2991 VP.t174 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2992 VP.t173 s1 fc1 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2993 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2994 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2995 fc1 s1 VP.t172 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2996 VP.t171 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2997 VP.t170 s1 fc1 VP.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2998 VN.t61 s4 fc2.t536 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2999 fc1 s1 VP.t168 VP.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3000 VP.t166 s1 fc1 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3001 fc2.t426 s4 VN.t60 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3002 fc2.t606 s4 VN.t59 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3003 fc2.t57 s3 out fc2.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3004 out s3 fc2.t55 fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3005 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3007 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3008 fc1 s1 VP.t165 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3009 fc2.t54 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3010 fc1 s1 VP.t164 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3011 fc2.t651 s4 VN.t58 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3012 VP.t163 s1 fc1 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3013 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3014 fc1 s1 VP.t162 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3015 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3016 fc2.t53 s3 out fc2.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3017 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3018 VP.t161 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3019 VP.t160 s1 fc1 VP.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3020 VP.t158 s1 fc1 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3021 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3022 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3023 VP.t157 s1 fc1 VP.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3024 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3025 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3026 VP.t155 s1 fc1 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3027 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3028 fc1 s1 VP.t154 VP.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3029 VP.t152 s1 fc1 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3030 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3031 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3032 fc1 s1 VP.t151 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3033 VP.t150 s1 fc1 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3034 VP.t149 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3035 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3036 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3037 fc2.t531 s4 VN.t57 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3038 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3039 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3040 fc2.t51 s3 out fc2.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3041 fc2.t578 s4 VN.t56 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3042 fc2.t615 s4 VN.t55 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3043 fc1 s1 VP.t148 VP.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3044 fc1 s1 VP.t146 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3045 fc1 s1 VP.t145 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3047 fc2.t612 s4 VN.t54 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3048 fc1 s1 VP.t144 VP.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3049 VP.t142 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3050 fc1 s1 VP.t141 VP.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3051 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3052 fc2.t603 s4 VN.t53 VN.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3053 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3054 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3055 fc1 s1 VP.t139 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3056 out s3 fc2.t49 fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3057 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3058 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3059 fc1 s1 VP.t138 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3060 fc1 s1 VP.t137 VP.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3061 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3062 VP.t135 s1 fc1 VP.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3063 fc1 s1 VP.t133 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3064 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3065 VP.t132 s1 fc1 VP.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3066 out s3 fc2.t48 fc2.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3068 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3069 fc1 s1 VP.t130 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3070 fc1 s1 VP.t129 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3071 out s3 fc2.t46 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3072 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3073 VN.t51 s4 fc2.t695 VN.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3074 VP.t128 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3075 VP.t127 s1 fc1 VP.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3076 out s3 fc2.t45 fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3077 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3078 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3079 VP.t125 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3080 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3081 fc1 s1 VP.t124 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3082 fc2.t736 s4 VN.t49 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3083 fc2.t596 s4 VN.t48 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3084 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3085 VP.t123 s1 fc1 VP.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3086 fc1 s1 VP.t121 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3088 VN.t46 s4 fc2.t428 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3089 fc2.t404 s4 VN.t44 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3090 fc2.t44 s3 out fc2.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3091 out s3 fc2.t42 fc2.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3092 fc1 s1 VP.t120 VP.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3093 VP.t118 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3094 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3095 VP.t117 s1 fc1 VP.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3096 fc1 s1 VP.t115 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3097 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3098 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3099 fc2.t40 s3 out fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3101 VP.t114 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3102 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3103 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3104 VP.t113 s1 fc1 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3105 fc1 s1 VP.t112 VP.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3106 VP.t110 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3107 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3108 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3109 VP.t109 s1 fc1 VP.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3110 VP.t107 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3111 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3112 fc1 s1 VP.t106 VP.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3113 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3114 fc2.t611 s4 VN.t43 VN.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3115 out s3 fc2.t39 fc2.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3116 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3117 VP.t104 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3118 fc2.t485 s4 VN.t41 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3119 fc2.t37 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3120 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3121 fc1 s1 VP.t103 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3122 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3123 fc2.t673 s4 VN.t40 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3124 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3125 fc2.t36 s3 out fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3126 fc1 s1 VP.t102 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3127 VP.t101 s1 fc1 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3128 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3129 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3130 fc2.t623 s4 VN.t38 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3131 fc1 s1 VP.t100 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3132 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3133 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3134 VP.t99 s1 fc1 VP.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3135 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3136 out s3 fc2.t35 fc2.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3137 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3138 VN.t36 s4 fc2.t431 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3139 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3140 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3141 fc1 s1 VP.t97 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3142 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3143 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3144 out s3 fc2.t33 fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3145 fc1 s1 VP.t96 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3146 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3147 VN.t35 s4 fc2.t618 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3148 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3149 fc2.t712 s4 VN.t34 VN.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3150 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3151 VP.t95 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3152 VP.t94 s1 fc1 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X3153 fc2.t558 s4 VN.t32 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X3154 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3156 fc1 s1 VP.t93 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3157 fc2.t678 s4 VN.t31 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3158 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3159 fc1 s1 VP.t92 VP.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3160 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3161 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3162 fc1 s1 VP.t90 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3163 fc1 s1 VP.t89 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3164 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3165 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3166 VP.t88 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3167 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3168 VN.t29 s4 fc2.t617 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3169 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3170 fc1 s1 VP.t87 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3171 out s3 fc2.t32 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3172 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3173 fc1 s1 VP.t86 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3174 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3175 VP.t85 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3176 VP.t84 s1 fc1 VP.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3177 fc1 s1 VP.t82 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3178 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3179 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3180 VN.t28 s4 fc2.t752 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3181 fc1 s1 VP.t81 VP.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3182 out s3 fc2.t31 fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3183 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3184 fc1 s1 VP.t79 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3185 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3186 VN.t27 s4 fc2.t738 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3187 fc1 s1 VP.t78 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3188 VP.t77 s1 fc1 VP.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3189 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3190 VP.t75 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3191 fc2.t540 s4 VN.t25 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3192 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3193 out s3 fc2.t30 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3194 fc2.t29 s3 out fc2.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3195 fc2.t27 s3 out fc2.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3196 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3197 fc1 s1 VP.t74 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3198 fc2.t707 s4 VN.t23 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3199 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X3200 fc1 s1 VP.t73 VP.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3201 VP.t71 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3202 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3203 VN.t21 s4 fc2.t519 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3205 fc1 s1 VP.t70 VP.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3206 VP.t68 s1 fc1 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3207 VP.t67 s1 fc1 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3208 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3209 VP.t66 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3210 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3211 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3212 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3213 VP.t65 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3214 VP.t64 s1 fc1 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3215 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3216 VP.t63 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3217 out s3 fc2.t25 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3218 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3219 VP.t62 s1 fc1 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3220 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3221 out s3 fc2.t24 fc2.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3222 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3223 fc1 s1 VP.t61 VP.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3224 VP.t59 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3225 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3226 fc1 s1 VP.t58 VP.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3227 out s3 fc2.t22 fc2.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X3228 VP.t56 s1 fc1 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3229 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3230 fc2.t20 s3 out fc2.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3231 fc2.t18 s3 out fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3232 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3234 fc1 s1 VP.t55 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3235 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3236 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3237 fc1 s1 VP.t54 VP.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3238 VN.t19 s4 fc2.t505 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3239 VP.t52 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3240 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3241 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3242 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3243 out s3 fc2.t17 fc2.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3244 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3246 fc1 s1 VP.t51 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3247 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3248 VP.t50 s1 fc1 VP.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3249 VP.t48 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3250 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3251 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3252 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3253 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3254 VN.t18 s4 fc2.t739 VN.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3255 out s3 fc2.t15 fc2.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3256 fc1 s1 VP.t47 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3257 out s3 fc2.t13 fc2.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3258 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3259 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3260 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3261 fc1 s1 VP.t46 VP.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3262 fc1 s1 VP.t44 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3263 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3264 fc1 s1 VP.t43 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3265 VP.t42 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3266 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3267 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3268 VP.t41 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3269 fc1 s1 VP.t40 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3270 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3271 VN.t16 s4 fc2.t737 VN.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3272 VN.t14 s4 fc2.t569 VN.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3273 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3274 fc1 s1 VP.t39 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3275 fc2.t11 s3 out fc2.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3276 fc1 s1 VP.t38 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3278 VN.t12 s4 fc2.t600 VN.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3279 VP.t37 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3280 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3281 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3282 VN.t10 s4 fc2.t676 VN.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3283 VN.t8 s4 fc2.t602 VN.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3284 out s3 fc2.t9 fc2.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3285 fc1 s1 VP.t36 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3286 out s3 fc2.t7 fc2.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3287 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3288 VP.t35 s1 fc1 VP.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3289 fc1 s1 VP.t33 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3290 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3291 VP.t32 s1 fc1 VP.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3292 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3293 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3294 VN.t6 s4 fc2.t522 VN.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3295 fc2.t523 s4 VN.t4 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3296 fc1 s1 VP.t30 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3297 fc1 s1 VP.t29 VP.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3298 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3299 VP.t27 s1 fc1 VP.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3300 fc2.t723 s4 VN.t3 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3301 VP.t25 s1 fc1 VP.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3302 VN.t1 s4 fc2.t677 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3303 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3304 fc1 s1 VP.t23 VP.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3305 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3306 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3307 VP.t21 s1 fc1 VP.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3308 VP.t19 s1 fc1 VP.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3309 fc1 s1 VP.t17 VP.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3310 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3311 VP.t15 s1 fc1 VP.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3312 VP.t13 s1 fc1 VP.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3313 fc1 s1 VP.t11 VP.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3314 fc2.t5 s3 out fc2.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3315 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3316 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3317 out s3 fc2.t3 fc2.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3318 VP.t9 s1 fc1 VP.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3319 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3320 VP.t7 s1 fc1 VP.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3321 VP.t5 s1 fc1 VP.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3322 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3323 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3324 fc2.t1 s3 out fc2.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3325 VP.t3 s1 fc1 VP.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3326 fc1 s1 VP.t1 VP.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3327 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
R0 VP.n10125 VP.n10124 153.554
R1 VP.n776 VP.n775 153.554
R2 VP.n1765 VP.n1764 153.554
R3 VP.n2726 VP.n2725 153.554
R4 VP.n3666 VP.n3665 153.554
R5 VP.n4572 VP.n4571 153.554
R6 VP.n5467 VP.n5466 153.554
R7 VP.n6323 VP.n6322 153.554
R8 VP.n7182 VP.n7181 153.554
R9 VP.n8010 VP.n8009 153.554
R10 VP.n9685 VP.n9684 153.554
R11 VP.n8844 VP.n8843 153.554
R12 VP.n2690 VP.n2689 153.118
R13 VP.n1446 VP.n1445 153.118
R14 VP.n10974 VP.n10973 153.118
R15 VP.n9609 VP.n9608 153.118
R16 VP.n8803 VP.n8802 153.118
R17 VP.n7912 VP.n7911 153.118
R18 VP.n7080 VP.n7079 153.118
R19 VP.n6161 VP.n6160 153.118
R20 VP.n5301 VP.n5300 153.118
R21 VP.n4341 VP.n4340 153.118
R22 VP.n3424 VP.n3423 153.118
R23 VP.n349 VP.n348 153.118
R24 VP.n10206 VP.n10205 146.135
R25 VP.n10204 VP.n10203 146.135
R26 VP.n10336 VP.n10335 146.135
R27 VP.n10324 VP.n10323 146.135
R28 VP.n10306 VP.n10305 146.135
R29 VP.n10290 VP.n10289 146.135
R30 VP.n10278 VP.n10277 146.135
R31 VP.n10262 VP.n10261 146.135
R32 VP.n10250 VP.n10249 146.135
R33 VP.n10234 VP.n10233 146.135
R34 VP.n10222 VP.n10221 146.135
R35 VP.n10339 VP.n10338 146.135
R36 VP.n201 VP.n200 145.699
R37 VP.n205 VP.n204 145.699
R38 VP.n209 VP.n208 145.699
R39 VP.n213 VP.n212 145.699
R40 VP.n217 VP.n216 145.699
R41 VP.n221 VP.n220 145.699
R42 VP.n225 VP.n224 145.699
R43 VP.n229 VP.n228 145.699
R44 VP.n233 VP.n232 145.699
R45 VP.n237 VP.n236 145.699
R46 VP.n142 VP.n141 145.699
R47 VP.n241 VP.n240 145.699
R48 VP.n10960 VP.n10959 101.08
R49 VP.n9585 VP.n9584 101.08
R50 VP.n8781 VP.n8780 101.08
R51 VP.n7894 VP.n7893 101.08
R52 VP.n7058 VP.n7057 101.08
R53 VP.n6143 VP.n6142 101.08
R54 VP.n5279 VP.n5278 101.08
R55 VP.n4323 VP.n4322 101.08
R56 VP.n3402 VP.n3401 101.08
R57 VP.n2597 VP.n2596 101.08
R58 VP.n1431 VP.n1430 101.08
R59 VP.n332 VP.n331 101.08
R60 VP.n10663 VP.n10662 98.123
R61 VP.n321 VP.n320 88.439
R62 VP.n10962 VP.n10961 65.312
R63 VP.n9587 VP.n9586 65.312
R64 VP.n8783 VP.n8782 65.312
R65 VP.n7896 VP.n7895 65.312
R66 VP.n7060 VP.n7059 65.312
R67 VP.n6145 VP.n6144 65.312
R68 VP.n5281 VP.n5280 65.312
R69 VP.n4325 VP.n4324 65.312
R70 VP.n3404 VP.n3403 65.312
R71 VP.n2599 VP.n2598 65.312
R72 VP.n1433 VP.n1432 65.312
R73 VP.n334 VP.n333 65.312
R74 VP.n10666 VP.n10665 62.872
R75 VP.n9666 VP.n9665 62.872
R76 VP.n9287 VP.n9286 62.872
R77 VP.n8460 VP.n8459 62.872
R78 VP.n7621 VP.n7620 62.872
R79 VP.n6782 VP.n6781 62.872
R80 VP.n5918 VP.n5917 62.872
R81 VP.n5054 VP.n5053 62.872
R82 VP.n4148 VP.n4147 62.872
R83 VP.n3227 VP.n3226 62.872
R84 VP.n2277 VP.n2276 62.872
R85 VP.n1300 VP.n1299 62.872
R86 VP.n10670 VP.t0 14.709
R87 VP.n10964 VP.t167 14.709
R88 VP.n9670 VP.t31 14.709
R89 VP.n9589 VP.t153 14.709
R90 VP.n9291 VP.t156 14.709
R91 VP.n8785 VP.t4 14.709
R92 VP.n8464 VP.t200 14.709
R93 VP.n7898 VP.t10 14.709
R94 VP.n7625 VP.t2 14.709
R95 VP.n7062 VP.t136 14.709
R96 VP.n6786 VP.t122 14.709
R97 VP.n6147 VP.t186 14.709
R98 VP.n5922 VP.t14 14.709
R99 VP.n5283 VP.t22 14.709
R100 VP.n5058 VP.t131 14.709
R101 VP.n4327 VP.t105 14.709
R102 VP.n4152 VP.t20 14.709
R103 VP.n3406 VP.t12 14.709
R104 VP.n3231 VP.t83 14.709
R105 VP.n2601 VP.t60 14.709
R106 VP.n2281 VP.t98 14.709
R107 VP.n1435 VP.t80 14.709
R108 VP.n1304 VP.t45 14.709
R109 VP.n337 VP.t69 14.709
R110 VP.t6 VP.n10436 14.219
R111 VP.t16 VP.n10976 14.219
R112 VP.t126 VP.n9814 14.219
R113 VP.t143 VP.n9611 14.219
R114 VP.t207 VP.n9050 14.219
R115 VP.t28 VP.n8805 14.219
R116 VP.t18 VP.n8212 14.219
R117 VP.t111 VP.n7914 14.219
R118 VP.t134 VP.n7355 14.219
R119 VP.t195 VP.n7082 14.219
R120 VP.t159 VP.n6502 14.219
R121 VP.t24 VP.n6163 14.219
R122 VP.t26 VP.n5617 14.219
R123 VP.t119 VP.n5303 14.219
R124 VP.t169 VP.n4728 14.219
R125 VP.t140 VP.n4343 14.219
R126 VP.t76 VP.n3793 14.219
R127 VP.t72 VP.n3426 14.219
R128 VP.t108 VP.n2848 14.219
R129 VP.t91 VP.n2587 14.219
R130 VP.t53 VP.n1867 14.219
R131 VP.t34 VP.n1448 14.219
R132 VP.t49 VP.n880 14.219
R133 VP.t57 VP.n351 14.219
R134 VP.t116 VP.n202 14.219
R135 VP.n322 VP.n321 10.138
R136 VP.n2690 VP.t385 6.541
R137 VP.n2588 VP.t103 6.541
R138 VP.n2843 VP.n2842 6.541
R139 VP.n2846 VP.t596 6.541
R140 VP.n2838 VP.n2837 6.541
R141 VP.n2821 VP.t1114 6.541
R142 VP.n3393 VP.n3392 6.541
R143 VP.n3396 VP.t277 6.541
R144 VP.n3388 VP.n3387 6.541
R145 VP.n3372 VP.t1332 6.541
R146 VP.n3788 VP.n3787 6.541
R147 VP.n3791 VP.t1194 6.541
R148 VP.n3783 VP.n3782 6.541
R149 VP.n3761 VP.t770 6.541
R150 VP.n4312 VP.n4311 6.541
R151 VP.n4315 VP.t632 6.541
R152 VP.n4307 VP.n4306 6.541
R153 VP.n4293 VP.t372 6.541
R154 VP.n4687 VP.n4686 6.541
R155 VP.n4690 VP.t229 6.541
R156 VP.n4682 VP.n4681 6.541
R157 VP.n4667 VP.t23 6.541
R158 VP.n5217 VP.n5216 6.541
R159 VP.n5220 VP.t1224 6.541
R160 VP.n5212 VP.n5211 6.541
R161 VP.n5199 VP.t965 6.541
R162 VP.n5582 VP.n5581 6.541
R163 VP.n5585 VP.t974 6.541
R164 VP.n5577 VP.n5576 6.541
R165 VP.n5562 VP.t587 6.541
R166 VP.n6082 VP.n6081 6.541
R167 VP.n6085 VP.t450 6.541
R168 VP.n6077 VP.n6076 6.541
R169 VP.n6064 VP.t406 6.541
R170 VP.n6438 VP.n6437 6.541
R171 VP.n6441 VP.t261 6.541
R172 VP.n6433 VP.n6432 6.541
R173 VP.n6418 VP.t1184 6.541
R174 VP.n6946 VP.n6945 6.541
R175 VP.n6949 VP.t1049 6.541
R176 VP.n6941 VP.n6940 6.541
R177 VP.n6928 VP.t996 6.541
R178 VP.n7297 VP.n7296 6.541
R179 VP.n7300 VP.t861 6.541
R180 VP.n7292 VP.n7291 6.541
R181 VP.n7277 VP.t485 6.541
R182 VP.n7784 VP.n7783 6.541
R183 VP.n7787 VP.t348 6.541
R184 VP.n7779 VP.n7778 6.541
R185 VP.n7766 VP.t289 6.541
R186 VP.n8125 VP.n8124 6.541
R187 VP.n8128 VP.t145 6.541
R188 VP.n8120 VP.n8119 6.541
R189 VP.n8105 VP.t1076 6.541
R190 VP.n8623 VP.n8622 6.541
R191 VP.n8626 VP.t938 6.541
R192 VP.n8618 VP.n8617 6.541
R193 VP.n8605 VP.t892 6.541
R194 VP.n8969 VP.n8968 6.541
R195 VP.n8972 VP.t755 6.541
R196 VP.n8964 VP.n8963 6.541
R197 VP.n8949 VP.t371 6.541
R198 VP.n9422 VP.n9421 6.541
R199 VP.n9425 VP.t378 6.541
R200 VP.n9417 VP.n9416 6.541
R201 VP.n9402 VP.t189 6.541
R202 VP.n10760 VP.n10759 6.541
R203 VP.n10763 VP.t971 6.541
R204 VP.n10755 VP.n10754 6.541
R205 VP.n10747 VP.t707 6.541
R206 VP.n10166 VP.n10165 6.541
R207 VP.n10169 VP.t1182 6.541
R208 VP.n10161 VP.n10160 6.541
R209 VP.n10152 VP.t405 6.541
R210 VP.n10354 VP.t868 6.541
R211 VP.n1446 VP.t234 6.541
R212 VP.n2245 VP.n2244 6.541
R213 VP.n2265 VP.t449 6.541
R214 VP.n2268 VP.t972 6.541
R215 VP.n2248 VP.n2247 6.541
R216 VP.n2332 VP.n2331 6.541
R217 VP.n2343 VP.t115 6.541
R218 VP.n2340 VP.t1183 6.541
R219 VP.n2335 VP.n2334 6.541
R220 VP.n3196 VP.n3195 6.541
R221 VP.n3215 VP.t1047 6.541
R222 VP.n3218 VP.t869 6.541
R223 VP.n3199 VP.n3198 6.541
R224 VP.n3359 VP.n3358 6.541
R225 VP.n3369 VP.t727 6.541
R226 VP.n3366 VP.t484 6.541
R227 VP.n3362 VP.n3361 6.541
R228 VP.n4087 VP.n4086 6.541
R229 VP.n4107 VP.t346 6.541
R230 VP.n4110 VP.t1216 6.541
R231 VP.n4090 VP.n4089 6.541
R232 VP.n4280 VP.n4279 6.541
R233 VP.n4290 VP.t1075 6.541
R234 VP.n4287 VP.t823 6.541
R235 VP.n4283 VP.n4282 6.541
R236 VP.n4970 VP.n4969 6.541
R237 VP.n4990 VP.t675 6.541
R238 VP.n4993 VP.t439 6.541
R239 VP.n4973 VP.n4972 6.541
R240 VP.n5186 VP.n5185 6.541
R241 VP.n5196 VP.t297 6.541
R242 VP.n5193 VP.t87 6.541
R243 VP.n5189 VP.n5188 6.541
R244 VP.n5807 VP.n5806 6.541
R245 VP.n5827 VP.t97 6.541
R246 VP.n5830 VP.t1036 6.541
R247 VP.n5810 VP.n5809 6.541
R248 VP.n6050 VP.n6049 6.541
R249 VP.n6061 VP.t902 6.541
R250 VP.n6058 VP.t855 6.541
R251 VP.n6053 VP.n6052 6.541
R252 VP.n6651 VP.n6650 6.541
R253 VP.n6670 VP.t705 6.541
R254 VP.n6673 VP.t338 6.541
R255 VP.n6654 VP.n6653 6.541
R256 VP.n6914 VP.n6913 6.541
R257 VP.n6925 VP.t196 6.541
R258 VP.n6922 VP.t129 6.541
R259 VP.n6917 VP.n6916 6.541
R260 VP.n7463 VP.n7462 6.541
R261 VP.n7482 VP.t1308 6.541
R262 VP.n7485 VP.t930 6.541
R263 VP.n7466 VP.n7465 6.541
R264 VP.n7753 VP.n7752 6.541
R265 VP.n7763 VP.t794 6.541
R266 VP.n7760 VP.t742 6.541
R267 VP.n7756 VP.n7755 6.541
R268 VP.n8279 VP.n8278 6.541
R269 VP.n8299 VP.t610 6.541
R270 VP.n8302 VP.t221 6.541
R271 VP.n8282 VP.n8281 6.541
R272 VP.n8592 VP.n8591 6.541
R273 VP.n8602 VP.t51 6.541
R274 VP.n8599 VP.t1341 6.541
R275 VP.n8595 VP.n8594 6.541
R276 VP.n9076 VP.n9075 6.541
R277 VP.n9096 VP.t1203 6.541
R278 VP.n9099 VP.t822 6.541
R279 VP.n9079 VP.n9078 6.541
R280 VP.n9388 VP.n9387 6.541
R281 VP.n9399 VP.t828 6.541
R282 VP.n9396 VP.t566 6.541
R283 VP.n9391 VP.n9390 6.541
R284 VP.n9839 VP.n9838 6.541
R285 VP.n9858 VP.t1034 6.541
R286 VP.n9861 VP.t253 6.541
R287 VP.n9842 VP.n9841 6.541
R288 VP.n10733 VP.n10732 6.541
R289 VP.n10744 VP.t714 6.541
R290 VP.n10741 VP.t475 6.541
R291 VP.n10736 VP.n10735 6.541
R292 VP.n10458 VP.n10457 6.541
R293 VP.n10466 VP.t336 6.541
R294 VP.n10469 VP.t148 6.541
R295 VP.n10461 VP.n10460 6.541
R296 VP.n10192 VP.t1317 6.541
R297 VP.n10341 VP.t451 6.541
R298 VP.n10328 VP.t206 6.541
R299 VP.n10423 VP.n10422 6.541
R300 VP.n10434 VP.t515 6.541
R301 VP.n10431 VP.t1037 6.541
R302 VP.n10426 VP.n10425 6.541
R303 VP.n10974 VP.t300 6.541
R304 VP.n10971 VP.t1 6.541
R305 VP.n9609 VP.t144 6.541
R306 VP.n9606 VP.t1205 6.541
R307 VP.n10053 VP.n10052 6.541
R308 VP.n10073 VP.t369 6.541
R309 VP.n10076 VP.t891 6.541
R310 VP.n10050 VP.n10049 6.541
R311 VP.n10983 VP.n10982 6.541
R312 VP.n11007 VP.t17 6.541
R313 VP.n11010 VP.t1097 6.541
R314 VP.n10980 VP.n10979 6.541
R315 VP.n10620 VP.n10619 6.541
R316 VP.n10644 VP.t962 6.541
R317 VP.n10647 VP.t795 6.541
R318 VP.n10617 VP.n10616 6.541
R319 VP.n10312 VP.t654 6.541
R320 VP.n8803 VP.t1153 6.541
R321 VP.n8800 VP.t1060 6.541
R322 VP.n9257 VP.n9256 6.541
R323 VP.n9275 VP.t220 6.541
R324 VP.n9278 VP.t595 6.541
R325 VP.n9254 VP.n9253 6.541
R326 VP.n9618 VP.n9617 6.541
R327 VP.n9635 VP.t1213 6.541
R328 VP.n9638 VP.t956 6.541
R329 VP.n9615 VP.n9614 6.541
R330 VP.n10013 VP.n10012 6.541
R331 VP.n10042 VP.t819 6.541
R332 VP.n10045 VP.t646 6.541
R333 VP.n10010 VP.n10009 6.541
R334 VP.n10924 VP.n10923 6.541
R335 VP.n10951 VP.t507 6.541
R336 VP.n10948 VP.t243 6.541
R337 VP.n10921 VP.n10920 6.541
R338 VP.n10582 VP.n10581 6.541
R339 VP.n10606 VP.t82 6.541
R340 VP.n10609 VP.t1241 6.541
R341 VP.n10579 VP.n10578 6.541
R342 VP.n10296 VP.t1095 6.541
R343 VP.n8756 VP.n8755 6.541
R344 VP.n8775 VP.t922 6.541
R345 VP.n8772 VP.t812 6.541
R346 VP.n8753 VP.n8752 6.541
R347 VP.n9036 VP.n9035 6.541
R348 VP.n9048 VP.t666 6.541
R349 VP.n9045 VP.t352 6.541
R350 VP.n9039 VP.n9038 6.541
R351 VP.n9568 VP.n9567 6.541
R352 VP.n9579 VP.t360 6.541
R353 VP.n9576 VP.t74 6.541
R354 VP.n9571 VP.n9570 6.541
R355 VP.n9801 VP.n9800 6.541
R356 VP.n9812 VP.t1263 6.541
R357 VP.n9809 VP.t1089 6.541
R358 VP.n9804 VP.n9803 6.541
R359 VP.n10905 VP.n10904 6.541
R360 VP.n10916 VP.t953 6.541
R361 VP.n10913 VP.t687 6.541
R362 VP.n10908 VP.n10907 6.541
R363 VP.n10400 VP.n10399 6.541
R364 VP.n10408 VP.t554 6.541
R365 VP.n10405 VP.t324 6.541
R366 VP.n10397 VP.n10396 6.541
R367 VP.n10284 VP.t181 6.541
R368 VP.n8199 VP.n8198 6.541
R369 VP.n8210 VP.t39 6.541
R370 VP.n8207 VP.t447 6.541
R371 VP.n8202 VP.n8201 6.541
R372 VP.n7912 VP.t1008 6.541
R373 VP.n7909 VP.t912 6.541
R374 VP.n7080 VP.t865 6.541
R375 VP.n7077 VP.t763 6.541
R376 VP.n7591 VP.n7590 6.541
R377 VP.n7609 VP.t1230 6.541
R378 VP.n7612 VP.t295 6.541
R379 VP.n7588 VP.n7587 6.541
R380 VP.n7953 VP.n7952 6.541
R381 VP.n7970 VP.t773 6.541
R382 VP.n7973 VP.t660 6.541
R383 VP.n7950 VP.n7949 6.541
R384 VP.n8419 VP.n8418 6.541
R385 VP.n8448 VP.t519 6.541
R386 VP.n8451 VP.t205 6.541
R387 VP.n8416 VP.n8415 6.541
R388 VP.n8729 VP.n8728 6.541
R389 VP.n8749 VP.t29 6.541
R390 VP.n8746 VP.t1256 6.541
R391 VP.n8726 VP.n8725 6.541
R392 VP.n9219 VP.n9218 6.541
R393 VP.n9246 VP.t1110 6.541
R394 VP.n9249 VP.t800 6.541
R395 VP.n9216 VP.n9215 6.541
R396 VP.n9535 VP.n9534 6.541
R397 VP.n9556 VP.t809 6.541
R398 VP.n9553 VP.t548 6.541
R399 VP.n9532 VP.n9531 6.541
R400 VP.n9976 VP.n9975 6.541
R401 VP.n10002 VP.t409 6.541
R402 VP.n10005 VP.t168 6.541
R403 VP.n9973 VP.n9972 6.541
R404 VP.n10873 VP.n10872 6.541
R405 VP.n10900 VP.t1334 6.541
R406 VP.n10897 VP.t1136 6.541
R407 VP.n10870 VP.n10869 6.541
R408 VP.n10547 VP.n10546 6.541
R409 VP.n10571 VP.t999 6.541
R410 VP.n10574 VP.t775 6.541
R411 VP.n10544 VP.n10543 6.541
R412 VP.n10268 VP.t635 6.541
R413 VP.n7033 VP.n7032 6.541
R414 VP.n7052 VP.t625 6.541
R415 VP.n7049 VP.t513 6.541
R416 VP.n7030 VP.n7029 6.541
R417 VP.n7341 VP.n7340 6.541
R418 VP.n7353 VP.t374 6.541
R419 VP.n7350 VP.t11 6.541
R420 VP.n7344 VP.n7343 6.541
R421 VP.n7876 VP.n7875 6.541
R422 VP.n7886 VP.t1220 6.541
R423 VP.n7883 VP.t1102 6.541
R424 VP.n7879 VP.n7878 6.541
R425 VP.n8162 VP.n8161 6.541
R426 VP.n8174 VP.t967 6.541
R427 VP.n8171 VP.t652 6.541
R428 VP.n8165 VP.n8164 6.541
R429 VP.n8712 VP.n8711 6.541
R430 VP.n8722 VP.t511 6.541
R431 VP.n8719 VP.t399 6.541
R432 VP.n8715 VP.n8714 6.541
R433 VP.n9006 VP.n9005 6.541
R434 VP.n9018 VP.t257 6.541
R435 VP.n9015 VP.t1176 6.541
R436 VP.n9009 VP.n9008 6.541
R437 VP.n9516 VP.n9515 6.541
R438 VP.n9527 VP.t1187 6.541
R439 VP.n9524 VP.t993 6.541
R440 VP.n9519 VP.n9518 6.541
R441 VP.n9779 VP.n9778 6.541
R442 VP.n9790 VP.t856 6.541
R443 VP.n9787 VP.t624 6.541
R444 VP.n9782 VP.n9781 6.541
R445 VP.n10854 VP.n10853 6.541
R446 VP.n10865 VP.t486 6.541
R447 VP.n10862 VP.t282 6.541
R448 VP.n10857 VP.n10856 6.541
R449 VP.n10383 VP.n10382 6.541
R450 VP.n10391 VP.t133 6.541
R451 VP.n10388 VP.t1219 6.541
R452 VP.n10380 VP.n10379 6.541
R453 VP.n10256 VP.t1077 6.541
R454 VP.n6489 VP.n6488 6.541
R455 VP.n6500 VP.t1078 6.541
R456 VP.n6497 VP.t137 6.541
R457 VP.n6492 VP.n6491 6.541
R458 VP.n6161 VP.t709 6.541
R459 VP.n6158 VP.t618 6.541
R460 VP.n5301 VP.t568 6.541
R461 VP.n5298 VP.t320 6.541
R462 VP.n5888 VP.n5887 6.541
R463 VP.n5906 VP.t933 6.541
R464 VP.n5909 VP.t1305 6.541
R465 VP.n5885 VP.n5884 6.541
R466 VP.n6266 VP.n6265 6.541
R467 VP.n6283 VP.t477 6.541
R468 VP.n6286 VP.t367 6.541
R469 VP.n6263 VP.n6262 6.541
R470 VP.n6741 VP.n6740 6.541
R471 VP.n6770 VP.t223 6.541
R472 VP.n6773 VP.t1210 6.541
R473 VP.n6738 VP.n6737 6.541
R474 VP.n7006 VP.n7005 6.541
R475 VP.n7026 VP.t1069 6.541
R476 VP.n7023 VP.t960 6.541
R477 VP.n7003 VP.n7002 6.541
R478 VP.n7553 VP.n7552 6.541
R479 VP.n7580 VP.t824 6.541
R480 VP.n7583 VP.t502 6.541
R481 VP.n7550 VP.n7549 6.541
R482 VP.n7844 VP.n7843 6.541
R483 VP.n7864 VP.t364 6.541
R484 VP.n7861 VP.t247 6.541
R485 VP.n7841 VP.n7840 6.541
R486 VP.n8370 VP.n8369 6.541
R487 VP.n8397 VP.t89 6.541
R488 VP.n8400 VP.t1027 6.541
R489 VP.n8367 VP.n8366 6.541
R490 VP.n8681 VP.n8680 6.541
R491 VP.n8701 VP.t894 6.541
R492 VP.n8698 VP.t849 6.541
R493 VP.n8678 VP.n8677 6.541
R494 VP.n9169 VP.n9168 6.541
R495 VP.n9196 VP.t700 6.541
R496 VP.n9199 VP.t332 6.541
R497 VP.n9166 VP.n9165 6.541
R498 VP.n9484 VP.n9483 6.541
R499 VP.n9505 VP.t341 6.541
R500 VP.n9502 VP.t121 6.541
R501 VP.n9481 VP.n9480 6.541
R502 VP.n9928 VP.n9927 6.541
R503 VP.n9954 VP.t1303 6.541
R504 VP.n9957 VP.t1070 6.541
R505 VP.n9925 VP.n9924 6.541
R506 VP.n10822 VP.n10821 6.541
R507 VP.n10849 VP.t932 6.541
R508 VP.n10846 VP.t734 6.541
R509 VP.n10819 VP.n10818 6.541
R510 VP.n10512 VP.n10511 6.541
R511 VP.n10536 VP.t601 6.541
R512 VP.n10539 VP.t365 6.541
R513 VP.n10509 VP.n10508 6.541
R514 VP.n10240 VP.t222 6.541
R515 VP.n5254 VP.n5253 6.541
R516 VP.n5273 VP.t330 6.541
R517 VP.n5270 VP.t36 6.541
R518 VP.n5251 VP.n5250 6.541
R519 VP.n5603 VP.n5602 6.541
R520 VP.n5615 VP.t44 6.541
R521 VP.n5612 VP.t1064 6.541
R522 VP.n5606 VP.n5605 6.541
R523 VP.n6125 VP.n6124 6.541
R524 VP.n6135 VP.t925 6.541
R525 VP.n6132 VP.t817 6.541
R526 VP.n6128 VP.n6127 6.541
R527 VP.n6452 VP.n6451 6.541
R528 VP.n6464 VP.t670 6.541
R529 VP.n6461 VP.t356 6.541
R530 VP.n6455 VP.n6454 6.541
R531 VP.n6988 VP.n6987 6.541
R532 VP.n6998 VP.t215 6.541
R533 VP.n6995 VP.t79 6.541
R534 VP.n6991 VP.n6990 6.541
R535 VP.n7311 VP.n7310 6.541
R536 VP.n7323 VP.t1270 6.541
R537 VP.n7320 VP.t882 6.541
R538 VP.n7314 VP.n7313 6.541
R539 VP.n7826 VP.n7825 6.541
R540 VP.n7836 VP.t745 6.541
R541 VP.n7833 VP.t691 6.541
R542 VP.n7829 VP.n7828 6.541
R543 VP.n8139 VP.n8138 6.541
R544 VP.n8151 VP.t560 6.541
R545 VP.n8148 VP.t177 6.541
R546 VP.n8142 VP.n8141 6.541
R547 VP.n8664 VP.n8663 6.541
R548 VP.n8674 VP.t1343 6.541
R549 VP.n8671 VP.t1295 6.541
R550 VP.n8667 VP.n8666 6.541
R551 VP.n8983 VP.n8982 6.541
R552 VP.n8995 VP.t1148 6.541
R553 VP.n8992 VP.t781 6.541
R554 VP.n8986 VP.n8985 6.541
R555 VP.n9465 VP.n9464 6.541
R556 VP.n9476 VP.t788 6.541
R557 VP.n9473 VP.t589 6.541
R558 VP.n9468 VP.n9467 6.541
R559 VP.n9757 VP.n9756 6.541
R560 VP.n9768 VP.t453 6.541
R561 VP.n9765 VP.t217 6.541
R562 VP.n9760 VP.n9759 6.541
R563 VP.n10803 VP.n10802 6.541
R564 VP.n10814 VP.t43 6.541
R565 VP.n10811 VP.t1186 6.541
R566 VP.n10806 VP.n10805 6.541
R567 VP.n10366 VP.n10365 6.541
R568 VP.n10374 VP.t1051 6.541
R569 VP.n10371 VP.t816 6.541
R570 VP.n10363 VP.n10362 6.541
R571 VP.n10228 VP.t669 6.541
R572 VP.n4715 VP.n4714 6.541
R573 VP.n4726 VP.t640 6.541
R574 VP.n4723 VP.t1151 6.541
R575 VP.n4718 VP.n4717 6.541
R576 VP.n4341 VP.t423 6.541
R577 VP.n4338 VP.t164 6.541
R578 VP.n3424 VP.t530 6.541
R579 VP.n3421 VP.t269 6.541
R580 VP.n4118 VP.n4117 6.541
R581 VP.n4136 VP.t741 6.541
R582 VP.n4139 VP.t1006 6.541
R583 VP.n4115 VP.n4114 6.541
R584 VP.n4515 VP.n4514 6.541
R585 VP.n4532 VP.t176 6.541
R586 VP.n4535 VP.t1227 6.541
R587 VP.n4512 VP.n4511 6.541
R588 VP.n5013 VP.n5012 6.541
R589 VP.n5042 VP.t1083 6.541
R590 VP.n5045 VP.t920 6.541
R591 VP.n5010 VP.n5009 6.541
R592 VP.n5227 VP.n5226 6.541
R593 VP.n5247 VP.t779 6.541
R594 VP.n5244 VP.t517 6.541
R595 VP.n5224 VP.n5223 6.541
R596 VP.n5850 VP.n5849 6.541
R597 VP.n5877 VP.t525 6.541
R598 VP.n5880 VP.t209 6.541
R599 VP.n5847 VP.n5846 6.541
R600 VP.n6093 VP.n6092 6.541
R601 VP.n6113 VP.t33 6.541
R602 VP.n6110 VP.t1262 6.541
R603 VP.n6090 VP.n6089 6.541
R604 VP.n6692 VP.n6691 6.541
R605 VP.n6719 VP.t1116 6.541
R606 VP.n6722 VP.t731 6.541
R607 VP.n6689 VP.n6688 6.541
R608 VP.n6957 VP.n6956 6.541
R609 VP.n6977 VP.t600 6.541
R610 VP.n6974 VP.t551 6.541
R611 VP.n6954 VP.n6953 6.541
R612 VP.n7504 VP.n7503 6.541
R613 VP.n7531 VP.t414 6.541
R614 VP.n7534 VP.t1333 6.541
R615 VP.n7501 VP.n7500 6.541
R616 VP.n7795 VP.n7794 6.541
R617 VP.n7815 VP.t1197 6.541
R618 VP.n7812 VP.t1140 6.541
R619 VP.n7792 VP.n7791 6.541
R620 VP.n8321 VP.n8320 6.541
R621 VP.n8348 VP.t1004 6.541
R622 VP.n8351 VP.t633 6.541
R623 VP.n8318 VP.n8317 6.541
R624 VP.n8633 VP.n8632 6.541
R625 VP.n8653 VP.t493 6.541
R626 VP.n8650 VP.t441 6.541
R627 VP.n8630 VP.n8629 6.541
R628 VP.n9119 VP.n9118 6.541
R629 VP.n9146 VP.t301 6.541
R630 VP.n9149 VP.t1226 6.541
R631 VP.n9116 VP.n9115 6.541
R632 VP.n9433 VP.n9432 6.541
R633 VP.n9454 VP.t1234 6.541
R634 VP.n9451 VP.t1039 6.541
R635 VP.n9430 VP.n9429 6.541
R636 VP.n9880 VP.n9879 6.541
R637 VP.n9906 VP.t905 6.541
R638 VP.n9909 VP.t664 6.541
R639 VP.n9877 VP.n9876 6.541
R640 VP.n10771 VP.n10770 6.541
R641 VP.n10798 VP.t523 6.541
R642 VP.n10795 VP.t340 6.541
R643 VP.n10768 VP.n10767 6.541
R644 VP.n10477 VP.n10476 6.541
R645 VP.n10501 VP.t198 6.541
R646 VP.n10504 VP.t1261 6.541
R647 VP.n10474 VP.n10473 6.541
R648 VP.n10212 VP.t1113 6.541
R649 VP.n349 VP.t58 6.541
R650 VP.n346 VP.t1130 6.541
R651 VP.n867 VP.n866 6.541
R652 VP.n878 VP.t296 6.541
R653 VP.n875 VP.t830 6.541
R654 VP.n870 VP.n869 6.541
R655 VP.n1409 VP.n1408 6.541
R656 VP.n1419 VP.t1290 6.541
R657 VP.n1416 VP.t1035 6.541
R658 VP.n1412 VP.n1411 6.541
R659 VP.n1853 VP.n1852 6.541
R660 VP.n1865 VP.t899 6.541
R661 VP.n1862 VP.t715 6.541
R662 VP.n1856 VP.n1855 6.541
R663 VP.n2621 VP.n2620 6.541
R664 VP.n2628 VP.t582 6.541
R665 VP.n2631 VP.t337 6.541
R666 VP.n2624 VP.n2623 6.541
R667 VP.n2806 VP.n2805 6.541
R668 VP.n2818 VP.t192 6.541
R669 VP.n2815 VP.t1319 6.541
R670 VP.n2809 VP.n2808 6.541
R671 VP.n3332 VP.n3331 6.541
R672 VP.n3342 VP.t1179 6.541
R673 VP.n3339 VP.t929 6.541
R674 VP.n3335 VP.n3334 6.541
R675 VP.n3746 VP.n3745 6.541
R676 VP.n3758 VP.t793 6.541
R677 VP.n3755 VP.t286 6.541
R678 VP.n3749 VP.n3748 6.541
R679 VP.n4253 VP.n4252 6.541
R680 VP.n4263 VP.t141 6.541
R681 VP.n4260 VP.t1268 6.541
R682 VP.n4256 VP.n4255 6.541
R683 VP.n4652 VP.n4651 6.541
R684 VP.n4664 VP.t1121 6.541
R685 VP.n4661 VP.t889 6.541
R686 VP.n4655 VP.n4654 6.541
R687 VP.n5159 VP.n5158 6.541
R688 VP.n5169 VP.t752 6.541
R689 VP.n5166 VP.t559 6.541
R690 VP.n5162 VP.n5161 6.541
R691 VP.n5547 VP.n5546 6.541
R692 VP.n5559 VP.t565 6.541
R693 VP.n5556 VP.t187 6.541
R694 VP.n5550 VP.n5549 6.541
R695 VP.n6023 VP.n6022 6.541
R696 VP.n6033 VP.t1348 6.541
R697 VP.n6030 VP.t1301 6.541
R698 VP.n6026 VP.n6025 6.541
R699 VP.n6403 VP.n6402 6.541
R700 VP.n6415 VP.t1154 6.541
R701 VP.n6412 VP.t786 6.541
R702 VP.n6406 VP.n6405 6.541
R703 VP.n6887 VP.n6886 6.541
R704 VP.n6897 VP.t644 6.541
R705 VP.n6894 VP.t597 6.541
R706 VP.n6890 VP.n6889 6.541
R707 VP.n7262 VP.n7261 6.541
R708 VP.n7274 VP.t459 6.541
R709 VP.n7271 VP.t40 6.541
R710 VP.n7265 VP.n7264 6.541
R711 VP.n7726 VP.n7725 6.541
R712 VP.n7736 VP.t1239 6.541
R713 VP.n7733 VP.t1195 6.541
R714 VP.n7729 VP.n7728 6.541
R715 VP.n8090 VP.n8089 6.541
R716 VP.n8102 VP.t1057 6.541
R717 VP.n8099 VP.t668 6.541
R718 VP.n8093 VP.n8092 6.541
R719 VP.n8565 VP.n8564 6.541
R720 VP.n8575 VP.t528 6.541
R721 VP.n8572 VP.t421 6.541
R722 VP.n8568 VP.n8567 6.541
R723 VP.n8934 VP.n8933 6.541
R724 VP.n8946 VP.t887 6.541
R725 VP.n8943 VP.t1266 6.541
R726 VP.n8937 VP.n8936 6.541
R727 VP.n9359 VP.n9358 6.541
R728 VP.n9370 VP.t571 6.541
R729 VP.n9367 VP.t326 6.541
R730 VP.n9362 VP.n9361 6.541
R731 VP.n9735 VP.n9734 6.541
R732 VP.n9746 VP.t183 6.541
R733 VP.n9743 VP.t1310 6.541
R734 VP.n9738 VP.n9737 6.541
R735 VP.n10704 VP.n10703 6.541
R736 VP.n10715 VP.t1164 6.541
R737 VP.n10712 VP.t924 6.541
R738 VP.n10707 VP.n10706 6.541
R739 VP.n10138 VP.n10137 6.541
R740 VP.n10149 VP.t784 6.541
R741 VP.n10146 VP.t612 6.541
R742 VP.n10141 VP.n10140 6.541
R743 VP.n10337 VP.t471 6.541
R744 VP.n243 VP.t546 6.541
R745 VP.n10126 VP.t1059 6.541
R746 VP.n10689 VP.n10688 6.541
R747 VP.n11013 VP.t322 6.541
R748 VP.n11016 VP.t30 6.541
R749 VP.n11019 VP.n11018 6.541
R750 VP.n9702 VP.n9701 6.541
R751 VP.n9724 VP.t636 6.541
R752 VP.n9721 VP.t461 6.541
R753 VP.n9705 VP.n9704 6.541
R754 VP.n9337 VP.n9336 6.541
R755 VP.n9348 VP.t1016 6.541
R756 VP.n9345 VP.t776 6.541
R757 VP.n9340 VP.n9339 6.541
R758 VP.n8911 VP.n8910 6.541
R759 VP.n8923 VP.t1337 6.541
R760 VP.n8920 VP.t1010 6.541
R761 VP.n8914 VP.n8913 6.541
R762 VP.n8544 VP.n8543 6.541
R763 VP.n8554 VP.t274 6.541
R764 VP.n8551 VP.t172 6.541
R765 VP.n8547 VP.n8546 6.541
R766 VP.n8067 VP.n8066 6.541
R767 VP.n8079 VP.t737 6.541
R768 VP.n8076 VP.t1111 6.541
R769 VP.n8070 VP.n8069 6.541
R770 VP.n7705 VP.n7704 6.541
R771 VP.n7715 VP.t383 6.541
R772 VP.n7712 VP.t266 6.541
R773 VP.n7708 VP.n7707 6.541
R774 VP.n7239 VP.n7238 6.541
R775 VP.n7251 VP.t909 6.541
R776 VP.n7248 VP.t520 6.541
R777 VP.n7242 VP.n7241 6.541
R778 VP.n6866 VP.n6865 6.541
R779 VP.n6876 VP.t1087 6.541
R780 VP.n6873 VP.t1046 6.541
R781 VP.n6869 VP.n6868 6.541
R782 VP.n6380 VP.n6379 6.541
R783 VP.n6392 VP.t307 6.541
R784 VP.n6389 VP.t1231 6.541
R785 VP.n6383 VP.n6382 6.541
R786 VP.n6002 VP.n6001 6.541
R787 VP.n6012 VP.t497 6.541
R788 VP.n6009 VP.t448 6.541
R789 VP.n6005 VP.n6004 6.541
R790 VP.n5524 VP.n5523 6.541
R791 VP.n5536 VP.t1009 6.541
R792 VP.n5533 VP.t638 6.541
R793 VP.n5527 VP.n5526 6.541
R794 VP.n5138 VP.n5137 6.541
R795 VP.n5148 VP.t1202 6.541
R796 VP.n5145 VP.t1002 6.541
R797 VP.n5141 VP.n5140 6.541
R798 VP.n4629 VP.n4628 6.541
R799 VP.n4641 VP.t265 6.541
R800 VP.n4638 VP.t1340 6.541
R801 VP.n4632 VP.n4631 6.541
R802 VP.n4232 VP.n4231 6.541
R803 VP.n4242 VP.t607 6.541
R804 VP.n4239 VP.t413 6.541
R805 VP.n4235 VP.n4234 6.541
R806 VP.n3723 VP.n3722 6.541
R807 VP.n3735 VP.t1237 6.541
R808 VP.n3732 VP.t738 6.541
R809 VP.n3726 VP.n3725 6.541
R810 VP.n3311 VP.n3310 6.541
R811 VP.n3321 VP.t258 6.541
R812 VP.n3318 VP.t38 6.541
R813 VP.n3314 VP.n3313 6.541
R814 VP.n2783 VP.n2782 6.541
R815 VP.n2795 VP.t642 6.541
R816 VP.n2792 VP.t400 6.541
R817 VP.n2786 VP.n2785 6.541
R818 VP.n2646 VP.n2645 6.541
R819 VP.n2653 VP.t1030 6.541
R820 VP.n2656 VP.t785 6.541
R821 VP.n2649 VP.n2648 6.541
R822 VP.n1823 VP.n1822 6.541
R823 VP.n1835 VP.t1346 6.541
R824 VP.n1832 VP.t1166 6.541
R825 VP.n1826 VP.n1825 6.541
R826 VP.n1385 VP.n1384 6.541
R827 VP.n1395 VP.t435 6.541
R828 VP.n1392 VP.t184 6.541
R829 VP.n1388 VP.n1387 6.541
R830 VP.n839 VP.n838 6.541
R831 VP.n849 VP.t750 6.541
R832 VP.n820 VP.t572 6.541
R833 VP.n842 VP.n841 6.541
R834 VP.n296 VP.n295 6.541
R835 VP.n318 VP.t1135 6.541
R836 VP.n315 VP.t888 6.541
R837 VP.n299 VP.n298 6.541
R838 VP.n201 VP.t529 6.541
R839 VP.n147 VP.t138 6.541
R840 VP.n205 VP.t70 6.541
R841 VP.n203 VP.t418 6.541
R842 VP.n267 VP.n266 6.541
R843 VP.n730 VP.t78 6.541
R844 VP.n733 VP.t1144 6.541
R845 VP.n736 VP.n735 6.541
R846 VP.n777 VP.t843 6.541
R847 VP.n209 VP.t952 6.541
R848 VP.n207 VP.t1273 6.541
R849 VP.n370 VP.n369 6.541
R850 VP.n394 VP.t959 6.541
R851 VP.n397 VP.t694 6.541
R852 VP.n373 VP.n372 6.541
R853 VP.n906 VP.n905 6.541
R854 VP.n926 VP.t563 6.541
R855 VP.n929 VP.t391 6.541
R856 VP.n909 VP.n908 6.541
R857 VP.n1339 VP.n1338 6.541
R858 VP.n1731 VP.t246 6.541
R859 VP.n1734 VP.t1298 6.541
R860 VP.n1737 VP.n1736 6.541
R861 VP.n1766 VP.t985 6.541
R862 VP.n213 VP.t1201 6.541
R863 VP.n211 VP.t827 6.541
R864 VP.n417 VP.n416 6.541
R865 VP.n441 VP.t512 6.541
R866 VP.n444 VP.t249 6.541
R867 VP.n420 VP.n419 6.541
R868 VP.n956 VP.n955 6.541
R869 VP.n976 VP.t93 6.541
R870 VP.n979 VP.t1248 6.541
R871 VP.n959 VP.n958 6.541
R872 VP.n1468 VP.n1467 6.541
R873 VP.n1482 VP.t1101 6.541
R874 VP.n1485 VP.t851 6.541
R875 VP.n1471 VP.n1470 6.541
R876 VP.n1893 VP.n1892 6.541
R877 VP.n1915 VP.t703 6.541
R878 VP.n1918 VP.t537 6.541
R879 VP.n1896 VP.n1895 6.541
R880 VP.n2315 VP.n2314 6.541
R881 VP.n2692 VP.t398 6.541
R882 VP.n2695 VP.t124 6.541
R883 VP.n2698 VP.n2697 6.541
R884 VP.n2727 VP.t1128 6.541
R885 VP.n217 VP.t753 6.541
R886 VP.n215 VP.t1127 6.541
R887 VP.n464 VP.n463 6.541
R888 VP.n488 VP.t761 6.541
R889 VP.n491 VP.t506 6.541
R890 VP.n467 VP.n466 6.541
R891 VP.n1006 VP.n1005 6.541
R892 VP.n1026 VP.t969 6.541
R893 VP.n1029 VP.t194 6.541
R894 VP.n1009 VP.n1008 6.541
R895 VP.n1506 VP.n1505 6.541
R896 VP.n1520 VP.t659 6.541
R897 VP.n1523 VP.t402 6.541
R898 VP.n1509 VP.n1508 6.541
R899 VP.n1945 VP.n1944 6.541
R900 VP.n1967 VP.t259 6.541
R901 VP.n1970 VP.t61 6.541
R902 VP.n1948 VP.n1947 6.541
R903 VP.n2568 VP.n2567 6.541
R904 VP.n2585 VP.t1255 6.541
R905 VP.n2582 VP.t994 6.541
R906 VP.n2571 VP.n2570 6.541
R907 VP.n2874 VP.n2873 6.541
R908 VP.n2896 VP.t858 6.541
R909 VP.n2899 VP.t681 6.541
R910 VP.n2877 VP.n2876 6.541
R911 VP.n3265 VP.n3264 6.541
R912 VP.n3632 VP.t547 6.541
R913 VP.n3635 VP.t284 6.541
R914 VP.n3638 VP.n3637 6.541
R915 VP.n3667 VP.t1021 6.541
R916 VP.n221 VP.t298 6.541
R917 VP.n219 VP.t679 6.541
R918 VP.n511 VP.n510 6.541
R919 VP.n535 VP.t308 6.541
R920 VP.n538 VP.t96 6.541
R921 VP.n514 VP.n513 6.541
R922 VP.n1056 VP.n1055 6.541
R923 VP.n1076 VP.t1282 6.541
R924 VP.n1079 VP.t1048 6.541
R925 VP.n1059 VP.n1058 6.541
R926 VP.n1544 VP.n1543 6.541
R927 VP.n1558 VP.t910 6.541
R928 VP.n1561 VP.t653 6.541
R929 VP.n1547 VP.n1546 6.541
R930 VP.n1997 VP.n1996 6.541
R931 VP.n2019 VP.t1112 6.541
R932 VP.n2022 VP.t347 6.541
R933 VP.n2000 VP.n1999 6.541
R934 VP.n2530 VP.n2529 6.541
R935 VP.n2547 VP.t811 6.541
R936 VP.n2544 VP.t550 6.541
R937 VP.n2533 VP.n2532 6.541
R938 VP.n2926 VP.n2925 6.541
R939 VP.n2948 VP.t411 6.541
R940 VP.n2951 VP.t238 6.541
R941 VP.n2929 VP.n2928 6.541
R942 VP.n3446 VP.n3445 6.541
R943 VP.n3460 VP.t73 6.541
R944 VP.n3463 VP.t1139 6.541
R945 VP.n3449 VP.n3448 6.541
R946 VP.n3819 VP.n3818 6.541
R947 VP.n3841 VP.t1001 6.541
R948 VP.n3844 VP.t574 6.541
R949 VP.n3822 VP.n3821 6.541
R950 VP.n4186 VP.n4185 6.541
R951 VP.n4538 VP.t438 6.541
R952 VP.n4541 VP.t188 6.541
R953 VP.n4544 VP.n4543 6.541
R954 VP.n4573 VP.t1169 6.541
R955 VP.n225 VP.t1146 6.541
R956 VP.n223 VP.t235 6.541
R957 VP.n558 VP.n557 6.541
R958 VP.n582 VP.t1155 6.541
R959 VP.n585 VP.t973 6.541
R960 VP.n561 VP.n560 6.541
R961 VP.n1106 VP.n1105 6.541
R962 VP.n1126 VP.t837 6.541
R963 VP.n1129 VP.t598 6.541
R964 VP.n1109 VP.n1108 6.541
R965 VP.n1582 VP.n1581 6.541
R966 VP.n1596 VP.t460 6.541
R967 VP.n1599 VP.t260 6.541
R968 VP.n1585 VP.n1584 6.541
R969 VP.n2049 VP.n2048 6.541
R970 VP.n2071 VP.t102 6.541
R971 VP.n2074 VP.t1196 6.541
R972 VP.n2052 VP.n2051 6.541
R973 VP.n2492 VP.n2491 6.541
R974 VP.n2509 VP.t1058 6.541
R975 VP.n2506 VP.t803 6.541
R976 VP.n2495 VP.n2494 6.541
R977 VP.n2978 VP.n2977 6.541
R978 VP.n3000 VP.t1267 6.541
R979 VP.n3003 VP.t492 6.541
R980 VP.n2981 VP.n2980 6.541
R981 VP.n3484 VP.n3483 6.541
R982 VP.n3498 VP.t955 6.541
R983 VP.n3501 VP.t690 6.541
R984 VP.n3487 VP.n3486 6.541
R985 VP.n3871 VP.n3870 6.541
R986 VP.n3893 VP.t557 6.541
R987 VP.n3896 VP.t106 6.541
R988 VP.n3874 VP.n3873 6.541
R989 VP.n4363 VP.n4362 6.541
R990 VP.n4377 VP.t1293 6.541
R991 VP.n4380 VP.t1038 6.541
R992 VP.n4366 VP.n4365 6.541
R993 VP.n4754 VP.n4753 6.541
R994 VP.n4776 VP.t904 6.541
R995 VP.n4779 VP.t717 6.541
R996 VP.n4757 VP.n4756 6.541
R997 VP.n5092 VP.n5091 6.541
R998 VP.n5433 VP.t586 6.541
R999 VP.n5436 VP.t339 6.541
R1000 VP.n5439 VP.n5438 6.541
R1001 VP.n5468 VP.t1323 6.541
R1002 VP.n229 VP.t699 6.541
R1003 VP.n227 VP.t1090 6.541
R1004 VP.n605 VP.n604 6.541
R1005 VP.n622 VP.t706 6.541
R1006 VP.n625 VP.t524 6.541
R1007 VP.n608 VP.n607 6.541
R1008 VP.n1156 VP.n1155 6.541
R1009 VP.n1164 VP.t386 6.541
R1010 VP.n1167 VP.t130 6.541
R1011 VP.n1159 VP.n1158 6.541
R1012 VP.n1620 VP.n1619 6.541
R1013 VP.n1628 VP.t1309 6.541
R1014 VP.n1631 VP.t1115 6.541
R1015 VP.n1623 VP.n1622 6.541
R1016 VP.n2101 VP.n2100 6.541
R1017 VP.n2112 VP.t978 6.541
R1018 VP.n2115 VP.t743 6.541
R1019 VP.n2104 VP.n2103 6.541
R1020 VP.n2460 VP.n2459 6.541
R1021 VP.n2471 VP.t611 6.541
R1022 VP.n2468 VP.t416 6.541
R1023 VP.n2463 VP.n2462 6.541
R1024 VP.n3030 VP.n3029 6.541
R1025 VP.n3041 VP.t268 6.541
R1026 VP.n3044 VP.t1342 6.541
R1027 VP.n3033 VP.n3032 6.541
R1028 VP.n3522 VP.n3521 6.541
R1029 VP.n3530 VP.t1204 6.541
R1030 VP.n3533 VP.t946 6.541
R1031 VP.n3525 VP.n3524 6.541
R1032 VP.n3923 VP.n3922 6.541
R1033 VP.n3934 VP.t86 6.541
R1034 VP.n3937 VP.t380 6.541
R1035 VP.n3926 VP.n3925 6.541
R1036 VP.n4401 VP.n4400 6.541
R1037 VP.n4409 VP.t848 6.541
R1038 VP.n4412 VP.t588 6.541
R1039 VP.n4404 VP.n4403 6.541
R1040 VP.n4806 VP.n4805 6.541
R1041 VP.n4817 VP.t452 6.541
R1042 VP.n4820 VP.t271 6.541
R1043 VP.n4809 VP.n4808 6.541
R1044 VP.n5323 VP.n5322 6.541
R1045 VP.n5331 VP.t120 6.541
R1046 VP.n5334 VP.t1185 6.541
R1047 VP.n5326 VP.n5325 6.541
R1048 VP.n5643 VP.n5642 6.541
R1049 VP.n5654 VP.t1198 6.541
R1050 VP.n5657 VP.t872 6.541
R1051 VP.n5646 VP.n5645 6.541
R1052 VP.n5956 VP.n5955 6.541
R1053 VP.n6289 VP.t730 6.541
R1054 VP.n6292 VP.t634 6.541
R1055 VP.n6295 VP.n6294 6.541
R1056 VP.n6324 VP.t162 6.541
R1057 VP.n233 VP.t254 6.541
R1058 VP.n231 VP.t648 6.541
R1059 VP.n645 VP.n644 6.541
R1060 VP.n652 VP.t262 6.541
R1061 VP.n655 VP.t46 6.541
R1062 VP.n648 VP.n647 6.541
R1063 VP.n1194 VP.n1193 6.541
R1064 VP.n1204 VP.t1242 6.541
R1065 VP.n1207 VP.t997 6.541
R1066 VP.n1197 VP.n1196 6.541
R1067 VP.n1652 VP.n1651 6.541
R1068 VP.n1660 VP.t862 6.541
R1069 VP.n1663 VP.t671 6.541
R1070 VP.n1655 VP.n1654 6.541
R1071 VP.n2142 VP.n2141 6.541
R1072 VP.n2153 VP.t532 6.541
R1073 VP.n2156 VP.t290 6.541
R1074 VP.n2145 VP.n2144 6.541
R1075 VP.n2428 VP.n2427 6.541
R1076 VP.n2439 VP.t146 6.541
R1077 VP.n2436 VP.t1271 6.541
R1078 VP.n2431 VP.n2430 6.541
R1079 VP.n3071 VP.n3070 6.541
R1080 VP.n3082 VP.t1124 6.541
R1081 VP.n3085 VP.t893 6.541
R1082 VP.n3074 VP.n3073 6.541
R1083 VP.n3554 VP.n3553 6.541
R1084 VP.n3562 VP.t756 6.541
R1085 VP.n3565 VP.t561 6.541
R1086 VP.n3557 VP.n3556 6.541
R1087 VP.n3964 VP.n3963 6.541
R1088 VP.n3975 VP.t422 6.541
R1089 VP.n3978 VP.t1235 6.541
R1090 VP.n3967 VP.n3966 6.541
R1091 VP.n4433 VP.n4432 6.541
R1092 VP.n4441 VP.t1093 6.541
R1093 VP.n4444 VP.t840 6.541
R1094 VP.n4436 VP.n4435 6.541
R1095 VP.n4847 VP.n4846 6.541
R1096 VP.n4858 VP.t1302 6.541
R1097 VP.n4861 VP.t526 6.541
R1098 VP.n4850 VP.n4849 6.541
R1099 VP.n5355 VP.n5354 6.541
R1100 VP.n5363 VP.t991 6.541
R1101 VP.n5366 VP.t732 6.541
R1102 VP.n5358 VP.n5357 6.541
R1103 VP.n5684 VP.n5683 6.541
R1104 VP.n5695 VP.t747 6.541
R1105 VP.n5698 VP.t426 6.541
R1106 VP.n5687 VP.n5686 6.541
R1107 VP.n6183 VP.n6182 6.541
R1108 VP.n6191 VP.t279 6.541
R1109 VP.n6194 VP.t178 6.541
R1110 VP.n6186 VP.n6185 6.541
R1111 VP.n6528 VP.n6527 6.541
R1112 VP.n6539 VP.t1344 6.541
R1113 VP.n6542 VP.t1013 6.541
R1114 VP.n6531 VP.n6530 6.541
R1115 VP.n6820 VP.n6819 6.541
R1116 VP.n7148 VP.t881 6.541
R1117 VP.n7151 VP.t782 6.541
R1118 VP.n7154 VP.n7153 6.541
R1119 VP.n7183 VP.t318 6.541
R1120 VP.n237 VP.t1108 6.541
R1121 VP.n235 VP.t202 6.541
R1122 VP.n675 VP.n674 6.541
R1123 VP.n684 VP.t1117 6.541
R1124 VP.n687 VP.t935 6.541
R1125 VP.n678 VP.n677 6.541
R1126 VP.n1234 VP.n1233 6.541
R1127 VP.n1245 VP.t797 6.541
R1128 VP.n1248 VP.t552 6.541
R1129 VP.n1237 VP.n1236 6.541
R1130 VP.n1684 VP.n1683 6.541
R1131 VP.n1692 VP.t415 6.541
R1132 VP.n1695 VP.t224 6.541
R1133 VP.n1687 VP.n1686 6.541
R1134 VP.n2183 VP.n2182 6.541
R1135 VP.n2194 VP.t54 6.541
R1136 VP.n2197 VP.t1141 6.541
R1137 VP.n2186 VP.n2185 6.541
R1138 VP.n2396 VP.n2395 6.541
R1139 VP.n2407 VP.t1005 6.541
R1140 VP.n2404 VP.t825 6.541
R1141 VP.n2399 VP.n2398 6.541
R1142 VP.n3112 VP.n3111 6.541
R1143 VP.n3123 VP.t677 6.541
R1144 VP.n3126 VP.t442 6.541
R1145 VP.n3115 VP.n3114 6.541
R1146 VP.n3586 VP.n3585 6.541
R1147 VP.n3594 VP.t302 6.541
R1148 VP.n3597 VP.t90 6.541
R1149 VP.n3589 VP.n3588 6.541
R1150 VP.n4005 VP.n4004 6.541
R1151 VP.n4016 VP.t1277 6.541
R1152 VP.n4019 VP.t790 6.541
R1153 VP.n4008 VP.n4007 6.541
R1154 VP.n4465 VP.n4464 6.541
R1155 VP.n4473 VP.t650 6.541
R1156 VP.n4476 VP.t456 6.541
R1157 VP.n4468 VP.n4467 6.541
R1158 VP.n4888 VP.n4887 6.541
R1159 VP.n4899 VP.t317 6.541
R1160 VP.n4902 VP.t47 6.541
R1161 VP.n4891 VP.n4890 6.541
R1162 VP.n5387 VP.n5386 6.541
R1163 VP.n5395 VP.t1244 6.541
R1164 VP.n5398 VP.t981 6.541
R1165 VP.n5390 VP.n5389 6.541
R1166 VP.n5725 VP.n5724 6.541
R1167 VP.n5736 VP.t293 6.541
R1168 VP.n5739 VP.t672 6.541
R1169 VP.n5728 VP.n5727 6.541
R1170 VP.n6215 VP.n6214 6.541
R1171 VP.n6223 VP.t1133 6.541
R1172 VP.n6226 VP.t1029 6.541
R1173 VP.n6218 VP.n6217 6.541
R1174 VP.n6569 VP.n6568 6.541
R1175 VP.n6580 VP.t896 6.541
R1176 VP.n6583 VP.t569 6.541
R1177 VP.n6572 VP.n6571 6.541
R1178 VP.n7102 VP.n7101 6.541
R1179 VP.n7110 VP.t432 6.541
R1180 VP.n7113 VP.t333 6.541
R1181 VP.n7105 VP.n7104 6.541
R1182 VP.n7381 VP.n7380 6.541
R1183 VP.n7392 VP.t190 6.541
R1184 VP.n7395 VP.t1161 6.541
R1185 VP.n7384 VP.n7383 6.541
R1186 VP.n7659 VP.n7658 6.541
R1187 VP.n7976 VP.t1026 6.541
R1188 VP.n7979 VP.t927 6.541
R1189 VP.n7982 VP.n7981 6.541
R1190 VP.n8011 VP.t470 6.541
R1191 VP.n142 VP.t275 6.541
R1192 VP.n140 VP.t604 6.541
R1193 VP.n274 VP.n273 6.541
R1194 VP.n292 VP.t281 6.541
R1195 VP.n289 VP.t1338 6.541
R1196 VP.n271 VP.n270 6.541
R1197 VP.n790 VP.n789 6.541
R1198 VP.n787 VP.t1199 6.541
R1199 VP.n817 VP.t1017 6.541
R1200 VP.n784 VP.n783 6.541
R1201 VP.n1346 VP.n1345 6.541
R1202 VP.n1370 VP.t884 6.541
R1203 VP.n1367 VP.t637 6.541
R1204 VP.n1343 VP.n1342 6.541
R1205 VP.n1776 VP.n1775 6.541
R1206 VP.n1806 VP.t495 6.541
R1207 VP.n1803 VP.t248 6.541
R1208 VP.n1773 VP.n1772 6.541
R1209 VP.n2663 VP.n2662 6.541
R1210 VP.n2684 VP.t92 6.541
R1211 VP.n2687 VP.t1229 6.541
R1212 VP.n2660 VP.n2659 6.541
R1213 VP.n2736 VP.n2735 6.541
R1214 VP.n2766 VP.t1085 6.541
R1215 VP.n2763 VP.t850 6.541
R1216 VP.n2733 VP.n2732 6.541
R1217 VP.n3272 VP.n3271 6.541
R1218 VP.n3296 VP.t701 6.541
R1219 VP.n3293 VP.t518 6.541
R1220 VP.n3269 VP.n3268 6.541
R1221 VP.n3676 VP.n3675 6.541
R1222 VP.n3706 VP.t381 6.541
R1223 VP.n3703 VP.t1193 6.541
R1224 VP.n3673 VP.n3672 6.541
R1225 VP.n4193 VP.n4192 6.541
R1226 VP.n4217 VP.t1055 6.541
R1227 VP.n4214 VP.t859 6.541
R1228 VP.n4190 VP.n4189 6.541
R1229 VP.n4585 VP.n4584 6.541
R1230 VP.n4582 VP.t711 6.541
R1231 VP.n4612 VP.t490 6.541
R1232 VP.n4579 VP.n4578 6.541
R1233 VP.n5099 VP.n5098 6.541
R1234 VP.n5123 VP.t351 6.541
R1235 VP.n5120 VP.t139 6.541
R1236 VP.n5096 VP.n5095 6.541
R1237 VP.n5477 VP.n5476 6.541
R1238 VP.n5507 VP.t151 6.541
R1239 VP.n5504 VP.t1080 6.541
R1240 VP.n5474 VP.n5473 6.541
R1241 VP.n5963 VP.n5962 6.541
R1242 VP.n5987 VP.t942 6.541
R1243 VP.n5984 VP.t901 6.541
R1244 VP.n5960 VP.n5959 6.541
R1245 VP.n6333 VP.n6332 6.541
R1246 VP.n6363 VP.t760 6.541
R1247 VP.n6360 VP.t375 6.541
R1248 VP.n6330 VP.n6329 6.541
R1249 VP.n6827 VP.n6826 6.541
R1250 VP.n6851 VP.t232 6.541
R1251 VP.n6848 VP.t100 6.541
R1252 VP.n6824 VP.n6823 6.541
R1253 VP.n7192 VP.n7191 6.541
R1254 VP.n7222 VP.t591 6.541
R1255 VP.n7219 VP.t968 6.541
R1256 VP.n7189 VP.n7188 6.541
R1257 VP.n7666 VP.n7665 6.541
R1258 VP.n7690 VP.t112 6.541
R1259 VP.n7687 VP.t1327 6.541
R1260 VP.n7663 VP.n7662 6.541
R1261 VP.n8020 VP.n8019 6.541
R1262 VP.n8050 VP.t1189 6.541
R1263 VP.n8047 VP.t867 6.541
R1264 VP.n8017 VP.n8016 6.541
R1265 VP.n8505 VP.n8504 6.541
R1266 VP.n8529 VP.t721 6.541
R1267 VP.n8526 VP.t628 6.541
R1268 VP.n8502 VP.n8501 6.541
R1269 VP.n8866 VP.n8865 6.541
R1270 VP.n8894 VP.t487 6.541
R1271 VP.n8891 VP.t154 6.541
R1272 VP.n8863 VP.n8862 6.541
R1273 VP.n9322 VP.n9321 6.541
R1274 VP.n9641 VP.t165 6.541
R1275 VP.n9644 VP.t1222 6.541
R1276 VP.n9647 VP.n9646 6.541
R1277 VP.n9686 VP.t911 6.541
R1278 VP.n2224 VP.n2223 6.541
R1279 VP.n2235 VP.t940 6.541
R1280 VP.n2238 VP.t692 6.541
R1281 VP.n2227 VP.n2226 6.541
R1282 VP.n2364 VP.n2363 6.541
R1283 VP.n2375 VP.t562 6.541
R1284 VP.n2372 VP.t373 6.541
R1285 VP.n2367 VP.n2366 6.541
R1286 VP.n3153 VP.n3152 6.541
R1287 VP.n3164 VP.t230 6.541
R1288 VP.n3167 VP.t1296 6.541
R1289 VP.n3156 VP.n3155 6.541
R1290 VP.n3618 VP.n3617 6.541
R1291 VP.n3626 VP.t1150 6.541
R1292 VP.n3629 VP.t966 6.541
R1293 VP.n3621 VP.n3620 6.541
R1294 VP.n4046 VP.n4045 6.541
R1295 VP.n4057 VP.t832 6.541
R1296 VP.n4060 VP.t344 6.541
R1297 VP.n4049 VP.n4048 6.541
R1298 VP.n4497 VP.n4496 6.541
R1299 VP.n4505 VP.t203 6.541
R1300 VP.n4508 VP.t1306 6.541
R1301 VP.n4500 VP.n4499 6.541
R1302 VP.n4929 VP.n4928 6.541
R1303 VP.n4940 VP.t1160 6.541
R1304 VP.n4943 VP.t936 6.541
R1305 VP.n4932 VP.n4931 6.541
R1306 VP.n5419 VP.n5418 6.541
R1307 VP.n5427 VP.t798 6.541
R1308 VP.n5430 VP.t606 6.541
R1309 VP.n5422 VP.n5421 6.541
R1310 VP.n5766 VP.n5765 6.541
R1311 VP.n5777 VP.t615 6.541
R1312 VP.n5780 VP.t225 6.541
R1313 VP.n5769 VP.n5768 6.541
R1314 VP.n6247 VP.n6246 6.541
R1315 VP.n6255 VP.t55 6.541
R1316 VP.n6258 VP.t1280 6.541
R1317 VP.n6250 VP.n6249 6.541
R1318 VP.n6610 VP.n6609 6.541
R1319 VP.n6621 VP.t444 6.541
R1320 VP.n6624 VP.t826 6.541
R1321 VP.n6613 VP.n6612 6.541
R1322 VP.n7134 VP.n7133 6.541
R1323 VP.n7142 VP.t1287 6.541
R1324 VP.n7145 VP.t1178 6.541
R1325 VP.n7137 VP.n7136 6.541
R1326 VP.n7422 VP.n7421 6.541
R1327 VP.n7433 VP.t1042 6.541
R1328 VP.n7436 VP.t712 6.541
R1329 VP.n7425 VP.n7424 6.541
R1330 VP.n7934 VP.n7933 6.541
R1331 VP.n7942 VP.t578 6.541
R1332 VP.n7945 VP.t479 6.541
R1333 VP.n7937 VP.n7936 6.541
R1334 VP.n8238 VP.n8237 6.541
R1335 VP.n8249 VP.t342 6.541
R1336 VP.n8252 VP.t1316 6.541
R1337 VP.n8241 VP.n8240 6.541
R1338 VP.n8498 VP.n8497 6.541
R1339 VP.n8807 VP.t1174 6.541
R1340 VP.n8810 VP.t1073 6.541
R1341 VP.n8813 VP.n8812 6.541
R1342 VP.n8845 VP.t616 6.541
R1343 VP.n241 VP.t723 6.541
R1344 VP.n239 VP.t1053 6.541
R1345 VP.n707 VP.n706 6.541
R1346 VP.n724 VP.t733 6.541
R1347 VP.n727 VP.t489 6.541
R1348 VP.n710 VP.n709 6.541
R1349 VP.n1275 VP.n1274 6.541
R1350 VP.n1286 VP.t349 6.541
R1351 VP.n1289 VP.t81 6.541
R1352 VP.n1278 VP.n1277 6.541
R1353 VP.n1716 VP.n1715 6.541
R1354 VP.n1725 VP.t1272 6.541
R1355 VP.n1728 VP.t1079 6.541
R1356 VP.n1719 VP.n1718 6.541
R1357 VP.n1443 VP.t1283 6.541
R1358 VP.n10094 VP.n10093 6.541
R1359 VP.n10098 VP.t1107 6.541
R1360 VP.n10079 VP.n10078 6.541
R1361 VP.n10081 VP.t1350 6.541
R1362 VP.n2590 VP.t558 6.105
R1363 VP.n2843 VP.t1259 6.105
R1364 VP.n2846 VP.n2845 6.105
R1365 VP.n2838 VP.t541 6.105
R1366 VP.n2821 VP.n2820 6.105
R1367 VP.n3393 VP.t1167 6.105
R1368 VP.n3396 VP.n3395 6.105
R1369 VP.n3388 VP.t463 6.105
R1370 VP.n3372 VP.n3371 6.105
R1371 VP.n3788 VP.t1147 6.105
R1372 VP.n3791 VP.n3790 6.105
R1373 VP.n3783 VP.t440 6.105
R1374 VP.n3761 VP.n3760 6.105
R1375 VP.n4312 VP.t213 6.105
R1376 VP.n4315 VP.n4314 6.105
R1377 VP.n4307 VP.t805 6.105
R1378 VP.n4293 VP.n4292 6.105
R1379 VP.n4687 VP.t199 6.105
R1380 VP.n4690 VP.n4689 6.105
R1381 VP.n4682 VP.t789 6.105
R1382 VP.n4667 VP.n4666 6.105
R1383 VP.n5217 VP.t813 6.105
R1384 VP.n5220 VP.n5219 6.105
R1385 VP.n5212 VP.t64 6.105
R1386 VP.n5199 VP.n5198 6.105
R1387 VP.n5582 VP.t939 6.105
R1388 VP.n5585 VP.n5584 6.105
R1389 VP.n5577 VP.t1312 6.105
R1390 VP.n5562 VP.n5561 6.105
R1391 VP.n6082 VP.t75 6.105
R1392 VP.n6085 VP.n6084 6.105
R1393 VP.n6077 VP.t683 6.105
R1394 VP.n6064 VP.n6063 6.105
R1395 VP.n6438 VP.t160 6.105
R1396 VP.n6441 VP.n6440 6.105
R1397 VP.n6433 VP.t757 6.105
R1398 VP.n6418 VP.n6417 6.105
R1399 VP.n6946 VP.t689 6.105
R1400 VP.n6949 VP.n6948 6.105
R1401 VP.n6941 VP.t1284 6.105
R1402 VP.n6928 VP.n6927 6.105
R1403 VP.n7297 VP.t767 6.105
R1404 VP.n7300 VP.n7299 6.105
R1405 VP.n7292 VP.t3 6.105
R1406 VP.n7277 VP.n7276 6.105
R1407 VP.n7784 VP.t1291 6.105
R1408 VP.n7787 VP.n7786 6.105
R1409 VP.n7779 VP.t573 6.105
R1410 VP.n7766 VP.n7765 6.105
R1411 VP.n8125 VP.t19 6.105
R1412 VP.n8128 VP.n8127 6.105
R1413 VP.n8120 VP.t649 6.105
R1414 VP.n8105 VP.n8104 6.105
R1415 VP.n8623 VP.t585 6.105
R1416 VP.n8626 VP.n8625 6.105
R1417 VP.n8618 VP.t1168 6.105
R1418 VP.n8605 VP.n8604 6.105
R1419 VP.n8969 VP.t655 6.105
R1420 VP.n8972 VP.n8971 6.105
R1421 VP.n8964 VP.t1243 6.105
R1422 VP.n8949 VP.n8948 6.105
R1423 VP.n9422 VP.t1329 6.105
R1424 VP.n9425 VP.n9424 6.105
R1425 VP.n9417 VP.t474 6.105
R1426 VP.n9402 VP.n9401 6.105
R1427 VP.n10760 VP.t629 6.105
R1428 VP.n10763 VP.n10762 6.105
R1429 VP.n10755 VP.t1138 6.105
R1430 VP.n10747 VP.n10746 6.105
R1431 VP.n10166 VP.t539 6.105
R1432 VP.n10169 VP.n10168 6.105
R1433 VP.n10161 VP.t1123 6.105
R1434 VP.n10152 VP.n10151 6.105
R1435 VP.n10206 VP.t1050 6.105
R1436 VP.n10353 VP.t462 6.105
R1437 VP.n2245 VP.t1104 6.105
R1438 VP.n2265 VP.n2264 6.105
R1439 VP.n2268 VP.n2267 6.105
R1440 VP.n2248 VP.t395 6.105
R1441 VP.n2332 VP.t1018 6.105
R1442 VP.n2343 VP.n2342 6.105
R1443 VP.n2340 VP.n2339 6.105
R1444 VP.n2335 VP.t310 6.105
R1445 VP.n3196 VP.t1003 6.105
R1446 VP.n3215 VP.n3214 6.105
R1447 VP.n3218 VP.n3217 6.105
R1448 VP.n3199 VP.t288 6.105
R1449 VP.n3359 VP.t323 6.105
R1450 VP.n3369 VP.n3368 6.105
R1451 VP.n3366 VP.n3365 6.105
R1452 VP.n3362 VP.t914 6.105
R1453 VP.n4087 VP.t299 6.105
R1454 VP.n4107 VP.n4106 6.105
R1455 VP.n4110 VP.n4109 6.105
R1456 VP.n4090 VP.t890 6.105
R1457 VP.n4280 VP.t661 6.105
R1458 VP.n4290 VP.n4289 6.105
R1459 VP.n4287 VP.n4286 6.105
R1460 VP.n4283 VP.t1250 6.105
R1461 VP.n4970 VP.t647 6.105
R1462 VP.n4990 VP.n4989 6.105
R1463 VP.n4993 VP.n4992 6.105
R1464 VP.n4973 VP.t1156 6.105
R1465 VP.n5186 VP.t1257 6.105
R1466 VP.n5196 VP.n5195 6.105
R1467 VP.n5193 VP.n5192 6.105
R1468 VP.n5189 VP.t540 6.105
R1469 VP.n5807 VP.t1321 6.105
R1470 VP.n5827 VP.n5826 6.105
R1471 VP.n5830 VP.n5829 6.105
R1472 VP.n5810 VP.t464 6.105
R1473 VP.n6050 VP.t549 6.105
R1474 VP.n6061 VP.n6060 6.105
R1475 VP.n6058 VP.n6057 6.105
R1476 VP.n6053 VP.t1131 6.105
R1477 VP.n6651 VP.t622 6.105
R1478 VP.n6670 VP.n6669 6.105
R1479 VP.n6673 VP.n6672 6.105
R1480 VP.n6654 VP.t1206 6.105
R1481 VP.n6914 VP.t1137 6.105
R1482 VP.n6925 VP.n6924 6.105
R1483 VP.n6922 VP.n6921 6.105
R1484 VP.n6917 VP.t428 6.105
R1485 VP.n7463 VP.t1214 6.105
R1486 VP.n7482 VP.n7481 6.105
R1487 VP.n7485 VP.n7484 6.105
R1488 VP.n7466 VP.t499 6.105
R1489 VP.n7753 VP.t437 6.105
R1490 VP.n7763 VP.n7762 6.105
R1491 VP.n7760 VP.n7759 6.105
R1492 VP.n7756 VP.t1020 6.105
R1493 VP.n8279 VP.t508 6.105
R1494 VP.n8299 VP.n8298 6.105
R1495 VP.n8302 VP.n8301 6.105
R1496 VP.n8282 VP.t1091 6.105
R1497 VP.n8592 VP.t1033 6.105
R1498 VP.n8602 VP.n8601 6.105
R1499 VP.n8599 VP.n8598 6.105
R1500 VP.n8595 VP.t325 6.105
R1501 VP.n9076 VP.t1096 6.105
R1502 VP.n9096 VP.n9095 6.105
R1503 VP.n9099 VP.n9098 6.105
R1504 VP.n9079 VP.t387 6.105
R1505 VP.n9388 VP.t482 6.105
R1506 VP.n9399 VP.n9398 6.105
R1507 VP.n9396 VP.n9395 6.105
R1508 VP.n9391 VP.t853 6.105
R1509 VP.n9839 VP.t393 6.105
R1510 VP.n9858 VP.n9857 6.105
R1511 VP.n9861 VP.n9860 6.105
R1512 VP.n9842 VP.t979 6.105
R1513 VP.n10733 VP.t309 6.105
R1514 VP.n10744 VP.n10743 6.105
R1515 VP.n10741 VP.n10740 6.105
R1516 VP.n10736 VP.t903 6.105
R1517 VP.n10458 VP.t287 6.105
R1518 VP.n10466 VP.n10465 6.105
R1519 VP.n10469 VP.n10468 6.105
R1520 VP.n10461 VP.t879 6.105
R1521 VP.n10204 VP.t197 6.105
R1522 VP.n10191 VP.t913 6.105
R1523 VP.n10342 VP.t631 6.105
R1524 VP.n10336 VP.t379 6.105
R1525 VP.n10327 VP.t1092 6.105
R1526 VP.n10423 VP.t1170 6.105
R1527 VP.n10434 VP.n10433 6.105
R1528 VP.n10431 VP.n10430 6.105
R1529 VP.n10426 VP.t465 6.105
R1530 VP.n10954 VP.t483 6.105
R1531 VP.n9602 VP.t185 6.105
R1532 VP.n10053 VP.t1022 6.105
R1533 VP.n10073 VP.n10072 6.105
R1534 VP.n10076 VP.n10075 6.105
R1535 VP.n10050 VP.t312 6.105
R1536 VP.n10983 VP.t945 6.105
R1537 VP.n11007 VP.n11006 6.105
R1538 VP.n11010 VP.n11009 6.105
R1539 VP.n10980 VP.t228 6.105
R1540 VP.n10620 VP.t931 6.105
R1541 VP.n10644 VP.n10643 6.105
R1542 VP.n10647 VP.n10646 6.105
R1543 VP.n10617 VP.t214 6.105
R1544 VP.n10324 VP.t831 6.105
R1545 VP.n10311 VP.t237 6.105
R1546 VP.n8796 VP.t1339 6.105
R1547 VP.n9257 VP.t876 6.105
R1548 VP.n9275 VP.n9274 6.105
R1549 VP.n9278 VP.n9277 6.105
R1550 VP.n9254 VP.t157 6.105
R1551 VP.n9618 VP.t802 6.105
R1552 VP.n9635 VP.n9634 6.105
R1553 VP.n9638 VP.n9637 6.105
R1554 VP.n9615 VP.t1240 6.105
R1555 VP.n10013 VP.t787 6.105
R1556 VP.n10042 VP.n10041 6.105
R1557 VP.n10045 VP.n10044 6.105
R1558 VP.n10010 VP.t32 6.105
R1559 VP.n10924 VP.t62 6.105
R1560 VP.n10951 VP.n10950 6.105
R1561 VP.n10948 VP.n10947 6.105
R1562 VP.n10921 VP.t674 6.105
R1563 VP.n10582 VP.t42 6.105
R1564 VP.n10606 VP.n10605 6.105
R1565 VP.n10609 VP.n10608 6.105
R1566 VP.n10579 VP.t662 6.105
R1567 VP.n10306 VP.t1276 6.105
R1568 VP.n10295 VP.t682 6.105
R1569 VP.n8756 VP.t505 6.105
R1570 VP.n8775 VP.n8774 6.105
R1571 VP.n8772 VP.n8771 6.105
R1572 VP.n8753 VP.t1088 6.105
R1573 VP.n9036 VP.t639 6.105
R1574 VP.n9048 VP.n9047 6.105
R1575 VP.n9045 VP.n9044 6.105
R1576 VP.n9039 VP.t1223 6.105
R1577 VP.n9568 VP.t1247 6.105
R1578 VP.n9579 VP.n9578 6.105
R1579 VP.n9576 VP.n9575 6.105
R1580 VP.n9571 VP.t384 6.105
R1581 VP.n9801 VP.t1233 6.105
R1582 VP.n9812 VP.n9811 6.105
R1583 VP.n9809 VP.n9808 6.105
R1584 VP.n9804 VP.t514 6.105
R1585 VP.n10905 VP.t536 6.105
R1586 VP.n10916 VP.n10915 6.105
R1587 VP.n10913 VP.n10912 6.105
R1588 VP.n10908 VP.t1119 6.105
R1589 VP.n10400 VP.t521 6.105
R1590 VP.n10408 VP.n10407 6.105
R1591 VP.n10405 VP.n10404 6.105
R1592 VP.n10397 VP.t1045 6.105
R1593 VP.n10290 VP.t419 6.105
R1594 VP.n10283 VP.t1129 6.105
R1595 VP.n8199 VP.t726 6.105
R1596 VP.n8210 VP.n8209 6.105
R1597 VP.n8207 VP.n8206 6.105
R1598 VP.n8202 VP.t1318 6.105
R1599 VP.n7905 VP.t1192 6.105
R1600 VP.n7073 VP.t1043 6.105
R1601 VP.n7591 VP.t581 6.105
R1602 VP.n7609 VP.n7608 6.105
R1603 VP.n7612 VP.n7611 6.105
R1604 VP.n7588 VP.t1165 6.105
R1605 VP.n7953 VP.t359 6.105
R1606 VP.n7970 VP.n7969 6.105
R1607 VP.n7973 VP.n7972 6.105
R1608 VP.n7950 VP.t943 6.105
R1609 VP.n8419 VP.t491 6.105
R1610 VP.n8448 VP.n8447 6.105
R1611 VP.n8451 VP.n8450 6.105
R1612 VP.n8416 VP.t1074 6.105
R1613 VP.n8729 VP.t951 6.105
R1614 VP.n8749 VP.n8748 6.105
R1615 VP.n8746 VP.n8745 6.105
R1616 VP.n8726 VP.t233 6.105
R1617 VP.n9219 VP.t1082 6.105
R1618 VP.n9246 VP.n9245 6.105
R1619 VP.n9249 VP.n9248 6.105
R1620 VP.n9216 VP.t368 6.105
R1621 VP.n9535 VP.t390 6.105
R1622 VP.n9556 VP.n9555 6.105
R1623 VP.n9553 VP.n9552 6.105
R1624 VP.n9532 VP.t835 6.105
R1625 VP.n9976 VP.t376 6.105
R1626 VP.n10002 VP.n10001 6.105
R1627 VP.n10005 VP.n10004 6.105
R1628 VP.n9973 VP.t900 6.105
R1629 VP.n10873 VP.t984 6.105
R1630 VP.n10900 VP.n10899 6.105
R1631 VP.n10897 VP.n10896 6.105
R1632 VP.n10870 VP.t264 6.105
R1633 VP.n10547 VP.t908 6.105
R1634 VP.n10571 VP.n10570 6.105
R1635 VP.n10574 VP.n10573 6.105
R1636 VP.n10544 VP.t193 6.105
R1637 VP.n10278 VP.t866 6.105
R1638 VP.n10267 VP.t273 6.105
R1639 VP.n7033 VP.t211 6.105
R1640 VP.n7052 VP.n7051 6.105
R1641 VP.n7049 VP.n7048 6.105
R1642 VP.n7030 VP.t799 6.105
R1643 VP.n7341 VP.t345 6.105
R1644 VP.n7353 VP.n7352 6.105
R1645 VP.n7350 VP.n7349 6.105
R1646 VP.n7344 VP.t928 6.105
R1647 VP.n7876 VP.t808 6.105
R1648 VP.n7886 VP.n7885 6.105
R1649 VP.n7883 VP.n7882 6.105
R1650 VP.n7879 VP.t56 6.105
R1651 VP.n8162 VP.t937 6.105
R1652 VP.n8174 VP.n8173 6.105
R1653 VP.n8171 VP.n8170 6.105
R1654 VP.n8165 VP.t219 6.105
R1655 VP.n8712 VP.t67 6.105
R1656 VP.n8722 VP.n8721 6.105
R1657 VP.n8719 VP.n8718 6.105
R1658 VP.n8715 VP.t678 6.105
R1659 VP.n9006 VP.t226 6.105
R1660 VP.n9018 VP.n9017 6.105
R1661 VP.n9015 VP.n9014 6.105
R1662 VP.n9009 VP.t751 6.105
R1663 VP.n9516 VP.t842 6.105
R1664 VP.n9527 VP.n9526 6.105
R1665 VP.n9524 VP.n9523 6.105
R1666 VP.n9519 VP.t1279 6.105
R1667 VP.n9779 VP.t759 6.105
R1668 VP.n9790 VP.n9789 6.105
R1669 VP.n9787 VP.n9786 6.105
R1670 VP.n9782 VP.t1347 6.105
R1671 VP.n10854 VP.t110 6.105
R1672 VP.n10865 VP.n10864 6.105
R1673 VP.n10862 VP.n10861 6.105
R1674 VP.n10857 VP.t710 6.105
R1675 VP.n10383 VP.t7 6.105
R1676 VP.n10391 VP.n10390 6.105
R1677 VP.n10388 VP.n10387 6.105
R1678 VP.n10380 VP.t643 6.105
R1679 VP.n10262 VP.t1315 6.105
R1680 VP.n10255 VP.t720 6.105
R1681 VP.n6489 VP.t434 6.105
R1682 VP.n6500 VP.n6499 6.105
R1683 VP.n6497 VP.n6496 6.105
R1684 VP.n6492 VP.t1015 6.105
R1685 VP.n6154 VP.t897 6.105
R1686 VP.n5294 VP.t748 6.105
R1687 VP.n5888 VP.t280 6.105
R1688 VP.n5906 VP.n5905 6.105
R1689 VP.n5909 VP.n5908 6.105
R1690 VP.n5885 VP.t722 6.105
R1691 VP.n6266 VP.t25 6.105
R1692 VP.n6283 VP.n6282 6.105
R1693 VP.n6286 VP.n6285 6.105
R1694 VP.n6263 VP.t651 6.105
R1695 VP.n6741 VP.t191 6.105
R1696 VP.n6770 VP.n6769 6.105
R1697 VP.n6773 VP.n6772 6.105
R1698 VP.n6738 VP.t783 6.105
R1699 VP.n7006 VP.t657 6.105
R1700 VP.n7026 VP.n7025 6.105
R1701 VP.n7023 VP.n7022 6.105
R1702 VP.n7003 VP.t1245 6.105
R1703 VP.n7553 VP.t791 6.105
R1704 VP.n7580 VP.n7579 6.105
R1705 VP.n7583 VP.n7582 6.105
R1706 VP.n7550 VP.t37 6.105
R1707 VP.n7844 VP.t1253 6.105
R1708 VP.n7864 VP.n7863 6.105
R1709 VP.n7861 VP.n7860 6.105
R1710 VP.n7841 VP.t533 6.105
R1711 VP.n8370 VP.t48 6.105
R1712 VP.n8397 VP.n8396 6.105
R1713 VP.n8400 VP.n8399 6.105
R1714 VP.n8367 VP.t605 6.105
R1715 VP.n8681 VP.t544 6.105
R1716 VP.n8701 VP.n8700 6.105
R1717 VP.n8698 VP.n8697 6.105
R1718 VP.n8678 VP.t1125 6.105
R1719 VP.n9169 VP.t614 6.105
R1720 VP.n9196 VP.n9195 6.105
R1721 VP.n9199 VP.n9198 6.105
R1722 VP.n9166 VP.t1200 6.105
R1723 VP.n9484 VP.t1286 6.105
R1724 VP.n9505 VP.n9504 6.105
R1725 VP.n9502 VP.n9501 6.105
R1726 VP.n9481 VP.t425 6.105
R1727 VP.n9928 VP.t1208 6.105
R1728 VP.n9954 VP.n9953 6.105
R1729 VP.n9957 VP.n9956 6.105
R1730 VP.n9925 VP.t496 6.105
R1731 VP.n10822 VP.t577 6.105
R1732 VP.n10849 VP.n10848 6.105
R1733 VP.n10846 VP.n10845 6.105
R1734 VP.n10819 VP.t1159 6.105
R1735 VP.n10512 VP.t500 6.105
R1736 VP.n10536 VP.n10535 6.105
R1737 VP.n10539 VP.n10538 6.105
R1738 VP.n10509 VP.t1086 6.105
R1739 VP.n10250 VP.t469 6.105
R1740 VP.n10239 VP.t1173 6.105
R1741 VP.n5254 VP.t1218 6.105
R1742 VP.n5273 VP.n5272 6.105
R1743 VP.n5270 VP.n5269 6.105
R1744 VP.n5251 VP.t501 6.105
R1745 VP.n5603 VP.t1345 6.105
R1746 VP.n5615 VP.n5614 6.105
R1747 VP.n5612 VP.n5611 6.105
R1748 VP.n5606 VP.t488 6.105
R1749 VP.n6125 VP.t509 6.105
R1750 VP.n6135 VP.n6134 6.105
R1751 VP.n6132 VP.n6131 6.105
R1752 VP.n6128 VP.t1094 6.105
R1753 VP.n6452 VP.t641 6.105
R1754 VP.n6464 VP.n6463 6.105
R1755 VP.n6461 VP.n6460 6.105
R1756 VP.n6455 VP.t1228 6.105
R1757 VP.n6988 VP.t1099 6.105
R1758 VP.n6998 VP.n6997 6.105
R1759 VP.n6995 VP.n6994 6.105
R1760 VP.n6991 VP.t388 6.105
R1761 VP.n7311 VP.t1236 6.105
R1762 VP.n7323 VP.n7322 6.105
R1763 VP.n7320 VP.n7319 6.105
R1764 VP.n7314 VP.t455 6.105
R1765 VP.n7826 VP.t397 6.105
R1766 VP.n7836 VP.n7835 6.105
R1767 VP.n7833 VP.n7832 6.105
R1768 VP.n7829 VP.t980 6.105
R1769 VP.n8139 VP.t468 6.105
R1770 VP.n8151 VP.n8150 6.105
R1771 VP.n8148 VP.n8147 6.105
R1772 VP.n8142 VP.t1054 6.105
R1773 VP.n8664 VP.t990 6.105
R1774 VP.n8674 VP.n8673 6.105
R1775 VP.n8671 VP.n8670 6.105
R1776 VP.n8667 VP.t270 6.105
R1777 VP.n8983 VP.t1062 6.105
R1778 VP.n8995 VP.n8994 6.105
R1779 VP.n8992 VP.n8991 6.105
R1780 VP.n8986 VP.t350 6.105
R1781 VP.n9465 VP.t431 6.105
R1782 VP.n9476 VP.n9475 6.105
R1783 VP.n9473 VP.n9472 6.105
R1784 VP.n9468 VP.t871 6.105
R1785 VP.n9757 VP.t355 6.105
R1786 VP.n9768 VP.n9767 6.105
R1787 VP.n9765 VP.n9764 6.105
R1788 VP.n9760 VP.t941 6.105
R1789 VP.n10803 VP.t1025 6.105
R1790 VP.n10814 VP.n10813 6.105
R1791 VP.n10811 VP.n10810 6.105
R1792 VP.n10806 VP.t316 6.105
R1793 VP.n10366 VP.t948 6.105
R1794 VP.n10374 VP.n10373 6.105
R1795 VP.n10371 VP.n10370 6.105
R1796 VP.n10363 VP.t231 6.105
R1797 VP.n10234 VP.t919 6.105
R1798 VP.n10227 VP.t329 6.105
R1799 VP.n4715 VP.t1294 6.105
R1800 VP.n4726 VP.n4725 6.105
R1801 VP.n4723 VP.n4722 6.105
R1802 VP.n4718 VP.t579 6.105
R1803 VP.n4334 VP.t602 6.105
R1804 VP.n3417 VP.t698 6.105
R1805 VP.n4118 VP.t77 6.105
R1806 VP.n4136 VP.n4135 6.105
R1807 VP.n4139 VP.n4138 6.105
R1808 VP.n4115 VP.t684 6.105
R1809 VP.n4515 VP.t1068 6.105
R1810 VP.n4532 VP.n4531 6.105
R1811 VP.n4535 VP.n4534 6.105
R1812 VP.n4512 VP.t354 6.105
R1813 VP.n5013 VP.t1052 6.105
R1814 VP.n5042 VP.n5041 6.105
R1815 VP.n5045 VP.n5044 6.105
R1816 VP.n5010 VP.t343 6.105
R1817 VP.n5227 VP.t362 6.105
R1818 VP.n5247 VP.n5246 6.105
R1819 VP.n5244 VP.n5243 6.105
R1820 VP.n5224 VP.t947 6.105
R1821 VP.n5850 VP.t494 6.105
R1822 VP.n5877 VP.n5876 6.105
R1823 VP.n5880 VP.n5879 6.105
R1824 VP.n5847 VP.t934 6.105
R1825 VP.n6093 VP.t957 6.105
R1826 VP.n6113 VP.n6112 6.105
R1827 VP.n6110 VP.n6109 6.105
R1828 VP.n6090 VP.t239 6.105
R1829 VP.n6692 VP.t1084 6.105
R1830 VP.n6719 VP.n6718 6.105
R1831 VP.n6722 VP.n6721 6.105
R1832 VP.n6689 VP.t304 6.105
R1833 VP.n6957 VP.t245 6.105
R1834 VP.n6977 VP.n6976 6.105
R1835 VP.n6974 VP.n6973 6.105
R1836 VP.n6954 VP.t839 6.105
R1837 VP.n7504 VP.t314 6.105
R1838 VP.n7531 VP.n7530 6.105
R1839 VP.n7534 VP.n7533 6.105
R1840 VP.n7501 VP.t906 6.105
R1841 VP.n7795 VP.t847 6.105
R1842 VP.n7815 VP.n7814 6.105
R1843 VP.n7812 VP.n7811 6.105
R1844 VP.n7792 VP.t104 6.105
R1845 VP.n8321 VP.t917 6.105
R1846 VP.n8348 VP.n8347 6.105
R1847 VP.n8351 VP.n8350 6.105
R1848 VP.n8318 VP.t201 6.105
R1849 VP.n8633 VP.t118 6.105
R1850 VP.n8653 VP.n8652 6.105
R1851 VP.n8650 VP.n8649 6.105
R1852 VP.n8630 VP.t716 6.105
R1853 VP.n9119 VP.t208 6.105
R1854 VP.n9146 VP.n9145 6.105
R1855 VP.n9149 VP.n9148 6.105
R1856 VP.n9116 VP.t796 6.105
R1857 VP.n9433 VP.t880 6.105
R1858 VP.n9454 VP.n9453 6.105
R1859 VP.n9451 VP.n9450 6.105
R1860 VP.n9430 VP.t1322 6.105
R1861 VP.n9880 VP.t804 6.105
R1862 VP.n9906 VP.n9905 6.105
R1863 VP.n9909 VP.n9908 6.105
R1864 VP.n9877 VP.t52 6.105
R1865 VP.n10771 VP.t175 6.105
R1866 VP.n10798 VP.n10797 6.105
R1867 VP.n10795 VP.n10794 6.105
R1868 VP.n10768 VP.t769 6.105
R1869 VP.n10477 VP.t63 6.105
R1870 VP.n10501 VP.n10500 6.105
R1871 VP.n10504 VP.n10503 6.105
R1872 VP.n10474 VP.t676 6.105
R1873 VP.n10222 VP.t1292 6.105
R1874 VP.n10211 VP.t778 6.105
R1875 VP.n342 VP.t94 6.105
R1876 VP.n867 VP.t961 6.105
R1877 VP.n878 VP.n877 6.105
R1878 VP.n875 VP.n874 6.105
R1879 VP.n870 VP.t242 6.105
R1880 VP.n1409 VP.t874 6.105
R1881 VP.n1419 VP.n1418 6.105
R1882 VP.n1416 VP.n1415 6.105
R1883 VP.n1412 VP.t155 6.105
R1884 VP.n1853 VP.t860 6.105
R1885 VP.n1865 VP.n1864 6.105
R1886 VP.n1862 VP.n1861 6.105
R1887 VP.n1856 VP.t128 6.105
R1888 VP.n2621 VP.t166 6.105
R1889 VP.n2628 VP.n2627 6.105
R1890 VP.n2631 VP.n2630 6.105
R1891 VP.n2624 VP.t764 6.105
R1892 VP.n2806 VP.t142 6.105
R1893 VP.n2818 VP.n2817 6.105
R1894 VP.n2815 VP.n2814 6.105
R1895 VP.n2809 VP.t740 6.105
R1896 VP.n3332 VP.t774 6.105
R1897 VP.n3342 VP.n3341 6.105
R1898 VP.n3339 VP.n3338 6.105
R1899 VP.n3335 VP.t13 6.105
R1900 VP.n3746 VP.t754 6.105
R1901 VP.n3758 VP.n3757 6.105
R1902 VP.n3755 VP.n3754 6.105
R1903 VP.n3749 VP.t1275 6.105
R1904 VP.n4253 VP.t1103 6.105
R1905 VP.n4263 VP.n4262 6.105
R1906 VP.n4260 VP.n4259 6.105
R1907 VP.n4256 VP.t394 6.105
R1908 VP.n4652 VP.t1019 6.105
R1909 VP.n4664 VP.n4663 6.105
R1910 VP.n4661 VP.n4660 6.105
R1911 VP.n4655 VP.t311 6.105
R1912 VP.n5159 VP.t403 6.105
R1913 VP.n5169 VP.n5168 6.105
R1914 VP.n5166 VP.n5165 6.105
R1915 VP.n5162 VP.t987 6.105
R1916 VP.n5547 VP.t473 6.105
R1917 VP.n5559 VP.n5558 6.105
R1918 VP.n5556 VP.n5555 6.105
R1919 VP.n5550 VP.t915 6.105
R1920 VP.n6023 VP.t995 6.105
R1921 VP.n6033 VP.n6032 6.105
R1922 VP.n6030 VP.n6029 6.105
R1923 VP.n6026 VP.t276 6.105
R1924 VP.n6403 VP.t1067 6.105
R1925 VP.n6415 VP.n6414 6.105
R1926 VP.n6412 VP.n6411 6.105
R1927 VP.n6406 VP.t353 6.105
R1928 VP.n6887 VP.t285 6.105
R1929 VP.n6897 VP.n6896 6.105
R1930 VP.n6894 VP.n6893 6.105
R1931 VP.n6890 VP.t875 6.105
R1932 VP.n7262 VP.t361 6.105
R1933 VP.n7274 VP.n7273 6.105
R1934 VP.n7271 VP.n7270 6.105
R1935 VP.n7265 VP.t944 6.105
R1936 VP.n7726 VP.t886 6.105
R1937 VP.n7736 VP.n7735 6.105
R1938 VP.n7733 VP.n7732 6.105
R1939 VP.n7729 VP.t171 6.105
R1940 VP.n8090 VP.t954 6.105
R1941 VP.n8102 VP.n8101 6.105
R1942 VP.n8099 VP.n8098 6.105
R1943 VP.n8093 VP.t236 6.105
R1944 VP.n8565 VP.t182 6.105
R1945 VP.n8575 VP.n8574 6.105
R1946 VP.n8572 VP.n8571 6.105
R1947 VP.n8568 VP.t695 6.105
R1948 VP.n8934 VP.t241 6.105
R1949 VP.n8946 VP.n8945 6.105
R1950 VP.n8943 VP.n8942 6.105
R1951 VP.n8937 VP.t838 6.105
R1952 VP.n9359 VP.t152 6.105
R1953 VP.n9370 VP.n9369 6.105
R1954 VP.n9367 VP.n9366 6.105
R1955 VP.n9362 VP.t609 6.105
R1956 VP.n9735 VP.t127 6.105
R1957 VP.n9746 VP.n9745 6.105
R1958 VP.n9743 VP.n9742 6.105
R1959 VP.n9738 VP.t729 6.105
R1960 VP.n10704 VP.t762 6.105
R1961 VP.n10715 VP.n10714 6.105
R1962 VP.n10712 VP.n10711 6.105
R1963 VP.n10707 VP.t1349 6.105
R1964 VP.n10138 VP.t739 6.105
R1965 VP.n10149 VP.n10148 6.105
R1966 VP.n10146 VP.n10145 6.105
R1967 VP.n10141 VP.t1331 6.105
R1968 VP.n10339 VP.t645 6.105
R1969 VP.n10340 VP.t9 6.105
R1970 VP.n129 VP.t833 6.105
R1971 VP.n10125 VP.t1191 6.105
R1972 VP.n10649 VP.t481 6.105
R1973 VP.n10689 VP.t1209 6.105
R1974 VP.n11013 VP.n11012 6.105
R1975 VP.n11016 VP.n11015 6.105
R1976 VP.n11019 VP.t498 6.105
R1977 VP.n9702 VP.t593 6.105
R1978 VP.n9724 VP.n9723 6.105
R1979 VP.n9721 VP.n9720 6.105
R1980 VP.n9705 VP.t1181 6.105
R1981 VP.n9337 VP.t617 6.105
R1982 VP.n9348 VP.n9347 6.105
R1983 VP.n9345 VP.n9344 6.105
R1984 VP.n9340 VP.t1056 6.105
R1985 VP.n8911 VP.t1299 6.105
R1986 VP.n8923 VP.n8922 6.105
R1987 VP.n8920 VP.n8919 6.105
R1988 VP.n8914 VP.t584 6.105
R1989 VP.n8544 VP.t1162 6.105
R1990 VP.n8554 VP.n8553 6.105
R1991 VP.n8551 VP.n8550 6.105
R1992 VP.n8547 VP.t458 6.105
R1993 VP.n8067 VP.t71 6.105
R1994 VP.n8079 VP.n8078 6.105
R1995 VP.n8076 VP.n8075 6.105
R1996 VP.n8070 VP.t680 6.105
R1997 VP.n7705 VP.t1336 6.105
R1998 VP.n7715 VP.n7714 6.105
R1999 VP.n7712 VP.n7711 6.105
R2000 VP.n7708 VP.t553 6.105
R2001 VP.n7239 VP.t810 6.105
R2002 VP.n7251 VP.n7250 6.105
R2003 VP.n7248 VP.n7247 6.105
R2004 VP.n7242 VP.t59 6.105
R2005 VP.n6866 VP.t736 6.105
R2006 VP.n6876 VP.n6875 6.105
R2007 VP.n6873 VP.n6872 6.105
R2008 VP.n6869 VP.t1326 6.105
R2009 VP.n6380 VP.t212 6.105
R2010 VP.n6392 VP.n6391 6.105
R2011 VP.n6389 VP.n6388 6.105
R2012 VP.n6383 VP.t801 6.105
R2013 VP.n6002 VP.t125 6.105
R2014 VP.n6012 VP.n6011 6.105
R2015 VP.n6009 VP.n6008 6.105
R2016 VP.n6005 VP.t725 6.105
R2017 VP.n5524 VP.t923 6.105
R2018 VP.n5536 VP.n5535 6.105
R2019 VP.n5533 VP.n5532 6.105
R2020 VP.n5527 VP.t15 6.105
R2021 VP.n5138 VP.t852 6.105
R2022 VP.n5148 VP.n5147 6.105
R2023 VP.n5145 VP.n5144 6.105
R2024 VP.n5141 VP.t114 6.105
R2025 VP.n4629 VP.t170 6.105
R2026 VP.n4641 VP.n4640 6.105
R2027 VP.n4638 VP.n4637 6.105
R2028 VP.n4632 VP.t765 6.105
R2029 VP.n4232 VP.t250 6.105
R2030 VP.n4242 VP.n4241 6.105
R2031 VP.n4239 VP.n4238 6.105
R2032 VP.n4235 VP.t845 6.105
R2033 VP.n3723 VP.t1126 6.105
R2034 VP.n3735 VP.n3734 6.105
R2035 VP.n3732 VP.n3731 6.105
R2036 VP.n3726 VP.t420 6.105
R2037 VP.n3311 VP.t1221 6.105
R2038 VP.n3321 VP.n3320 6.105
R2039 VP.n3318 VP.n3317 6.105
R2040 VP.n3314 VP.t503 6.105
R2041 VP.n2783 VP.t608 6.105
R2042 VP.n2795 VP.n2794 6.105
R2043 VP.n2792 VP.n2791 6.105
R2044 VP.n2786 VP.t1120 6.105
R2045 VP.n2646 VP.t626 6.105
R2046 VP.n2653 VP.n2652 6.105
R2047 VP.n2656 VP.n2655 6.105
R2048 VP.n2649 VP.t1211 6.105
R2049 VP.n1823 VP.t1307 6.105
R2050 VP.n1835 VP.n1834 6.105
R2051 VP.n1832 VP.n1831 6.105
R2052 VP.n1826 VP.t594 6.105
R2053 VP.n1385 VP.t1325 6.105
R2054 VP.n1395 VP.n1394 6.105
R2055 VP.n1392 VP.n1391 6.105
R2056 VP.n1388 VP.t619 6.105
R2057 VP.n839 VP.t704 6.105
R2058 VP.n849 VP.n848 6.105
R2059 VP.n820 VP.n819 6.105
R2060 VP.n842 VP.t1300 6.105
R2061 VP.n296 VP.t724 6.105
R2062 VP.n318 VP.n317 6.105
R2063 VP.n315 VP.n314 6.105
R2064 VP.n299 VP.t1163 6.105
R2065 VP.n146 VP.t818 6.105
R2066 VP.n206 VP.t382 6.105
R2067 VP.n267 VP.t992 6.105
R2068 VP.n730 VP.n729 6.105
R2069 VP.n733 VP.n732 6.105
R2070 VP.n736 VP.t107 6.105
R2071 VP.n776 VP.t975 6.105
R2072 VP.n1291 VP.t256 6.105
R2073 VP.n210 VP.t1238 6.105
R2074 VP.n370 VP.t545 6.105
R2075 VP.n394 VP.n393 6.105
R2076 VP.n397 VP.n396 6.105
R2077 VP.n373 VP.t982 6.105
R2078 VP.n906 VP.t527 6.105
R2079 VP.n926 VP.n925 6.105
R2080 VP.n929 VP.n928 6.105
R2081 VP.n909 VP.t1109 6.105
R2082 VP.n1339 VP.t1134 6.105
R2083 VP.n1731 VP.n1730 6.105
R2084 VP.n1734 VP.n1733 6.105
R2085 VP.n1737 VP.t427 6.105
R2086 VP.n1765 VP.t1118 6.105
R2087 VP.n2270 VP.t408 6.105
R2088 VP.n214 VP.t179 6.105
R2089 VP.n417 VP.t68 6.105
R2090 VP.n441 VP.n440 6.105
R2091 VP.n444 VP.n443 6.105
R2092 VP.n420 VP.t534 6.105
R2093 VP.n956 VP.t50 6.105
R2094 VP.n976 VP.n975 6.105
R2095 VP.n979 VP.n978 6.105
R2096 VP.n959 VP.t667 6.105
R2097 VP.n1468 VP.t686 6.105
R2098 VP.n1482 VP.n1481 6.105
R2099 VP.n1485 VP.n1484 6.105
R2100 VP.n1471 VP.t1281 6.105
R2101 VP.n1893 VP.t673 6.105
R2102 VP.n1915 VP.n1914 6.105
R2103 VP.n1918 VP.n1917 6.105
R2104 VP.n1896 VP.t1265 6.105
R2105 VP.n2315 VP.t1288 6.105
R2106 VP.n2692 VP.n2691 6.105
R2107 VP.n2695 VP.n2694 6.105
R2108 VP.n2698 VP.t570 6.105
R2109 VP.n2726 VP.t1274 6.105
R2110 VP.n3220 VP.t556 6.105
R2111 VP.n218 VP.t1031 6.105
R2112 VP.n464 VP.t410 6.105
R2113 VP.n488 VP.n487 6.105
R2114 VP.n491 VP.n490 6.105
R2115 VP.n467 VP.t792 6.105
R2116 VP.n1006 VP.t334 6.105
R2117 VP.n1026 VP.n1025 6.105
R2118 VP.n1029 VP.n1028 6.105
R2119 VP.n1009 VP.t921 6.105
R2120 VP.n1506 VP.t240 6.105
R2121 VP.n1520 VP.n1519 6.105
R2122 VP.n1523 VP.n1522 6.105
R2123 VP.n1509 VP.t836 6.105
R2124 VP.n1945 VP.t227 6.105
R2125 VP.n1967 VP.n1966 6.105
R2126 VP.n1970 VP.n1969 6.105
R2127 VP.n1948 VP.t820 6.105
R2128 VP.n2568 VP.t844 6.105
R2129 VP.n2585 VP.n2584 6.105
R2130 VP.n2582 VP.n2581 6.105
R2131 VP.n2571 VP.t101 6.105
R2132 VP.n2874 VP.t829 6.105
R2133 VP.n2896 VP.n2895 6.105
R2134 VP.n2899 VP.n2898 6.105
R2135 VP.n2877 VP.t84 6.105
R2136 VP.n3265 VP.t113 6.105
R2137 VP.n3632 VP.n3631 6.105
R2138 VP.n3635 VP.n3634 6.105
R2139 VP.n3638 VP.t713 6.105
R2140 VP.n3666 VP.t95 6.105
R2141 VP.n4141 VP.t696 6.105
R2142 VP.n222 VP.t583 6.105
R2143 VP.n511 VP.t1264 6.105
R2144 VP.n535 VP.n534 6.105
R2145 VP.n538 VP.n537 6.105
R2146 VP.n514 VP.t401 6.105
R2147 VP.n1056 VP.t1180 6.105
R2148 VP.n1076 VP.n1075 6.105
R2149 VP.n1079 VP.n1078 6.105
R2150 VP.n1059 VP.t472 6.105
R2151 VP.n1544 VP.t555 6.105
R2152 VP.n1558 VP.n1557 6.105
R2153 VP.n1561 VP.n1560 6.105
R2154 VP.n1547 VP.t1081 6.105
R2155 VP.n1997 VP.t480 6.105
R2156 VP.n2019 VP.n2018 6.105
R2157 VP.n2022 VP.n2021 6.105
R2158 VP.n2000 VP.t1066 6.105
R2159 VP.n2530 VP.t392 6.105
R2160 VP.n2547 VP.n2546 6.105
R2161 VP.n2544 VP.n2543 6.105
R2162 VP.n2533 VP.t977 6.105
R2163 VP.n2926 VP.t377 6.105
R2164 VP.n2948 VP.n2947 6.105
R2165 VP.n2951 VP.n2950 6.105
R2166 VP.n2929 VP.t963 6.105
R2167 VP.n3446 VP.t986 6.105
R2168 VP.n3460 VP.n3459 6.105
R2169 VP.n3463 VP.n3462 6.105
R2170 VP.n3449 VP.t267 6.105
R2171 VP.n3819 VP.t970 6.105
R2172 VP.n3841 VP.n3840 6.105
R2173 VP.n3844 VP.n3843 6.105
R2174 VP.n3822 VP.t251 6.105
R2175 VP.n4186 VP.t1328 6.105
R2176 VP.n4538 VP.n4537 6.105
R2177 VP.n4541 VP.n4540 6.105
R2178 VP.n4544 VP.t621 6.105
R2179 VP.n4572 VP.t1311 6.105
R2180 VP.n5047 VP.t599 6.105
R2181 VP.n226 VP.t117 6.105
R2182 VP.n558 VP.t821 6.105
R2183 VP.n582 VP.n581 6.105
R2184 VP.n585 VP.n584 6.105
R2185 VP.n561 VP.t1258 6.105
R2186 VP.n1106 VP.t728 6.105
R2187 VP.n1126 VP.n1125 6.105
R2188 VP.n1129 VP.n1128 6.105
R2189 VP.n1109 VP.t1320 6.105
R2190 VP.n1582 VP.t85 6.105
R2191 VP.n1596 VP.n1595 6.105
R2192 VP.n1599 VP.n1598 6.105
R2193 VP.n1585 VP.t688 6.105
R2194 VP.n2049 VP.t1330 6.105
R2195 VP.n2071 VP.n2070 6.105
R2196 VP.n2074 VP.n2073 6.105
R2197 VP.n2052 VP.t620 6.105
R2198 VP.n2492 VP.t697 6.105
R2199 VP.n2509 VP.n2508 6.105
R2200 VP.n2506 VP.n2505 6.105
R2201 VP.n2495 VP.t1232 6.105
R2202 VP.n2978 VP.t630 6.105
R2203 VP.n3000 VP.n2999 6.105
R2204 VP.n3003 VP.n3002 6.105
R2205 VP.n2981 VP.t1215 6.105
R2206 VP.n3484 VP.t538 6.105
R2207 VP.n3498 VP.n3497 6.105
R2208 VP.n3501 VP.n3500 6.105
R2209 VP.n3487 VP.t1122 6.105
R2210 VP.n3871 VP.t522 6.105
R2211 VP.n3893 VP.n3892 6.105
R2212 VP.n3896 VP.n3895 6.105
R2213 VP.n3874 VP.t1105 6.105
R2214 VP.n4363 VP.t877 6.105
R2215 VP.n4377 VP.n4376 6.105
R2216 VP.n4380 VP.n4379 6.105
R2217 VP.n4366 VP.t158 6.105
R2218 VP.n4754 VP.t863 6.105
R2219 VP.n4776 VP.n4775 6.105
R2220 VP.n4779 VP.n4778 6.105
R2221 VP.n4757 VP.t132 6.105
R2222 VP.n5092 VP.t173 6.105
R2223 VP.n5433 VP.n5432 6.105
R2224 VP.n5436 VP.n5435 6.105
R2225 VP.n5439 VP.t766 6.105
R2226 VP.n5467 VP.t303 6.105
R2227 VP.n5911 VP.t744 6.105
R2228 VP.n230 VP.t988 6.105
R2229 VP.n605 VP.t370 6.105
R2230 VP.n622 VP.n621 6.105
R2231 VP.n625 VP.n624 6.105
R2232 VP.n608 VP.t814 6.105
R2233 VP.n1156 VP.t278 6.105
R2234 VP.n1164 VP.n1163 6.105
R2235 VP.n1167 VP.n1166 6.105
R2236 VP.n1159 VP.t870 6.105
R2237 VP.n1620 VP.t964 6.105
R2238 VP.n1628 VP.n1627 6.105
R2239 VP.n1631 VP.n1630 6.105
R2240 VP.n1623 VP.t244 6.105
R2241 VP.n2101 VP.t878 6.105
R2242 VP.n2112 VP.n2111 6.105
R2243 VP.n2115 VP.n2114 6.105
R2244 VP.n2104 VP.t161 6.105
R2245 VP.n2460 VP.t252 6.105
R2246 VP.n2471 VP.n2470 6.105
R2247 VP.n2468 VP.n2467 6.105
R2248 VP.n2463 VP.t846 6.105
R2249 VP.n3030 VP.t174 6.105
R2250 VP.n3041 VP.n3040 6.105
R2251 VP.n3044 VP.n3043 6.105
R2252 VP.n3033 VP.t768 6.105
R2253 VP.n3522 VP.t854 6.105
R2254 VP.n3530 VP.n3529 6.105
R2255 VP.n3533 VP.n3532 6.105
R2256 VP.n3525 VP.t41 6.105
R2257 VP.n3923 VP.t777 6.105
R2258 VP.n3934 VP.n3933 6.105
R2259 VP.n3937 VP.n3936 6.105
R2260 VP.n3926 VP.t21 6.105
R2261 VP.n4401 VP.t429 6.105
R2262 VP.n4409 VP.n4408 6.105
R2263 VP.n4412 VP.n4411 6.105
R2264 VP.n4404 VP.t1011 6.105
R2265 VP.n4806 VP.t417 6.105
R2266 VP.n4817 VP.n4816 6.105
R2267 VP.n4820 VP.n4819 6.105
R2268 VP.n4809 VP.t998 6.105
R2269 VP.n5323 VP.t1023 6.105
R2270 VP.n5331 VP.n5330 6.105
R2271 VP.n5334 VP.n5333 6.105
R2272 VP.n5326 VP.t313 6.105
R2273 VP.n5643 VP.t1149 6.105
R2274 VP.n5654 VP.n5653 6.105
R2275 VP.n5657 VP.n5656 6.105
R2276 VP.n5646 VP.t291 6.105
R2277 VP.n5956 VP.t327 6.105
R2278 VP.n6289 VP.n6288 6.105
R2279 VP.n6292 VP.n6291 6.105
R2280 VP.n6295 VP.t916 6.105
R2281 VP.n6323 VP.t454 6.105
R2282 VP.n6775 VP.t1040 6.105
R2283 VP.n234 VP.t542 6.105
R2284 VP.n645 VP.t1225 6.105
R2285 VP.n652 VP.n651 6.105
R2286 VP.n655 VP.n654 6.105
R2287 VP.n648 VP.t363 6.105
R2288 VP.n1194 VP.t1132 6.105
R2289 VP.n1204 VP.n1203 6.105
R2290 VP.n1207 VP.n1206 6.105
R2291 VP.n1197 VP.t424 6.105
R2292 VP.n1652 VP.t516 6.105
R2293 VP.n1660 VP.n1659 6.105
R2294 VP.n1663 VP.n1662 6.105
R2295 VP.n1655 VP.t1098 6.105
R2296 VP.n2142 VP.t430 6.105
R2297 VP.n2153 VP.n2152 6.105
R2298 VP.n2156 VP.n2155 6.105
R2299 VP.n2145 VP.t1012 6.105
R2300 VP.n2428 VP.t1106 6.105
R2301 VP.n2439 VP.n2438 6.105
R2302 VP.n2436 VP.n2435 6.105
R2303 VP.n2431 VP.t396 6.105
R2304 VP.n3071 VP.t1024 6.105
R2305 VP.n3082 VP.n3081 6.105
R2306 VP.n3085 VP.n3084 6.105
R2307 VP.n3074 VP.t315 6.105
R2308 VP.n3554 VP.t404 6.105
R2309 VP.n3562 VP.n3561 6.105
R2310 VP.n3565 VP.n3564 6.105
R2311 VP.n3557 VP.t989 6.105
R2312 VP.n3964 VP.t328 6.105
R2313 VP.n3975 VP.n3974 6.105
R2314 VP.n3978 VP.n3977 6.105
R2315 VP.n3967 VP.t918 6.105
R2316 VP.n4433 VP.t746 6.105
R2317 VP.n4441 VP.n4440 6.105
R2318 VP.n4444 VP.n4443 6.105
R2319 VP.n4436 VP.t1269 6.105
R2320 VP.n4847 VP.t665 6.105
R2321 VP.n4858 VP.n4857 6.105
R2322 VP.n4861 VP.n4860 6.105
R2323 VP.n4850 VP.t1252 6.105
R2324 VP.n5355 VP.t575 6.105
R2325 VP.n5363 VP.n5362 6.105
R2326 VP.n5366 VP.n5365 6.105
R2327 VP.n5358 VP.t1157 6.105
R2328 VP.n5684 VP.t702 6.105
R2329 VP.n5695 VP.n5694 6.105
R2330 VP.n5698 VP.n5697 6.105
R2331 VP.n5687 VP.t1142 6.105
R2332 VP.n6183 VP.t1171 6.105
R2333 VP.n6191 VP.n6190 6.105
R2334 VP.n6194 VP.n6193 6.105
R2335 VP.n6186 VP.t466 6.105
R2336 VP.n6528 VP.t1304 6.105
R2337 VP.n6539 VP.n6538 6.105
R2338 VP.n6542 VP.n6541 6.105
R2339 VP.n6531 VP.t590 6.105
R2340 VP.n6820 VP.t476 6.105
R2341 VP.n7148 VP.n7147 6.105
R2342 VP.n7151 VP.n7150 6.105
R2343 VP.n7154 VP.t1061 6.105
R2344 VP.n7182 VP.t603 6.105
R2345 VP.n7614 VP.t1188 6.105
R2346 VP.n238 VP.t149 6.105
R2347 VP.n675 VP.t780 6.105
R2348 VP.n684 VP.n683 6.105
R2349 VP.n687 VP.n686 6.105
R2350 VP.n678 VP.t1217 6.105
R2351 VP.n1234 VP.t685 6.105
R2352 VP.n1245 VP.n1244 6.105
R2353 VP.n1248 VP.n1247 6.105
R2354 VP.n1237 VP.t1278 6.105
R2355 VP.n1684 VP.t35 6.105
R2356 VP.n1692 VP.n1691 6.105
R2357 VP.n1695 VP.n1694 6.105
R2358 VP.n1687 VP.t656 6.105
R2359 VP.n2183 VP.t1285 6.105
R2360 VP.n2194 VP.n2193 6.105
R2361 VP.n2197 VP.n2196 6.105
R2362 VP.n2186 VP.t567 6.105
R2363 VP.n2396 VP.t663 6.105
R2364 VP.n2407 VP.n2406 6.105
R2365 VP.n2404 VP.n2403 6.105
R2366 VP.n2399 VP.t1251 6.105
R2367 VP.n3112 VP.t576 6.105
R2368 VP.n3123 VP.n3122 6.105
R2369 VP.n3126 VP.n3125 6.105
R2370 VP.n3115 VP.t1158 6.105
R2371 VP.n3586 VP.t1260 6.105
R2372 VP.n3594 VP.n3593 6.105
R2373 VP.n3597 VP.n3596 6.105
R2374 VP.n3589 VP.t543 6.105
R2375 VP.n4005 VP.t1172 6.105
R2376 VP.n4016 VP.n4015 6.105
R2377 VP.n4019 VP.n4018 6.105
R2378 VP.n4008 VP.t467 6.105
R2379 VP.n4465 VP.t292 6.105
R2380 VP.n4473 VP.n4472 6.105
R2381 VP.n4476 VP.n4475 6.105
R2382 VP.n4468 VP.t883 6.105
R2383 VP.n4888 VP.t218 6.105
R2384 VP.n4899 VP.n4898 6.105
R2385 VP.n4902 VP.n4901 6.105
R2386 VP.n4891 VP.t807 6.105
R2387 VP.n5387 VP.t895 6.105
R2388 VP.n5395 VP.n5394 6.105
R2389 VP.n5398 VP.n5397 6.105
R2390 VP.n5390 VP.t88 6.105
R2391 VP.n5725 VP.t958 6.105
R2392 VP.n5736 VP.n5735 6.105
R2393 VP.n5739 VP.n5738 6.105
R2394 VP.n5728 VP.t66 6.105
R2395 VP.n6215 VP.t719 6.105
R2396 VP.n6223 VP.n6222 6.105
R2397 VP.n6226 VP.n6225 6.105
R2398 VP.n6218 VP.t1313 6.105
R2399 VP.n6569 VP.t857 6.105
R2400 VP.n6580 VP.n6579 6.105
R2401 VP.n6583 VP.n6582 6.105
R2402 VP.n6572 VP.t123 6.105
R2403 VP.n7102 VP.t1324 6.105
R2404 VP.n7110 VP.n7109 6.105
R2405 VP.n7113 VP.n7112 6.105
R2406 VP.n7105 VP.t613 6.105
R2407 VP.n7381 VP.t135 6.105
R2408 VP.n7392 VP.n7391 6.105
R2409 VP.n7395 VP.n7394 6.105
R2410 VP.n7384 VP.t735 6.105
R2411 VP.n7659 VP.t623 6.105
R2412 VP.n7976 VP.n7975 6.105
R2413 VP.n7979 VP.n7978 6.105
R2414 VP.n7982 VP.t1207 6.105
R2415 VP.n8010 VP.t749 6.105
R2416 VP.n8453 VP.t1335 6.105
R2417 VP.n139 VP.t564 6.105
R2418 VP.n274 VP.t1175 6.105
R2419 VP.n292 VP.n291 6.105
R2420 VP.n289 VP.n288 6.105
R2421 VP.n271 VP.t321 6.105
R2422 VP.n790 VP.t1152 6.105
R2423 VP.n787 VP.n786 6.105
R2424 VP.n817 VP.n816 6.105
R2425 VP.n784 VP.t446 6.105
R2426 VP.n1346 VP.t478 6.105
R2427 VP.n1370 VP.n1369 6.105
R2428 VP.n1367 VP.n1366 6.105
R2429 VP.n1343 VP.t1065 6.105
R2430 VP.n1776 VP.t457 6.105
R2431 VP.n1806 VP.n1805 6.105
R2432 VP.n1803 VP.n1802 6.105
R2433 VP.n1773 VP.t976 6.105
R2434 VP.n2663 VP.t1071 6.105
R2435 VP.n2684 VP.n2683 6.105
R2436 VP.n2687 VP.n2686 6.105
R2437 VP.n2660 VP.t357 6.105
R2438 VP.n2736 VP.t983 6.105
R2439 VP.n2766 VP.n2765 6.105
R2440 VP.n2763 VP.n2762 6.105
R2441 VP.n2733 VP.t263 6.105
R2442 VP.n3272 VP.t366 6.105
R2443 VP.n3296 VP.n3295 6.105
R2444 VP.n3293 VP.n3292 6.105
R2445 VP.n3269 VP.t949 6.105
R2446 VP.n3676 VP.t272 6.105
R2447 VP.n3706 VP.n3705 6.105
R2448 VP.n3703 VP.n3702 6.105
R2449 VP.n3673 VP.t864 6.105
R2450 VP.n4193 VP.t693 6.105
R2451 VP.n4217 VP.n4216 6.105
R2452 VP.n4214 VP.n4213 6.105
R2453 VP.n4190 VP.t1289 6.105
R2454 VP.n4585 VP.t627 6.105
R2455 VP.n4582 VP.n4581 6.105
R2456 VP.n4612 VP.n4611 6.105
R2457 VP.n4579 VP.t1212 6.105
R2458 VP.n5099 VP.t1297 6.105
R2459 VP.n5123 VP.n5122 6.105
R2460 VP.n5120 VP.n5119 6.105
R2461 VP.n5096 VP.t580 6.105
R2462 VP.n5477 VP.t27 6.105
R2463 VP.n5507 VP.n5506 6.105
R2464 VP.n5504 VP.n5503 6.105
R2465 VP.n5474 VP.t504 6.105
R2466 VP.n5963 VP.t592 6.105
R2467 VP.n5987 VP.n5986 6.105
R2468 VP.n5984 VP.n5983 6.105
R2469 VP.n5960 VP.t1177 6.105
R2470 VP.n6333 VP.t658 6.105
R2471 VP.n6363 VP.n6362 6.105
R2472 VP.n6360 VP.n6359 6.105
R2473 VP.n6330 VP.t1246 6.105
R2474 VP.n6827 VP.t1190 6.105
R2475 VP.n6851 VP.n6850 6.105
R2476 VP.n6848 VP.n6847 6.105
R2477 VP.n6824 VP.t407 6.105
R2478 VP.n7192 VP.t1254 6.105
R2479 VP.n7222 VP.n7221 6.105
R2480 VP.n7219 VP.n7218 6.105
R2481 VP.n7189 VP.t535 6.105
R2482 VP.n7666 VP.t1014 6.105
R2483 VP.n7690 VP.n7689 6.105
R2484 VP.n7687 VP.n7686 6.105
R2485 VP.n7663 VP.t306 6.105
R2486 VP.n8020 VP.t1145 6.105
R2487 VP.n8050 VP.n8049 6.105
R2488 VP.n8047 VP.n8046 6.105
R2489 VP.n8017 VP.t436 6.105
R2490 VP.n8505 VP.t319 6.105
R2491 VP.n8529 VP.n8528 6.105
R2492 VP.n8526 VP.n8525 6.105
R2493 VP.n8502 VP.t907 6.105
R2494 VP.n8866 VP.t445 6.105
R2495 VP.n8894 VP.n8893 6.105
R2496 VP.n8891 VP.n8890 6.105
R2497 VP.n8863 VP.t1032 6.105
R2498 VP.n9322 VP.t1063 6.105
R2499 VP.n9641 VP.n9640 6.105
R2500 VP.n9644 VP.n9643 6.105
R2501 VP.n9647 VP.t204 6.105
R2502 VP.n9685 VP.t1044 6.105
R2503 VP.n10100 VP.t335 6.105
R2504 VP.n2224 VP.t841 6.105
R2505 VP.n2235 VP.n2234 6.105
R2506 VP.n2238 VP.n2237 6.105
R2507 VP.n2227 VP.t99 6.105
R2508 VP.n2364 VP.t216 6.105
R2509 VP.n2375 VP.n2374 6.105
R2510 VP.n2372 VP.n2371 6.105
R2511 VP.n2367 VP.t806 6.105
R2512 VP.n3153 VP.t109 6.105
R2513 VP.n3164 VP.n3163 6.105
R2514 VP.n3167 VP.n3166 6.105
R2515 VP.n3156 VP.t708 6.105
R2516 VP.n3618 VP.t815 6.105
R2517 VP.n3626 VP.n3625 6.105
R2518 VP.n3629 VP.n3628 6.105
R2519 VP.n3621 VP.t65 6.105
R2520 VP.n4046 VP.t718 6.105
R2521 VP.n4057 VP.n4056 6.105
R2522 VP.n4060 VP.n4059 6.105
R2523 VP.n4049 VP.t1314 6.105
R2524 VP.n4497 VP.t1143 6.105
R2525 VP.n4505 VP.n4504 6.105
R2526 VP.n4508 VP.n4507 6.105
R2527 VP.n4500 VP.t433 6.105
R2528 VP.n4929 VP.t1072 6.105
R2529 VP.n4940 VP.n4939 6.105
R2530 VP.n4943 VP.n4942 6.105
R2531 VP.n4932 VP.t358 6.105
R2532 VP.n5419 VP.t443 6.105
R2533 VP.n5427 VP.n5426 6.105
R2534 VP.n5430 VP.n5429 6.105
R2535 VP.n5422 VP.t1028 6.105
R2536 VP.n5766 VP.t510 6.105
R2537 VP.n5777 VP.n5776 6.105
R2538 VP.n5780 VP.n5779 6.105
R2539 VP.n5769 VP.t950 6.105
R2540 VP.n6247 VP.t1041 6.105
R2541 VP.n6255 VP.n6254 6.105
R2542 VP.n6258 VP.n6257 6.105
R2543 VP.n6250 VP.t255 6.105
R2544 VP.n6610 VP.t1100 6.105
R2545 VP.n6621 VP.n6620 6.105
R2546 VP.n6624 VP.n6623 6.105
R2547 VP.n6613 VP.t389 6.105
R2548 VP.n7134 VP.t873 6.105
R2549 VP.n7142 VP.n7141 6.105
R2550 VP.n7145 VP.n7144 6.105
R2551 VP.n7137 VP.t150 6.105
R2552 VP.n7422 VP.t1000 6.105
R2553 VP.n7433 VP.n7432 6.105
R2554 VP.n7436 VP.n7435 6.105
R2555 VP.n7425 VP.t283 6.105
R2556 VP.n7934 VP.t163 6.105
R2557 VP.n7942 VP.n7941 6.105
R2558 VP.n7945 VP.n7944 6.105
R2559 VP.n7937 VP.t758 6.105
R2560 VP.n8238 VP.t294 6.105
R2561 VP.n8249 VP.n8248 6.105
R2562 VP.n8252 VP.n8251 6.105
R2563 VP.n8241 VP.t885 6.105
R2564 VP.n8498 VP.t771 6.105
R2565 VP.n8807 VP.n8806 6.105
R2566 VP.n8810 VP.n8809 6.105
R2567 VP.n8813 VP.t5 6.105
R2568 VP.n8844 VP.t898 6.105
R2569 VP.n9280 VP.t180 6.105
R2570 VP.n242 VP.t1007 6.105
R2571 VP.n707 VP.t331 6.105
R2572 VP.n724 VP.n723 6.105
R2573 VP.n727 VP.n726 6.105
R2574 VP.n710 VP.t772 6.105
R2575 VP.n1275 VP.t305 6.105
R2576 VP.n1286 VP.n1285 6.105
R2577 VP.n1289 VP.n1288 6.105
R2578 VP.n1278 VP.t834 6.105
R2579 VP.n1716 VP.t926 6.105
R2580 VP.n1725 VP.n1724 6.105
R2581 VP.n1728 VP.n1727 6.105
R2582 VP.n1719 VP.t210 6.105
R2583 VP.n1440 VP.t412 6.105
R2584 VP.n10094 VP.t531 6.105
R2585 VP.n10098 VP.n10097 6.105
R2586 VP.n10079 VP.t1249 6.105
R2587 VP.n10081 VP.n10080 6.105
R2588 VP.n10964 VP.n10962 4.263
R2589 VP.n9589 VP.n9587 4.263
R2590 VP.n8785 VP.n8783 4.263
R2591 VP.n7898 VP.n7896 4.263
R2592 VP.n7062 VP.n7060 4.263
R2593 VP.n6147 VP.n6145 4.263
R2594 VP.n5283 VP.n5281 4.263
R2595 VP.n4327 VP.n4325 4.263
R2596 VP.n3406 VP.n3404 4.263
R2597 VP.n2601 VP.n2599 4.263
R2598 VP.n1435 VP.n1433 4.263
R2599 VP.n337 VP.n334 4.263
R2600 VP.n10667 VP.n10666 3.857
R2601 VP.n9667 VP.n9666 3.857
R2602 VP.n9288 VP.n9287 3.857
R2603 VP.n8461 VP.n8460 3.857
R2604 VP.n7622 VP.n7621 3.857
R2605 VP.n6783 VP.n6782 3.857
R2606 VP.n5919 VP.n5918 3.857
R2607 VP.n5055 VP.n5054 3.857
R2608 VP.n4149 VP.n4148 3.857
R2609 VP.n3228 VP.n3227 3.857
R2610 VP.n2278 VP.n2277 3.857
R2611 VP.n1301 VP.n1300 3.857
R2612 VP.n10436 VP.t147 2.635
R2613 VP.n328 VP.n327 0.233
R2614 VP.n248 VP.n247 0.184
R2615 VP.n4 VP.n3 0.173
R2616 VP.n135 VP.n134 0.169
R2617 VP.n10347 VP.n10346 0.163
R2618 VP.n10326 VP.n10325 0.158
R2619 VP VP.n249 0.157
R2620 VP.n10064 VP.n10063 0.156
R2621 VP.n10994 VP.n10993 0.156
R2622 VP.n10020 VP.n10019 0.156
R2623 VP.n10935 VP.n10934 0.156
R2624 VP.n8426 VP.n8425 0.156
R2625 VP.n9226 VP.n9225 0.156
R2626 VP.n9983 VP.n9982 0.156
R2627 VP.n10884 VP.n10883 0.156
R2628 VP.n6748 VP.n6747 0.156
R2629 VP.n7560 VP.n7559 0.156
R2630 VP.n8377 VP.n8376 0.156
R2631 VP.n9176 VP.n9175 0.156
R2632 VP.n9935 VP.n9934 0.156
R2633 VP.n10833 VP.n10832 0.156
R2634 VP.n5020 VP.n5019 0.156
R2635 VP.n5857 VP.n5856 0.156
R2636 VP.n6699 VP.n6698 0.156
R2637 VP.n7511 VP.n7510 0.156
R2638 VP.n8328 VP.n8327 0.156
R2639 VP.n9126 VP.n9125 0.156
R2640 VP.n9887 VP.n9886 0.156
R2641 VP.n10782 VP.n10781 0.156
R2642 VP.n9820 VP.n9817 0.156
R2643 VP.n9056 VP.n9053 0.156
R2644 VP.n8259 VP.n8256 0.156
R2645 VP.n7443 VP.n7440 0.156
R2646 VP.n6631 VP.n6628 0.156
R2647 VP.n5787 VP.n5784 0.156
R2648 VP.n4950 VP.n4947 0.156
R2649 VP.n4067 VP.n4064 0.156
R2650 VP.n3174 VP.n3171 0.156
R2651 VP.n886 VP.n885 0.156
R2652 VP.n936 VP.n935 0.156
R2653 VP.n1873 VP.n1872 0.156
R2654 VP.n986 VP.n985 0.156
R2655 VP.n1925 VP.n1924 0.156
R2656 VP.n2854 VP.n2853 0.156
R2657 VP.n1036 VP.n1035 0.156
R2658 VP.n1977 VP.n1976 0.156
R2659 VP.n2906 VP.n2905 0.156
R2660 VP.n3799 VP.n3798 0.156
R2661 VP.n1086 VP.n1085 0.156
R2662 VP.n2029 VP.n2028 0.156
R2663 VP.n2958 VP.n2957 0.156
R2664 VP.n3851 VP.n3850 0.156
R2665 VP.n4734 VP.n4733 0.156
R2666 VP.n1136 VP.n1135 0.156
R2667 VP.n2081 VP.n2080 0.156
R2668 VP.n3010 VP.n3009 0.156
R2669 VP.n3903 VP.n3902 0.156
R2670 VP.n4786 VP.n4785 0.156
R2671 VP.n5623 VP.n5622 0.156
R2672 VP.n1174 VP.n1173 0.156
R2673 VP.n2122 VP.n2121 0.156
R2674 VP.n3051 VP.n3050 0.156
R2675 VP.n3944 VP.n3943 0.156
R2676 VP.n4827 VP.n4826 0.156
R2677 VP.n5664 VP.n5663 0.156
R2678 VP.n6508 VP.n6507 0.156
R2679 VP.n1214 VP.n1213 0.156
R2680 VP.n2163 VP.n2162 0.156
R2681 VP.n3092 VP.n3091 0.156
R2682 VP.n3985 VP.n3984 0.156
R2683 VP.n4868 VP.n4867 0.156
R2684 VP.n5705 VP.n5704 0.156
R2685 VP.n6549 VP.n6548 0.156
R2686 VP.n7361 VP.n7360 0.156
R2687 VP.n1255 VP.n1254 0.156
R2688 VP.n2204 VP.n2203 0.156
R2689 VP.n3133 VP.n3132 0.156
R2690 VP.n4026 VP.n4025 0.156
R2691 VP.n4909 VP.n4908 0.156
R2692 VP.n5746 VP.n5745 0.156
R2693 VP.n6590 VP.n6589 0.156
R2694 VP.n7402 VP.n7401 0.156
R2695 VP.n8218 VP.n8217 0.156
R2696 VP.n801 VP.n800 0.156
R2697 VP.n1787 VP.n1786 0.156
R2698 VP.n2747 VP.n2746 0.156
R2699 VP.n3687 VP.n3686 0.156
R2700 VP.n4596 VP.n4595 0.156
R2701 VP.n5488 VP.n5487 0.156
R2702 VP.n6344 VP.n6343 0.156
R2703 VP.n7203 VP.n7202 0.156
R2704 VP.n8031 VP.n8030 0.156
R2705 VP.n8875 VP.n8874 0.156
R2706 VP.n884 VP.n883 0.152
R2707 VP.n934 VP.n933 0.152
R2708 VP.n1871 VP.n1870 0.152
R2709 VP.n1975 VP.n1974 0.152
R2710 VP.n3797 VP.n3796 0.152
R2711 VP.n1084 VP.n1083 0.152
R2712 VP.n2027 VP.n2026 0.152
R2713 VP.n1134 VP.n1133 0.152
R2714 VP.n3901 VP.n3900 0.152
R2715 VP.n4784 VP.n4783 0.152
R2716 VP.n2120 VP.n2119 0.152
R2717 VP.n3942 VP.n3941 0.152
R2718 VP.n4825 VP.n4824 0.152
R2719 VP.n5662 VP.n5661 0.152
R2720 VP.n2161 VP.n2160 0.152
R2721 VP.n7359 VP.n7358 0.152
R2722 VP.n2202 VP.n2201 0.152
R2723 VP.n4907 VP.n4906 0.152
R2724 VP.n5744 VP.n5743 0.152
R2725 VP.n1785 VP.n1784 0.152
R2726 VP.n3685 VP.n3684 0.152
R2727 VP.n8029 VP.n8028 0.152
R2728 VP.n8873 VP.n8872 0.152
R2729 VP.n10350 VP.n10344 0.144
R2730 VP.n10109 VP.n10108 0.138
R2731 VP.n10119 VP.n10116 0.138
R2732 VP.n10664 VP.n10663 0.136
R2733 VP.n845 VP.n844 0.134
R2734 VP.n1745 VP.n1743 0.128
R2735 VP.n2706 VP.n2704 0.128
R2736 VP.n3646 VP.n3644 0.128
R2737 VP.n4552 VP.n4550 0.128
R2738 VP.n5447 VP.n5445 0.128
R2739 VP.n6303 VP.n6301 0.128
R2740 VP.n7162 VP.n7160 0.128
R2741 VP.n7990 VP.n7988 0.128
R2742 VP.n336 VP.n335 0.123
R2743 VP.n10333 VP.n10330 0.12
R2744 VP.n11047 VP.n11034 0.12
R2745 VP.n11058 VP.n1320 0.12
R2746 VP.n11057 VP.n2296 0.12
R2747 VP.n11056 VP.n3246 0.12
R2748 VP.n11055 VP.n4167 0.12
R2749 VP.n11054 VP.n5073 0.12
R2750 VP.n11053 VP.n5937 0.12
R2751 VP.n11052 VP.n6801 0.12
R2752 VP.n11051 VP.n7640 0.12
R2753 VP.n11050 VP.n8479 0.12
R2754 VP.n11048 VP.n10113 0.12
R2755 VP.n11049 VP.n9306 0.119
R2756 VP.n8765 VP.n8764 0.117
R2757 VP.n7042 VP.n7041 0.117
R2758 VP.n5263 VP.n5262 0.117
R2759 VP.n1406 VP.n1405 0.117
R2760 VP.n3384 VP.n3383 0.117
R2761 VP.n1316 VP.n1311 0.117
R2762 VP.n10057 VP.n10055 0.116
R2763 VP.n10987 VP.n10985 0.116
R2764 VP.n10037 VP.n10035 0.116
R2765 VP.n10928 VP.n10926 0.116
R2766 VP.n8443 VP.n8441 0.116
R2767 VP.n9241 VP.n9239 0.116
R2768 VP.n9997 VP.n9995 0.116
R2769 VP.n10877 VP.n10875 0.116
R2770 VP.n6765 VP.n6763 0.116
R2771 VP.n7575 VP.n7573 0.116
R2772 VP.n8392 VP.n8390 0.116
R2773 VP.n9191 VP.n9189 0.116
R2774 VP.n9949 VP.n9947 0.116
R2775 VP.n10826 VP.n10824 0.116
R2776 VP.n5037 VP.n5035 0.116
R2777 VP.n5872 VP.n5870 0.116
R2778 VP.n6714 VP.n6712 0.116
R2779 VP.n7526 VP.n7524 0.116
R2780 VP.n8343 VP.n8341 0.116
R2781 VP.n9141 VP.n9139 0.116
R2782 VP.n9901 VP.n9899 0.116
R2783 VP.n10775 VP.n10773 0.116
R2784 VP.n9824 VP.n9823 0.116
R2785 VP.n9060 VP.n9059 0.116
R2786 VP.n8263 VP.n8262 0.116
R2787 VP.n7447 VP.n7446 0.116
R2788 VP.n6635 VP.n6634 0.116
R2789 VP.n5791 VP.n5790 0.116
R2790 VP.n4954 VP.n4953 0.116
R2791 VP.n4071 VP.n4070 0.116
R2792 VP.n3178 VP.n3177 0.116
R2793 VP.n10700 VP.n10698 0.116
R2794 VP.n263 VP.n261 0.116
R2795 VP.n1740 VP.n1739 0.116
R2796 VP.n365 VP.n363 0.116
R2797 VP.n902 VP.n900 0.116
R2798 VP.n1336 VP.n1334 0.116
R2799 VP.n2701 VP.n2700 0.116
R2800 VP.n412 VP.n410 0.116
R2801 VP.n952 VP.n950 0.116
R2802 VP.n1464 VP.n1462 0.116
R2803 VP.n1889 VP.n1887 0.116
R2804 VP.n2312 VP.n2310 0.116
R2805 VP.n3641 VP.n3640 0.116
R2806 VP.n459 VP.n457 0.116
R2807 VP.n1002 VP.n1000 0.116
R2808 VP.n1502 VP.n1500 0.116
R2809 VP.n1941 VP.n1939 0.116
R2810 VP.n2564 VP.n2562 0.116
R2811 VP.n2870 VP.n2868 0.116
R2812 VP.n3262 VP.n3260 0.116
R2813 VP.n4547 VP.n4546 0.116
R2814 VP.n506 VP.n504 0.116
R2815 VP.n1052 VP.n1050 0.116
R2816 VP.n1540 VP.n1538 0.116
R2817 VP.n1993 VP.n1991 0.116
R2818 VP.n2526 VP.n2524 0.116
R2819 VP.n2922 VP.n2920 0.116
R2820 VP.n3442 VP.n3440 0.116
R2821 VP.n3815 VP.n3813 0.116
R2822 VP.n4183 VP.n4181 0.116
R2823 VP.n5442 VP.n5441 0.116
R2824 VP.n553 VP.n551 0.116
R2825 VP.n1102 VP.n1100 0.116
R2826 VP.n1578 VP.n1576 0.116
R2827 VP.n2045 VP.n2043 0.116
R2828 VP.n2488 VP.n2486 0.116
R2829 VP.n2974 VP.n2972 0.116
R2830 VP.n3480 VP.n3478 0.116
R2831 VP.n3867 VP.n3865 0.116
R2832 VP.n4359 VP.n4357 0.116
R2833 VP.n4750 VP.n4748 0.116
R2834 VP.n5089 VP.n5087 0.116
R2835 VP.n6298 VP.n6297 0.116
R2836 VP.n600 VP.n598 0.116
R2837 VP.n1152 VP.n1150 0.116
R2838 VP.n1616 VP.n1614 0.116
R2839 VP.n2097 VP.n2095 0.116
R2840 VP.n2456 VP.n2454 0.116
R2841 VP.n3026 VP.n3024 0.116
R2842 VP.n3518 VP.n3516 0.116
R2843 VP.n3919 VP.n3917 0.116
R2844 VP.n4397 VP.n4395 0.116
R2845 VP.n4802 VP.n4800 0.116
R2846 VP.n5319 VP.n5317 0.116
R2847 VP.n5639 VP.n5637 0.116
R2848 VP.n5953 VP.n5951 0.116
R2849 VP.n7157 VP.n7156 0.116
R2850 VP.n640 VP.n638 0.116
R2851 VP.n1190 VP.n1188 0.116
R2852 VP.n1648 VP.n1646 0.116
R2853 VP.n2138 VP.n2136 0.116
R2854 VP.n2424 VP.n2422 0.116
R2855 VP.n3067 VP.n3065 0.116
R2856 VP.n3550 VP.n3548 0.116
R2857 VP.n3960 VP.n3958 0.116
R2858 VP.n4429 VP.n4427 0.116
R2859 VP.n4843 VP.n4841 0.116
R2860 VP.n5351 VP.n5349 0.116
R2861 VP.n5680 VP.n5678 0.116
R2862 VP.n6179 VP.n6177 0.116
R2863 VP.n6524 VP.n6522 0.116
R2864 VP.n6817 VP.n6815 0.116
R2865 VP.n7985 VP.n7984 0.116
R2866 VP.n670 VP.n668 0.116
R2867 VP.n1230 VP.n1228 0.116
R2868 VP.n1680 VP.n1678 0.116
R2869 VP.n2179 VP.n2177 0.116
R2870 VP.n2392 VP.n2390 0.116
R2871 VP.n3108 VP.n3106 0.116
R2872 VP.n3582 VP.n3580 0.116
R2873 VP.n4001 VP.n3999 0.116
R2874 VP.n4461 VP.n4459 0.116
R2875 VP.n4884 VP.n4882 0.116
R2876 VP.n5383 VP.n5381 0.116
R2877 VP.n5721 VP.n5719 0.116
R2878 VP.n6211 VP.n6209 0.116
R2879 VP.n6565 VP.n6563 0.116
R2880 VP.n7098 VP.n7096 0.116
R2881 VP.n7377 VP.n7375 0.116
R2882 VP.n7656 VP.n7654 0.116
R2883 VP.n9651 VP.n9650 0.116
R2884 VP.n702 VP.n700 0.116
R2885 VP.n1271 VP.n1269 0.116
R2886 VP.n1712 VP.n1710 0.116
R2887 VP.n2220 VP.n2218 0.116
R2888 VP.n2360 VP.n2358 0.116
R2889 VP.n3149 VP.n3147 0.116
R2890 VP.n3614 VP.n3612 0.116
R2891 VP.n4042 VP.n4040 0.116
R2892 VP.n4493 VP.n4491 0.116
R2893 VP.n4925 VP.n4923 0.116
R2894 VP.n5415 VP.n5413 0.116
R2895 VP.n5762 VP.n5760 0.116
R2896 VP.n6243 VP.n6241 0.116
R2897 VP.n6606 VP.n6604 0.116
R2898 VP.n7130 VP.n7128 0.116
R2899 VP.n7418 VP.n7416 0.116
R2900 VP.n7930 VP.n7928 0.116
R2901 VP.n8234 VP.n8232 0.116
R2902 VP.n8495 VP.n8493 0.116
R2903 VP.n8817 VP.n8816 0.116
R2904 VP.n278 VP.n276 0.116
R2905 VP.n794 VP.n792 0.116
R2906 VP.n1350 VP.n1348 0.116
R2907 VP.n1780 VP.n1778 0.116
R2908 VP.n2667 VP.n2665 0.116
R2909 VP.n2740 VP.n2738 0.116
R2910 VP.n3276 VP.n3274 0.116
R2911 VP.n3680 VP.n3678 0.116
R2912 VP.n4197 VP.n4195 0.116
R2913 VP.n4589 VP.n4587 0.116
R2914 VP.n5103 VP.n5101 0.116
R2915 VP.n5481 VP.n5479 0.116
R2916 VP.n5967 VP.n5965 0.116
R2917 VP.n6337 VP.n6335 0.116
R2918 VP.n6831 VP.n6829 0.116
R2919 VP.n7196 VP.n7194 0.116
R2920 VP.n7670 VP.n7668 0.116
R2921 VP.n8024 VP.n8022 0.116
R2922 VP.n8509 VP.n8507 0.116
R2923 VP.n8870 VP.n8868 0.116
R2924 VP.n11023 VP.n11021 0.116
R2925 VP.n128 VP.n127 0.114
R2926 VP.n120 VP.n119 0.114
R2927 VP.n115 VP.n114 0.114
R2928 VP.n107 VP.n106 0.114
R2929 VP.n102 VP.n101 0.114
R2930 VP.n96 VP.n95 0.114
R2931 VP.n89 VP.n88 0.114
R2932 VP.n81 VP.n80 0.114
R2933 VP.n76 VP.n75 0.114
R2934 VP.n70 VP.n69 0.114
R2935 VP.n63 VP.n62 0.114
R2936 VP.n55 VP.n54 0.114
R2937 VP.n50 VP.n49 0.114
R2938 VP.n44 VP.n43 0.114
R2939 VP.n34 VP.n33 0.114
R2940 VP.n24 VP.n23 0.114
R2941 VP.n17 VP.n16 0.114
R2942 VP.n2833 VP.n2825 0.113
R2943 VP.n259 VP.n258 0.11
R2944 VP.n361 VP.n360 0.11
R2945 VP.n408 VP.n407 0.11
R2946 VP.n455 VP.n454 0.11
R2947 VP.n502 VP.n501 0.11
R2948 VP.n549 VP.n548 0.11
R2949 VP.n596 VP.n595 0.11
R2950 VP.n636 VP.n635 0.11
R2951 VP.n666 VP.n665 0.11
R2952 VP.n698 VP.n697 0.11
R2953 VP.n10639 VP.n10638 0.11
R2954 VP.n1295 VP.n1294 0.108
R2955 VP.n9 VP.n8 0.106
R2956 VP.n11002 VP.n11001 0.106
R2957 VP.n10943 VP.n10942 0.106
R2958 VP.n8741 VP.n8740 0.106
R2959 VP.n9548 VP.n9547 0.106
R2960 VP.n10892 VP.n10891 0.106
R2961 VP.n7018 VP.n7017 0.106
R2962 VP.n7856 VP.n7855 0.106
R2963 VP.n8693 VP.n8692 0.106
R2964 VP.n9497 VP.n9496 0.106
R2965 VP.n10841 VP.n10840 0.106
R2966 VP.n5239 VP.n5238 0.106
R2967 VP.n6105 VP.n6104 0.106
R2968 VP.n6969 VP.n6968 0.106
R2969 VP.n7807 VP.n7806 0.106
R2970 VP.n8645 VP.n8644 0.106
R2971 VP.n9446 VP.n9445 0.106
R2972 VP.n10790 VP.n10789 0.106
R2973 VP.n10725 VP.n10722 0.106
R2974 VP.n9380 VP.n9377 0.106
R2975 VP.n8585 VP.n8582 0.106
R2976 VP.n7746 VP.n7743 0.106
R2977 VP.n6907 VP.n6904 0.106
R2978 VP.n6043 VP.n6040 0.106
R2979 VP.n5179 VP.n5176 0.106
R2980 VP.n4273 VP.n4270 0.106
R2981 VP.n3352 VP.n3349 0.106
R2982 VP.n897 VP.n896 0.106
R2983 VP.n1331 VP.n1330 0.106
R2984 VP.n947 VP.n946 0.106
R2985 VP.n1459 VP.n1458 0.106
R2986 VP.n1884 VP.n1883 0.106
R2987 VP.n2307 VP.n2306 0.106
R2988 VP.n997 VP.n996 0.106
R2989 VP.n1497 VP.n1496 0.106
R2990 VP.n1936 VP.n1935 0.106
R2991 VP.n2559 VP.n2558 0.106
R2992 VP.n2865 VP.n2864 0.106
R2993 VP.n3257 VP.n3256 0.106
R2994 VP.n1047 VP.n1046 0.106
R2995 VP.n1535 VP.n1534 0.106
R2996 VP.n1988 VP.n1987 0.106
R2997 VP.n2521 VP.n2520 0.106
R2998 VP.n2917 VP.n2916 0.106
R2999 VP.n3437 VP.n3436 0.106
R3000 VP.n3810 VP.n3809 0.106
R3001 VP.n4178 VP.n4177 0.106
R3002 VP.n1097 VP.n1096 0.106
R3003 VP.n1573 VP.n1572 0.106
R3004 VP.n2040 VP.n2039 0.106
R3005 VP.n2483 VP.n2482 0.106
R3006 VP.n2969 VP.n2968 0.106
R3007 VP.n3475 VP.n3474 0.106
R3008 VP.n3862 VP.n3861 0.106
R3009 VP.n4354 VP.n4353 0.106
R3010 VP.n4745 VP.n4744 0.106
R3011 VP.n5084 VP.n5083 0.106
R3012 VP.n1147 VP.n1146 0.106
R3013 VP.n1611 VP.n1610 0.106
R3014 VP.n2092 VP.n2091 0.106
R3015 VP.n2451 VP.n2450 0.106
R3016 VP.n3021 VP.n3020 0.106
R3017 VP.n3513 VP.n3512 0.106
R3018 VP.n3914 VP.n3913 0.106
R3019 VP.n4392 VP.n4391 0.106
R3020 VP.n4797 VP.n4796 0.106
R3021 VP.n5314 VP.n5313 0.106
R3022 VP.n5634 VP.n5633 0.106
R3023 VP.n5948 VP.n5947 0.106
R3024 VP.n1185 VP.n1184 0.106
R3025 VP.n1643 VP.n1642 0.106
R3026 VP.n2133 VP.n2132 0.106
R3027 VP.n2419 VP.n2418 0.106
R3028 VP.n3062 VP.n3061 0.106
R3029 VP.n3545 VP.n3544 0.106
R3030 VP.n3955 VP.n3954 0.106
R3031 VP.n4424 VP.n4423 0.106
R3032 VP.n4838 VP.n4837 0.106
R3033 VP.n5346 VP.n5345 0.106
R3034 VP.n5675 VP.n5674 0.106
R3035 VP.n6174 VP.n6173 0.106
R3036 VP.n6519 VP.n6518 0.106
R3037 VP.n6812 VP.n6811 0.106
R3038 VP.n1225 VP.n1224 0.106
R3039 VP.n1675 VP.n1674 0.106
R3040 VP.n2174 VP.n2173 0.106
R3041 VP.n2387 VP.n2386 0.106
R3042 VP.n3103 VP.n3102 0.106
R3043 VP.n3577 VP.n3576 0.106
R3044 VP.n3996 VP.n3995 0.106
R3045 VP.n4456 VP.n4455 0.106
R3046 VP.n4879 VP.n4878 0.106
R3047 VP.n5378 VP.n5377 0.106
R3048 VP.n5716 VP.n5715 0.106
R3049 VP.n6206 VP.n6205 0.106
R3050 VP.n6560 VP.n6559 0.106
R3051 VP.n7093 VP.n7092 0.106
R3052 VP.n7372 VP.n7371 0.106
R3053 VP.n7651 VP.n7650 0.106
R3054 VP.n1266 VP.n1265 0.106
R3055 VP.n1707 VP.n1706 0.106
R3056 VP.n2215 VP.n2214 0.106
R3057 VP.n2355 VP.n2354 0.106
R3058 VP.n3144 VP.n3143 0.106
R3059 VP.n3609 VP.n3608 0.106
R3060 VP.n4037 VP.n4036 0.106
R3061 VP.n4488 VP.n4487 0.106
R3062 VP.n4920 VP.n4919 0.106
R3063 VP.n5410 VP.n5409 0.106
R3064 VP.n5757 VP.n5756 0.106
R3065 VP.n6238 VP.n6237 0.106
R3066 VP.n6601 VP.n6600 0.106
R3067 VP.n7125 VP.n7124 0.106
R3068 VP.n7413 VP.n7412 0.106
R3069 VP.n7925 VP.n7924 0.106
R3070 VP.n8229 VP.n8228 0.106
R3071 VP.n8490 VP.n8489 0.106
R3072 VP.n812 VP.n811 0.106
R3073 VP.n1362 VP.n1361 0.106
R3074 VP.n1798 VP.n1797 0.106
R3075 VP.n2679 VP.n2678 0.106
R3076 VP.n2758 VP.n2757 0.106
R3077 VP.n3288 VP.n3287 0.106
R3078 VP.n3698 VP.n3697 0.106
R3079 VP.n4209 VP.n4208 0.106
R3080 VP.n4607 VP.n4606 0.106
R3081 VP.n5115 VP.n5114 0.106
R3082 VP.n5499 VP.n5498 0.106
R3083 VP.n5979 VP.n5978 0.106
R3084 VP.n6355 VP.n6354 0.106
R3085 VP.n6843 VP.n6842 0.106
R3086 VP.n7214 VP.n7213 0.106
R3087 VP.n7682 VP.n7681 0.106
R3088 VP.n8042 VP.n8041 0.106
R3089 VP.n8521 VP.n8520 0.106
R3090 VP.n8886 VP.n8885 0.106
R3091 VP.n747 VP.n740 0.104
R3092 VP.n390 VP.n383 0.104
R3093 VP.n437 VP.n430 0.104
R3094 VP.n484 VP.n477 0.104
R3095 VP.n531 VP.n524 0.104
R3096 VP.n578 VP.n571 0.104
R3097 VP.n618 VP.n611 0.104
R3098 VP.n720 VP.n713 0.104
R3099 VP.n9316 VP.n9315 0.104
R3100 VP.n10133 VP.n10132 0.101
R3101 VP.n1317 VP.n1310 0.101
R3102 VP.n770 VP.n769 0.101
R3103 VP.n2293 VP.n2287 0.101
R3104 VP.n1759 VP.n1758 0.101
R3105 VP.n3243 VP.n3237 0.101
R3106 VP.n2720 VP.n2719 0.101
R3107 VP.n4164 VP.n4158 0.101
R3108 VP.n3660 VP.n3659 0.101
R3109 VP.n5070 VP.n5064 0.101
R3110 VP.n4566 VP.n4565 0.101
R3111 VP.n5934 VP.n5928 0.101
R3112 VP.n5461 VP.n5460 0.101
R3113 VP.n6798 VP.n6792 0.101
R3114 VP.n6317 VP.n6316 0.101
R3115 VP.n7637 VP.n7631 0.101
R3116 VP.n7176 VP.n7175 0.101
R3117 VP.n8476 VP.n8470 0.101
R3118 VP.n8004 VP.n8003 0.101
R3119 VP.n9682 VP.n9676 0.101
R3120 VP.n8838 VP.n8837 0.101
R3121 VP.n9303 VP.n9297 0.101
R3122 VP.n10659 VP.n10658 0.101
R3123 VP.n746 VP.n742 0.098
R3124 VP.n389 VP.n385 0.098
R3125 VP.n436 VP.n432 0.098
R3126 VP.n483 VP.n479 0.098
R3127 VP.n530 VP.n526 0.098
R3128 VP.n577 VP.n573 0.098
R3129 VP.n617 VP.n613 0.098
R3130 VP.n719 VP.n715 0.098
R3131 VP.n10030 VP.n10027 0.097
R3132 VP.n8436 VP.n8433 0.097
R3133 VP.n6758 VP.n6755 0.097
R3134 VP.n5030 VP.n5027 0.097
R3135 VP.n3182 VP.n3179 0.097
R3136 VP.n10322 VP.n10318 0.092
R3137 VP.n10304 VP.n10300 0.092
R3138 VP.n10276 VP.n10272 0.092
R3139 VP.n10248 VP.n10244 0.092
R3140 VP.n10220 VP.n10216 0.092
R3141 VP.n10202 VP.n10201 0.092
R3142 VP.n125 VP.n122 0.091
R3143 VP.n118 VP.n117 0.091
R3144 VP.n112 VP.n109 0.091
R3145 VP.n105 VP.n104 0.091
R3146 VP.n99 VP.n98 0.091
R3147 VP.n94 VP.n93 0.091
R3148 VP.n86 VP.n83 0.091
R3149 VP.n79 VP.n78 0.091
R3150 VP.n73 VP.n72 0.091
R3151 VP.n68 VP.n67 0.091
R3152 VP.n60 VP.n57 0.091
R3153 VP.n53 VP.n52 0.091
R3154 VP.n47 VP.n46 0.091
R3155 VP.n42 VP.n41 0.091
R3156 VP.n32 VP.n31 0.091
R3157 VP.n22 VP.n21 0.091
R3158 VP.n14 VP.n11 0.091
R3159 VP.n133 VP.n132 0.091
R3160 VP.n246 VP.n245 0.091
R3161 VP.n2 VP.n1 0.091
R3162 VP.n751 VP.n750 0.09
R3163 VP.n1200 VP.n1199 0.09
R3164 VP.n681 VP.n680 0.09
R3165 VP.n781 VP.n780 0.089
R3166 VP.n10115 VP.n10114 0.088
R3167 VP.n10601 VP.n10596 0.084
R3168 VP.n10566 VP.n10561 0.084
R3169 VP.n10531 VP.n10526 0.084
R3170 VP.n10496 VP.n10491 0.084
R3171 VP.n10598 VP.n10597 0.084
R3172 VP.n10563 VP.n10562 0.084
R3173 VP.n10528 VP.n10527 0.084
R3174 VP.n10493 VP.n10492 0.084
R3175 VP.n1315 VP.n1314 0.084
R3176 VP.n765 VP.n764 0.084
R3177 VP.n2291 VP.n2290 0.084
R3178 VP.n892 VP.n891 0.084
R3179 VP.n1754 VP.n1753 0.084
R3180 VP.n3241 VP.n3240 0.084
R3181 VP.n942 VP.n941 0.084
R3182 VP.n1879 VP.n1878 0.084
R3183 VP.n2715 VP.n2714 0.084
R3184 VP.n4162 VP.n4161 0.084
R3185 VP.n992 VP.n991 0.084
R3186 VP.n1931 VP.n1930 0.084
R3187 VP.n2860 VP.n2859 0.084
R3188 VP.n3655 VP.n3654 0.084
R3189 VP.n5068 VP.n5067 0.084
R3190 VP.n1042 VP.n1041 0.084
R3191 VP.n1983 VP.n1982 0.084
R3192 VP.n2912 VP.n2911 0.084
R3193 VP.n3805 VP.n3804 0.084
R3194 VP.n4561 VP.n4560 0.084
R3195 VP.n5932 VP.n5931 0.084
R3196 VP.n1092 VP.n1091 0.084
R3197 VP.n2035 VP.n2034 0.084
R3198 VP.n2964 VP.n2963 0.084
R3199 VP.n3857 VP.n3856 0.084
R3200 VP.n4740 VP.n4739 0.084
R3201 VP.n5456 VP.n5455 0.084
R3202 VP.n6796 VP.n6795 0.084
R3203 VP.n1142 VP.n1141 0.084
R3204 VP.n2087 VP.n2086 0.084
R3205 VP.n3016 VP.n3015 0.084
R3206 VP.n3909 VP.n3908 0.084
R3207 VP.n4792 VP.n4791 0.084
R3208 VP.n5629 VP.n5628 0.084
R3209 VP.n6312 VP.n6311 0.084
R3210 VP.n7635 VP.n7634 0.084
R3211 VP.n1180 VP.n1179 0.084
R3212 VP.n2128 VP.n2127 0.084
R3213 VP.n3057 VP.n3056 0.084
R3214 VP.n3950 VP.n3949 0.084
R3215 VP.n4833 VP.n4832 0.084
R3216 VP.n5670 VP.n5669 0.084
R3217 VP.n6514 VP.n6513 0.084
R3218 VP.n7171 VP.n7170 0.084
R3219 VP.n8474 VP.n8473 0.084
R3220 VP.n1220 VP.n1219 0.084
R3221 VP.n2169 VP.n2168 0.084
R3222 VP.n3098 VP.n3097 0.084
R3223 VP.n3991 VP.n3990 0.084
R3224 VP.n4874 VP.n4873 0.084
R3225 VP.n5711 VP.n5710 0.084
R3226 VP.n6555 VP.n6554 0.084
R3227 VP.n7367 VP.n7366 0.084
R3228 VP.n7999 VP.n7998 0.084
R3229 VP.n9680 VP.n9679 0.084
R3230 VP.n1261 VP.n1260 0.084
R3231 VP.n2210 VP.n2209 0.084
R3232 VP.n3139 VP.n3138 0.084
R3233 VP.n4032 VP.n4031 0.084
R3234 VP.n4915 VP.n4914 0.084
R3235 VP.n5752 VP.n5751 0.084
R3236 VP.n6596 VP.n6595 0.084
R3237 VP.n7408 VP.n7407 0.084
R3238 VP.n8224 VP.n8223 0.084
R3239 VP.n8833 VP.n8832 0.084
R3240 VP.n9301 VP.n9300 0.084
R3241 VP.n807 VP.n806 0.084
R3242 VP.n1793 VP.n1792 0.084
R3243 VP.n2753 VP.n2752 0.084
R3244 VP.n3693 VP.n3692 0.084
R3245 VP.n4602 VP.n4601 0.084
R3246 VP.n5494 VP.n5493 0.084
R3247 VP.n6350 VP.n6349 0.084
R3248 VP.n7209 VP.n7208 0.084
R3249 VP.n8037 VP.n8036 0.084
R3250 VP.n8881 VP.n8880 0.084
R3251 VP.n10654 VP.n10653 0.084
R3252 VP.n7 VP.n6 0.084
R3253 VP.t8 VP.n10334 0.083
R3254 VP.n10673 VP.n10672 0.082
R3255 VP.n9673 VP.n9672 0.082
R3256 VP.n9294 VP.n9293 0.082
R3257 VP.n8467 VP.n8466 0.082
R3258 VP.n7628 VP.n7627 0.082
R3259 VP.n6789 VP.n6788 0.082
R3260 VP.n5925 VP.n5924 0.082
R3261 VP.n5061 VP.n5060 0.082
R3262 VP.n4155 VP.n4154 0.082
R3263 VP.n3234 VP.n3233 0.082
R3264 VP.n2284 VP.n2283 0.082
R3265 VP.n1307 VP.n1306 0.082
R3266 VP.n10181 VP.n10180 0.08
R3267 VP.n10633 VP.n10632 0.079
R3268 VP.n10697 VP.n10695 0.077
R3269 VP.n750 VP.n749 0.077
R3270 VP.n127 VP.n126 0.077
R3271 VP.n114 VP.n113 0.077
R3272 VP.n101 VP.n100 0.077
R3273 VP.n88 VP.n87 0.077
R3274 VP.n75 VP.n74 0.077
R3275 VP.n62 VP.n61 0.077
R3276 VP.n49 VP.n48 0.077
R3277 VP.n16 VP.n15 0.077
R3278 VP.n1318 VP.n1307 0.075
R3279 VP.n2294 VP.n2284 0.075
R3280 VP.n3244 VP.n3234 0.075
R3281 VP.n4165 VP.n4155 0.075
R3282 VP.n5071 VP.n5061 0.075
R3283 VP.n5935 VP.n5925 0.075
R3284 VP.n6799 VP.n6789 0.075
R3285 VP.n7638 VP.n7628 0.075
R3286 VP.n8477 VP.n8467 0.075
R3287 VP.n9683 VP.n9673 0.075
R3288 VP.n9304 VP.n9294 0.075
R3289 VP.n10674 VP.n10673 0.075
R3290 VP.n9022 VP.n9020 0.075
R3291 VP.n7327 VP.n7325 0.075
R3292 VP.n5589 VP.n5587 0.075
R3293 VP.n1839 VP.n1838 0.075
R3294 VP.n3766 VP.n3765 0.075
R3295 VP.n10288 VP.n10287 0.075
R3296 VP.n10260 VP.n10259 0.075
R3297 VP.n10232 VP.n10231 0.075
R3298 VP.n10453 VP.n10452 0.075
R3299 VP.n9834 VP.n9833 0.075
R3300 VP.n9071 VP.n9070 0.075
R3301 VP.n8274 VP.n8273 0.075
R3302 VP.n7458 VP.n7457 0.075
R3303 VP.n6646 VP.n6645 0.075
R3304 VP.n5802 VP.n5801 0.075
R3305 VP.n4965 VP.n4964 0.075
R3306 VP.n4082 VP.n4081 0.075
R3307 VP.n2327 VP.n2326 0.075
R3308 VP.n9627 VP.n9626 0.074
R3309 VP.n7962 VP.n7961 0.074
R3310 VP.n9238 VP.n9237 0.074
R3311 VP.n9994 VP.n9993 0.074
R3312 VP.n6275 VP.n6274 0.074
R3313 VP.n7572 VP.n7571 0.074
R3314 VP.n8389 VP.n8388 0.074
R3315 VP.n9188 VP.n9187 0.074
R3316 VP.n9946 VP.n9945 0.074
R3317 VP.n4524 VP.n4523 0.074
R3318 VP.n5869 VP.n5868 0.074
R3319 VP.n6711 VP.n6710 0.074
R3320 VP.n7523 VP.n7522 0.074
R3321 VP.n8340 VP.n8339 0.074
R3322 VP.n9138 VP.n9137 0.074
R3323 VP.n9898 VP.n9897 0.074
R3324 VP.n10177 VP.n10176 0.074
R3325 VP.n3191 VP.n3190 0.072
R3326 VP.n10958 VP.n10957 0.072
R3327 VP.n9583 VP.n9582 0.072
R3328 VP.n8779 VP.n8778 0.072
R3329 VP.n7892 VP.n7891 0.072
R3330 VP.n7056 VP.n7055 0.072
R3331 VP.n6141 VP.n6140 0.072
R3332 VP.n5277 VP.n5276 0.072
R3333 VP.n4321 VP.n4320 0.072
R3334 VP.n3400 VP.n3399 0.072
R3335 VP.n2595 VP.n2594 0.072
R3336 VP.n1429 VP.n1428 0.072
R3337 VP.n330 VP.n329 0.072
R3338 VP.n10034 VP.n10033 0.072
R3339 VP.n8440 VP.n8439 0.072
R3340 VP.n6762 VP.n6761 0.072
R3341 VP.n5034 VP.n5033 0.072
R3342 VP.n10310 VP.n10309 0.069
R3343 VP.n10294 VP.n10293 0.069
R3344 VP.n10282 VP.n10281 0.069
R3345 VP.n10266 VP.n10265 0.069
R3346 VP.n10254 VP.n10253 0.069
R3347 VP.n10238 VP.n10237 0.069
R3348 VP.n10226 VP.n10225 0.069
R3349 VP.n10210 VP.n10209 0.069
R3350 VP.n10190 VP.n10189 0.069
R3351 VP.n10356 VP.n10355 0.069
R3352 VP.n10184 VP.n10183 0.069
R3353 VP.n9 VP.n7 0.069
R3354 VP.n10624 VP.n10623 0.068
R3355 VP.n10586 VP.n10585 0.068
R3356 VP.n10551 VP.n10550 0.068
R3357 VP.n10516 VP.n10515 0.068
R3358 VP.n10481 VP.n10480 0.068
R3359 VP.n10441 VP.n10440 0.068
R3360 VP.n10684 VP.n10683 0.068
R3361 VP.n10990 VP.n10989 0.067
R3362 VP.n10318 VP.n10317 0.067
R3363 VP.n10318 VP.n10315 0.067
R3364 VP.n9621 VP.n9620 0.067
R3365 VP.n10300 VP.n10299 0.067
R3366 VP.n10300 VP.n10298 0.067
R3367 VP.n10287 VP.n10286 0.067
R3368 VP.n10287 VP.n10285 0.067
R3369 VP.n7956 VP.n7955 0.067
R3370 VP.n10272 VP.n10271 0.067
R3371 VP.n10272 VP.n10270 0.067
R3372 VP.n10259 VP.n10258 0.067
R3373 VP.n10259 VP.n10257 0.067
R3374 VP.n6269 VP.n6268 0.067
R3375 VP.n10244 VP.n10243 0.067
R3376 VP.n10244 VP.n10242 0.067
R3377 VP.n10231 VP.n10230 0.067
R3378 VP.n10231 VP.n10229 0.067
R3379 VP.n4518 VP.n4517 0.067
R3380 VP.n10216 VP.n10215 0.067
R3381 VP.n10216 VP.n10214 0.067
R3382 VP.n10176 VP.n10171 0.067
R3383 VP.n2318 VP.n2317 0.067
R3384 VP.n1307 VP.n1295 0.067
R3385 VP.n1307 VP.n1296 0.067
R3386 VP.n2284 VP.n2272 0.067
R3387 VP.n2284 VP.n2273 0.067
R3388 VP.n3234 VP.n3222 0.067
R3389 VP.n3234 VP.n3223 0.067
R3390 VP.n4155 VP.n4143 0.067
R3391 VP.n4155 VP.n4144 0.067
R3392 VP.n5061 VP.n5049 0.067
R3393 VP.n5061 VP.n5050 0.067
R3394 VP.n5925 VP.n5913 0.067
R3395 VP.n5925 VP.n5914 0.067
R3396 VP.n6789 VP.n6777 0.067
R3397 VP.n6789 VP.n6778 0.067
R3398 VP.n7628 VP.n7616 0.067
R3399 VP.n7628 VP.n7617 0.067
R3400 VP.n8467 VP.n8455 0.067
R3401 VP.n8467 VP.n8456 0.067
R3402 VP.n9673 VP.n9661 0.067
R3403 VP.n9294 VP.n9283 0.067
R3404 VP.n9294 VP.n9282 0.067
R3405 VP.n9673 VP.n9662 0.067
R3406 VP.n10673 VP.n10661 0.067
R3407 VP.n10673 VP.n10660 0.067
R3408 VP.n10201 VP.n10200 0.067
R3409 VP.n10201 VP.n10198 0.067
R3410 VP.n10176 VP.n10175 0.067
R3411 VP.n2243 VP.n2242 0.066
R3412 VP.n8178 VP.n8177 0.066
R3413 VP.n6468 VP.n6467 0.066
R3414 VP.n4694 VP.n4693 0.066
R3415 VP.n128 VP.n125 0.066
R3416 VP.n120 VP.n118 0.066
R3417 VP.n381 VP.n376 0.066
R3418 VP.n115 VP.n112 0.066
R3419 VP.n107 VP.n105 0.066
R3420 VP.n428 VP.n423 0.066
R3421 VP.n102 VP.n99 0.066
R3422 VP.n96 VP.n94 0.066
R3423 VP.n475 VP.n470 0.066
R3424 VP.n89 VP.n86 0.066
R3425 VP.n81 VP.n79 0.066
R3426 VP.n522 VP.n517 0.066
R3427 VP.n76 VP.n73 0.066
R3428 VP.n70 VP.n68 0.066
R3429 VP.n569 VP.n564 0.066
R3430 VP.n63 VP.n60 0.066
R3431 VP.n55 VP.n53 0.066
R3432 VP.n50 VP.n47 0.066
R3433 VP.n44 VP.n42 0.066
R3434 VP.n34 VP.n32 0.066
R3435 VP.n24 VP.n22 0.066
R3436 VP.n17 VP.n14 0.066
R3437 VP.n135 VP.n133 0.066
R3438 VP.n149 VP.n148 0.066
R3439 VP.n248 VP.n246 0.066
R3440 VP.n4 VP.n2 0.066
R3441 VP.n9308 VP.n9307 0.065
R3442 VP.n199 VP.n198 0.064
R3443 VP.n772 VP.n761 0.063
R3444 VP.n1761 VP.n1750 0.063
R3445 VP.n2722 VP.n2711 0.063
R3446 VP.n3662 VP.n3651 0.063
R3447 VP.n4568 VP.n4557 0.063
R3448 VP.n5463 VP.n5452 0.063
R3449 VP.n6319 VP.n6308 0.063
R3450 VP.n7178 VP.n7167 0.063
R3451 VP.n8006 VP.n7995 0.063
R3452 VP.n8840 VP.n8829 0.063
R3453 VP.n10111 VP.n10105 0.063
R3454 VP.n10638 VP.n10637 0.062
R3455 VP.n10596 VP.n10595 0.062
R3456 VP.n10561 VP.n10560 0.062
R3457 VP.n10526 VP.n10525 0.062
R3458 VP.n10491 VP.n10490 0.062
R3459 VP.n199 VP.n158 0.062
R3460 VP.n758 VP.n757 0.062
R3461 VP.n10068 VP.n10067 0.061
R3462 VP.t8 VP.n10181 0.061
R3463 VP.n2609 VP.n2607 0.06
R3464 VP.n921 VP.n920 0.059
R3465 VP.n971 VP.n970 0.059
R3466 VP.n1021 VP.n1020 0.059
R3467 VP.n1071 VP.n1070 0.059
R3468 VP.n1121 VP.n1120 0.059
R3469 VP.n10033 VP.n10032 0.058
R3470 VP.n8439 VP.n8438 0.058
R3471 VP.n6761 VP.n6760 0.058
R3472 VP.n5033 VP.n5032 0.058
R3473 VP.n3190 VP.n3189 0.058
R3474 VP.n308 VP.n307 0.058
R3475 VP.n1905 VP.n1901 0.058
R3476 VP.n1957 VP.n1953 0.058
R3477 VP.n3831 VP.n3827 0.058
R3478 VP.n2009 VP.n2005 0.058
R3479 VP.n1068 VP.n1064 0.058
R3480 VP.n2061 VP.n2057 0.058
R3481 VP.n9598 VP.n9593 0.057
R3482 VP.n8791 VP.n8789 0.057
R3483 VP.n7068 VP.n7066 0.057
R3484 VP.n5289 VP.n5287 0.057
R3485 VP.n3412 VP.n3410 0.057
R3486 VP.n10438 VP.n10437 0.056
R3487 VP.n10677 VP.n10676 0.056
R3488 VP.n244 VP.n243 0.056
R3489 VP.n10099 VP.n10098 0.055
R3490 VP.n10176 VP.n10174 0.055
R3491 VP.n10352 VP.n10342 0.055
R3492 VP.n10135 VP.n10134 0.055
R3493 VP.n10972 VP.n10971 0.055
R3494 VP.n9607 VP.n9606 0.055
R3495 VP.n8801 VP.n8800 0.055
R3496 VP.n7910 VP.n7909 0.055
R3497 VP.n7078 VP.n7077 0.055
R3498 VP.n6159 VP.n6158 0.055
R3499 VP.n5299 VP.n5298 0.055
R3500 VP.n4339 VP.n4338 0.055
R3501 VP.n3422 VP.n3421 0.055
R3502 VP.n347 VP.n346 0.055
R3503 VP.n1444 VP.n1443 0.055
R3504 VP.n2610 VP.n2590 0.054
R3505 VP.n10650 VP.n10649 0.054
R3506 VP.n1292 VP.n1291 0.054
R3507 VP.n2271 VP.n2270 0.054
R3508 VP.n3221 VP.n3220 0.054
R3509 VP.n4142 VP.n4141 0.054
R3510 VP.n5048 VP.n5047 0.054
R3511 VP.n5912 VP.n5911 0.054
R3512 VP.n6776 VP.n6775 0.054
R3513 VP.n7615 VP.n7614 0.054
R3514 VP.n8454 VP.n8453 0.054
R3515 VP.n10101 VP.n10100 0.054
R3516 VP.n9281 VP.n9280 0.054
R3517 VP.n8769 VP.n8767 0.054
R3518 VP.n7046 VP.n7044 0.054
R3519 VP.n5267 VP.n5265 0.054
R3520 VP.n10632 VP.n10631 0.054
R3521 VP.n8765 VP.n8763 0.054
R3522 VP.n7042 VP.n7040 0.054
R3523 VP.n5263 VP.n5261 0.054
R3524 VP.n752 VP.n738 0.054
R3525 VP.n122 VP.n121 0.054
R3526 VP.n117 VP.n116 0.054
R3527 VP.n109 VP.n108 0.054
R3528 VP.n104 VP.n103 0.054
R3529 VP.n98 VP.n97 0.054
R3530 VP.n93 VP.n92 0.054
R3531 VP.n83 VP.n82 0.054
R3532 VP.n78 VP.n77 0.054
R3533 VP.n72 VP.n71 0.054
R3534 VP.n67 VP.n66 0.054
R3535 VP.n57 VP.n56 0.054
R3536 VP.n52 VP.n51 0.054
R3537 VP.n46 VP.n45 0.054
R3538 VP.n41 VP.n40 0.054
R3539 VP.n31 VP.n30 0.054
R3540 VP.n21 VP.n20 0.054
R3541 VP.n11 VP.n10 0.054
R3542 VP.n6 VP.n5 0.054
R3543 VP.n9696 VP.n9695 0.054
R3544 VP.n9691 VP.n9690 0.054
R3545 VP.n9328 VP.n9327 0.054
R3546 VP.n8901 VP.n8900 0.054
R3547 VP.n8535 VP.n8534 0.054
R3548 VP.n8057 VP.n8056 0.054
R3549 VP.n7696 VP.n7695 0.054
R3550 VP.n7229 VP.n7228 0.054
R3551 VP.n6857 VP.n6856 0.054
R3552 VP.n6370 VP.n6369 0.054
R3553 VP.n5993 VP.n5992 0.054
R3554 VP.n5514 VP.n5513 0.054
R3555 VP.n5129 VP.n5128 0.054
R3556 VP.n4619 VP.n4618 0.054
R3557 VP.n4223 VP.n4222 0.054
R3558 VP.n3713 VP.n3712 0.054
R3559 VP.n3302 VP.n3301 0.054
R3560 VP.n2773 VP.n2772 0.054
R3561 VP.n2637 VP.n2636 0.054
R3562 VP.n1813 VP.n1812 0.054
R3563 VP.n1376 VP.n1375 0.054
R3564 VP.n827 VP.n826 0.054
R3565 VP.n10417 VP.n10416 0.054
R3566 VP.n2269 VP.n2268 0.054
R3567 VP.n2341 VP.n2340 0.054
R3568 VP.n3219 VP.n3218 0.054
R3569 VP.n3367 VP.n3366 0.054
R3570 VP.n4111 VP.n4110 0.054
R3571 VP.n4288 VP.n4287 0.054
R3572 VP.n4994 VP.n4993 0.054
R3573 VP.n5194 VP.n5193 0.054
R3574 VP.n5831 VP.n5830 0.054
R3575 VP.n6059 VP.n6058 0.054
R3576 VP.n6674 VP.n6673 0.054
R3577 VP.n6923 VP.n6922 0.054
R3578 VP.n7486 VP.n7485 0.054
R3579 VP.n7761 VP.n7760 0.054
R3580 VP.n8303 VP.n8302 0.054
R3581 VP.n8600 VP.n8599 0.054
R3582 VP.n9100 VP.n9099 0.054
R3583 VP.n9397 VP.n9396 0.054
R3584 VP.n9862 VP.n9861 0.054
R3585 VP.n10742 VP.n10741 0.054
R3586 VP.n10470 VP.n10469 0.054
R3587 VP.n10432 VP.n10431 0.054
R3588 VP.n10077 VP.n10076 0.054
R3589 VP.n11011 VP.n11010 0.054
R3590 VP.n10648 VP.n10647 0.054
R3591 VP.n9279 VP.n9278 0.054
R3592 VP.n9639 VP.n9638 0.054
R3593 VP.n10046 VP.n10045 0.054
R3594 VP.n10949 VP.n10948 0.054
R3595 VP.n10610 VP.n10609 0.054
R3596 VP.n8773 VP.n8772 0.054
R3597 VP.n9046 VP.n9045 0.054
R3598 VP.n9577 VP.n9576 0.054
R3599 VP.n9810 VP.n9809 0.054
R3600 VP.n10914 VP.n10913 0.054
R3601 VP.n10406 VP.n10405 0.054
R3602 VP.n8208 VP.n8207 0.054
R3603 VP.n7613 VP.n7612 0.054
R3604 VP.n7974 VP.n7973 0.054
R3605 VP.n8452 VP.n8451 0.054
R3606 VP.n8747 VP.n8746 0.054
R3607 VP.n9250 VP.n9249 0.054
R3608 VP.n9554 VP.n9553 0.054
R3609 VP.n10006 VP.n10005 0.054
R3610 VP.n10898 VP.n10897 0.054
R3611 VP.n10575 VP.n10574 0.054
R3612 VP.n7050 VP.n7049 0.054
R3613 VP.n7351 VP.n7350 0.054
R3614 VP.n7884 VP.n7883 0.054
R3615 VP.n8172 VP.n8171 0.054
R3616 VP.n8720 VP.n8719 0.054
R3617 VP.n9016 VP.n9015 0.054
R3618 VP.n9525 VP.n9524 0.054
R3619 VP.n9788 VP.n9787 0.054
R3620 VP.n10863 VP.n10862 0.054
R3621 VP.n10389 VP.n10388 0.054
R3622 VP.n6498 VP.n6497 0.054
R3623 VP.n5910 VP.n5909 0.054
R3624 VP.n6287 VP.n6286 0.054
R3625 VP.n6774 VP.n6773 0.054
R3626 VP.n7024 VP.n7023 0.054
R3627 VP.n7584 VP.n7583 0.054
R3628 VP.n7862 VP.n7861 0.054
R3629 VP.n8401 VP.n8400 0.054
R3630 VP.n8699 VP.n8698 0.054
R3631 VP.n9200 VP.n9199 0.054
R3632 VP.n9503 VP.n9502 0.054
R3633 VP.n9958 VP.n9957 0.054
R3634 VP.n10847 VP.n10846 0.054
R3635 VP.n10540 VP.n10539 0.054
R3636 VP.n5271 VP.n5270 0.054
R3637 VP.n5613 VP.n5612 0.054
R3638 VP.n6133 VP.n6132 0.054
R3639 VP.n6462 VP.n6461 0.054
R3640 VP.n6996 VP.n6995 0.054
R3641 VP.n7321 VP.n7320 0.054
R3642 VP.n7834 VP.n7833 0.054
R3643 VP.n8149 VP.n8148 0.054
R3644 VP.n8672 VP.n8671 0.054
R3645 VP.n8993 VP.n8992 0.054
R3646 VP.n9474 VP.n9473 0.054
R3647 VP.n9766 VP.n9765 0.054
R3648 VP.n10812 VP.n10811 0.054
R3649 VP.n10372 VP.n10371 0.054
R3650 VP.n4724 VP.n4723 0.054
R3651 VP.n4140 VP.n4139 0.054
R3652 VP.n4536 VP.n4535 0.054
R3653 VP.n5046 VP.n5045 0.054
R3654 VP.n5245 VP.n5244 0.054
R3655 VP.n5881 VP.n5880 0.054
R3656 VP.n6111 VP.n6110 0.054
R3657 VP.n6723 VP.n6722 0.054
R3658 VP.n6975 VP.n6974 0.054
R3659 VP.n7535 VP.n7534 0.054
R3660 VP.n7813 VP.n7812 0.054
R3661 VP.n8352 VP.n8351 0.054
R3662 VP.n8651 VP.n8650 0.054
R3663 VP.n9150 VP.n9149 0.054
R3664 VP.n9452 VP.n9451 0.054
R3665 VP.n9910 VP.n9909 0.054
R3666 VP.n10796 VP.n10795 0.054
R3667 VP.n10505 VP.n10504 0.054
R3668 VP.n876 VP.n875 0.054
R3669 VP.n1417 VP.n1416 0.054
R3670 VP.n1863 VP.n1862 0.054
R3671 VP.n2632 VP.n2631 0.054
R3672 VP.n2816 VP.n2815 0.054
R3673 VP.n3340 VP.n3339 0.054
R3674 VP.n3756 VP.n3755 0.054
R3675 VP.n4261 VP.n4260 0.054
R3676 VP.n4662 VP.n4661 0.054
R3677 VP.n5167 VP.n5166 0.054
R3678 VP.n5557 VP.n5556 0.054
R3679 VP.n6031 VP.n6030 0.054
R3680 VP.n6413 VP.n6412 0.054
R3681 VP.n6895 VP.n6894 0.054
R3682 VP.n7272 VP.n7271 0.054
R3683 VP.n7734 VP.n7733 0.054
R3684 VP.n8100 VP.n8099 0.054
R3685 VP.n8573 VP.n8572 0.054
R3686 VP.n8944 VP.n8943 0.054
R3687 VP.n9368 VP.n9367 0.054
R3688 VP.n9744 VP.n9743 0.054
R3689 VP.n10713 VP.n10712 0.054
R3690 VP.n10147 VP.n10146 0.054
R3691 VP.n11017 VP.n11016 0.054
R3692 VP.n9722 VP.n9721 0.054
R3693 VP.n9346 VP.n9345 0.054
R3694 VP.n8921 VP.n8920 0.054
R3695 VP.n8552 VP.n8551 0.054
R3696 VP.n8077 VP.n8076 0.054
R3697 VP.n7713 VP.n7712 0.054
R3698 VP.n7249 VP.n7248 0.054
R3699 VP.n6874 VP.n6873 0.054
R3700 VP.n6390 VP.n6389 0.054
R3701 VP.n6010 VP.n6009 0.054
R3702 VP.n5534 VP.n5533 0.054
R3703 VP.n5146 VP.n5145 0.054
R3704 VP.n4639 VP.n4638 0.054
R3705 VP.n4240 VP.n4239 0.054
R3706 VP.n3733 VP.n3732 0.054
R3707 VP.n3319 VP.n3318 0.054
R3708 VP.n2793 VP.n2792 0.054
R3709 VP.n2657 VP.n2656 0.054
R3710 VP.n1833 VP.n1832 0.054
R3711 VP.n1393 VP.n1392 0.054
R3712 VP.n821 VP.n820 0.054
R3713 VP.n316 VP.n315 0.054
R3714 VP.n734 VP.n733 0.054
R3715 VP.n398 VP.n397 0.054
R3716 VP.n930 VP.n929 0.054
R3717 VP.n1735 VP.n1734 0.054
R3718 VP.n445 VP.n444 0.054
R3719 VP.n980 VP.n979 0.054
R3720 VP.n1486 VP.n1485 0.054
R3721 VP.n1919 VP.n1918 0.054
R3722 VP.n2696 VP.n2695 0.054
R3723 VP.n492 VP.n491 0.054
R3724 VP.n1030 VP.n1029 0.054
R3725 VP.n1524 VP.n1523 0.054
R3726 VP.n1971 VP.n1970 0.054
R3727 VP.n2583 VP.n2582 0.054
R3728 VP.n2900 VP.n2899 0.054
R3729 VP.n3636 VP.n3635 0.054
R3730 VP.n539 VP.n538 0.054
R3731 VP.n1080 VP.n1079 0.054
R3732 VP.n1562 VP.n1561 0.054
R3733 VP.n2023 VP.n2022 0.054
R3734 VP.n2545 VP.n2544 0.054
R3735 VP.n2952 VP.n2951 0.054
R3736 VP.n3464 VP.n3463 0.054
R3737 VP.n3845 VP.n3844 0.054
R3738 VP.n4542 VP.n4541 0.054
R3739 VP.n586 VP.n585 0.054
R3740 VP.n1130 VP.n1129 0.054
R3741 VP.n1600 VP.n1599 0.054
R3742 VP.n2075 VP.n2074 0.054
R3743 VP.n2507 VP.n2506 0.054
R3744 VP.n3004 VP.n3003 0.054
R3745 VP.n3502 VP.n3501 0.054
R3746 VP.n3897 VP.n3896 0.054
R3747 VP.n4381 VP.n4380 0.054
R3748 VP.n4780 VP.n4779 0.054
R3749 VP.n5437 VP.n5436 0.054
R3750 VP.n626 VP.n625 0.054
R3751 VP.n1168 VP.n1167 0.054
R3752 VP.n1632 VP.n1631 0.054
R3753 VP.n2116 VP.n2115 0.054
R3754 VP.n2469 VP.n2468 0.054
R3755 VP.n3045 VP.n3044 0.054
R3756 VP.n3534 VP.n3533 0.054
R3757 VP.n3938 VP.n3937 0.054
R3758 VP.n4413 VP.n4412 0.054
R3759 VP.n4821 VP.n4820 0.054
R3760 VP.n5335 VP.n5334 0.054
R3761 VP.n5658 VP.n5657 0.054
R3762 VP.n6293 VP.n6292 0.054
R3763 VP.n656 VP.n655 0.054
R3764 VP.n1208 VP.n1207 0.054
R3765 VP.n1664 VP.n1663 0.054
R3766 VP.n2157 VP.n2156 0.054
R3767 VP.n2437 VP.n2436 0.054
R3768 VP.n3086 VP.n3085 0.054
R3769 VP.n3566 VP.n3565 0.054
R3770 VP.n3979 VP.n3978 0.054
R3771 VP.n4445 VP.n4444 0.054
R3772 VP.n4862 VP.n4861 0.054
R3773 VP.n5367 VP.n5366 0.054
R3774 VP.n5699 VP.n5698 0.054
R3775 VP.n6195 VP.n6194 0.054
R3776 VP.n6543 VP.n6542 0.054
R3777 VP.n7152 VP.n7151 0.054
R3778 VP.n688 VP.n687 0.054
R3779 VP.n1249 VP.n1248 0.054
R3780 VP.n1696 VP.n1695 0.054
R3781 VP.n2198 VP.n2197 0.054
R3782 VP.n2405 VP.n2404 0.054
R3783 VP.n3127 VP.n3126 0.054
R3784 VP.n3598 VP.n3597 0.054
R3785 VP.n4020 VP.n4019 0.054
R3786 VP.n4477 VP.n4476 0.054
R3787 VP.n4903 VP.n4902 0.054
R3788 VP.n5399 VP.n5398 0.054
R3789 VP.n5740 VP.n5739 0.054
R3790 VP.n6227 VP.n6226 0.054
R3791 VP.n6584 VP.n6583 0.054
R3792 VP.n7114 VP.n7113 0.054
R3793 VP.n7396 VP.n7395 0.054
R3794 VP.n7980 VP.n7979 0.054
R3795 VP.n290 VP.n289 0.054
R3796 VP.n818 VP.n817 0.054
R3797 VP.n1368 VP.n1367 0.054
R3798 VP.n1804 VP.n1803 0.054
R3799 VP.n2688 VP.n2687 0.054
R3800 VP.n2764 VP.n2763 0.054
R3801 VP.n3294 VP.n3293 0.054
R3802 VP.n3704 VP.n3703 0.054
R3803 VP.n4215 VP.n4214 0.054
R3804 VP.n4613 VP.n4612 0.054
R3805 VP.n5121 VP.n5120 0.054
R3806 VP.n5505 VP.n5504 0.054
R3807 VP.n5985 VP.n5984 0.054
R3808 VP.n6361 VP.n6360 0.054
R3809 VP.n6849 VP.n6848 0.054
R3810 VP.n7220 VP.n7219 0.054
R3811 VP.n7688 VP.n7687 0.054
R3812 VP.n8048 VP.n8047 0.054
R3813 VP.n8527 VP.n8526 0.054
R3814 VP.n8892 VP.n8891 0.054
R3815 VP.n9645 VP.n9644 0.054
R3816 VP.n2239 VP.n2238 0.054
R3817 VP.n2373 VP.n2372 0.054
R3818 VP.n3168 VP.n3167 0.054
R3819 VP.n3630 VP.n3629 0.054
R3820 VP.n4061 VP.n4060 0.054
R3821 VP.n4509 VP.n4508 0.054
R3822 VP.n4944 VP.n4943 0.054
R3823 VP.n5431 VP.n5430 0.054
R3824 VP.n5781 VP.n5780 0.054
R3825 VP.n6259 VP.n6258 0.054
R3826 VP.n6625 VP.n6624 0.054
R3827 VP.n7146 VP.n7145 0.054
R3828 VP.n7437 VP.n7436 0.054
R3829 VP.n7946 VP.n7945 0.054
R3830 VP.n8253 VP.n8252 0.054
R3831 VP.n8811 VP.n8810 0.054
R3832 VP.n728 VP.n727 0.054
R3833 VP.n1290 VP.n1289 0.054
R3834 VP.n1729 VP.n1728 0.054
R3835 VP.n10967 VP.n10966 0.053
R3836 VP.n7901 VP.n7900 0.053
R3837 VP.n6150 VP.n6149 0.053
R3838 VP.n4330 VP.n4329 0.053
R3839 VP.n2604 VP.n2603 0.053
R3840 VP.n3409 VP.n3408 0.053
R3841 VP.n5286 VP.n5285 0.053
R3842 VP.n7065 VP.n7064 0.053
R3843 VP.n8788 VP.n8787 0.053
R3844 VP.n9592 VP.n9591 0.053
R3845 VP.n10591 VP.n10590 0.053
R3846 VP.n10556 VP.n10555 0.053
R3847 VP.n10521 VP.n10520 0.053
R3848 VP.n10486 VP.n10485 0.053
R3849 VP.n10096 VP.n10085 0.053
R3850 VP.n10969 VP.n10968 0.052
R3851 VP.n1438 VP.n1437 0.052
R3852 VP.n340 VP.n339 0.052
R3853 VP.n10016 VP.n10015 0.052
R3854 VP.n8422 VP.n8421 0.052
R3855 VP.n9222 VP.n9221 0.052
R3856 VP.n9979 VP.n9978 0.052
R3857 VP.n6744 VP.n6743 0.052
R3858 VP.n7556 VP.n7555 0.052
R3859 VP.n8373 VP.n8372 0.052
R3860 VP.n9172 VP.n9171 0.052
R3861 VP.n9931 VP.n9930 0.052
R3862 VP.n5016 VP.n5015 0.052
R3863 VP.n5853 VP.n5852 0.052
R3864 VP.n6695 VP.n6694 0.052
R3865 VP.n7507 VP.n7506 0.052
R3866 VP.n8324 VP.n8323 0.052
R3867 VP.n9122 VP.n9121 0.052
R3868 VP.n9883 VP.n9882 0.052
R3869 VP.n9819 VP.n9818 0.052
R3870 VP.n9055 VP.n9054 0.052
R3871 VP.n8258 VP.n8257 0.052
R3872 VP.n7442 VP.n7441 0.052
R3873 VP.n6630 VP.n6629 0.052
R3874 VP.n5786 VP.n5785 0.052
R3875 VP.n4949 VP.n4948 0.052
R3876 VP.n4066 VP.n4065 0.052
R3877 VP.n3173 VP.n3172 0.052
R3878 VP.n251 VP.n250 0.052
R3879 VP.n353 VP.n352 0.052
R3880 VP.n400 VP.n399 0.052
R3881 VP.n447 VP.n446 0.052
R3882 VP.n494 VP.n493 0.052
R3883 VP.n541 VP.n540 0.052
R3884 VP.n588 VP.n587 0.052
R3885 VP.n628 VP.n627 0.052
R3886 VP.n658 VP.n657 0.052
R3887 VP.n9654 VP.n9653 0.052
R3888 VP.n690 VP.n689 0.052
R3889 VP.n8820 VP.n8819 0.052
R3890 VP.n11026 VP.n11025 0.052
R3891 VP.n831 VP.n830 0.052
R3892 VP.n1439 VP.n1438 0.051
R3893 VP.n10629 VP.n10628 0.051
R3894 VP.t8 VP.n10310 0.051
R3895 VP.t8 VP.n10308 0.051
R3896 VP.t8 VP.n10294 0.051
R3897 VP.t8 VP.n10292 0.051
R3898 VP.t8 VP.n10282 0.051
R3899 VP.t8 VP.n10280 0.051
R3900 VP.t8 VP.n10266 0.051
R3901 VP.t8 VP.n10264 0.051
R3902 VP.t8 VP.n10254 0.051
R3903 VP.t8 VP.n10252 0.051
R3904 VP.t8 VP.n10238 0.051
R3905 VP.t8 VP.n10236 0.051
R3906 VP.t8 VP.n10226 0.051
R3907 VP.t8 VP.n10224 0.051
R3908 VP.t8 VP.n10210 0.051
R3909 VP.t8 VP.n10208 0.051
R3910 VP.t8 VP.n10184 0.051
R3911 VP.t8 VP.n10186 0.051
R3912 VP.t8 VP.n10190 0.051
R3913 VP.t8 VP.n10188 0.051
R3914 VP.t8 VP.n10356 0.051
R3915 VP.t8 VP.n10358 0.051
R3916 VP.n341 VP.n340 0.051
R3917 VP.n260 VP.n259 0.05
R3918 VP.n362 VP.n361 0.05
R3919 VP.n409 VP.n408 0.05
R3920 VP.n456 VP.n455 0.05
R3921 VP.n503 VP.n502 0.05
R3922 VP.n550 VP.n549 0.05
R3923 VP.n597 VP.n596 0.05
R3924 VP.n637 VP.n636 0.05
R3925 VP.n667 VP.n666 0.05
R3926 VP.n699 VP.n698 0.05
R3927 VP.n2840 VP.n2839 0.05
R3928 VP.n3390 VP.n3389 0.05
R3929 VP.n3785 VP.n3784 0.05
R3930 VP.n4309 VP.n4308 0.05
R3931 VP.n4684 VP.n4683 0.05
R3932 VP.n5214 VP.n5213 0.05
R3933 VP.n5579 VP.n5578 0.05
R3934 VP.n6079 VP.n6078 0.05
R3935 VP.n6435 VP.n6434 0.05
R3936 VP.n6943 VP.n6942 0.05
R3937 VP.n7294 VP.n7293 0.05
R3938 VP.n7781 VP.n7780 0.05
R3939 VP.n8122 VP.n8121 0.05
R3940 VP.n8620 VP.n8619 0.05
R3941 VP.n8966 VP.n8965 0.05
R3942 VP.n9419 VP.n9418 0.05
R3943 VP.n10757 VP.n10756 0.05
R3944 VP.n10163 VP.n10162 0.05
R3945 VP.n10060 VP.n10059 0.049
R3946 VP.n10932 VP.n10931 0.049
R3947 VP.n9031 VP.n9023 0.049
R3948 VP.n8194 VP.n8186 0.049
R3949 VP.n10881 VP.n10880 0.049
R3950 VP.n7336 VP.n7328 0.049
R3951 VP.n6484 VP.n6476 0.049
R3952 VP.n10830 VP.n10829 0.049
R3953 VP.n5598 VP.n5590 0.049
R3954 VP.n4710 VP.n4702 0.049
R3955 VP.n10779 VP.n10778 0.049
R3956 VP.n862 VP.n851 0.049
R3957 VP.n1848 VP.n1840 0.049
R3958 VP.n884 VP.n881 0.049
R3959 VP.n1322 VP.n1321 0.049
R3960 VP.n934 VP.n931 0.049
R3961 VP.n1450 VP.n1449 0.049
R3962 VP.n1871 VP.n1868 0.049
R3963 VP.n2298 VP.n2297 0.049
R3964 VP.n982 VP.n981 0.049
R3965 VP.n1488 VP.n1487 0.049
R3966 VP.n1921 VP.n1920 0.049
R3967 VP.n2550 VP.n2549 0.049
R3968 VP.n2850 VP.n2849 0.049
R3969 VP.n3248 VP.n3247 0.049
R3970 VP.n1032 VP.n1031 0.049
R3971 VP.n1526 VP.n1525 0.049
R3972 VP.n1975 VP.n1972 0.049
R3973 VP.n2512 VP.n2511 0.049
R3974 VP.n2902 VP.n2901 0.049
R3975 VP.n3428 VP.n3427 0.049
R3976 VP.n3797 VP.n3794 0.049
R3977 VP.n4169 VP.n4168 0.049
R3978 VP.n1084 VP.n1081 0.049
R3979 VP.n1564 VP.n1563 0.049
R3980 VP.n2027 VP.n2024 0.049
R3981 VP.n2474 VP.n2473 0.049
R3982 VP.n2954 VP.n2953 0.049
R3983 VP.n3466 VP.n3465 0.049
R3984 VP.n3847 VP.n3846 0.049
R3985 VP.n4345 VP.n4344 0.049
R3986 VP.n4730 VP.n4729 0.049
R3987 VP.n5075 VP.n5074 0.049
R3988 VP.n1134 VP.n1131 0.049
R3989 VP.n1602 VP.n1601 0.049
R3990 VP.n2077 VP.n2076 0.049
R3991 VP.n2442 VP.n2441 0.049
R3992 VP.n3006 VP.n3005 0.049
R3993 VP.n3504 VP.n3503 0.049
R3994 VP.n3901 VP.n3898 0.049
R3995 VP.n4383 VP.n4382 0.049
R3996 VP.n4784 VP.n4781 0.049
R3997 VP.n5305 VP.n5304 0.049
R3998 VP.n5619 VP.n5618 0.049
R3999 VP.n5939 VP.n5938 0.049
R4000 VP.n1170 VP.n1169 0.049
R4001 VP.n1634 VP.n1633 0.049
R4002 VP.n2120 VP.n2117 0.049
R4003 VP.n2410 VP.n2409 0.049
R4004 VP.n3047 VP.n3046 0.049
R4005 VP.n3536 VP.n3535 0.049
R4006 VP.n3942 VP.n3939 0.049
R4007 VP.n4415 VP.n4414 0.049
R4008 VP.n4825 VP.n4822 0.049
R4009 VP.n5337 VP.n5336 0.049
R4010 VP.n5662 VP.n5659 0.049
R4011 VP.n6165 VP.n6164 0.049
R4012 VP.n6504 VP.n6503 0.049
R4013 VP.n6803 VP.n6802 0.049
R4014 VP.n1210 VP.n1209 0.049
R4015 VP.n1666 VP.n1665 0.049
R4016 VP.n2161 VP.n2158 0.049
R4017 VP.n2378 VP.n2377 0.049
R4018 VP.n3088 VP.n3087 0.049
R4019 VP.n3568 VP.n3567 0.049
R4020 VP.n3981 VP.n3980 0.049
R4021 VP.n4447 VP.n4446 0.049
R4022 VP.n4864 VP.n4863 0.049
R4023 VP.n5369 VP.n5368 0.049
R4024 VP.n5701 VP.n5700 0.049
R4025 VP.n6197 VP.n6196 0.049
R4026 VP.n6545 VP.n6544 0.049
R4027 VP.n7084 VP.n7083 0.049
R4028 VP.n7359 VP.n7356 0.049
R4029 VP.n7642 VP.n7641 0.049
R4030 VP.n1251 VP.n1250 0.049
R4031 VP.n1698 VP.n1697 0.049
R4032 VP.n2202 VP.n2199 0.049
R4033 VP.n2346 VP.n2345 0.049
R4034 VP.n3129 VP.n3128 0.049
R4035 VP.n3600 VP.n3599 0.049
R4036 VP.n4022 VP.n4021 0.049
R4037 VP.n4479 VP.n4478 0.049
R4038 VP.n4907 VP.n4904 0.049
R4039 VP.n5401 VP.n5400 0.049
R4040 VP.n5744 VP.n5741 0.049
R4041 VP.n6229 VP.n6228 0.049
R4042 VP.n6586 VP.n6585 0.049
R4043 VP.n7116 VP.n7115 0.049
R4044 VP.n7398 VP.n7397 0.049
R4045 VP.n7916 VP.n7915 0.049
R4046 VP.n8214 VP.n8213 0.049
R4047 VP.n8481 VP.n8480 0.049
R4048 VP.n281 VP.n280 0.049
R4049 VP.n797 VP.n796 0.049
R4050 VP.n1353 VP.n1352 0.049
R4051 VP.n1785 VP.n1782 0.049
R4052 VP.n2670 VP.n2669 0.049
R4053 VP.n2743 VP.n2742 0.049
R4054 VP.n3279 VP.n3278 0.049
R4055 VP.n3685 VP.n3682 0.049
R4056 VP.n4200 VP.n4199 0.049
R4057 VP.n4592 VP.n4591 0.049
R4058 VP.n5106 VP.n5105 0.049
R4059 VP.n5484 VP.n5483 0.049
R4060 VP.n5970 VP.n5969 0.049
R4061 VP.n6340 VP.n6339 0.049
R4062 VP.n6834 VP.n6833 0.049
R4063 VP.n7199 VP.n7198 0.049
R4064 VP.n7673 VP.n7672 0.049
R4065 VP.n8029 VP.n8026 0.049
R4066 VP.n8512 VP.n8511 0.049
R4067 VP.n10418 VP.n10410 0.049
R4068 VP.n3775 VP.n3767 0.049
R4069 VP.n9793 VP.n9792 0.048
R4070 VP.n8154 VP.n8153 0.048
R4071 VP.n8998 VP.n8997 0.048
R4072 VP.n9771 VP.n9770 0.048
R4073 VP.n6444 VP.n6443 0.048
R4074 VP.n7303 VP.n7302 0.048
R4075 VP.n8131 VP.n8130 0.048
R4076 VP.n8975 VP.n8974 0.048
R4077 VP.n9749 VP.n9748 0.048
R4078 VP.n2798 VP.n2797 0.048
R4079 VP.n3738 VP.n3737 0.048
R4080 VP.n4644 VP.n4643 0.048
R4081 VP.n5539 VP.n5538 0.048
R4082 VP.n6395 VP.n6394 0.048
R4083 VP.n7254 VP.n7253 0.048
R4084 VP.n8082 VP.n8081 0.048
R4085 VP.n8926 VP.n8925 0.048
R4086 VP.n9727 VP.n9726 0.048
R4087 VP.n4671 VP.n4670 0.048
R4088 VP.n5566 VP.n5565 0.048
R4089 VP.n6422 VP.n6421 0.048
R4090 VP.n7281 VP.n7280 0.048
R4091 VP.n8109 VP.n8108 0.048
R4092 VP.n8953 VP.n8952 0.048
R4093 VP.n10087 VP.n10086 0.048
R4094 VP.n7903 VP.n7902 0.048
R4095 VP.n6152 VP.n6151 0.048
R4096 VP.n4332 VP.n4331 0.048
R4097 VP.n10180 VP.n10179 0.048
R4098 VP.n10349 VP.n10348 0.048
R4099 VP.n2606 VP.n2605 0.048
R4100 VP.n10096 VP.n10092 0.048
R4101 VP.n3380 VP.n3379 0.047
R4102 VP.n8762 VP.n8761 0.047
R4103 VP.n7039 VP.n7038 0.047
R4104 VP.n5260 VP.n5259 0.047
R4105 VP.n1402 VP.n1401 0.047
R4106 VP.t8 VP.n10178 0.047
R4107 VP.n311 VP.n310 0.047
R4108 VP.n150 VP.n149 0.047
R4109 VP.n2263 VP.n2249 0.047
R4110 VP.n2338 VP.n2336 0.047
R4111 VP.n3213 VP.n3200 0.047
R4112 VP.n3364 VP.n3363 0.047
R4113 VP.n4105 VP.n4091 0.047
R4114 VP.n4285 VP.n4284 0.047
R4115 VP.n4988 VP.n4974 0.047
R4116 VP.n5191 VP.n5190 0.047
R4117 VP.n5825 VP.n5811 0.047
R4118 VP.n6056 VP.n6054 0.047
R4119 VP.n6668 VP.n6655 0.047
R4120 VP.n6920 VP.n6918 0.047
R4121 VP.n7480 VP.n7467 0.047
R4122 VP.n7758 VP.n7757 0.047
R4123 VP.n8297 VP.n8283 0.047
R4124 VP.n8597 VP.n8596 0.047
R4125 VP.n9094 VP.n9080 0.047
R4126 VP.n9394 VP.n9392 0.047
R4127 VP.n9856 VP.n9843 0.047
R4128 VP.n10739 VP.n10737 0.047
R4129 VP.n10464 VP.n10462 0.047
R4130 VP.n10429 VP.n10427 0.047
R4131 VP.n10970 VP.n10955 0.047
R4132 VP.n9605 VP.n9603 0.047
R4133 VP.n10071 VP.n10051 0.047
R4134 VP.n11005 VP.n10981 0.047
R4135 VP.n10642 VP.n10618 0.047
R4136 VP.n8799 VP.n8797 0.047
R4137 VP.n9273 VP.n9255 0.047
R4138 VP.n9633 VP.n9616 0.047
R4139 VP.n10040 VP.n10011 0.047
R4140 VP.n10946 VP.n10922 0.047
R4141 VP.n10604 VP.n10580 0.047
R4142 VP.n8770 VP.n8754 0.047
R4143 VP.n9043 VP.n9040 0.047
R4144 VP.n9574 VP.n9572 0.047
R4145 VP.n9807 VP.n9805 0.047
R4146 VP.n10911 VP.n10909 0.047
R4147 VP.n10403 VP.n10398 0.047
R4148 VP.n8205 VP.n8203 0.047
R4149 VP.n7908 VP.n7906 0.047
R4150 VP.n7076 VP.n7074 0.047
R4151 VP.n7607 VP.n7589 0.047
R4152 VP.n7968 VP.n7951 0.047
R4153 VP.n8446 VP.n8417 0.047
R4154 VP.n8744 VP.n8727 0.047
R4155 VP.n9244 VP.n9217 0.047
R4156 VP.n9551 VP.n9533 0.047
R4157 VP.n10000 VP.n9974 0.047
R4158 VP.n10895 VP.n10871 0.047
R4159 VP.n10569 VP.n10545 0.047
R4160 VP.n7047 VP.n7031 0.047
R4161 VP.n7348 VP.n7345 0.047
R4162 VP.n7881 VP.n7880 0.047
R4163 VP.n8169 VP.n8166 0.047
R4164 VP.n8717 VP.n8716 0.047
R4165 VP.n9013 VP.n9010 0.047
R4166 VP.n9522 VP.n9520 0.047
R4167 VP.n9785 VP.n9783 0.047
R4168 VP.n10860 VP.n10858 0.047
R4169 VP.n10386 VP.n10381 0.047
R4170 VP.n6495 VP.n6493 0.047
R4171 VP.n6157 VP.n6155 0.047
R4172 VP.n5297 VP.n5295 0.047
R4173 VP.n5904 VP.n5886 0.047
R4174 VP.n6281 VP.n6264 0.047
R4175 VP.n6768 VP.n6739 0.047
R4176 VP.n7021 VP.n7004 0.047
R4177 VP.n7578 VP.n7551 0.047
R4178 VP.n7859 VP.n7842 0.047
R4179 VP.n8395 VP.n8368 0.047
R4180 VP.n8696 VP.n8679 0.047
R4181 VP.n9194 VP.n9167 0.047
R4182 VP.n9500 VP.n9482 0.047
R4183 VP.n9952 VP.n9926 0.047
R4184 VP.n10844 VP.n10820 0.047
R4185 VP.n10534 VP.n10510 0.047
R4186 VP.n5268 VP.n5252 0.047
R4187 VP.n5610 VP.n5607 0.047
R4188 VP.n6130 VP.n6129 0.047
R4189 VP.n6459 VP.n6456 0.047
R4190 VP.n6993 VP.n6992 0.047
R4191 VP.n7318 VP.n7315 0.047
R4192 VP.n7831 VP.n7830 0.047
R4193 VP.n8146 VP.n8143 0.047
R4194 VP.n8669 VP.n8668 0.047
R4195 VP.n8990 VP.n8987 0.047
R4196 VP.n9471 VP.n9469 0.047
R4197 VP.n9763 VP.n9761 0.047
R4198 VP.n10809 VP.n10807 0.047
R4199 VP.n10369 VP.n10364 0.047
R4200 VP.n4721 VP.n4719 0.047
R4201 VP.n4337 VP.n4335 0.047
R4202 VP.n3420 VP.n3418 0.047
R4203 VP.n4134 VP.n4116 0.047
R4204 VP.n4530 VP.n4513 0.047
R4205 VP.n5040 VP.n5011 0.047
R4206 VP.n5242 VP.n5225 0.047
R4207 VP.n5875 VP.n5848 0.047
R4208 VP.n6108 VP.n6091 0.047
R4209 VP.n6717 VP.n6690 0.047
R4210 VP.n6972 VP.n6955 0.047
R4211 VP.n7529 VP.n7502 0.047
R4212 VP.n7810 VP.n7793 0.047
R4213 VP.n8346 VP.n8319 0.047
R4214 VP.n8648 VP.n8631 0.047
R4215 VP.n9144 VP.n9117 0.047
R4216 VP.n9449 VP.n9431 0.047
R4217 VP.n9904 VP.n9878 0.047
R4218 VP.n10793 VP.n10769 0.047
R4219 VP.n10499 VP.n10475 0.047
R4220 VP.n345 VP.n343 0.047
R4221 VP.n873 VP.n871 0.047
R4222 VP.n1414 VP.n1413 0.047
R4223 VP.n1860 VP.n1857 0.047
R4224 VP.n2626 VP.n2625 0.047
R4225 VP.n2813 VP.n2810 0.047
R4226 VP.n3337 VP.n3336 0.047
R4227 VP.n3753 VP.n3750 0.047
R4228 VP.n4258 VP.n4257 0.047
R4229 VP.n4659 VP.n4656 0.047
R4230 VP.n5164 VP.n5163 0.047
R4231 VP.n5554 VP.n5551 0.047
R4232 VP.n6028 VP.n6027 0.047
R4233 VP.n6410 VP.n6407 0.047
R4234 VP.n6892 VP.n6891 0.047
R4235 VP.n7269 VP.n7266 0.047
R4236 VP.n7731 VP.n7730 0.047
R4237 VP.n8097 VP.n8094 0.047
R4238 VP.n8570 VP.n8569 0.047
R4239 VP.n8941 VP.n8938 0.047
R4240 VP.n9365 VP.n9363 0.047
R4241 VP.n9741 VP.n9739 0.047
R4242 VP.n10710 VP.n10708 0.047
R4243 VP.n10144 VP.n10142 0.047
R4244 VP.n11032 VP.n11020 0.047
R4245 VP.n9719 VP.n9706 0.047
R4246 VP.n9343 VP.n9341 0.047
R4247 VP.n8918 VP.n8915 0.047
R4248 VP.n8549 VP.n8548 0.047
R4249 VP.n8074 VP.n8071 0.047
R4250 VP.n7710 VP.n7709 0.047
R4251 VP.n7246 VP.n7243 0.047
R4252 VP.n6871 VP.n6870 0.047
R4253 VP.n6387 VP.n6384 0.047
R4254 VP.n6007 VP.n6006 0.047
R4255 VP.n5531 VP.n5528 0.047
R4256 VP.n5143 VP.n5142 0.047
R4257 VP.n4636 VP.n4633 0.047
R4258 VP.n4237 VP.n4236 0.047
R4259 VP.n3730 VP.n3727 0.047
R4260 VP.n3316 VP.n3315 0.047
R4261 VP.n2790 VP.n2787 0.047
R4262 VP.n2651 VP.n2650 0.047
R4263 VP.n1830 VP.n1827 0.047
R4264 VP.n1390 VP.n1389 0.047
R4265 VP.n847 VP.n843 0.047
R4266 VP.n313 VP.n300 0.047
R4267 VP.n758 VP.n737 0.047
R4268 VP.n392 VP.n374 0.047
R4269 VP.n924 VP.n910 0.047
R4270 VP.n1747 VP.n1738 0.047
R4271 VP.n439 VP.n421 0.047
R4272 VP.n974 VP.n960 0.047
R4273 VP.n1480 VP.n1472 0.047
R4274 VP.n1913 VP.n1897 0.047
R4275 VP.n2708 VP.n2699 0.047
R4276 VP.n486 VP.n468 0.047
R4277 VP.n1024 VP.n1010 0.047
R4278 VP.n1518 VP.n1510 0.047
R4279 VP.n1965 VP.n1949 0.047
R4280 VP.n2580 VP.n2572 0.047
R4281 VP.n2894 VP.n2878 0.047
R4282 VP.n3648 VP.n3639 0.047
R4283 VP.n533 VP.n515 0.047
R4284 VP.n1074 VP.n1060 0.047
R4285 VP.n1556 VP.n1548 0.047
R4286 VP.n2017 VP.n2001 0.047
R4287 VP.n2542 VP.n2534 0.047
R4288 VP.n2946 VP.n2930 0.047
R4289 VP.n3458 VP.n3450 0.047
R4290 VP.n3839 VP.n3823 0.047
R4291 VP.n4554 VP.n4545 0.047
R4292 VP.n580 VP.n562 0.047
R4293 VP.n1124 VP.n1110 0.047
R4294 VP.n1594 VP.n1586 0.047
R4295 VP.n2069 VP.n2053 0.047
R4296 VP.n2504 VP.n2496 0.047
R4297 VP.n2998 VP.n2982 0.047
R4298 VP.n3496 VP.n3488 0.047
R4299 VP.n3891 VP.n3875 0.047
R4300 VP.n4375 VP.n4367 0.047
R4301 VP.n4774 VP.n4758 0.047
R4302 VP.n5449 VP.n5440 0.047
R4303 VP.n620 VP.n609 0.047
R4304 VP.n1162 VP.n1160 0.047
R4305 VP.n1626 VP.n1624 0.047
R4306 VP.n2110 VP.n2105 0.047
R4307 VP.n2466 VP.n2464 0.047
R4308 VP.n3039 VP.n3034 0.047
R4309 VP.n3528 VP.n3526 0.047
R4310 VP.n3932 VP.n3927 0.047
R4311 VP.n4407 VP.n4405 0.047
R4312 VP.n4815 VP.n4810 0.047
R4313 VP.n5329 VP.n5327 0.047
R4314 VP.n5652 VP.n5647 0.047
R4315 VP.n6305 VP.n6296 0.047
R4316 VP.n650 VP.n649 0.047
R4317 VP.n1202 VP.n1198 0.047
R4318 VP.n1658 VP.n1656 0.047
R4319 VP.n2151 VP.n2146 0.047
R4320 VP.n2434 VP.n2432 0.047
R4321 VP.n3080 VP.n3075 0.047
R4322 VP.n3560 VP.n3558 0.047
R4323 VP.n3973 VP.n3968 0.047
R4324 VP.n4439 VP.n4437 0.047
R4325 VP.n4856 VP.n4851 0.047
R4326 VP.n5361 VP.n5359 0.047
R4327 VP.n5693 VP.n5688 0.047
R4328 VP.n6189 VP.n6187 0.047
R4329 VP.n6537 VP.n6532 0.047
R4330 VP.n7164 VP.n7155 0.047
R4331 VP.n682 VP.n679 0.047
R4332 VP.n1243 VP.n1238 0.047
R4333 VP.n1690 VP.n1688 0.047
R4334 VP.n2192 VP.n2187 0.047
R4335 VP.n2402 VP.n2400 0.047
R4336 VP.n3121 VP.n3116 0.047
R4337 VP.n3592 VP.n3590 0.047
R4338 VP.n4014 VP.n4009 0.047
R4339 VP.n4471 VP.n4469 0.047
R4340 VP.n4897 VP.n4892 0.047
R4341 VP.n5393 VP.n5391 0.047
R4342 VP.n5734 VP.n5729 0.047
R4343 VP.n6221 VP.n6219 0.047
R4344 VP.n6578 VP.n6573 0.047
R4345 VP.n7108 VP.n7106 0.047
R4346 VP.n7390 VP.n7385 0.047
R4347 VP.n7992 VP.n7983 0.047
R4348 VP.n287 VP.n272 0.047
R4349 VP.n815 VP.n785 0.047
R4350 VP.n1365 VP.n1344 0.047
R4351 VP.n1801 VP.n1774 0.047
R4352 VP.n2682 VP.n2661 0.047
R4353 VP.n2761 VP.n2734 0.047
R4354 VP.n3291 VP.n3270 0.047
R4355 VP.n3701 VP.n3674 0.047
R4356 VP.n4212 VP.n4191 0.047
R4357 VP.n4610 VP.n4580 0.047
R4358 VP.n5118 VP.n5097 0.047
R4359 VP.n5502 VP.n5475 0.047
R4360 VP.n5982 VP.n5961 0.047
R4361 VP.n6358 VP.n6331 0.047
R4362 VP.n6846 VP.n6825 0.047
R4363 VP.n7217 VP.n7190 0.047
R4364 VP.n7685 VP.n7664 0.047
R4365 VP.n8045 VP.n8018 0.047
R4366 VP.n8524 VP.n8503 0.047
R4367 VP.n8889 VP.n8864 0.047
R4368 VP.n9659 VP.n9648 0.047
R4369 VP.n2233 VP.n2228 0.047
R4370 VP.n2370 VP.n2368 0.047
R4371 VP.n3162 VP.n3157 0.047
R4372 VP.n3624 VP.n3622 0.047
R4373 VP.n4055 VP.n4050 0.047
R4374 VP.n4503 VP.n4501 0.047
R4375 VP.n4938 VP.n4933 0.047
R4376 VP.n5425 VP.n5423 0.047
R4377 VP.n5775 VP.n5770 0.047
R4378 VP.n6253 VP.n6251 0.047
R4379 VP.n6619 VP.n6614 0.047
R4380 VP.n7140 VP.n7138 0.047
R4381 VP.n7431 VP.n7426 0.047
R4382 VP.n7940 VP.n7938 0.047
R4383 VP.n8247 VP.n8242 0.047
R4384 VP.n8826 VP.n8814 0.047
R4385 VP.n722 VP.n711 0.047
R4386 VP.n1284 VP.n1279 0.047
R4387 VP.n1723 VP.n1720 0.047
R4388 VP.n1442 VP.n1441 0.047
R4389 VP.n10096 VP.n10095 0.047
R4390 VP.n856 VP.n855 0.046
R4391 VP.n1839 VP.n1837 0.046
R4392 VP.n3766 VP.n3764 0.046
R4393 VP.n9022 VP.n9021 0.046
R4394 VP.n7327 VP.n7326 0.046
R4395 VP.n5589 VP.n5588 0.046
R4396 VP.n9693 VP.n9692 0.046
R4397 VP.n8903 VP.n8902 0.046
R4398 VP.n8059 VP.n8058 0.046
R4399 VP.n7231 VP.n7230 0.046
R4400 VP.n6372 VP.n6371 0.046
R4401 VP.n5516 VP.n5515 0.046
R4402 VP.n4621 VP.n4620 0.046
R4403 VP.n3715 VP.n3714 0.046
R4404 VP.n2775 VP.n2774 0.046
R4405 VP.n1815 VP.n1814 0.046
R4406 VP.n9309 VP.n9308 0.045
R4407 VP.n11001 VP.n11000 0.045
R4408 VP.n10637 VP.n10636 0.045
R4409 VP.n10942 VP.n10941 0.045
R4410 VP.n10595 VP.n10594 0.045
R4411 VP.n8740 VP.n8739 0.045
R4412 VP.n9547 VP.n9546 0.045
R4413 VP.n10891 VP.n10890 0.045
R4414 VP.n10560 VP.n10559 0.045
R4415 VP.n7017 VP.n7016 0.045
R4416 VP.n7855 VP.n7854 0.045
R4417 VP.n8692 VP.n8691 0.045
R4418 VP.n9496 VP.n9495 0.045
R4419 VP.n10840 VP.n10839 0.045
R4420 VP.n10525 VP.n10524 0.045
R4421 VP.n5238 VP.n5237 0.045
R4422 VP.n6104 VP.n6103 0.045
R4423 VP.n6968 VP.n6967 0.045
R4424 VP.n7806 VP.n7805 0.045
R4425 VP.n8644 VP.n8643 0.045
R4426 VP.n9445 VP.n9444 0.045
R4427 VP.n10789 VP.n10788 0.045
R4428 VP.n10490 VP.n10489 0.045
R4429 VP.n10722 VP.n10721 0.045
R4430 VP.n9377 VP.n9376 0.045
R4431 VP.n8582 VP.n8581 0.045
R4432 VP.n7743 VP.n7742 0.045
R4433 VP.n6904 VP.n6903 0.045
R4434 VP.n6040 VP.n6039 0.045
R4435 VP.n5176 VP.n5175 0.045
R4436 VP.n4270 VP.n4269 0.045
R4437 VP.n3349 VP.n3348 0.045
R4438 VP.n10132 VP.n10131 0.045
R4439 VP.n10697 VP.n10691 0.045
R4440 VP.n1310 VP.n1309 0.045
R4441 VP.n769 VP.n768 0.045
R4442 VP.n2287 VP.n2286 0.045
R4443 VP.n1745 VP.n1742 0.045
R4444 VP.n896 VP.n895 0.045
R4445 VP.n1330 VP.n1329 0.045
R4446 VP.n1758 VP.n1757 0.045
R4447 VP.n3237 VP.n3236 0.045
R4448 VP.n2706 VP.n2703 0.045
R4449 VP.n946 VP.n945 0.045
R4450 VP.n1458 VP.n1457 0.045
R4451 VP.n1883 VP.n1882 0.045
R4452 VP.n2306 VP.n2305 0.045
R4453 VP.n2719 VP.n2718 0.045
R4454 VP.n4158 VP.n4157 0.045
R4455 VP.n3646 VP.n3643 0.045
R4456 VP.n996 VP.n995 0.045
R4457 VP.n1496 VP.n1495 0.045
R4458 VP.n1935 VP.n1934 0.045
R4459 VP.n2558 VP.n2557 0.045
R4460 VP.n2864 VP.n2863 0.045
R4461 VP.n3256 VP.n3255 0.045
R4462 VP.n3659 VP.n3658 0.045
R4463 VP.n5064 VP.n5063 0.045
R4464 VP.n4552 VP.n4549 0.045
R4465 VP.n1046 VP.n1045 0.045
R4466 VP.n1534 VP.n1533 0.045
R4467 VP.n1987 VP.n1986 0.045
R4468 VP.n2520 VP.n2519 0.045
R4469 VP.n2916 VP.n2915 0.045
R4470 VP.n3436 VP.n3435 0.045
R4471 VP.n3809 VP.n3808 0.045
R4472 VP.n4177 VP.n4176 0.045
R4473 VP.n4565 VP.n4564 0.045
R4474 VP.n5928 VP.n5927 0.045
R4475 VP.n5447 VP.n5444 0.045
R4476 VP.n1096 VP.n1095 0.045
R4477 VP.n1572 VP.n1571 0.045
R4478 VP.n2039 VP.n2038 0.045
R4479 VP.n2482 VP.n2481 0.045
R4480 VP.n2968 VP.n2967 0.045
R4481 VP.n3474 VP.n3473 0.045
R4482 VP.n3861 VP.n3860 0.045
R4483 VP.n4353 VP.n4352 0.045
R4484 VP.n4744 VP.n4743 0.045
R4485 VP.n5083 VP.n5082 0.045
R4486 VP.n5460 VP.n5459 0.045
R4487 VP.n6792 VP.n6791 0.045
R4488 VP.n6303 VP.n6300 0.045
R4489 VP.n1146 VP.n1145 0.045
R4490 VP.n1610 VP.n1609 0.045
R4491 VP.n2091 VP.n2090 0.045
R4492 VP.n2450 VP.n2449 0.045
R4493 VP.n3020 VP.n3019 0.045
R4494 VP.n3512 VP.n3511 0.045
R4495 VP.n3913 VP.n3912 0.045
R4496 VP.n4391 VP.n4390 0.045
R4497 VP.n4796 VP.n4795 0.045
R4498 VP.n5313 VP.n5312 0.045
R4499 VP.n5633 VP.n5632 0.045
R4500 VP.n5947 VP.n5946 0.045
R4501 VP.n6316 VP.n6315 0.045
R4502 VP.n7631 VP.n7630 0.045
R4503 VP.n7162 VP.n7159 0.045
R4504 VP.n1184 VP.n1183 0.045
R4505 VP.n1642 VP.n1641 0.045
R4506 VP.n2132 VP.n2131 0.045
R4507 VP.n2418 VP.n2417 0.045
R4508 VP.n3061 VP.n3060 0.045
R4509 VP.n3544 VP.n3543 0.045
R4510 VP.n3954 VP.n3953 0.045
R4511 VP.n4423 VP.n4422 0.045
R4512 VP.n4837 VP.n4836 0.045
R4513 VP.n5345 VP.n5344 0.045
R4514 VP.n5674 VP.n5673 0.045
R4515 VP.n6173 VP.n6172 0.045
R4516 VP.n6518 VP.n6517 0.045
R4517 VP.n6811 VP.n6810 0.045
R4518 VP.n7175 VP.n7174 0.045
R4519 VP.n8470 VP.n8469 0.045
R4520 VP.n7990 VP.n7987 0.045
R4521 VP.n1224 VP.n1223 0.045
R4522 VP.n1674 VP.n1673 0.045
R4523 VP.n2173 VP.n2172 0.045
R4524 VP.n2386 VP.n2385 0.045
R4525 VP.n3102 VP.n3101 0.045
R4526 VP.n3576 VP.n3575 0.045
R4527 VP.n3995 VP.n3994 0.045
R4528 VP.n4455 VP.n4454 0.045
R4529 VP.n4878 VP.n4877 0.045
R4530 VP.n5377 VP.n5376 0.045
R4531 VP.n5715 VP.n5714 0.045
R4532 VP.n6205 VP.n6204 0.045
R4533 VP.n6559 VP.n6558 0.045
R4534 VP.n7092 VP.n7091 0.045
R4535 VP.n7371 VP.n7370 0.045
R4536 VP.n7650 VP.n7649 0.045
R4537 VP.n8003 VP.n8002 0.045
R4538 VP.n9676 VP.n9675 0.045
R4539 VP.n1265 VP.n1264 0.045
R4540 VP.n1706 VP.n1705 0.045
R4541 VP.n2214 VP.n2213 0.045
R4542 VP.n2354 VP.n2353 0.045
R4543 VP.n3143 VP.n3142 0.045
R4544 VP.n3608 VP.n3607 0.045
R4545 VP.n4036 VP.n4035 0.045
R4546 VP.n4487 VP.n4486 0.045
R4547 VP.n4919 VP.n4918 0.045
R4548 VP.n5409 VP.n5408 0.045
R4549 VP.n5756 VP.n5755 0.045
R4550 VP.n6237 VP.n6236 0.045
R4551 VP.n6600 VP.n6599 0.045
R4552 VP.n7124 VP.n7123 0.045
R4553 VP.n7412 VP.n7411 0.045
R4554 VP.n7924 VP.n7923 0.045
R4555 VP.n8228 VP.n8227 0.045
R4556 VP.n8489 VP.n8488 0.045
R4557 VP.n8837 VP.n8836 0.045
R4558 VP.n9297 VP.n9296 0.045
R4559 VP.n811 VP.n810 0.045
R4560 VP.n1361 VP.n1360 0.045
R4561 VP.n1797 VP.n1796 0.045
R4562 VP.n2678 VP.n2677 0.045
R4563 VP.n2757 VP.n2756 0.045
R4564 VP.n3287 VP.n3286 0.045
R4565 VP.n3697 VP.n3696 0.045
R4566 VP.n4208 VP.n4207 0.045
R4567 VP.n4606 VP.n4605 0.045
R4568 VP.n5114 VP.n5113 0.045
R4569 VP.n5498 VP.n5497 0.045
R4570 VP.n5978 VP.n5977 0.045
R4571 VP.n6354 VP.n6353 0.045
R4572 VP.n6842 VP.n6841 0.045
R4573 VP.n7213 VP.n7212 0.045
R4574 VP.n7681 VP.n7680 0.045
R4575 VP.n8041 VP.n8040 0.045
R4576 VP.n8520 VP.n8519 0.045
R4577 VP.n8885 VP.n8884 0.045
R4578 VP.n10658 VP.n10657 0.045
R4579 VP.n260 VP.n257 0.045
R4580 VP.n362 VP.n359 0.045
R4581 VP.n409 VP.n406 0.045
R4582 VP.n456 VP.n453 0.045
R4583 VP.n503 VP.n500 0.045
R4584 VP.n550 VP.n547 0.045
R4585 VP.n597 VP.n594 0.045
R4586 VP.n637 VP.n634 0.045
R4587 VP.n667 VP.n664 0.045
R4588 VP.n699 VP.n696 0.045
R4589 VP.n10031 VP.n10030 0.044
R4590 VP.n8437 VP.n8436 0.044
R4591 VP.n6759 VP.n6758 0.044
R4592 VP.n5031 VP.n5030 0.044
R4593 VP.n3188 VP.n3182 0.044
R4594 VP.n721 VP.n720 0.044
R4595 VP.n10321 VP.n10320 0.044
R4596 VP.n10303 VP.n10302 0.044
R4597 VP.n10275 VP.n10274 0.044
R4598 VP.n10247 VP.n10246 0.044
R4599 VP.n10219 VP.n10218 0.044
R4600 VP.n10196 VP.n10195 0.044
R4601 VP.n9306 VP.n8827 0.043
R4602 VP.n11047 VP.n11046 0.043
R4603 VP.n8185 VP.n8184 0.043
R4604 VP.n6475 VP.n6474 0.043
R4605 VP.n4701 VP.n4700 0.043
R4606 VP.n9264 VP.n9261 0.043
R4607 VP.n7598 VP.n7595 0.043
R4608 VP.n5895 VP.n5892 0.043
R4609 VP.n4125 VP.n4122 0.043
R4610 VP.n1320 VP.n759 0.043
R4611 VP.n2296 VP.n1748 0.043
R4612 VP.n3246 VP.n2709 0.043
R4613 VP.n4167 VP.n3649 0.043
R4614 VP.n5073 VP.n4555 0.043
R4615 VP.n5937 VP.n5450 0.043
R4616 VP.n6801 VP.n6306 0.043
R4617 VP.n7640 VP.n7165 0.043
R4618 VP.n8479 VP.n7993 0.043
R4619 VP.n9992 VP.n9991 0.042
R4620 VP.n9236 VP.n9235 0.042
R4621 VP.n9944 VP.n9943 0.042
R4622 VP.n9186 VP.n9185 0.042
R4623 VP.n8387 VP.n8386 0.042
R4624 VP.n7570 VP.n7569 0.042
R4625 VP.n9896 VP.n9895 0.042
R4626 VP.n9136 VP.n9135 0.042
R4627 VP.n8338 VP.n8337 0.042
R4628 VP.n7521 VP.n7520 0.042
R4629 VP.n6709 VP.n6708 0.042
R4630 VP.n5867 VP.n5866 0.042
R4631 VP.n10451 VP.n10446 0.042
R4632 VP.n9832 VP.n9827 0.042
R4633 VP.n9069 VP.n9064 0.042
R4634 VP.n8272 VP.n8267 0.042
R4635 VP.n7456 VP.n7451 0.042
R4636 VP.n6644 VP.n6639 0.042
R4637 VP.n5800 VP.n5795 0.042
R4638 VP.n4963 VP.n4958 0.042
R4639 VP.n4080 VP.n4075 0.042
R4640 VP.n10615 VP.n10614 0.042
R4641 VP.n1282 VP.n1281 0.042
R4642 VP.n5650 VP.n5649 0.042
R4643 VP.n4813 VP.n4812 0.042
R4644 VP.n3930 VP.n3929 0.042
R4645 VP.n3037 VP.n3036 0.042
R4646 VP.n2108 VP.n2107 0.042
R4647 VP.n6535 VP.n6534 0.042
R4648 VP.n5691 VP.n5690 0.042
R4649 VP.n4854 VP.n4853 0.042
R4650 VP.n3971 VP.n3970 0.042
R4651 VP.n3078 VP.n3077 0.042
R4652 VP.n2149 VP.n2148 0.042
R4653 VP.n7388 VP.n7387 0.042
R4654 VP.n6576 VP.n6575 0.042
R4655 VP.n5732 VP.n5731 0.042
R4656 VP.n4895 VP.n4894 0.042
R4657 VP.n4012 VP.n4011 0.042
R4658 VP.n3119 VP.n3118 0.042
R4659 VP.n2190 VP.n2189 0.042
R4660 VP.n1241 VP.n1240 0.042
R4661 VP.n8245 VP.n8244 0.042
R4662 VP.n7429 VP.n7428 0.042
R4663 VP.n6617 VP.n6616 0.042
R4664 VP.n5773 VP.n5772 0.042
R4665 VP.n4936 VP.n4935 0.042
R4666 VP.n4053 VP.n4052 0.042
R4667 VP.n3160 VP.n3159 0.042
R4668 VP.n2231 VP.n2230 0.042
R4669 VP.t116 VP.n37 0.042
R4670 VP.t116 VP.n27 0.042
R4671 VP.t116 VP.n138 0.042
R4672 VP.n198 VP.n197 0.042
R4673 VP.n9313 VP.n9312 0.042
R4674 VP.n1313 VP.n1312 0.041
R4675 VP.n755 VP.n754 0.041
R4676 VP.n2257 VP.n2256 0.041
R4677 VP.n154 VP.n153 0.041
R4678 VP.n9042 VP.n9041 0.041
R4679 VP.n9012 VP.n9011 0.041
R4680 VP.n8168 VP.n8167 0.041
R4681 VP.n7347 VP.n7346 0.041
R4682 VP.n8989 VP.n8988 0.041
R4683 VP.n8145 VP.n8144 0.041
R4684 VP.n7317 VP.n7316 0.041
R4685 VP.n6458 VP.n6457 0.041
R4686 VP.n5609 VP.n5608 0.041
R4687 VP.n8940 VP.n8939 0.041
R4688 VP.n8096 VP.n8095 0.041
R4689 VP.n7268 VP.n7267 0.041
R4690 VP.n6409 VP.n6408 0.041
R4691 VP.n5553 VP.n5552 0.041
R4692 VP.n4658 VP.n4657 0.041
R4693 VP.n3752 VP.n3751 0.041
R4694 VP.n2812 VP.n2811 0.041
R4695 VP.n1859 VP.n1858 0.041
R4696 VP.n8015 VP.n8014 0.041
R4697 VP.n7187 VP.n7186 0.041
R4698 VP.n6328 VP.n6327 0.041
R4699 VP.n5472 VP.n5471 0.041
R4700 VP.n4577 VP.n4576 0.041
R4701 VP.n3671 VP.n3670 0.041
R4702 VP.n2731 VP.n2730 0.041
R4703 VP.n1771 VP.n1770 0.041
R4704 VP.n782 VP.n781 0.041
R4705 VP.n8961 VP.n8960 0.041
R4706 VP.n8117 VP.n8116 0.041
R4707 VP.n7289 VP.n7288 0.041
R4708 VP.n6430 VP.n6429 0.041
R4709 VP.n5574 VP.n5573 0.041
R4710 VP.n4679 VP.n4678 0.041
R4711 VP.n3780 VP.n3779 0.041
R4712 VP.n846 VP.n845 0.041
R4713 VP.n1829 VP.n1828 0.041
R4714 VP.n2789 VP.n2788 0.041
R4715 VP.n3729 VP.n3728 0.041
R4716 VP.n4635 VP.n4634 0.041
R4717 VP.n5530 VP.n5529 0.041
R4718 VP.n6386 VP.n6385 0.041
R4719 VP.n7245 VP.n7244 0.041
R4720 VP.n8073 VP.n8072 0.041
R4721 VP.n8917 VP.n8916 0.041
R4722 VP.n10600 VP.n10599 0.041
R4723 VP.n10565 VP.n10564 0.041
R4724 VP.n10530 VP.n10529 0.041
R4725 VP.n10495 VP.n10494 0.041
R4726 VP.n9697 VP.n9694 0.041
R4727 VP.n9332 VP.n9330 0.041
R4728 VP.n8906 VP.n8904 0.041
R4729 VP.n8539 VP.n8537 0.041
R4730 VP.n8062 VP.n8060 0.041
R4731 VP.n7700 VP.n7698 0.041
R4732 VP.n7234 VP.n7232 0.041
R4733 VP.n6861 VP.n6859 0.041
R4734 VP.n6375 VP.n6373 0.041
R4735 VP.n5997 VP.n5995 0.041
R4736 VP.n5519 VP.n5517 0.041
R4737 VP.n5133 VP.n5131 0.041
R4738 VP.n4624 VP.n4622 0.041
R4739 VP.n4227 VP.n4225 0.041
R4740 VP.n3718 VP.n3716 0.041
R4741 VP.n3306 VP.n3304 0.041
R4742 VP.n2778 VP.n2776 0.041
R4743 VP.n2641 VP.n2639 0.041
R4744 VP.n1818 VP.n1816 0.041
R4745 VP.n1380 VP.n1378 0.041
R4746 VP.n834 VP.n832 0.041
R4747 VP.n1201 VP.n1200 0.04
R4748 VP.n9214 VP.n9202 0.04
R4749 VP.n9164 VP.n9152 0.04
R4750 VP.n9114 VP.n9102 0.04
R4751 VP.n5845 VP.n5833 0.04
R4752 VP.n9093 VP.n9081 0.04
R4753 VP.n8296 VP.n8284 0.04
R4754 VP.n5824 VP.n5812 0.04
R4755 VP.n4987 VP.n4975 0.04
R4756 VP.n4104 VP.n4092 0.04
R4757 VP.n197 VP.n159 0.04
R4758 VP.n619 VP.n618 0.04
R4759 VP.n9268 VP.n9267 0.04
R4760 VP.n9560 VP.n9559 0.04
R4761 VP.n7602 VP.n7601 0.04
R4762 VP.n7868 VP.n7867 0.04
R4763 VP.n8705 VP.n8704 0.04
R4764 VP.n9509 VP.n9508 0.04
R4765 VP.n5899 VP.n5898 0.04
R4766 VP.n6117 VP.n6116 0.04
R4767 VP.n6981 VP.n6980 0.04
R4768 VP.n7819 VP.n7818 0.04
R4769 VP.n8657 VP.n8656 0.04
R4770 VP.n9458 VP.n9457 0.04
R4771 VP.n4129 VP.n4128 0.04
R4772 VP.n2259 VP.n2258 0.04
R4773 VP.n2613 VP.n2612 0.04
R4774 VP.n3325 VP.n3324 0.04
R4775 VP.n4246 VP.n4245 0.04
R4776 VP.n5152 VP.n5151 0.04
R4777 VP.n6016 VP.n6015 0.04
R4778 VP.n6880 VP.n6879 0.04
R4779 VP.n7719 VP.n7718 0.04
R4780 VP.n8558 VP.n8557 0.04
R4781 VP.n9352 VP.n9351 0.04
R4782 VP.n381 VP.n380 0.04
R4783 VP.n428 VP.n427 0.04
R4784 VP.n475 VP.n474 0.04
R4785 VP.n522 VP.n521 0.04
R4786 VP.n569 VP.n568 0.04
R4787 VP.n4298 VP.n4297 0.04
R4788 VP.n5204 VP.n5203 0.04
R4789 VP.n6069 VP.n6068 0.04
R4790 VP.n6933 VP.n6932 0.04
R4791 VP.n7771 VP.n7770 0.04
R4792 VP.n8610 VP.n8609 0.04
R4793 VP.n9408 VP.n9407 0.04
R4794 VP.n303 VP.n302 0.04
R4795 VP.t8 VP.n10326 0.04
R4796 VP.n131 VP.n130 0.039
R4797 VP.n124 VP.n123 0.039
R4798 VP.n111 VP.n110 0.039
R4799 VP.n91 VP.n90 0.039
R4800 VP.n85 VP.n84 0.039
R4801 VP.n65 VP.n64 0.039
R4802 VP.n59 VP.n58 0.039
R4803 VP.n39 VP.n38 0.039
R4804 VP.n29 VP.n28 0.039
R4805 VP.n19 VP.n18 0.039
R4806 VP.n13 VP.n12 0.039
R4807 VP.n1438 VP.n1427 0.039
R4808 VP.n10347 VP.n10345 0.039
R4809 VP.n10967 VP.n10956 0.039
R4810 VP.n9592 VP.n9581 0.039
R4811 VP.n8788 VP.n8777 0.039
R4812 VP.n7901 VP.n7890 0.039
R4813 VP.n7065 VP.n7054 0.039
R4814 VP.n6150 VP.n6139 0.039
R4815 VP.n5286 VP.n5275 0.039
R4816 VP.n4330 VP.n4319 0.039
R4817 VP.n3409 VP.n3398 0.039
R4818 VP.n2604 VP.n2593 0.039
R4819 VP.n9408 VP.n9405 0.039
R4820 VP.n8610 VP.n8608 0.039
R4821 VP.n7771 VP.n7769 0.039
R4822 VP.n6933 VP.n6931 0.039
R4823 VP.n6069 VP.n6067 0.039
R4824 VP.n5204 VP.n5202 0.039
R4825 VP.n4298 VP.n4296 0.039
R4826 VP.n10931 VP.n10930 0.039
R4827 VP.n9260 VP.n9259 0.039
R4828 VP.n9560 VP.n9558 0.039
R4829 VP.n10880 VP.n10879 0.039
R4830 VP.n9541 VP.n9540 0.039
R4831 VP.n8734 VP.n8733 0.039
R4832 VP.n7594 VP.n7593 0.039
R4833 VP.n9509 VP.n9507 0.039
R4834 VP.n8705 VP.n8703 0.039
R4835 VP.n7868 VP.n7866 0.039
R4836 VP.n10829 VP.n10828 0.039
R4837 VP.n9490 VP.n9489 0.039
R4838 VP.n8686 VP.n8685 0.039
R4839 VP.n7849 VP.n7848 0.039
R4840 VP.n7011 VP.n7010 0.039
R4841 VP.n5891 VP.n5890 0.039
R4842 VP.n9458 VP.n9456 0.039
R4843 VP.n8657 VP.n8655 0.039
R4844 VP.n7819 VP.n7817 0.039
R4845 VP.n6981 VP.n6979 0.039
R4846 VP.n6117 VP.n6115 0.039
R4847 VP.n10778 VP.n10777 0.039
R4848 VP.n9439 VP.n9438 0.039
R4849 VP.n8638 VP.n8637 0.039
R4850 VP.n7800 VP.n7799 0.039
R4851 VP.n6962 VP.n6961 0.039
R4852 VP.n6098 VP.n6097 0.039
R4853 VP.n5232 VP.n5231 0.039
R4854 VP.n4121 VP.n4120 0.039
R4855 VP.n10718 VP.n10717 0.039
R4856 VP.n9373 VP.n9372 0.039
R4857 VP.n8578 VP.n8577 0.039
R4858 VP.n7739 VP.n7738 0.039
R4859 VP.n6900 VP.n6899 0.039
R4860 VP.n6036 VP.n6035 0.039
R4861 VP.n5172 VP.n5171 0.039
R4862 VP.n4266 VP.n4265 0.039
R4863 VP.n3345 VP.n3344 0.039
R4864 VP.n2259 VP.n2253 0.039
R4865 VP.n9352 VP.n9350 0.039
R4866 VP.n8558 VP.n8556 0.039
R4867 VP.n7719 VP.n7717 0.039
R4868 VP.n6880 VP.n6878 0.039
R4869 VP.n6016 VP.n6014 0.039
R4870 VP.n5152 VP.n5150 0.039
R4871 VP.n4246 VP.n4244 0.039
R4872 VP.n3325 VP.n3323 0.039
R4873 VP.n2613 VP.n2611 0.039
R4874 VP.t116 VP.n145 0.039
R4875 VP.n10966 VP.n10958 0.039
R4876 VP.n9591 VP.n9583 0.039
R4877 VP.n8787 VP.n8779 0.039
R4878 VP.n7900 VP.n7892 0.039
R4879 VP.n7064 VP.n7056 0.039
R4880 VP.n6149 VP.n6141 0.039
R4881 VP.n5285 VP.n5277 0.039
R4882 VP.n4329 VP.n4321 0.039
R4883 VP.n3408 VP.n3400 0.039
R4884 VP.n2603 VP.n2595 0.039
R4885 VP.n1437 VP.n1429 0.039
R4886 VP.n339 VP.n330 0.039
R4887 VP.n340 VP.n328 0.039
R4888 VP.n9316 VP.n9313 0.038
R4889 VP.n5008 VP.n4996 0.038
R4890 VP.n8861 VP.n8848 0.038
R4891 VP.t8 VP.n10333 0.038
R4892 VP.n9272 VP.n9260 0.038
R4893 VP.n7606 VP.n7594 0.038
R4894 VP.n5903 VP.n5891 0.038
R4895 VP.n4133 VP.n4121 0.038
R4896 VP.n9264 VP.n9263 0.038
R4897 VP.n7598 VP.n7597 0.038
R4898 VP.n5895 VP.n5894 0.038
R4899 VP.n4125 VP.n4124 0.038
R4900 VP.n3211 VP.n3202 0.037
R4901 VP.n4103 VP.n4094 0.037
R4902 VP.n4986 VP.n4977 0.037
R4903 VP.n5823 VP.n5814 0.037
R4904 VP.n6666 VP.n6657 0.037
R4905 VP.n7478 VP.n7469 0.037
R4906 VP.n8295 VP.n8286 0.037
R4907 VP.n9092 VP.n9083 0.037
R4908 VP.n9854 VP.n9845 0.037
R4909 VP.n8413 VP.n8404 0.037
R4910 VP.n9213 VP.n9204 0.037
R4911 VP.n9970 VP.n9961 0.037
R4912 VP.n6735 VP.n6726 0.037
R4913 VP.n7547 VP.n7538 0.037
R4914 VP.n8364 VP.n8355 0.037
R4915 VP.n9163 VP.n9154 0.037
R4916 VP.n9922 VP.n9913 0.037
R4917 VP.n5007 VP.n4998 0.037
R4918 VP.n5844 VP.n5835 0.037
R4919 VP.n6686 VP.n6677 0.037
R4920 VP.n7498 VP.n7489 0.037
R4921 VP.n8315 VP.n8306 0.037
R4922 VP.n9113 VP.n9104 0.037
R4923 VP.n9874 VP.n9865 0.037
R4924 VP.n10133 VP.n10129 0.037
R4925 VP.n1317 VP.n1316 0.037
R4926 VP.n770 VP.n766 0.037
R4927 VP.n2293 VP.n2292 0.037
R4928 VP.n1759 VP.n1755 0.037
R4929 VP.n3243 VP.n3242 0.037
R4930 VP.n2720 VP.n2716 0.037
R4931 VP.n4164 VP.n4163 0.037
R4932 VP.n3660 VP.n3656 0.037
R4933 VP.n5070 VP.n5069 0.037
R4934 VP.n4566 VP.n4562 0.037
R4935 VP.n5934 VP.n5933 0.037
R4936 VP.n5461 VP.n5457 0.037
R4937 VP.n6798 VP.n6797 0.037
R4938 VP.n6317 VP.n6313 0.037
R4939 VP.n7637 VP.n7636 0.037
R4940 VP.n7176 VP.n7172 0.037
R4941 VP.n8476 VP.n8475 0.037
R4942 VP.n8004 VP.n8000 0.037
R4943 VP.n9682 VP.n9681 0.037
R4944 VP.n8838 VP.n8834 0.037
R4945 VP.n9303 VP.n9302 0.037
R4946 VP.n10109 VP.n10107 0.037
R4947 VP.n10119 VP.n10118 0.037
R4948 VP.n10659 VP.n10655 0.037
R4949 VP.n8860 VP.n8851 0.037
R4950 VP.n9717 VP.n9708 0.037
R4951 VP.n10071 VP.n10058 0.036
R4952 VP.n11005 VP.n10988 0.036
R4953 VP.n10642 VP.n10627 0.036
R4954 VP.n10946 VP.n10929 0.036
R4955 VP.n10604 VP.n10589 0.036
R4956 VP.n9574 VP.n9565 0.036
R4957 VP.n8744 VP.n8732 0.036
R4958 VP.n9551 VP.n9539 0.036
R4959 VP.n10895 VP.n10878 0.036
R4960 VP.n10569 VP.n10554 0.036
R4961 VP.n7881 VP.n7873 0.036
R4962 VP.n8717 VP.n8709 0.036
R4963 VP.n9522 VP.n9513 0.036
R4964 VP.n7021 VP.n7009 0.036
R4965 VP.n7859 VP.n7847 0.036
R4966 VP.n8696 VP.n8684 0.036
R4967 VP.n9500 VP.n9488 0.036
R4968 VP.n10844 VP.n10827 0.036
R4969 VP.n10534 VP.n10519 0.036
R4970 VP.n6130 VP.n6122 0.036
R4971 VP.n6993 VP.n6985 0.036
R4972 VP.n7831 VP.n7823 0.036
R4973 VP.n8669 VP.n8661 0.036
R4974 VP.n9471 VP.n9462 0.036
R4975 VP.n5242 VP.n5230 0.036
R4976 VP.n6108 VP.n6096 0.036
R4977 VP.n6972 VP.n6960 0.036
R4978 VP.n7810 VP.n7798 0.036
R4979 VP.n8648 VP.n8636 0.036
R4980 VP.n9449 VP.n9437 0.036
R4981 VP.n10793 VP.n10776 0.036
R4982 VP.n10499 VP.n10484 0.036
R4983 VP.n10739 VP.n10730 0.036
R4984 VP.n9394 VP.n9385 0.036
R4985 VP.n8597 VP.n8589 0.036
R4986 VP.n7758 VP.n7750 0.036
R4987 VP.n6920 VP.n6911 0.036
R4988 VP.n6056 VP.n6047 0.036
R4989 VP.n5191 VP.n5183 0.036
R4990 VP.n4285 VP.n4277 0.036
R4991 VP.n3364 VP.n3356 0.036
R4992 VP.n2626 VP.n2618 0.036
R4993 VP.n3337 VP.n3329 0.036
R4994 VP.n4258 VP.n4250 0.036
R4995 VP.n5164 VP.n5156 0.036
R4996 VP.n6028 VP.n6020 0.036
R4997 VP.n6892 VP.n6884 0.036
R4998 VP.n7731 VP.n7723 0.036
R4999 VP.n8570 VP.n8562 0.036
R5000 VP.n9365 VP.n9356 0.036
R5001 VP.n10710 VP.n10701 0.036
R5002 VP.n924 VP.n903 0.036
R5003 VP.n1747 VP.n1337 0.036
R5004 VP.n974 VP.n953 0.036
R5005 VP.n1480 VP.n1465 0.036
R5006 VP.n1913 VP.n1890 0.036
R5007 VP.n2708 VP.n2313 0.036
R5008 VP.n1024 VP.n1003 0.036
R5009 VP.n1518 VP.n1503 0.036
R5010 VP.n1965 VP.n1942 0.036
R5011 VP.n2580 VP.n2565 0.036
R5012 VP.n2894 VP.n2871 0.036
R5013 VP.n3648 VP.n3263 0.036
R5014 VP.n1074 VP.n1053 0.036
R5015 VP.n1556 VP.n1541 0.036
R5016 VP.n2017 VP.n1994 0.036
R5017 VP.n2542 VP.n2527 0.036
R5018 VP.n2946 VP.n2923 0.036
R5019 VP.n3458 VP.n3443 0.036
R5020 VP.n3839 VP.n3816 0.036
R5021 VP.n4554 VP.n4184 0.036
R5022 VP.n1124 VP.n1103 0.036
R5023 VP.n1594 VP.n1579 0.036
R5024 VP.n2069 VP.n2046 0.036
R5025 VP.n2504 VP.n2489 0.036
R5026 VP.n2998 VP.n2975 0.036
R5027 VP.n3496 VP.n3481 0.036
R5028 VP.n3891 VP.n3868 0.036
R5029 VP.n4375 VP.n4360 0.036
R5030 VP.n4774 VP.n4751 0.036
R5031 VP.n5449 VP.n5090 0.036
R5032 VP.n1162 VP.n1153 0.036
R5033 VP.n1626 VP.n1617 0.036
R5034 VP.n2110 VP.n2098 0.036
R5035 VP.n2466 VP.n2457 0.036
R5036 VP.n3039 VP.n3027 0.036
R5037 VP.n3528 VP.n3519 0.036
R5038 VP.n3932 VP.n3920 0.036
R5039 VP.n4407 VP.n4398 0.036
R5040 VP.n4815 VP.n4803 0.036
R5041 VP.n5329 VP.n5320 0.036
R5042 VP.n5652 VP.n5640 0.036
R5043 VP.n6305 VP.n5954 0.036
R5044 VP.n1202 VP.n1191 0.036
R5045 VP.n1658 VP.n1649 0.036
R5046 VP.n2151 VP.n2139 0.036
R5047 VP.n2434 VP.n2425 0.036
R5048 VP.n3080 VP.n3068 0.036
R5049 VP.n3560 VP.n3551 0.036
R5050 VP.n3973 VP.n3961 0.036
R5051 VP.n4439 VP.n4430 0.036
R5052 VP.n4856 VP.n4844 0.036
R5053 VP.n5361 VP.n5352 0.036
R5054 VP.n5693 VP.n5681 0.036
R5055 VP.n6189 VP.n6180 0.036
R5056 VP.n6537 VP.n6525 0.036
R5057 VP.n7164 VP.n6818 0.036
R5058 VP.n1243 VP.n1231 0.036
R5059 VP.n1690 VP.n1681 0.036
R5060 VP.n2192 VP.n2180 0.036
R5061 VP.n2402 VP.n2393 0.036
R5062 VP.n3121 VP.n3109 0.036
R5063 VP.n3592 VP.n3583 0.036
R5064 VP.n4014 VP.n4002 0.036
R5065 VP.n4471 VP.n4462 0.036
R5066 VP.n4897 VP.n4885 0.036
R5067 VP.n5393 VP.n5384 0.036
R5068 VP.n5734 VP.n5722 0.036
R5069 VP.n6221 VP.n6212 0.036
R5070 VP.n6578 VP.n6566 0.036
R5071 VP.n7108 VP.n7099 0.036
R5072 VP.n7390 VP.n7378 0.036
R5073 VP.n7992 VP.n7657 0.036
R5074 VP.n9659 VP.n9652 0.036
R5075 VP.n1284 VP.n1272 0.036
R5076 VP.n1723 VP.n1713 0.036
R5077 VP.n2233 VP.n2221 0.036
R5078 VP.n2370 VP.n2361 0.036
R5079 VP.n3162 VP.n3150 0.036
R5080 VP.n3624 VP.n3615 0.036
R5081 VP.n4055 VP.n4043 0.036
R5082 VP.n4503 VP.n4494 0.036
R5083 VP.n4938 VP.n4926 0.036
R5084 VP.n5425 VP.n5416 0.036
R5085 VP.n5775 VP.n5763 0.036
R5086 VP.n6253 VP.n6244 0.036
R5087 VP.n6619 VP.n6607 0.036
R5088 VP.n7140 VP.n7131 0.036
R5089 VP.n7431 VP.n7419 0.036
R5090 VP.n7940 VP.n7931 0.036
R5091 VP.n8247 VP.n8235 0.036
R5092 VP.n8826 VP.n8496 0.036
R5093 VP.n8826 VP.n8818 0.036
R5094 VP.n287 VP.n279 0.036
R5095 VP.n815 VP.n795 0.036
R5096 VP.n1365 VP.n1351 0.036
R5097 VP.n1801 VP.n1781 0.036
R5098 VP.n2682 VP.n2668 0.036
R5099 VP.n2761 VP.n2741 0.036
R5100 VP.n3291 VP.n3277 0.036
R5101 VP.n3701 VP.n3681 0.036
R5102 VP.n4212 VP.n4198 0.036
R5103 VP.n4610 VP.n4590 0.036
R5104 VP.n5118 VP.n5104 0.036
R5105 VP.n5502 VP.n5482 0.036
R5106 VP.n5982 VP.n5968 0.036
R5107 VP.n6358 VP.n6338 0.036
R5108 VP.n6846 VP.n6832 0.036
R5109 VP.n7217 VP.n7197 0.036
R5110 VP.n7685 VP.n7671 0.036
R5111 VP.n8045 VP.n8025 0.036
R5112 VP.n8524 VP.n8510 0.036
R5113 VP.n8889 VP.n8871 0.036
R5114 VP.n11032 VP.n10687 0.036
R5115 VP.n11032 VP.n11024 0.036
R5116 VP.n4305 VP.n4303 0.036
R5117 VP.n5210 VP.n5208 0.036
R5118 VP.n6075 VP.n6073 0.036
R5119 VP.n6939 VP.n6937 0.036
R5120 VP.n7777 VP.n7775 0.036
R5121 VP.n8616 VP.n8614 0.036
R5122 VP.n9415 VP.n9412 0.036
R5123 VP.n11002 VP.n10998 0.036
R5124 VP.n10943 VP.n10939 0.036
R5125 VP.n8741 VP.n8737 0.036
R5126 VP.n9548 VP.n9544 0.036
R5127 VP.n10892 VP.n10888 0.036
R5128 VP.n7018 VP.n7014 0.036
R5129 VP.n7856 VP.n7852 0.036
R5130 VP.n8693 VP.n8689 0.036
R5131 VP.n9497 VP.n9493 0.036
R5132 VP.n10841 VP.n10837 0.036
R5133 VP.n5239 VP.n5235 0.036
R5134 VP.n6105 VP.n6101 0.036
R5135 VP.n6969 VP.n6965 0.036
R5136 VP.n7807 VP.n7803 0.036
R5137 VP.n8645 VP.n8641 0.036
R5138 VP.n9446 VP.n9442 0.036
R5139 VP.n10790 VP.n10786 0.036
R5140 VP.n10725 VP.n10724 0.036
R5141 VP.n9380 VP.n9379 0.036
R5142 VP.n8585 VP.n8584 0.036
R5143 VP.n7746 VP.n7745 0.036
R5144 VP.n6907 VP.n6906 0.036
R5145 VP.n6043 VP.n6042 0.036
R5146 VP.n5179 VP.n5178 0.036
R5147 VP.n4273 VP.n4272 0.036
R5148 VP.n3352 VP.n3351 0.036
R5149 VP.n897 VP.n893 0.036
R5150 VP.n1331 VP.n1327 0.036
R5151 VP.n947 VP.n943 0.036
R5152 VP.n1459 VP.n1455 0.036
R5153 VP.n1884 VP.n1880 0.036
R5154 VP.n2307 VP.n2303 0.036
R5155 VP.n997 VP.n993 0.036
R5156 VP.n1497 VP.n1493 0.036
R5157 VP.n1936 VP.n1932 0.036
R5158 VP.n2559 VP.n2555 0.036
R5159 VP.n2865 VP.n2861 0.036
R5160 VP.n3257 VP.n3253 0.036
R5161 VP.n1047 VP.n1043 0.036
R5162 VP.n1535 VP.n1531 0.036
R5163 VP.n1988 VP.n1984 0.036
R5164 VP.n2521 VP.n2517 0.036
R5165 VP.n2917 VP.n2913 0.036
R5166 VP.n3437 VP.n3433 0.036
R5167 VP.n3810 VP.n3806 0.036
R5168 VP.n4178 VP.n4174 0.036
R5169 VP.n1097 VP.n1093 0.036
R5170 VP.n1573 VP.n1569 0.036
R5171 VP.n2040 VP.n2036 0.036
R5172 VP.n2483 VP.n2479 0.036
R5173 VP.n2969 VP.n2965 0.036
R5174 VP.n3475 VP.n3471 0.036
R5175 VP.n3862 VP.n3858 0.036
R5176 VP.n4354 VP.n4350 0.036
R5177 VP.n4745 VP.n4741 0.036
R5178 VP.n5084 VP.n5080 0.036
R5179 VP.n1147 VP.n1143 0.036
R5180 VP.n1611 VP.n1607 0.036
R5181 VP.n2092 VP.n2088 0.036
R5182 VP.n2451 VP.n2447 0.036
R5183 VP.n3021 VP.n3017 0.036
R5184 VP.n3513 VP.n3509 0.036
R5185 VP.n3914 VP.n3910 0.036
R5186 VP.n4392 VP.n4388 0.036
R5187 VP.n4797 VP.n4793 0.036
R5188 VP.n5314 VP.n5310 0.036
R5189 VP.n5634 VP.n5630 0.036
R5190 VP.n5948 VP.n5944 0.036
R5191 VP.n1185 VP.n1181 0.036
R5192 VP.n1643 VP.n1639 0.036
R5193 VP.n2133 VP.n2129 0.036
R5194 VP.n2419 VP.n2415 0.036
R5195 VP.n3062 VP.n3058 0.036
R5196 VP.n3545 VP.n3541 0.036
R5197 VP.n3955 VP.n3951 0.036
R5198 VP.n4424 VP.n4420 0.036
R5199 VP.n4838 VP.n4834 0.036
R5200 VP.n5346 VP.n5342 0.036
R5201 VP.n5675 VP.n5671 0.036
R5202 VP.n6174 VP.n6170 0.036
R5203 VP.n6519 VP.n6515 0.036
R5204 VP.n6812 VP.n6808 0.036
R5205 VP.n1225 VP.n1221 0.036
R5206 VP.n1675 VP.n1671 0.036
R5207 VP.n2174 VP.n2170 0.036
R5208 VP.n2387 VP.n2383 0.036
R5209 VP.n3103 VP.n3099 0.036
R5210 VP.n3577 VP.n3573 0.036
R5211 VP.n3996 VP.n3992 0.036
R5212 VP.n4456 VP.n4452 0.036
R5213 VP.n4879 VP.n4875 0.036
R5214 VP.n5378 VP.n5374 0.036
R5215 VP.n5716 VP.n5712 0.036
R5216 VP.n6206 VP.n6202 0.036
R5217 VP.n6560 VP.n6556 0.036
R5218 VP.n7093 VP.n7089 0.036
R5219 VP.n7372 VP.n7368 0.036
R5220 VP.n7651 VP.n7647 0.036
R5221 VP.n1266 VP.n1262 0.036
R5222 VP.n1707 VP.n1703 0.036
R5223 VP.n2215 VP.n2211 0.036
R5224 VP.n2355 VP.n2351 0.036
R5225 VP.n3144 VP.n3140 0.036
R5226 VP.n3609 VP.n3605 0.036
R5227 VP.n4037 VP.n4033 0.036
R5228 VP.n4488 VP.n4484 0.036
R5229 VP.n4920 VP.n4916 0.036
R5230 VP.n5410 VP.n5406 0.036
R5231 VP.n5757 VP.n5753 0.036
R5232 VP.n6238 VP.n6234 0.036
R5233 VP.n6601 VP.n6597 0.036
R5234 VP.n7125 VP.n7121 0.036
R5235 VP.n7413 VP.n7409 0.036
R5236 VP.n7925 VP.n7921 0.036
R5237 VP.n8229 VP.n8225 0.036
R5238 VP.n8490 VP.n8486 0.036
R5239 VP.n812 VP.n808 0.036
R5240 VP.n1362 VP.n1358 0.036
R5241 VP.n1798 VP.n1794 0.036
R5242 VP.n2679 VP.n2675 0.036
R5243 VP.n2758 VP.n2754 0.036
R5244 VP.n3288 VP.n3284 0.036
R5245 VP.n3698 VP.n3694 0.036
R5246 VP.n4209 VP.n4205 0.036
R5247 VP.n4607 VP.n4603 0.036
R5248 VP.n5115 VP.n5111 0.036
R5249 VP.n5499 VP.n5495 0.036
R5250 VP.n5979 VP.n5975 0.036
R5251 VP.n6355 VP.n6351 0.036
R5252 VP.n6843 VP.n6839 0.036
R5253 VP.n7214 VP.n7210 0.036
R5254 VP.n7682 VP.n7678 0.036
R5255 VP.n8042 VP.n8038 0.036
R5256 VP.n8521 VP.n8517 0.036
R5257 VP.n8886 VP.n8882 0.036
R5258 VP.n10601 VP.n10600 0.036
R5259 VP.n10566 VP.n10565 0.036
R5260 VP.n10531 VP.n10530 0.036
R5261 VP.n10496 VP.n10495 0.036
R5262 VP.n2589 VP.n2588 0.035
R5263 VP.n10127 VP.n10126 0.035
R5264 VP.n778 VP.n777 0.035
R5265 VP.n1767 VP.n1766 0.035
R5266 VP.n2728 VP.n2727 0.035
R5267 VP.n3668 VP.n3667 0.035
R5268 VP.n4574 VP.n4573 0.035
R5269 VP.n5469 VP.n5468 0.035
R5270 VP.n6325 VP.n6324 0.035
R5271 VP.n7184 VP.n7183 0.035
R5272 VP.n8012 VP.n8011 0.035
R5273 VP.n9687 VP.n9686 0.035
R5274 VP.n8846 VP.n8845 0.035
R5275 VP.n1910 VP.n1909 0.035
R5276 VP.n2891 VP.n2890 0.035
R5277 VP.n1962 VP.n1961 0.035
R5278 VP.n3836 VP.n3835 0.035
R5279 VP.n2943 VP.n2942 0.035
R5280 VP.n2014 VP.n2013 0.035
R5281 VP.n4771 VP.n4770 0.035
R5282 VP.n3888 VP.n3887 0.035
R5283 VP.n2995 VP.n2994 0.035
R5284 VP.n2066 VP.n2065 0.035
R5285 VP.n10069 VP.n10068 0.035
R5286 VP.n10025 VP.n10024 0.035
R5287 VP.n8431 VP.n8430 0.035
R5288 VP.n6753 VP.n6752 0.035
R5289 VP.n5025 VP.n5024 0.035
R5290 VP.n3186 VP.n3185 0.035
R5291 VP.n8760 VP.n8759 0.035
R5292 VP.n7037 VP.n7036 0.035
R5293 VP.n5258 VP.n5257 0.035
R5294 VP.t8 VP.n10354 0.035
R5295 VP.t8 VP.n10192 0.035
R5296 VP.t8 VP.n10328 0.035
R5297 VP.t8 VP.n10312 0.035
R5298 VP.t8 VP.n10296 0.035
R5299 VP.t8 VP.n10284 0.035
R5300 VP.t8 VP.n10268 0.035
R5301 VP.t8 VP.n10256 0.035
R5302 VP.t8 VP.n10240 0.035
R5303 VP.t8 VP.n10228 0.035
R5304 VP.t8 VP.n10212 0.035
R5305 VP.t8 VP.n10337 0.035
R5306 VP.t116 VP.n147 0.035
R5307 VP.t116 VP.n203 0.035
R5308 VP.t116 VP.n207 0.035
R5309 VP.t116 VP.n211 0.035
R5310 VP.t116 VP.n215 0.035
R5311 VP.t116 VP.n219 0.035
R5312 VP.t116 VP.n223 0.035
R5313 VP.t116 VP.n227 0.035
R5314 VP.t116 VP.n231 0.035
R5315 VP.t116 VP.n235 0.035
R5316 VP.t116 VP.n140 0.035
R5317 VP.t116 VP.n239 0.035
R5318 VP.n391 VP.n390 0.035
R5319 VP.n438 VP.n437 0.035
R5320 VP.n485 VP.n484 0.035
R5321 VP.n532 VP.n531 0.035
R5322 VP.n579 VP.n578 0.035
R5323 VP.n10639 VP.n10634 0.034
R5324 VP.n11034 VP.n11033 0.034
R5325 VP.n10113 VP.n9660 0.034
R5326 VP.n9043 VP.n9033 0.034
R5327 VP.n8763 VP.n8762 0.034
R5328 VP.n7348 VP.n7338 0.034
R5329 VP.n7040 VP.n7039 0.034
R5330 VP.n5610 VP.n5600 0.034
R5331 VP.n5261 VP.n5260 0.034
R5332 VP.n873 VP.n864 0.034
R5333 VP.n1400 VP.n1398 0.034
R5334 VP.n1403 VP.n1402 0.034
R5335 VP.n1860 VP.n1850 0.034
R5336 VP.n9719 VP.n9699 0.034
R5337 VP.n9343 VP.n9334 0.034
R5338 VP.n8918 VP.n8908 0.034
R5339 VP.n8549 VP.n8541 0.034
R5340 VP.n8074 VP.n8064 0.034
R5341 VP.n7710 VP.n7702 0.034
R5342 VP.n7246 VP.n7236 0.034
R5343 VP.n6871 VP.n6863 0.034
R5344 VP.n6387 VP.n6377 0.034
R5345 VP.n6007 VP.n5999 0.034
R5346 VP.n5531 VP.n5521 0.034
R5347 VP.n5143 VP.n5135 0.034
R5348 VP.n4636 VP.n4626 0.034
R5349 VP.n4237 VP.n4229 0.034
R5350 VP.n3730 VP.n3720 0.034
R5351 VP.n3316 VP.n3308 0.034
R5352 VP.n2790 VP.n2780 0.034
R5353 VP.n2651 VP.n2643 0.034
R5354 VP.n1830 VP.n1820 0.034
R5355 VP.n1390 VP.n1382 0.034
R5356 VP.n847 VP.n836 0.034
R5357 VP.n10429 VP.n10420 0.034
R5358 VP.n3378 VP.n3376 0.034
R5359 VP.n3381 VP.n3380 0.034
R5360 VP.n3781 VP.n3777 0.034
R5361 VP.n916 VP.n915 0.034
R5362 VP.n1903 VP.n1902 0.034
R5363 VP.n1907 VP.n1906 0.034
R5364 VP.n966 VP.n965 0.034
R5365 VP.n2884 VP.n2883 0.034
R5366 VP.n2888 VP.n2887 0.034
R5367 VP.n1955 VP.n1954 0.034
R5368 VP.n1959 VP.n1958 0.034
R5369 VP.n1016 VP.n1015 0.034
R5370 VP.n3829 VP.n3828 0.034
R5371 VP.n3833 VP.n3832 0.034
R5372 VP.n2936 VP.n2935 0.034
R5373 VP.n2940 VP.n2939 0.034
R5374 VP.n2007 VP.n2006 0.034
R5375 VP.n2011 VP.n2010 0.034
R5376 VP.n1066 VP.n1065 0.034
R5377 VP.n4764 VP.n4763 0.034
R5378 VP.n4768 VP.n4767 0.034
R5379 VP.n3881 VP.n3880 0.034
R5380 VP.n3885 VP.n3884 0.034
R5381 VP.n2988 VP.n2987 0.034
R5382 VP.n2992 VP.n2991 0.034
R5383 VP.n2059 VP.n2058 0.034
R5384 VP.n2063 VP.n2062 0.034
R5385 VP.n1116 VP.n1115 0.034
R5386 VP.n10394 VP.n10393 0.034
R5387 VP.n10377 VP.n10376 0.034
R5388 VP.n10360 VP.n10359 0.034
R5389 VP.n10157 VP.n10156 0.034
R5390 VP.t8 VP.n10353 0.034
R5391 VP.t8 VP.n10191 0.034
R5392 VP.t8 VP.n10327 0.034
R5393 VP.t8 VP.n10311 0.034
R5394 VP.t8 VP.n10295 0.034
R5395 VP.t8 VP.n10283 0.034
R5396 VP.t8 VP.n10267 0.034
R5397 VP.t8 VP.n10255 0.034
R5398 VP.t8 VP.n10239 0.034
R5399 VP.t8 VP.n10227 0.034
R5400 VP.t8 VP.n10211 0.034
R5401 VP.t8 VP.n10340 0.034
R5402 VP.t116 VP.n146 0.034
R5403 VP.t116 VP.n206 0.034
R5404 VP.t116 VP.n210 0.034
R5405 VP.t116 VP.n214 0.034
R5406 VP.t116 VP.n218 0.034
R5407 VP.t116 VP.n222 0.034
R5408 VP.t116 VP.n226 0.034
R5409 VP.t116 VP.n230 0.034
R5410 VP.t116 VP.n234 0.034
R5411 VP.t116 VP.n238 0.034
R5412 VP.t116 VP.n139 0.034
R5413 VP.t116 VP.n242 0.034
R5414 VP.n1424 VP.n1423 0.033
R5415 VP.n918 VP.n917 0.033
R5416 VP.n1905 VP.n1904 0.033
R5417 VP.n1476 VP.n1475 0.033
R5418 VP.n968 VP.n967 0.033
R5419 VP.n2886 VP.n2885 0.033
R5420 VP.n2576 VP.n2575 0.033
R5421 VP.n1957 VP.n1956 0.033
R5422 VP.n1514 VP.n1513 0.033
R5423 VP.n1018 VP.n1017 0.033
R5424 VP.n3831 VP.n3830 0.033
R5425 VP.n3454 VP.n3453 0.033
R5426 VP.n2938 VP.n2937 0.033
R5427 VP.n2538 VP.n2537 0.033
R5428 VP.n2009 VP.n2008 0.033
R5429 VP.n1552 VP.n1551 0.033
R5430 VP.n1068 VP.n1067 0.033
R5431 VP.n4766 VP.n4765 0.033
R5432 VP.n4371 VP.n4370 0.033
R5433 VP.n3883 VP.n3882 0.033
R5434 VP.n3492 VP.n3491 0.033
R5435 VP.n2990 VP.n2989 0.033
R5436 VP.n2500 VP.n2499 0.033
R5437 VP.n2061 VP.n2060 0.033
R5438 VP.n1590 VP.n1589 0.033
R5439 VP.n1118 VP.n1117 0.033
R5440 VP.n1318 VP.n1317 0.033
R5441 VP.n2294 VP.n2293 0.033
R5442 VP.n3244 VP.n3243 0.033
R5443 VP.n4165 VP.n4164 0.033
R5444 VP.n5071 VP.n5070 0.033
R5445 VP.n5935 VP.n5934 0.033
R5446 VP.n6799 VP.n6798 0.033
R5447 VP.n7638 VP.n7637 0.033
R5448 VP.n8477 VP.n8476 0.033
R5449 VP.n9683 VP.n9682 0.033
R5450 VP.n9304 VP.n9303 0.033
R5451 VP.n10674 VP.n10659 0.033
R5452 VP.n2833 VP.n2832 0.033
R5453 VP.n9319 VP.n9318 0.032
R5454 VP.n10135 VP.n10133 0.032
R5455 VP.n10623 VP.n10622 0.032
R5456 VP.n10585 VP.n10584 0.032
R5457 VP.n10550 VP.n10549 0.032
R5458 VP.n10515 VP.n10514 0.032
R5459 VP.n10480 VP.n10479 0.032
R5460 VP.n10440 VP.n10439 0.032
R5461 VP.n9968 VP.n9967 0.032
R5462 VP.n9211 VP.n9210 0.032
R5463 VP.n8411 VP.n8410 0.032
R5464 VP.n9920 VP.n9919 0.032
R5465 VP.n9161 VP.n9160 0.032
R5466 VP.n8362 VP.n8361 0.032
R5467 VP.n7545 VP.n7544 0.032
R5468 VP.n6733 VP.n6732 0.032
R5469 VP.n9872 VP.n9871 0.032
R5470 VP.n9111 VP.n9110 0.032
R5471 VP.n8313 VP.n8312 0.032
R5472 VP.n7496 VP.n7495 0.032
R5473 VP.n6684 VP.n6683 0.032
R5474 VP.n5842 VP.n5841 0.032
R5475 VP.n5005 VP.n5004 0.032
R5476 VP.n8858 VP.n8857 0.032
R5477 VP.n9711 VP.n9710 0.032
R5478 VP.n9852 VP.n9851 0.032
R5479 VP.n9090 VP.n9089 0.032
R5480 VP.n8293 VP.n8292 0.032
R5481 VP.n7476 VP.n7475 0.032
R5482 VP.n6664 VP.n6663 0.032
R5483 VP.n5821 VP.n5820 0.032
R5484 VP.n4984 VP.n4983 0.032
R5485 VP.n4101 VP.n4100 0.032
R5486 VP.n3209 VP.n3208 0.032
R5487 VP.n1404 VP.n1403 0.032
R5488 VP.n3382 VP.n3381 0.032
R5489 VP.t91 VP.n2589 0.031
R5490 VP.t6 VP.n10127 0.031
R5491 VP.t49 VP.n778 0.031
R5492 VP.t53 VP.n1767 0.031
R5493 VP.t108 VP.n2728 0.031
R5494 VP.t76 VP.n3668 0.031
R5495 VP.t169 VP.n4574 0.031
R5496 VP.t26 VP.n5469 0.031
R5497 VP.t159 VP.n6325 0.031
R5498 VP.t134 VP.n7184 0.031
R5499 VP.t18 VP.n8012 0.031
R5500 VP.t126 VP.n9687 0.031
R5501 VP.t207 VP.n8846 0.031
R5502 VP.n9317 VP.n9316 0.031
R5503 VP.n2841 VP.n2823 0.031
R5504 VP.n3391 VP.n3374 0.031
R5505 VP.n3786 VP.n3763 0.031
R5506 VP.n4310 VP.n4295 0.031
R5507 VP.n4685 VP.n4669 0.031
R5508 VP.n5215 VP.n5201 0.031
R5509 VP.n5580 VP.n5564 0.031
R5510 VP.n6080 VP.n6066 0.031
R5511 VP.n6436 VP.n6420 0.031
R5512 VP.n6944 VP.n6930 0.031
R5513 VP.n7295 VP.n7279 0.031
R5514 VP.n7782 VP.n7768 0.031
R5515 VP.n8123 VP.n8107 0.031
R5516 VP.n8621 VP.n8607 0.031
R5517 VP.n8967 VP.n8951 0.031
R5518 VP.n9420 VP.n9404 0.031
R5519 VP.n10758 VP.n10749 0.031
R5520 VP.n10164 VP.n10154 0.031
R5521 VP.n2329 VP.n2318 0.031
R5522 VP.n10202 VP.n10196 0.031
R5523 VP.n10322 VP.n10321 0.031
R5524 VP.n10304 VP.n10303 0.031
R5525 VP.n10276 VP.n10275 0.031
R5526 VP.n10248 VP.n10247 0.031
R5527 VP.n10220 VP.n10219 0.031
R5528 VP.n7903 VP.n7889 0.031
R5529 VP.n6152 VP.n6138 0.031
R5530 VP.n4332 VP.n4318 0.031
R5531 VP.n2606 VP.n2592 0.031
R5532 VP.n9632 VP.n9621 0.031
R5533 VP.n7967 VP.n7956 0.031
R5534 VP.n6280 VP.n6269 0.031
R5535 VP.n4529 VP.n4518 0.031
R5536 VP.n2823 VP.n2822 0.031
R5537 VP.n3374 VP.n3373 0.031
R5538 VP.n3763 VP.n3762 0.031
R5539 VP.n4295 VP.n4294 0.031
R5540 VP.n4669 VP.n4668 0.031
R5541 VP.n5201 VP.n5200 0.031
R5542 VP.n5564 VP.n5563 0.031
R5543 VP.n6066 VP.n6065 0.031
R5544 VP.n6420 VP.n6419 0.031
R5545 VP.n6930 VP.n6929 0.031
R5546 VP.n7279 VP.n7278 0.031
R5547 VP.n7768 VP.n7767 0.031
R5548 VP.n8107 VP.n8106 0.031
R5549 VP.n8607 VP.n8606 0.031
R5550 VP.n8951 VP.n8950 0.031
R5551 VP.n9404 VP.n9403 0.031
R5552 VP.n10749 VP.n10748 0.031
R5553 VP.n10154 VP.n10153 0.031
R5554 VP.n9310 VP.n9309 0.03
R5555 VP.n10642 VP.n10615 0.03
R5556 VP.n10642 VP.n10612 0.03
R5557 VP.n5652 VP.n5650 0.03
R5558 VP.n5652 VP.n5651 0.03
R5559 VP.n4815 VP.n4813 0.03
R5560 VP.n4815 VP.n4814 0.03
R5561 VP.n3932 VP.n3930 0.03
R5562 VP.n3932 VP.n3931 0.03
R5563 VP.n3039 VP.n3037 0.03
R5564 VP.n3039 VP.n3038 0.03
R5565 VP.n2110 VP.n2108 0.03
R5566 VP.n2110 VP.n2109 0.03
R5567 VP.n6537 VP.n6535 0.03
R5568 VP.n6537 VP.n6536 0.03
R5569 VP.n5693 VP.n5691 0.03
R5570 VP.n5693 VP.n5692 0.03
R5571 VP.n4856 VP.n4854 0.03
R5572 VP.n4856 VP.n4855 0.03
R5573 VP.n3973 VP.n3971 0.03
R5574 VP.n3973 VP.n3972 0.03
R5575 VP.n3080 VP.n3078 0.03
R5576 VP.n3080 VP.n3079 0.03
R5577 VP.n2151 VP.n2149 0.03
R5578 VP.n2151 VP.n2150 0.03
R5579 VP.n7390 VP.n7388 0.03
R5580 VP.n7390 VP.n7389 0.03
R5581 VP.n6578 VP.n6576 0.03
R5582 VP.n6578 VP.n6577 0.03
R5583 VP.n5734 VP.n5732 0.03
R5584 VP.n5734 VP.n5733 0.03
R5585 VP.n4897 VP.n4895 0.03
R5586 VP.n4897 VP.n4896 0.03
R5587 VP.n4014 VP.n4012 0.03
R5588 VP.n4014 VP.n4013 0.03
R5589 VP.n3121 VP.n3119 0.03
R5590 VP.n3121 VP.n3120 0.03
R5591 VP.n2192 VP.n2190 0.03
R5592 VP.n2192 VP.n2191 0.03
R5593 VP.n1243 VP.n1241 0.03
R5594 VP.n1243 VP.n1242 0.03
R5595 VP.n1284 VP.n1282 0.03
R5596 VP.n1284 VP.n1283 0.03
R5597 VP.n8247 VP.n8245 0.03
R5598 VP.n8247 VP.n8246 0.03
R5599 VP.n7431 VP.n7429 0.03
R5600 VP.n7431 VP.n7430 0.03
R5601 VP.n6619 VP.n6617 0.03
R5602 VP.n6619 VP.n6618 0.03
R5603 VP.n5775 VP.n5773 0.03
R5604 VP.n5775 VP.n5774 0.03
R5605 VP.n4938 VP.n4936 0.03
R5606 VP.n4938 VP.n4937 0.03
R5607 VP.n4055 VP.n4053 0.03
R5608 VP.n4055 VP.n4054 0.03
R5609 VP.n3162 VP.n3160 0.03
R5610 VP.n3162 VP.n3161 0.03
R5611 VP.n2233 VP.n2231 0.03
R5612 VP.n2233 VP.n2232 0.03
R5613 VP.n8957 VP.n8953 0.029
R5614 VP.n8113 VP.n8109 0.029
R5615 VP.n7285 VP.n7281 0.029
R5616 VP.n6426 VP.n6422 0.029
R5617 VP.n5570 VP.n5566 0.029
R5618 VP.n4675 VP.n4671 0.029
R5619 VP.n9797 VP.n9793 0.029
R5620 VP.n9775 VP.n9771 0.029
R5621 VP.n9002 VP.n8998 0.029
R5622 VP.n8158 VP.n8154 0.029
R5623 VP.n9753 VP.n9749 0.029
R5624 VP.n8979 VP.n8975 0.029
R5625 VP.n8135 VP.n8131 0.029
R5626 VP.n7307 VP.n7303 0.029
R5627 VP.n6448 VP.n6444 0.029
R5628 VP.n9731 VP.n9727 0.029
R5629 VP.n8930 VP.n8926 0.029
R5630 VP.n8086 VP.n8082 0.029
R5631 VP.n7258 VP.n7254 0.029
R5632 VP.n6399 VP.n6395 0.029
R5633 VP.n5543 VP.n5539 0.029
R5634 VP.n4648 VP.n4644 0.029
R5635 VP.n3742 VP.n3738 0.029
R5636 VP.n2802 VP.n2798 0.029
R5637 VP.n761 VP.n760 0.029
R5638 VP.n1750 VP.n1749 0.029
R5639 VP.n2711 VP.n2710 0.029
R5640 VP.n3651 VP.n3650 0.029
R5641 VP.n4557 VP.n4556 0.029
R5642 VP.n5452 VP.n5451 0.029
R5643 VP.n6308 VP.n6307 0.029
R5644 VP.n7167 VP.n7166 0.029
R5645 VP.n7995 VP.n7994 0.029
R5646 VP.n8829 VP.n8828 0.029
R5647 VP.n10105 VP.n10104 0.029
R5648 VP.n2832 VP.n2831 0.029
R5649 VP.n9798 VP.n9797 0.029
R5650 VP.n8159 VP.n8158 0.029
R5651 VP.n9003 VP.n9002 0.029
R5652 VP.n9776 VP.n9775 0.029
R5653 VP.n6449 VP.n6448 0.029
R5654 VP.n7308 VP.n7307 0.029
R5655 VP.n8136 VP.n8135 0.029
R5656 VP.n8980 VP.n8979 0.029
R5657 VP.n9754 VP.n9753 0.029
R5658 VP.n2803 VP.n2802 0.029
R5659 VP.n3743 VP.n3742 0.029
R5660 VP.n4649 VP.n4648 0.029
R5661 VP.n5544 VP.n5543 0.029
R5662 VP.n6400 VP.n6399 0.029
R5663 VP.n7259 VP.n7258 0.029
R5664 VP.n8087 VP.n8086 0.029
R5665 VP.n8931 VP.n8930 0.029
R5666 VP.n9732 VP.n9731 0.029
R5667 VP.n4676 VP.n4675 0.029
R5668 VP.n5571 VP.n5570 0.029
R5669 VP.n6427 VP.n6426 0.029
R5670 VP.n7286 VP.n7285 0.029
R5671 VP.n8114 VP.n8113 0.029
R5672 VP.n8958 VP.n8957 0.029
R5673 VP.n9029 VP.n9028 0.029
R5674 VP.n7334 VP.n7333 0.029
R5675 VP.n5596 VP.n5595 0.029
R5676 VP.n860 VP.n859 0.029
R5677 VP.n1846 VP.n1845 0.029
R5678 VP.n3773 VP.n3772 0.029
R5679 VP.n10599 VP.n10598 0.028
R5680 VP.n8185 VP.n8178 0.028
R5681 VP.n7908 VP.n7904 0.028
R5682 VP.n10564 VP.n10563 0.028
R5683 VP.n6475 VP.n6468 0.028
R5684 VP.n6157 VP.n6153 0.028
R5685 VP.n10529 VP.n10528 0.028
R5686 VP.n4701 VP.n4694 0.028
R5687 VP.n4337 VP.n4333 0.028
R5688 VP.n10494 VP.n10493 0.028
R5689 VP.n308 VP.n306 0.028
R5690 VP.n8182 VP.n8181 0.028
R5691 VP.n6472 VP.n6471 0.028
R5692 VP.n4698 VP.n4697 0.028
R5693 VP.n378 VP.n377 0.028
R5694 VP.n425 VP.n424 0.028
R5695 VP.n472 VP.n471 0.028
R5696 VP.n519 VP.n518 0.028
R5697 VP.n566 VP.n565 0.028
R5698 VP.n155 VP.n154 0.028
R5699 VP.n10090 VP.n10087 0.028
R5700 VP.n10057 VP.n10056 0.027
R5701 VP.n10987 VP.n10986 0.027
R5702 VP.n9270 VP.n9269 0.027
R5703 VP.n9630 VP.n9629 0.027
R5704 VP.n10037 VP.n10036 0.027
R5705 VP.n10928 VP.n10927 0.027
R5706 VP.n7604 VP.n7603 0.027
R5707 VP.n7965 VP.n7964 0.027
R5708 VP.n8443 VP.n8442 0.027
R5709 VP.n9241 VP.n9240 0.027
R5710 VP.n9538 VP.n9537 0.027
R5711 VP.n9997 VP.n9996 0.027
R5712 VP.n10877 VP.n10876 0.027
R5713 VP.n5901 VP.n5900 0.027
R5714 VP.n6278 VP.n6277 0.027
R5715 VP.n6765 VP.n6764 0.027
R5716 VP.n7575 VP.n7574 0.027
R5717 VP.n8392 VP.n8391 0.027
R5718 VP.n9191 VP.n9190 0.027
R5719 VP.n9487 VP.n9486 0.027
R5720 VP.n9949 VP.n9948 0.027
R5721 VP.n10826 VP.n10825 0.027
R5722 VP.n4131 VP.n4130 0.027
R5723 VP.n4527 VP.n4526 0.027
R5724 VP.n5037 VP.n5036 0.027
R5725 VP.n5872 VP.n5871 0.027
R5726 VP.n6714 VP.n6713 0.027
R5727 VP.n7526 VP.n7525 0.027
R5728 VP.n8343 VP.n8342 0.027
R5729 VP.n9141 VP.n9140 0.027
R5730 VP.n9436 VP.n9435 0.027
R5731 VP.n9901 VP.n9900 0.027
R5732 VP.n10775 VP.n10774 0.027
R5733 VP.n10729 VP.n10728 0.027
R5734 VP.n9824 VP.n9822 0.027
R5735 VP.n9384 VP.n9383 0.027
R5736 VP.n9060 VP.n9058 0.027
R5737 VP.n8263 VP.n8261 0.027
R5738 VP.n7447 VP.n7445 0.027
R5739 VP.n6635 VP.n6633 0.027
R5740 VP.n5791 VP.n5789 0.027
R5741 VP.n4954 VP.n4952 0.027
R5742 VP.n4071 VP.n4069 0.027
R5743 VP.n3178 VP.n3176 0.027
R5744 VP.n2321 VP.n2320 0.027
R5745 VP.n10700 VP.n10699 0.027
R5746 VP.n263 VP.n262 0.027
R5747 VP.n365 VP.n364 0.027
R5748 VP.n902 VP.n901 0.027
R5749 VP.n1336 VP.n1335 0.027
R5750 VP.n412 VP.n411 0.027
R5751 VP.n952 VP.n951 0.027
R5752 VP.n1464 VP.n1463 0.027
R5753 VP.n1889 VP.n1888 0.027
R5754 VP.n2312 VP.n2311 0.027
R5755 VP.n459 VP.n458 0.027
R5756 VP.n1002 VP.n1001 0.027
R5757 VP.n1502 VP.n1501 0.027
R5758 VP.n1941 VP.n1940 0.027
R5759 VP.n2564 VP.n2563 0.027
R5760 VP.n2870 VP.n2869 0.027
R5761 VP.n3262 VP.n3261 0.027
R5762 VP.n506 VP.n505 0.027
R5763 VP.n1052 VP.n1051 0.027
R5764 VP.n1540 VP.n1539 0.027
R5765 VP.n1993 VP.n1992 0.027
R5766 VP.n2526 VP.n2525 0.027
R5767 VP.n2922 VP.n2921 0.027
R5768 VP.n3442 VP.n3441 0.027
R5769 VP.n3815 VP.n3814 0.027
R5770 VP.n4183 VP.n4182 0.027
R5771 VP.n553 VP.n552 0.027
R5772 VP.n1102 VP.n1101 0.027
R5773 VP.n1578 VP.n1577 0.027
R5774 VP.n2045 VP.n2044 0.027
R5775 VP.n2488 VP.n2487 0.027
R5776 VP.n2974 VP.n2973 0.027
R5777 VP.n3480 VP.n3479 0.027
R5778 VP.n3867 VP.n3866 0.027
R5779 VP.n4359 VP.n4358 0.027
R5780 VP.n4750 VP.n4749 0.027
R5781 VP.n5089 VP.n5088 0.027
R5782 VP.n600 VP.n599 0.027
R5783 VP.n1152 VP.n1151 0.027
R5784 VP.n1616 VP.n1615 0.027
R5785 VP.n2097 VP.n2096 0.027
R5786 VP.n2456 VP.n2455 0.027
R5787 VP.n3026 VP.n3025 0.027
R5788 VP.n3518 VP.n3517 0.027
R5789 VP.n3919 VP.n3918 0.027
R5790 VP.n4397 VP.n4396 0.027
R5791 VP.n4802 VP.n4801 0.027
R5792 VP.n5319 VP.n5318 0.027
R5793 VP.n5639 VP.n5638 0.027
R5794 VP.n5953 VP.n5952 0.027
R5795 VP.n640 VP.n639 0.027
R5796 VP.n1190 VP.n1189 0.027
R5797 VP.n1648 VP.n1647 0.027
R5798 VP.n2138 VP.n2137 0.027
R5799 VP.n2424 VP.n2423 0.027
R5800 VP.n3067 VP.n3066 0.027
R5801 VP.n3550 VP.n3549 0.027
R5802 VP.n3960 VP.n3959 0.027
R5803 VP.n4429 VP.n4428 0.027
R5804 VP.n4843 VP.n4842 0.027
R5805 VP.n5351 VP.n5350 0.027
R5806 VP.n5680 VP.n5679 0.027
R5807 VP.n6179 VP.n6178 0.027
R5808 VP.n6524 VP.n6523 0.027
R5809 VP.n6817 VP.n6816 0.027
R5810 VP.n670 VP.n669 0.027
R5811 VP.n1230 VP.n1229 0.027
R5812 VP.n1680 VP.n1679 0.027
R5813 VP.n2179 VP.n2178 0.027
R5814 VP.n2392 VP.n2391 0.027
R5815 VP.n3108 VP.n3107 0.027
R5816 VP.n3582 VP.n3581 0.027
R5817 VP.n4001 VP.n4000 0.027
R5818 VP.n4461 VP.n4460 0.027
R5819 VP.n4884 VP.n4883 0.027
R5820 VP.n5383 VP.n5382 0.027
R5821 VP.n5721 VP.n5720 0.027
R5822 VP.n6211 VP.n6210 0.027
R5823 VP.n6565 VP.n6564 0.027
R5824 VP.n7098 VP.n7097 0.027
R5825 VP.n7377 VP.n7376 0.027
R5826 VP.n7656 VP.n7655 0.027
R5827 VP.n9651 VP.n9649 0.027
R5828 VP.n702 VP.n701 0.027
R5829 VP.n1271 VP.n1270 0.027
R5830 VP.n1712 VP.n1711 0.027
R5831 VP.n2220 VP.n2219 0.027
R5832 VP.n2360 VP.n2359 0.027
R5833 VP.n3149 VP.n3148 0.027
R5834 VP.n3614 VP.n3613 0.027
R5835 VP.n4042 VP.n4041 0.027
R5836 VP.n4493 VP.n4492 0.027
R5837 VP.n4925 VP.n4924 0.027
R5838 VP.n5415 VP.n5414 0.027
R5839 VP.n5762 VP.n5761 0.027
R5840 VP.n6243 VP.n6242 0.027
R5841 VP.n6606 VP.n6605 0.027
R5842 VP.n7130 VP.n7129 0.027
R5843 VP.n7418 VP.n7417 0.027
R5844 VP.n7930 VP.n7929 0.027
R5845 VP.n8234 VP.n8233 0.027
R5846 VP.n8495 VP.n8494 0.027
R5847 VP.n8817 VP.n8815 0.027
R5848 VP.n278 VP.n277 0.027
R5849 VP.n794 VP.n793 0.027
R5850 VP.n1350 VP.n1349 0.027
R5851 VP.n1780 VP.n1779 0.027
R5852 VP.n2667 VP.n2666 0.027
R5853 VP.n2740 VP.n2739 0.027
R5854 VP.n3276 VP.n3275 0.027
R5855 VP.n3680 VP.n3679 0.027
R5856 VP.n4197 VP.n4196 0.027
R5857 VP.n4589 VP.n4588 0.027
R5858 VP.n5103 VP.n5102 0.027
R5859 VP.n5481 VP.n5480 0.027
R5860 VP.n5967 VP.n5966 0.027
R5861 VP.n6337 VP.n6336 0.027
R5862 VP.n6831 VP.n6830 0.027
R5863 VP.n7196 VP.n7195 0.027
R5864 VP.n7670 VP.n7669 0.027
R5865 VP.n8024 VP.n8023 0.027
R5866 VP.n8509 VP.n8508 0.027
R5867 VP.n8870 VP.n8869 0.027
R5868 VP.n11023 VP.n11022 0.027
R5869 VP.n7940 VP.n7939 0.027
R5870 VP.n7140 VP.n7139 0.027
R5871 VP.n6253 VP.n6252 0.027
R5872 VP.n5425 VP.n5424 0.027
R5873 VP.n4503 VP.n4502 0.027
R5874 VP.n3624 VP.n3623 0.027
R5875 VP.n2370 VP.n2369 0.027
R5876 VP.n10680 VP.n10679 0.027
R5877 VP.n8184 VP.n8183 0.027
R5878 VP.n6474 VP.n6473 0.027
R5879 VP.n4700 VP.n4699 0.027
R5880 VP.n10090 VP.n10089 0.027
R5881 VP.t116 VP.n199 0.026
R5882 VP.n2261 VP.n2251 0.026
R5883 VP.n1746 VP.n1741 0.026
R5884 VP.n923 VP.n912 0.026
R5885 VP.n2707 VP.n2702 0.026
R5886 VP.n1912 VP.n1899 0.026
R5887 VP.n1479 VP.n1474 0.026
R5888 VP.n973 VP.n962 0.026
R5889 VP.n3647 VP.n3642 0.026
R5890 VP.n2893 VP.n2880 0.026
R5891 VP.n2579 VP.n2574 0.026
R5892 VP.n1964 VP.n1951 0.026
R5893 VP.n1517 VP.n1512 0.026
R5894 VP.n1023 VP.n1012 0.026
R5895 VP.n4553 VP.n4548 0.026
R5896 VP.n3838 VP.n3825 0.026
R5897 VP.n3457 VP.n3452 0.026
R5898 VP.n2945 VP.n2932 0.026
R5899 VP.n2541 VP.n2536 0.026
R5900 VP.n2016 VP.n2003 0.026
R5901 VP.n1555 VP.n1550 0.026
R5902 VP.n1073 VP.n1062 0.026
R5903 VP.n5448 VP.n5443 0.026
R5904 VP.n4773 VP.n4760 0.026
R5905 VP.n4374 VP.n4369 0.026
R5906 VP.n3890 VP.n3877 0.026
R5907 VP.n3495 VP.n3490 0.026
R5908 VP.n2997 VP.n2984 0.026
R5909 VP.n2503 VP.n2498 0.026
R5910 VP.n2068 VP.n2055 0.026
R5911 VP.n1593 VP.n1588 0.026
R5912 VP.n1123 VP.n1112 0.026
R5913 VP.n6304 VP.n6299 0.026
R5914 VP.n7163 VP.n7158 0.026
R5915 VP.n7991 VP.n7986 0.026
R5916 VP.n10023 VP.n10022 0.025
R5917 VP.n8429 VP.n8428 0.025
R5918 VP.n9229 VP.n9228 0.025
R5919 VP.n9986 VP.n9985 0.025
R5920 VP.n6751 VP.n6750 0.025
R5921 VP.n7563 VP.n7562 0.025
R5922 VP.n8380 VP.n8379 0.025
R5923 VP.n9179 VP.n9178 0.025
R5924 VP.n9938 VP.n9937 0.025
R5925 VP.n5023 VP.n5022 0.025
R5926 VP.n5860 VP.n5859 0.025
R5927 VP.n6702 VP.n6701 0.025
R5928 VP.n7514 VP.n7513 0.025
R5929 VP.n8331 VP.n8330 0.025
R5930 VP.n9129 VP.n9128 0.025
R5931 VP.n9890 VP.n9889 0.025
R5932 VP.n8205 VP.n8196 0.025
R5933 VP.n6495 VP.n6486 0.025
R5934 VP.n4721 VP.n4712 0.025
R5935 VP.n2836 VP.n2833 0.025
R5936 VP.n9797 VP.n9796 0.025
R5937 VP.n8158 VP.n8157 0.025
R5938 VP.n9002 VP.n9001 0.025
R5939 VP.n9775 VP.n9774 0.025
R5940 VP.n6448 VP.n6447 0.025
R5941 VP.n7307 VP.n7306 0.025
R5942 VP.n8135 VP.n8134 0.025
R5943 VP.n8979 VP.n8978 0.025
R5944 VP.n9753 VP.n9752 0.025
R5945 VP.n2802 VP.n2801 0.025
R5946 VP.n3742 VP.n3741 0.025
R5947 VP.n4648 VP.n4647 0.025
R5948 VP.n5543 VP.n5542 0.025
R5949 VP.n6399 VP.n6398 0.025
R5950 VP.n7258 VP.n7257 0.025
R5951 VP.n8086 VP.n8085 0.025
R5952 VP.n8930 VP.n8929 0.025
R5953 VP.n9731 VP.n9730 0.025
R5954 VP.n4675 VP.n4674 0.025
R5955 VP.n5570 VP.n5569 0.025
R5956 VP.n6426 VP.n6425 0.025
R5957 VP.n7285 VP.n7284 0.025
R5958 VP.n8113 VP.n8112 0.025
R5959 VP.n8957 VP.n8956 0.025
R5960 VP.n10455 VP.n10438 0.025
R5961 VP.n9664 VP.n9663 0.024
R5962 VP.n9285 VP.n9284 0.024
R5963 VP.n8458 VP.n8457 0.024
R5964 VP.n7619 VP.n7618 0.024
R5965 VP.n6780 VP.n6779 0.024
R5966 VP.n5916 VP.n5915 0.024
R5967 VP.n5052 VP.n5051 0.024
R5968 VP.n4146 VP.n4145 0.024
R5969 VP.n3225 VP.n3224 0.024
R5970 VP.n2275 VP.n2274 0.024
R5971 VP.n1298 VP.n1297 0.024
R5972 VP.n10448 VP.n10447 0.024
R5973 VP.n9829 VP.n9828 0.024
R5974 VP.n9066 VP.n9065 0.024
R5975 VP.n8269 VP.n8268 0.024
R5976 VP.n7453 VP.n7452 0.024
R5977 VP.n6641 VP.n6640 0.024
R5978 VP.n5797 VP.n5796 0.024
R5979 VP.n4960 VP.n4959 0.024
R5980 VP.n4077 VP.n4076 0.024
R5981 VP.n3184 VP.n3183 0.024
R5982 VP.n255 VP.n254 0.024
R5983 VP.n357 VP.n356 0.024
R5984 VP.n404 VP.n403 0.024
R5985 VP.n451 VP.n450 0.024
R5986 VP.n498 VP.n497 0.024
R5987 VP.n545 VP.n544 0.024
R5988 VP.n592 VP.n591 0.024
R5989 VP.n632 VP.n631 0.024
R5990 VP.n662 VP.n661 0.024
R5991 VP.n694 VP.n693 0.024
R5992 VP.n11000 VP.n10999 0.024
R5993 VP.n10636 VP.n10635 0.024
R5994 VP.n10029 VP.n10028 0.024
R5995 VP.n10941 VP.n10940 0.024
R5996 VP.n10594 VP.n10593 0.024
R5997 VP.n8760 VP.n8758 0.024
R5998 VP.n8435 VP.n8434 0.024
R5999 VP.n8739 VP.n8738 0.024
R6000 VP.n9546 VP.n9545 0.024
R6001 VP.n10890 VP.n10889 0.024
R6002 VP.n10559 VP.n10558 0.024
R6003 VP.n7037 VP.n7035 0.024
R6004 VP.n6757 VP.n6756 0.024
R6005 VP.n7016 VP.n7015 0.024
R6006 VP.n7854 VP.n7853 0.024
R6007 VP.n8691 VP.n8690 0.024
R6008 VP.n9495 VP.n9494 0.024
R6009 VP.n10839 VP.n10838 0.024
R6010 VP.n10524 VP.n10523 0.024
R6011 VP.n5258 VP.n5256 0.024
R6012 VP.n5029 VP.n5028 0.024
R6013 VP.n5237 VP.n5236 0.024
R6014 VP.n6103 VP.n6102 0.024
R6015 VP.n6967 VP.n6966 0.024
R6016 VP.n7805 VP.n7804 0.024
R6017 VP.n8643 VP.n8642 0.024
R6018 VP.n9444 VP.n9443 0.024
R6019 VP.n10788 VP.n10787 0.024
R6020 VP.n10489 VP.n10488 0.024
R6021 VP.n10721 VP.n10720 0.024
R6022 VP.n9376 VP.n9375 0.024
R6023 VP.n8581 VP.n8580 0.024
R6024 VP.n7742 VP.n7741 0.024
R6025 VP.n6903 VP.n6902 0.024
R6026 VP.n6039 VP.n6038 0.024
R6027 VP.n5175 VP.n5174 0.024
R6028 VP.n4269 VP.n4268 0.024
R6029 VP.n3348 VP.n3347 0.024
R6030 VP.n3181 VP.n3180 0.024
R6031 VP.n1400 VP.n1399 0.024
R6032 VP.n10131 VP.n10130 0.024
R6033 VP.n309 VP.n308 0.024
R6034 VP.n1309 VP.n1308 0.024
R6035 VP.n740 VP.n739 0.024
R6036 VP.n768 VP.n767 0.024
R6037 VP.n2286 VP.n2285 0.024
R6038 VP.n383 VP.n382 0.024
R6039 VP.n895 VP.n894 0.024
R6040 VP.n1329 VP.n1328 0.024
R6041 VP.n1757 VP.n1756 0.024
R6042 VP.n3236 VP.n3235 0.024
R6043 VP.n430 VP.n429 0.024
R6044 VP.n945 VP.n944 0.024
R6045 VP.n1457 VP.n1456 0.024
R6046 VP.n1882 VP.n1881 0.024
R6047 VP.n2305 VP.n2304 0.024
R6048 VP.n2718 VP.n2717 0.024
R6049 VP.n4157 VP.n4156 0.024
R6050 VP.n477 VP.n476 0.024
R6051 VP.n995 VP.n994 0.024
R6052 VP.n1495 VP.n1494 0.024
R6053 VP.n1934 VP.n1933 0.024
R6054 VP.n2557 VP.n2556 0.024
R6055 VP.n2863 VP.n2862 0.024
R6056 VP.n3255 VP.n3254 0.024
R6057 VP.n3658 VP.n3657 0.024
R6058 VP.n5063 VP.n5062 0.024
R6059 VP.n524 VP.n523 0.024
R6060 VP.n1045 VP.n1044 0.024
R6061 VP.n1533 VP.n1532 0.024
R6062 VP.n1986 VP.n1985 0.024
R6063 VP.n2519 VP.n2518 0.024
R6064 VP.n2915 VP.n2914 0.024
R6065 VP.n3435 VP.n3434 0.024
R6066 VP.n3808 VP.n3807 0.024
R6067 VP.n4176 VP.n4175 0.024
R6068 VP.n4564 VP.n4563 0.024
R6069 VP.n5927 VP.n5926 0.024
R6070 VP.n571 VP.n570 0.024
R6071 VP.n1095 VP.n1094 0.024
R6072 VP.n1571 VP.n1570 0.024
R6073 VP.n2038 VP.n2037 0.024
R6074 VP.n2481 VP.n2480 0.024
R6075 VP.n2967 VP.n2966 0.024
R6076 VP.n3473 VP.n3472 0.024
R6077 VP.n3860 VP.n3859 0.024
R6078 VP.n4352 VP.n4351 0.024
R6079 VP.n4743 VP.n4742 0.024
R6080 VP.n5082 VP.n5081 0.024
R6081 VP.n5459 VP.n5458 0.024
R6082 VP.n6791 VP.n6790 0.024
R6083 VP.n611 VP.n610 0.024
R6084 VP.n1145 VP.n1144 0.024
R6085 VP.n1609 VP.n1608 0.024
R6086 VP.n2090 VP.n2089 0.024
R6087 VP.n2449 VP.n2448 0.024
R6088 VP.n3019 VP.n3018 0.024
R6089 VP.n3511 VP.n3510 0.024
R6090 VP.n3912 VP.n3911 0.024
R6091 VP.n4390 VP.n4389 0.024
R6092 VP.n4795 VP.n4794 0.024
R6093 VP.n5312 VP.n5311 0.024
R6094 VP.n5632 VP.n5631 0.024
R6095 VP.n5946 VP.n5945 0.024
R6096 VP.n6315 VP.n6314 0.024
R6097 VP.n7630 VP.n7629 0.024
R6098 VP.n1183 VP.n1182 0.024
R6099 VP.n1641 VP.n1640 0.024
R6100 VP.n2131 VP.n2130 0.024
R6101 VP.n2417 VP.n2416 0.024
R6102 VP.n3060 VP.n3059 0.024
R6103 VP.n3543 VP.n3542 0.024
R6104 VP.n3953 VP.n3952 0.024
R6105 VP.n4422 VP.n4421 0.024
R6106 VP.n4836 VP.n4835 0.024
R6107 VP.n5344 VP.n5343 0.024
R6108 VP.n5673 VP.n5672 0.024
R6109 VP.n6172 VP.n6171 0.024
R6110 VP.n6517 VP.n6516 0.024
R6111 VP.n6810 VP.n6809 0.024
R6112 VP.n7174 VP.n7173 0.024
R6113 VP.n8469 VP.n8468 0.024
R6114 VP.n1223 VP.n1222 0.024
R6115 VP.n1673 VP.n1672 0.024
R6116 VP.n2172 VP.n2171 0.024
R6117 VP.n2385 VP.n2384 0.024
R6118 VP.n3101 VP.n3100 0.024
R6119 VP.n3575 VP.n3574 0.024
R6120 VP.n3994 VP.n3993 0.024
R6121 VP.n4454 VP.n4453 0.024
R6122 VP.n4877 VP.n4876 0.024
R6123 VP.n5376 VP.n5375 0.024
R6124 VP.n5714 VP.n5713 0.024
R6125 VP.n6204 VP.n6203 0.024
R6126 VP.n6558 VP.n6557 0.024
R6127 VP.n7091 VP.n7090 0.024
R6128 VP.n7370 VP.n7369 0.024
R6129 VP.n7649 VP.n7648 0.024
R6130 VP.n8002 VP.n8001 0.024
R6131 VP.n9675 VP.n9674 0.024
R6132 VP.n713 VP.n712 0.024
R6133 VP.n1264 VP.n1263 0.024
R6134 VP.n1705 VP.n1704 0.024
R6135 VP.n2213 VP.n2212 0.024
R6136 VP.n2353 VP.n2352 0.024
R6137 VP.n3142 VP.n3141 0.024
R6138 VP.n3607 VP.n3606 0.024
R6139 VP.n4035 VP.n4034 0.024
R6140 VP.n4486 VP.n4485 0.024
R6141 VP.n4918 VP.n4917 0.024
R6142 VP.n5408 VP.n5407 0.024
R6143 VP.n5755 VP.n5754 0.024
R6144 VP.n6236 VP.n6235 0.024
R6145 VP.n6599 VP.n6598 0.024
R6146 VP.n7123 VP.n7122 0.024
R6147 VP.n7411 VP.n7410 0.024
R6148 VP.n7923 VP.n7922 0.024
R6149 VP.n8227 VP.n8226 0.024
R6150 VP.n8488 VP.n8487 0.024
R6151 VP.n8836 VP.n8835 0.024
R6152 VP.n9296 VP.n9295 0.024
R6153 VP.n810 VP.n809 0.024
R6154 VP.n1360 VP.n1359 0.024
R6155 VP.n1796 VP.n1795 0.024
R6156 VP.n2677 VP.n2676 0.024
R6157 VP.n2756 VP.n2755 0.024
R6158 VP.n3286 VP.n3285 0.024
R6159 VP.n3696 VP.n3695 0.024
R6160 VP.n4207 VP.n4206 0.024
R6161 VP.n4605 VP.n4604 0.024
R6162 VP.n5113 VP.n5112 0.024
R6163 VP.n5497 VP.n5496 0.024
R6164 VP.n5977 VP.n5976 0.024
R6165 VP.n6353 VP.n6352 0.024
R6166 VP.n6841 VP.n6840 0.024
R6167 VP.n7212 VP.n7211 0.024
R6168 VP.n7680 VP.n7679 0.024
R6169 VP.n8040 VP.n8039 0.024
R6170 VP.n8519 VP.n8518 0.024
R6171 VP.n8884 VP.n8883 0.024
R6172 VP.n9315 VP.n9314 0.024
R6173 VP.n10657 VP.n10656 0.024
R6174 VP.n3378 VP.n3377 0.024
R6175 VP.n10626 VP.n10625 0.024
R6176 VP.n10588 VP.n10587 0.024
R6177 VP.n10553 VP.n10552 0.024
R6178 VP.n10518 VP.n10517 0.024
R6179 VP.n10483 VP.n10482 0.024
R6180 VP.n10443 VP.n10442 0.024
R6181 VP.n10686 VP.n10685 0.024
R6182 VP.n10965 VP.n10960 0.024
R6183 VP.n9590 VP.n9585 0.024
R6184 VP.n8786 VP.n8781 0.024
R6185 VP.n7899 VP.n7894 0.024
R6186 VP.n7063 VP.n7058 0.024
R6187 VP.n6148 VP.n6143 0.024
R6188 VP.n5284 VP.n5279 0.024
R6189 VP.n4328 VP.n4323 0.024
R6190 VP.n3407 VP.n3402 0.024
R6191 VP.n2602 VP.n2597 0.024
R6192 VP.n1436 VP.n1431 0.024
R6193 VP.n338 VP.n332 0.024
R6194 VP.n1319 VP.n772 0.024
R6195 VP.n2295 VP.n1761 0.024
R6196 VP.n3245 VP.n2722 0.024
R6197 VP.n4166 VP.n3662 0.024
R6198 VP.n5072 VP.n4568 0.024
R6199 VP.n5936 VP.n5463 0.024
R6200 VP.n6800 VP.n6319 0.024
R6201 VP.n7639 VP.n7178 0.024
R6202 VP.n8478 VP.n8006 0.024
R6203 VP.n9305 VP.n8840 0.024
R6204 VP.n10112 VP.n10111 0.024
R6205 VP.n10675 VP.n10121 0.024
R6206 VP.n10671 VP.n10667 0.024
R6207 VP.n9671 VP.n9667 0.024
R6208 VP.n9292 VP.n9288 0.024
R6209 VP.n8465 VP.n8461 0.024
R6210 VP.n7626 VP.n7622 0.024
R6211 VP.n6787 VP.n6783 0.024
R6212 VP.n5923 VP.n5919 0.024
R6213 VP.n5059 VP.n5055 0.024
R6214 VP.n4153 VP.n4149 0.024
R6215 VP.n3232 VP.n3228 0.024
R6216 VP.n2282 VP.n2278 0.024
R6217 VP.n1305 VP.n1301 0.024
R6218 VP.n324 VP.n322 0.024
R6219 VP.n9325 VP.n9324 0.024
R6220 VP.n8898 VP.n8897 0.024
R6221 VP.n8532 VP.n8531 0.024
R6222 VP.n8054 VP.n8053 0.024
R6223 VP.n7693 VP.n7692 0.024
R6224 VP.n7226 VP.n7225 0.024
R6225 VP.n6854 VP.n6853 0.024
R6226 VP.n6367 VP.n6366 0.024
R6227 VP.n5990 VP.n5989 0.024
R6228 VP.n5511 VP.n5510 0.024
R6229 VP.n5126 VP.n5125 0.024
R6230 VP.n4616 VP.n4615 0.024
R6231 VP.n4220 VP.n4219 0.024
R6232 VP.n3710 VP.n3709 0.024
R6233 VP.n3299 VP.n3298 0.024
R6234 VP.n2770 VP.n2769 0.024
R6235 VP.n2634 VP.n2633 0.024
R6236 VP.n1810 VP.n1809 0.024
R6237 VP.n1373 VP.n1372 0.024
R6238 VP.n824 VP.n823 0.024
R6239 VP.n10414 VP.n10413 0.024
R6240 VP.n747 VP.n746 0.024
R6241 VP.n390 VP.n389 0.024
R6242 VP.n437 VP.n436 0.024
R6243 VP.n484 VP.n483 0.024
R6244 VP.n531 VP.n530 0.024
R6245 VP.n578 VP.n577 0.024
R6246 VP.n618 VP.n617 0.024
R6247 VP.n720 VP.n719 0.024
R6248 VP.n9807 VP.n9798 0.024
R6249 VP.n8169 VP.n8159 0.024
R6250 VP.n9013 VP.n9003 0.024
R6251 VP.n9785 VP.n9776 0.024
R6252 VP.n6459 VP.n6449 0.024
R6253 VP.n7318 VP.n7308 0.024
R6254 VP.n8146 VP.n8136 0.024
R6255 VP.n8990 VP.n8980 0.024
R6256 VP.n9763 VP.n9754 0.024
R6257 VP.n2813 VP.n2803 0.024
R6258 VP.n3753 VP.n3743 0.024
R6259 VP.n4659 VP.n4649 0.024
R6260 VP.n5554 VP.n5544 0.024
R6261 VP.n6410 VP.n6400 0.024
R6262 VP.n7269 VP.n7259 0.024
R6263 VP.n8097 VP.n8087 0.024
R6264 VP.n8941 VP.n8931 0.024
R6265 VP.n9741 VP.n9732 0.024
R6266 VP.n1723 VP.n1722 0.024
R6267 VP.n4680 VP.n4676 0.024
R6268 VP.n5575 VP.n5571 0.024
R6269 VP.n6431 VP.n6427 0.024
R6270 VP.n7290 VP.n7286 0.024
R6271 VP.n8118 VP.n8114 0.024
R6272 VP.n8962 VP.n8958 0.024
R6273 VP.n9625 VP.n9624 0.024
R6274 VP.n9992 VP.n9988 0.024
R6275 VP.n9236 VP.n9231 0.024
R6276 VP.n7960 VP.n7959 0.024
R6277 VP.n9944 VP.n9940 0.024
R6278 VP.n9186 VP.n9181 0.024
R6279 VP.n8387 VP.n8382 0.024
R6280 VP.n7570 VP.n7565 0.024
R6281 VP.n6273 VP.n6272 0.024
R6282 VP.n9896 VP.n9892 0.024
R6283 VP.n9136 VP.n9131 0.024
R6284 VP.n8338 VP.n8333 0.024
R6285 VP.n7521 VP.n7516 0.024
R6286 VP.n6709 VP.n6704 0.024
R6287 VP.n5867 VP.n5862 0.024
R6288 VP.n4522 VP.n4521 0.024
R6289 VP.n10451 VP.n10450 0.024
R6290 VP.n9832 VP.n9831 0.024
R6291 VP.n9069 VP.n9068 0.024
R6292 VP.n8272 VP.n8271 0.024
R6293 VP.n7456 VP.n7455 0.024
R6294 VP.n6644 VP.n6643 0.024
R6295 VP.n5800 VP.n5799 0.024
R6296 VP.n4963 VP.n4962 0.024
R6297 VP.n4080 VP.n4079 0.024
R6298 VP.n2325 VP.n2324 0.024
R6299 VP.n8189 VP.n8187 0.023
R6300 VP.n6479 VP.n6477 0.023
R6301 VP.n4705 VP.n4703 0.023
R6302 VP.n2829 VP.n2827 0.023
R6303 VP.n9598 VP.n9597 0.023
R6304 VP.n9597 VP.n9596 0.023
R6305 VP.n9601 VP.n9599 0.023
R6306 VP.n8791 VP.n8790 0.023
R6307 VP.n8795 VP.n8792 0.023
R6308 VP.n9263 VP.n9262 0.023
R6309 VP.n8794 VP.n8793 0.023
R6310 VP.n8191 VP.n8190 0.023
R6311 VP.n9026 VP.n9024 0.023
R6312 VP.n9028 VP.n9027 0.023
R6313 VP.n8769 VP.n8768 0.023
R6314 VP.n8193 VP.n8192 0.023
R6315 VP.n7068 VP.n7067 0.023
R6316 VP.n7072 VP.n7069 0.023
R6317 VP.n7597 VP.n7596 0.023
R6318 VP.n7071 VP.n7070 0.023
R6319 VP.n9970 VP.n9962 0.023
R6320 VP.n9213 VP.n9205 0.023
R6321 VP.n8413 VP.n8405 0.023
R6322 VP.n6481 VP.n6480 0.023
R6323 VP.n7331 VP.n7329 0.023
R6324 VP.n7333 VP.n7332 0.023
R6325 VP.n7046 VP.n7045 0.023
R6326 VP.n6483 VP.n6482 0.023
R6327 VP.n5289 VP.n5288 0.023
R6328 VP.n5293 VP.n5290 0.023
R6329 VP.n5894 VP.n5893 0.023
R6330 VP.n5292 VP.n5291 0.023
R6331 VP.n9922 VP.n9914 0.023
R6332 VP.n9163 VP.n9155 0.023
R6333 VP.n8364 VP.n8356 0.023
R6334 VP.n7547 VP.n7539 0.023
R6335 VP.n6735 VP.n6727 0.023
R6336 VP.n4707 VP.n4706 0.023
R6337 VP.n5593 VP.n5591 0.023
R6338 VP.n5595 VP.n5594 0.023
R6339 VP.n5267 VP.n5266 0.023
R6340 VP.n4709 VP.n4708 0.023
R6341 VP.n3412 VP.n3411 0.023
R6342 VP.n3416 VP.n3413 0.023
R6343 VP.n4124 VP.n4123 0.023
R6344 VP.n3415 VP.n3414 0.023
R6345 VP.n9874 VP.n9866 0.023
R6346 VP.n9113 VP.n9105 0.023
R6347 VP.n8315 VP.n8307 0.023
R6348 VP.n7498 VP.n7490 0.023
R6349 VP.n6686 VP.n6678 0.023
R6350 VP.n5844 VP.n5836 0.023
R6351 VP.n5007 VP.n4999 0.023
R6352 VP.n1426 VP.n1425 0.023
R6353 VP.n857 VP.n852 0.023
R6354 VP.n859 VP.n858 0.023
R6355 VP.n1843 VP.n1841 0.023
R6356 VP.n1845 VP.n1844 0.023
R6357 VP.n751 VP.n748 0.023
R6358 VP.n36 VP.n35 0.023
R6359 VP.n26 VP.n25 0.023
R6360 VP.n137 VP.n136 0.023
R6361 VP.n8860 VP.n8852 0.023
R6362 VP.n9697 VP.n9696 0.023
R6363 VP.n9690 VP.n9689 0.023
R6364 VP.n9332 VP.n9331 0.023
R6365 VP.n9327 VP.n9326 0.023
R6366 VP.n8906 VP.n8905 0.023
R6367 VP.n8900 VP.n8899 0.023
R6368 VP.n8539 VP.n8538 0.023
R6369 VP.n8534 VP.n8533 0.023
R6370 VP.n8062 VP.n8061 0.023
R6371 VP.n8056 VP.n8055 0.023
R6372 VP.n7700 VP.n7699 0.023
R6373 VP.n7695 VP.n7694 0.023
R6374 VP.n7234 VP.n7233 0.023
R6375 VP.n7228 VP.n7227 0.023
R6376 VP.n6861 VP.n6860 0.023
R6377 VP.n6856 VP.n6855 0.023
R6378 VP.n6375 VP.n6374 0.023
R6379 VP.n6369 VP.n6368 0.023
R6380 VP.n5997 VP.n5996 0.023
R6381 VP.n5992 VP.n5991 0.023
R6382 VP.n5519 VP.n5518 0.023
R6383 VP.n5513 VP.n5512 0.023
R6384 VP.n5133 VP.n5132 0.023
R6385 VP.n5128 VP.n5127 0.023
R6386 VP.n4624 VP.n4623 0.023
R6387 VP.n4618 VP.n4617 0.023
R6388 VP.n4227 VP.n4226 0.023
R6389 VP.n4222 VP.n4221 0.023
R6390 VP.n3718 VP.n3717 0.023
R6391 VP.n3712 VP.n3711 0.023
R6392 VP.n3306 VP.n3305 0.023
R6393 VP.n3301 VP.n3300 0.023
R6394 VP.n2778 VP.n2777 0.023
R6395 VP.n2772 VP.n2771 0.023
R6396 VP.n2641 VP.n2640 0.023
R6397 VP.n2636 VP.n2635 0.023
R6398 VP.n1818 VP.n1817 0.023
R6399 VP.n1812 VP.n1811 0.023
R6400 VP.n1380 VP.n1379 0.023
R6401 VP.n1375 VP.n1374 0.023
R6402 VP.n834 VP.n833 0.023
R6403 VP.n826 VP.n825 0.023
R6404 VP.n199 VP.n157 0.023
R6405 VP.n144 VP.n143 0.023
R6406 VP.n9717 VP.n9709 0.023
R6407 VP.n10416 VP.n10415 0.023
R6408 VP.n10418 VP.n10411 0.023
R6409 VP.n9854 VP.n9846 0.023
R6410 VP.n9092 VP.n9084 0.023
R6411 VP.n8295 VP.n8287 0.023
R6412 VP.n7478 VP.n7470 0.023
R6413 VP.n6666 VP.n6658 0.023
R6414 VP.n5823 VP.n5815 0.023
R6415 VP.n4986 VP.n4978 0.023
R6416 VP.n4103 VP.n4095 0.023
R6417 VP.n3211 VP.n3203 0.023
R6418 VP.n2830 VP.n2826 0.023
R6419 VP.n3770 VP.n3768 0.023
R6420 VP.n3772 VP.n3771 0.023
R6421 VP.n10085 VP.n10084 0.023
R6422 VP.n914 VP.n913 0.023
R6423 VP.n1901 VP.n1900 0.023
R6424 VP.n1909 VP.n1908 0.023
R6425 VP.n964 VP.n963 0.023
R6426 VP.n2882 VP.n2881 0.023
R6427 VP.n2890 VP.n2889 0.023
R6428 VP.n1953 VP.n1952 0.023
R6429 VP.n1961 VP.n1960 0.023
R6430 VP.n1014 VP.n1013 0.023
R6431 VP.n3827 VP.n3826 0.023
R6432 VP.n3835 VP.n3834 0.023
R6433 VP.n2934 VP.n2933 0.023
R6434 VP.n2942 VP.n2941 0.023
R6435 VP.n2005 VP.n2004 0.023
R6436 VP.n2013 VP.n2012 0.023
R6437 VP.n1064 VP.n1063 0.023
R6438 VP.n4762 VP.n4761 0.023
R6439 VP.n4770 VP.n4769 0.023
R6440 VP.n3879 VP.n3878 0.023
R6441 VP.n3887 VP.n3886 0.023
R6442 VP.n2986 VP.n2985 0.023
R6443 VP.n2994 VP.n2993 0.023
R6444 VP.n2057 VP.n2056 0.023
R6445 VP.n2065 VP.n2064 0.023
R6446 VP.n1114 VP.n1113 0.023
R6447 VP.n746 VP.n745 0.022
R6448 VP.n389 VP.n388 0.022
R6449 VP.n436 VP.n435 0.022
R6450 VP.n483 VP.n482 0.022
R6451 VP.n530 VP.n529 0.022
R6452 VP.n577 VP.n576 0.022
R6453 VP.n617 VP.n616 0.022
R6454 VP.n719 VP.n718 0.022
R6455 VP.n10062 VP.n10061 0.022
R6456 VP.n10018 VP.n10017 0.022
R6457 VP.n8183 VP.n8182 0.022
R6458 VP.n8424 VP.n8423 0.022
R6459 VP.n9224 VP.n9223 0.022
R6460 VP.n9981 VP.n9980 0.022
R6461 VP.n9964 VP.n9963 0.022
R6462 VP.n9207 VP.n9206 0.022
R6463 VP.n8407 VP.n8406 0.022
R6464 VP.n6473 VP.n6472 0.022
R6465 VP.n6746 VP.n6745 0.022
R6466 VP.n7558 VP.n7557 0.022
R6467 VP.n8375 VP.n8374 0.022
R6468 VP.n9174 VP.n9173 0.022
R6469 VP.n9933 VP.n9932 0.022
R6470 VP.n9916 VP.n9915 0.022
R6471 VP.n9157 VP.n9156 0.022
R6472 VP.n8358 VP.n8357 0.022
R6473 VP.n7541 VP.n7540 0.022
R6474 VP.n6729 VP.n6728 0.022
R6475 VP.n4699 VP.n4698 0.022
R6476 VP.n5018 VP.n5017 0.022
R6477 VP.n5855 VP.n5854 0.022
R6478 VP.n6697 VP.n6696 0.022
R6479 VP.n7509 VP.n7508 0.022
R6480 VP.n8326 VP.n8325 0.022
R6481 VP.n9124 VP.n9123 0.022
R6482 VP.n9885 VP.n9884 0.022
R6483 VP.n9868 VP.n9867 0.022
R6484 VP.n9107 VP.n9106 0.022
R6485 VP.n8309 VP.n8308 0.022
R6486 VP.n7492 VP.n7491 0.022
R6487 VP.n6680 VP.n6679 0.022
R6488 VP.n5838 VP.n5837 0.022
R6489 VP.n5001 VP.n5000 0.022
R6490 VP.n9816 VP.n9815 0.022
R6491 VP.n9052 VP.n9051 0.022
R6492 VP.n8255 VP.n8254 0.022
R6493 VP.n7439 VP.n7438 0.022
R6494 VP.n6627 VP.n6626 0.022
R6495 VP.n5783 VP.n5782 0.022
R6496 VP.n4946 VP.n4945 0.022
R6497 VP.n4063 VP.n4062 0.022
R6498 VP.n3170 VP.n3169 0.022
R6499 VP.n10693 VP.n10692 0.022
R6500 VP.n1314 VP.n1313 0.022
R6501 VP.n745 VP.n744 0.022
R6502 VP.n125 VP.n124 0.022
R6503 VP.n764 VP.n763 0.022
R6504 VP.n2290 VP.n2289 0.022
R6505 VP.n388 VP.n387 0.022
R6506 VP.n112 VP.n111 0.022
R6507 VP.n891 VP.n890 0.022
R6508 VP.n883 VP.n882 0.022
R6509 VP.n1753 VP.n1752 0.022
R6510 VP.n3240 VP.n3239 0.022
R6511 VP.n435 VP.n434 0.022
R6512 VP.n94 VP.n91 0.022
R6513 VP.n941 VP.n940 0.022
R6514 VP.n933 VP.n932 0.022
R6515 VP.n1878 VP.n1877 0.022
R6516 VP.n1870 VP.n1869 0.022
R6517 VP.n2714 VP.n2713 0.022
R6518 VP.n4161 VP.n4160 0.022
R6519 VP.n482 VP.n481 0.022
R6520 VP.n86 VP.n85 0.022
R6521 VP.n991 VP.n990 0.022
R6522 VP.n984 VP.n983 0.022
R6523 VP.n1930 VP.n1929 0.022
R6524 VP.n1923 VP.n1922 0.022
R6525 VP.n2859 VP.n2858 0.022
R6526 VP.n2852 VP.n2851 0.022
R6527 VP.n3654 VP.n3653 0.022
R6528 VP.n5067 VP.n5066 0.022
R6529 VP.n529 VP.n528 0.022
R6530 VP.n68 VP.n65 0.022
R6531 VP.n1041 VP.n1040 0.022
R6532 VP.n1034 VP.n1033 0.022
R6533 VP.n1982 VP.n1981 0.022
R6534 VP.n1974 VP.n1973 0.022
R6535 VP.n2911 VP.n2910 0.022
R6536 VP.n2904 VP.n2903 0.022
R6537 VP.n3804 VP.n3803 0.022
R6538 VP.n3796 VP.n3795 0.022
R6539 VP.n4560 VP.n4559 0.022
R6540 VP.n5931 VP.n5930 0.022
R6541 VP.n576 VP.n575 0.022
R6542 VP.n60 VP.n59 0.022
R6543 VP.n1091 VP.n1090 0.022
R6544 VP.n1083 VP.n1082 0.022
R6545 VP.n2034 VP.n2033 0.022
R6546 VP.n2026 VP.n2025 0.022
R6547 VP.n2963 VP.n2962 0.022
R6548 VP.n2956 VP.n2955 0.022
R6549 VP.n3856 VP.n3855 0.022
R6550 VP.n3849 VP.n3848 0.022
R6551 VP.n4739 VP.n4738 0.022
R6552 VP.n4732 VP.n4731 0.022
R6553 VP.n5455 VP.n5454 0.022
R6554 VP.n6795 VP.n6794 0.022
R6555 VP.n616 VP.n615 0.022
R6556 VP.n42 VP.n39 0.022
R6557 VP.n1141 VP.n1140 0.022
R6558 VP.n1133 VP.n1132 0.022
R6559 VP.n2086 VP.n2085 0.022
R6560 VP.n2079 VP.n2078 0.022
R6561 VP.n3015 VP.n3014 0.022
R6562 VP.n3008 VP.n3007 0.022
R6563 VP.n3908 VP.n3907 0.022
R6564 VP.n3900 VP.n3899 0.022
R6565 VP.n4791 VP.n4790 0.022
R6566 VP.n4783 VP.n4782 0.022
R6567 VP.n5628 VP.n5627 0.022
R6568 VP.n5621 VP.n5620 0.022
R6569 VP.n6311 VP.n6310 0.022
R6570 VP.n7634 VP.n7633 0.022
R6571 VP.n32 VP.n29 0.022
R6572 VP.n1179 VP.n1178 0.022
R6573 VP.n1172 VP.n1171 0.022
R6574 VP.n2127 VP.n2126 0.022
R6575 VP.n2119 VP.n2118 0.022
R6576 VP.n3056 VP.n3055 0.022
R6577 VP.n3049 VP.n3048 0.022
R6578 VP.n3949 VP.n3948 0.022
R6579 VP.n3941 VP.n3940 0.022
R6580 VP.n4832 VP.n4831 0.022
R6581 VP.n4824 VP.n4823 0.022
R6582 VP.n5669 VP.n5668 0.022
R6583 VP.n5661 VP.n5660 0.022
R6584 VP.n6513 VP.n6512 0.022
R6585 VP.n6506 VP.n6505 0.022
R6586 VP.n7170 VP.n7169 0.022
R6587 VP.n8473 VP.n8472 0.022
R6588 VP.n22 VP.n19 0.022
R6589 VP.n1219 VP.n1218 0.022
R6590 VP.n1212 VP.n1211 0.022
R6591 VP.n2168 VP.n2167 0.022
R6592 VP.n2160 VP.n2159 0.022
R6593 VP.n3097 VP.n3096 0.022
R6594 VP.n3090 VP.n3089 0.022
R6595 VP.n3990 VP.n3989 0.022
R6596 VP.n3983 VP.n3982 0.022
R6597 VP.n4873 VP.n4872 0.022
R6598 VP.n4866 VP.n4865 0.022
R6599 VP.n5710 VP.n5709 0.022
R6600 VP.n5703 VP.n5702 0.022
R6601 VP.n6554 VP.n6553 0.022
R6602 VP.n6547 VP.n6546 0.022
R6603 VP.n7366 VP.n7365 0.022
R6604 VP.n7358 VP.n7357 0.022
R6605 VP.n7998 VP.n7997 0.022
R6606 VP.n9679 VP.n9678 0.022
R6607 VP.n8854 VP.n8853 0.022
R6608 VP.n718 VP.n717 0.022
R6609 VP.n14 VP.n13 0.022
R6610 VP.n1260 VP.n1259 0.022
R6611 VP.n1253 VP.n1252 0.022
R6612 VP.n2209 VP.n2208 0.022
R6613 VP.n2201 VP.n2200 0.022
R6614 VP.n3138 VP.n3137 0.022
R6615 VP.n3131 VP.n3130 0.022
R6616 VP.n4031 VP.n4030 0.022
R6617 VP.n4024 VP.n4023 0.022
R6618 VP.n4914 VP.n4913 0.022
R6619 VP.n4906 VP.n4905 0.022
R6620 VP.n5751 VP.n5750 0.022
R6621 VP.n5743 VP.n5742 0.022
R6622 VP.n6595 VP.n6594 0.022
R6623 VP.n6588 VP.n6587 0.022
R6624 VP.n7407 VP.n7406 0.022
R6625 VP.n7400 VP.n7399 0.022
R6626 VP.n8223 VP.n8222 0.022
R6627 VP.n8216 VP.n8215 0.022
R6628 VP.n8832 VP.n8831 0.022
R6629 VP.n9300 VP.n9299 0.022
R6630 VP.n133 VP.n131 0.022
R6631 VP.n806 VP.n805 0.022
R6632 VP.n799 VP.n798 0.022
R6633 VP.n1792 VP.n1791 0.022
R6634 VP.n1784 VP.n1783 0.022
R6635 VP.n2752 VP.n2751 0.022
R6636 VP.n2745 VP.n2744 0.022
R6637 VP.n3692 VP.n3691 0.022
R6638 VP.n3684 VP.n3683 0.022
R6639 VP.n4601 VP.n4600 0.022
R6640 VP.n4594 VP.n4593 0.022
R6641 VP.n5493 VP.n5492 0.022
R6642 VP.n5486 VP.n5485 0.022
R6643 VP.n6349 VP.n6348 0.022
R6644 VP.n6342 VP.n6341 0.022
R6645 VP.n7208 VP.n7207 0.022
R6646 VP.n7201 VP.n7200 0.022
R6647 VP.n8036 VP.n8035 0.022
R6648 VP.n8028 VP.n8027 0.022
R6649 VP.n8880 VP.n8879 0.022
R6650 VP.n156 VP.n155 0.022
R6651 VP.n9714 VP.n9713 0.022
R6652 VP.n10653 VP.n10652 0.022
R6653 VP.n2 VP.n0 0.022
R6654 VP.n9848 VP.n9847 0.022
R6655 VP.n9086 VP.n9085 0.022
R6656 VP.n8289 VP.n8288 0.022
R6657 VP.n7472 VP.n7471 0.022
R6658 VP.n6660 VP.n6659 0.022
R6659 VP.n5817 VP.n5816 0.022
R6660 VP.n4980 VP.n4979 0.022
R6661 VP.n4097 VP.n4096 0.022
R6662 VP.n3205 VP.n3204 0.022
R6663 VP.n11003 VP.n11002 0.022
R6664 VP.n10944 VP.n10943 0.022
R6665 VP.n8742 VP.n8741 0.022
R6666 VP.n9549 VP.n9548 0.022
R6667 VP.n10893 VP.n10892 0.022
R6668 VP.n7019 VP.n7018 0.022
R6669 VP.n7857 VP.n7856 0.022
R6670 VP.n8694 VP.n8693 0.022
R6671 VP.n9498 VP.n9497 0.022
R6672 VP.n10842 VP.n10841 0.022
R6673 VP.n5240 VP.n5239 0.022
R6674 VP.n6106 VP.n6105 0.022
R6675 VP.n6970 VP.n6969 0.022
R6676 VP.n7808 VP.n7807 0.022
R6677 VP.n8646 VP.n8645 0.022
R6678 VP.n9447 VP.n9446 0.022
R6679 VP.n10791 VP.n10790 0.022
R6680 VP.n10726 VP.n10725 0.022
R6681 VP.n9381 VP.n9380 0.022
R6682 VP.n8586 VP.n8585 0.022
R6683 VP.n7747 VP.n7746 0.022
R6684 VP.n6908 VP.n6907 0.022
R6685 VP.n6044 VP.n6043 0.022
R6686 VP.n5180 VP.n5179 0.022
R6687 VP.n4274 VP.n4273 0.022
R6688 VP.n3353 VP.n3352 0.022
R6689 VP.n898 VP.n897 0.022
R6690 VP.n1332 VP.n1331 0.022
R6691 VP.n948 VP.n947 0.022
R6692 VP.n1460 VP.n1459 0.022
R6693 VP.n1885 VP.n1884 0.022
R6694 VP.n2308 VP.n2307 0.022
R6695 VP.n998 VP.n997 0.022
R6696 VP.n1498 VP.n1497 0.022
R6697 VP.n1937 VP.n1936 0.022
R6698 VP.n2560 VP.n2559 0.022
R6699 VP.n2866 VP.n2865 0.022
R6700 VP.n3258 VP.n3257 0.022
R6701 VP.n1048 VP.n1047 0.022
R6702 VP.n1536 VP.n1535 0.022
R6703 VP.n1989 VP.n1988 0.022
R6704 VP.n2522 VP.n2521 0.022
R6705 VP.n2918 VP.n2917 0.022
R6706 VP.n3438 VP.n3437 0.022
R6707 VP.n3811 VP.n3810 0.022
R6708 VP.n4179 VP.n4178 0.022
R6709 VP.n1098 VP.n1097 0.022
R6710 VP.n1574 VP.n1573 0.022
R6711 VP.n2041 VP.n2040 0.022
R6712 VP.n2484 VP.n2483 0.022
R6713 VP.n2970 VP.n2969 0.022
R6714 VP.n3476 VP.n3475 0.022
R6715 VP.n3863 VP.n3862 0.022
R6716 VP.n4355 VP.n4354 0.022
R6717 VP.n4746 VP.n4745 0.022
R6718 VP.n5085 VP.n5084 0.022
R6719 VP.n1148 VP.n1147 0.022
R6720 VP.n1612 VP.n1611 0.022
R6721 VP.n2093 VP.n2092 0.022
R6722 VP.n2452 VP.n2451 0.022
R6723 VP.n3022 VP.n3021 0.022
R6724 VP.n3514 VP.n3513 0.022
R6725 VP.n3915 VP.n3914 0.022
R6726 VP.n4393 VP.n4392 0.022
R6727 VP.n4798 VP.n4797 0.022
R6728 VP.n5315 VP.n5314 0.022
R6729 VP.n5635 VP.n5634 0.022
R6730 VP.n5949 VP.n5948 0.022
R6731 VP.n1186 VP.n1185 0.022
R6732 VP.n1644 VP.n1643 0.022
R6733 VP.n2134 VP.n2133 0.022
R6734 VP.n2420 VP.n2419 0.022
R6735 VP.n3063 VP.n3062 0.022
R6736 VP.n3546 VP.n3545 0.022
R6737 VP.n3956 VP.n3955 0.022
R6738 VP.n4425 VP.n4424 0.022
R6739 VP.n4839 VP.n4838 0.022
R6740 VP.n5347 VP.n5346 0.022
R6741 VP.n5676 VP.n5675 0.022
R6742 VP.n6175 VP.n6174 0.022
R6743 VP.n6520 VP.n6519 0.022
R6744 VP.n6813 VP.n6812 0.022
R6745 VP.n1226 VP.n1225 0.022
R6746 VP.n1676 VP.n1675 0.022
R6747 VP.n2175 VP.n2174 0.022
R6748 VP.n2388 VP.n2387 0.022
R6749 VP.n3104 VP.n3103 0.022
R6750 VP.n3578 VP.n3577 0.022
R6751 VP.n3997 VP.n3996 0.022
R6752 VP.n4457 VP.n4456 0.022
R6753 VP.n4880 VP.n4879 0.022
R6754 VP.n5379 VP.n5378 0.022
R6755 VP.n5717 VP.n5716 0.022
R6756 VP.n6207 VP.n6206 0.022
R6757 VP.n6561 VP.n6560 0.022
R6758 VP.n7094 VP.n7093 0.022
R6759 VP.n7373 VP.n7372 0.022
R6760 VP.n7652 VP.n7651 0.022
R6761 VP.n1267 VP.n1266 0.022
R6762 VP.n1708 VP.n1707 0.022
R6763 VP.n2216 VP.n2215 0.022
R6764 VP.n2356 VP.n2355 0.022
R6765 VP.n3145 VP.n3144 0.022
R6766 VP.n3610 VP.n3609 0.022
R6767 VP.n4038 VP.n4037 0.022
R6768 VP.n4489 VP.n4488 0.022
R6769 VP.n4921 VP.n4920 0.022
R6770 VP.n5411 VP.n5410 0.022
R6771 VP.n5758 VP.n5757 0.022
R6772 VP.n6239 VP.n6238 0.022
R6773 VP.n6602 VP.n6601 0.022
R6774 VP.n7126 VP.n7125 0.022
R6775 VP.n7414 VP.n7413 0.022
R6776 VP.n7926 VP.n7925 0.022
R6777 VP.n8230 VP.n8229 0.022
R6778 VP.n8491 VP.n8490 0.022
R6779 VP.n813 VP.n812 0.022
R6780 VP.n1363 VP.n1362 0.022
R6781 VP.n1799 VP.n1798 0.022
R6782 VP.n2680 VP.n2679 0.022
R6783 VP.n2759 VP.n2758 0.022
R6784 VP.n3289 VP.n3288 0.022
R6785 VP.n3699 VP.n3698 0.022
R6786 VP.n4210 VP.n4209 0.022
R6787 VP.n4608 VP.n4607 0.022
R6788 VP.n5116 VP.n5115 0.022
R6789 VP.n5500 VP.n5499 0.022
R6790 VP.n5980 VP.n5979 0.022
R6791 VP.n6356 VP.n6355 0.022
R6792 VP.n6844 VP.n6843 0.022
R6793 VP.n7215 VP.n7214 0.022
R6794 VP.n7683 VP.n7682 0.022
R6795 VP.n8043 VP.n8042 0.022
R6796 VP.n8522 VP.n8521 0.022
R6797 VP.n8887 VP.n8886 0.022
R6798 VP.n8193 VP.n8189 0.022
R6799 VP.n6483 VP.n6479 0.022
R6800 VP.n4709 VP.n4705 0.022
R6801 VP.n2830 VP.n2829 0.022
R6802 VP.n9659 VP.n9317 0.021
R6803 VP.n8767 VP.n8766 0.021
R6804 VP.n7044 VP.n7043 0.021
R6805 VP.n5265 VP.n5264 0.021
R6806 VP.n2260 VP.n2252 0.021
R6807 VP.n854 VP.n853 0.021
R6808 VP.n1745 VP.n1744 0.021
R6809 VP.n922 VP.n921 0.021
R6810 VP.n2706 VP.n2705 0.021
R6811 VP.n1911 VP.n1910 0.021
R6812 VP.n1478 VP.n1477 0.021
R6813 VP.n972 VP.n971 0.021
R6814 VP.n3646 VP.n3645 0.021
R6815 VP.n2892 VP.n2891 0.021
R6816 VP.n2578 VP.n2577 0.021
R6817 VP.n1963 VP.n1962 0.021
R6818 VP.n1516 VP.n1515 0.021
R6819 VP.n1022 VP.n1021 0.021
R6820 VP.n4552 VP.n4551 0.021
R6821 VP.n3837 VP.n3836 0.021
R6822 VP.n3456 VP.n3455 0.021
R6823 VP.n2944 VP.n2943 0.021
R6824 VP.n2540 VP.n2539 0.021
R6825 VP.n2015 VP.n2014 0.021
R6826 VP.n1554 VP.n1553 0.021
R6827 VP.n1072 VP.n1071 0.021
R6828 VP.n5447 VP.n5446 0.021
R6829 VP.n4772 VP.n4771 0.021
R6830 VP.n4373 VP.n4372 0.021
R6831 VP.n3889 VP.n3888 0.021
R6832 VP.n3494 VP.n3493 0.021
R6833 VP.n2996 VP.n2995 0.021
R6834 VP.n2502 VP.n2501 0.021
R6835 VP.n2067 VP.n2066 0.021
R6836 VP.n1592 VP.n1591 0.021
R6837 VP.n1122 VP.n1121 0.021
R6838 VP.n6303 VP.n6302 0.021
R6839 VP.n7162 VP.n7161 0.021
R6840 VP.n7990 VP.n7989 0.021
R6841 VP.n2825 VP.n2824 0.021
R6842 VP.n10120 VP.n10119 0.021
R6843 VP.n771 VP.n770 0.021
R6844 VP.n1760 VP.n1759 0.021
R6845 VP.n2721 VP.n2720 0.021
R6846 VP.n3661 VP.n3660 0.021
R6847 VP.n4567 VP.n4566 0.021
R6848 VP.n5462 VP.n5461 0.021
R6849 VP.n6318 VP.n6317 0.021
R6850 VP.n7177 VP.n7176 0.021
R6851 VP.n8005 VP.n8004 0.021
R6852 VP.n8839 VP.n8838 0.021
R6853 VP.n10110 VP.n10109 0.021
R6854 VP.n10089 VP.n10088 0.021
R6855 VP.n8956 VP.n8955 0.021
R6856 VP.n8112 VP.n8111 0.021
R6857 VP.n7284 VP.n7283 0.021
R6858 VP.n6425 VP.n6424 0.021
R6859 VP.n5569 VP.n5568 0.021
R6860 VP.n4674 VP.n4673 0.021
R6861 VP.n10030 VP.n10029 0.021
R6862 VP.n9266 VP.n9265 0.021
R6863 VP.n9796 VP.n9795 0.021
R6864 VP.n9026 VP.n9025 0.021
R6865 VP.n9991 VP.n9990 0.021
R6866 VP.n9235 VP.n9234 0.021
R6867 VP.n8436 VP.n8435 0.021
R6868 VP.n7600 VP.n7599 0.021
R6869 VP.n9774 VP.n9773 0.021
R6870 VP.n9001 VP.n9000 0.021
R6871 VP.n8157 VP.n8156 0.021
R6872 VP.n7331 VP.n7330 0.021
R6873 VP.n9943 VP.n9942 0.021
R6874 VP.n9185 VP.n9184 0.021
R6875 VP.n8386 VP.n8385 0.021
R6876 VP.n7569 VP.n7568 0.021
R6877 VP.n6758 VP.n6757 0.021
R6878 VP.n5897 VP.n5896 0.021
R6879 VP.n9752 VP.n9751 0.021
R6880 VP.n8978 VP.n8977 0.021
R6881 VP.n8134 VP.n8133 0.021
R6882 VP.n7306 VP.n7305 0.021
R6883 VP.n6447 VP.n6446 0.021
R6884 VP.n5593 VP.n5592 0.021
R6885 VP.n9895 VP.n9894 0.021
R6886 VP.n9135 VP.n9134 0.021
R6887 VP.n8337 VP.n8336 0.021
R6888 VP.n7520 VP.n7519 0.021
R6889 VP.n6708 VP.n6707 0.021
R6890 VP.n5866 VP.n5865 0.021
R6891 VP.n5030 VP.n5029 0.021
R6892 VP.n4127 VP.n4126 0.021
R6893 VP.n10446 VP.n10445 0.021
R6894 VP.n9827 VP.n9826 0.021
R6895 VP.n9064 VP.n9063 0.021
R6896 VP.n8267 VP.n8266 0.021
R6897 VP.n7451 VP.n7450 0.021
R6898 VP.n6639 VP.n6638 0.021
R6899 VP.n5795 VP.n5794 0.021
R6900 VP.n4958 VP.n4957 0.021
R6901 VP.n4075 VP.n4074 0.021
R6902 VP.n3182 VP.n3181 0.021
R6903 VP.n2255 VP.n2254 0.021
R6904 VP.n9730 VP.n9729 0.021
R6905 VP.n8929 VP.n8928 0.021
R6906 VP.n8085 VP.n8084 0.021
R6907 VP.n7257 VP.n7256 0.021
R6908 VP.n6398 VP.n6397 0.021
R6909 VP.n5542 VP.n5541 0.021
R6910 VP.n4647 VP.n4646 0.021
R6911 VP.n3741 VP.n3740 0.021
R6912 VP.n2801 VP.n2800 0.021
R6913 VP.n857 VP.n856 0.021
R6914 VP.n1843 VP.n1842 0.021
R6915 VP.n824 VP.n822 0.021
R6916 VP.n1810 VP.n1808 0.021
R6917 VP.n2770 VP.n2768 0.021
R6918 VP.n3710 VP.n3708 0.021
R6919 VP.n4616 VP.n4614 0.021
R6920 VP.n5511 VP.n5509 0.021
R6921 VP.n6367 VP.n6365 0.021
R6922 VP.n7226 VP.n7224 0.021
R6923 VP.n8054 VP.n8052 0.021
R6924 VP.n8898 VP.n8896 0.021
R6925 VP.n257 VP.n256 0.021
R6926 VP.n359 VP.n358 0.021
R6927 VP.n406 VP.n405 0.021
R6928 VP.n453 VP.n452 0.021
R6929 VP.n500 VP.n499 0.021
R6930 VP.n547 VP.n546 0.021
R6931 VP.n594 VP.n593 0.021
R6932 VP.n634 VP.n633 0.021
R6933 VP.n664 VP.n663 0.021
R6934 VP.n696 VP.n695 0.021
R6935 VP.n10414 VP.n10412 0.021
R6936 VP.n3770 VP.n3769 0.021
R6937 VP.n830 VP.n828 0.02
R6938 VP.n8196 VP.n8195 0.02
R6939 VP.n6486 VP.n6485 0.02
R6940 VP.n4712 VP.n4711 0.02
R6941 VP.n10333 VP.n10332 0.019
R6942 VP.n10071 VP.n10070 0.019
R6943 VP.n10991 VP.n10990 0.019
R6944 VP.n11005 VP.n11004 0.019
R6945 VP.n10642 VP.n10641 0.019
R6946 VP.n10946 VP.n10945 0.019
R6947 VP.n10604 VP.n10603 0.019
R6948 VP.n9033 VP.n9032 0.019
R6949 VP.n9574 VP.n9563 0.019
R6950 VP.n8177 VP.n8176 0.019
R6951 VP.n8744 VP.n8743 0.019
R6952 VP.n9551 VP.n9550 0.019
R6953 VP.n10895 VP.n10894 0.019
R6954 VP.n10569 VP.n10568 0.019
R6955 VP.n9966 VP.n9965 0.019
R6956 VP.n9209 VP.n9208 0.019
R6957 VP.n8409 VP.n8408 0.019
R6958 VP.n7338 VP.n7337 0.019
R6959 VP.n7881 VP.n7871 0.019
R6960 VP.n8717 VP.n8707 0.019
R6961 VP.n9522 VP.n9511 0.019
R6962 VP.n6467 VP.n6466 0.019
R6963 VP.n7021 VP.n7020 0.019
R6964 VP.n7859 VP.n7858 0.019
R6965 VP.n8696 VP.n8695 0.019
R6966 VP.n9500 VP.n9499 0.019
R6967 VP.n10844 VP.n10843 0.019
R6968 VP.n10534 VP.n10533 0.019
R6969 VP.n9918 VP.n9917 0.019
R6970 VP.n9159 VP.n9158 0.019
R6971 VP.n8360 VP.n8359 0.019
R6972 VP.n7543 VP.n7542 0.019
R6973 VP.n6731 VP.n6730 0.019
R6974 VP.n5600 VP.n5599 0.019
R6975 VP.n6130 VP.n6120 0.019
R6976 VP.n6993 VP.n6983 0.019
R6977 VP.n7831 VP.n7821 0.019
R6978 VP.n8669 VP.n8659 0.019
R6979 VP.n9471 VP.n9460 0.019
R6980 VP.n4693 VP.n4692 0.019
R6981 VP.n5242 VP.n5241 0.019
R6982 VP.n6108 VP.n6107 0.019
R6983 VP.n6972 VP.n6971 0.019
R6984 VP.n7810 VP.n7809 0.019
R6985 VP.n8648 VP.n8647 0.019
R6986 VP.n9449 VP.n9448 0.019
R6987 VP.n10793 VP.n10792 0.019
R6988 VP.n10499 VP.n10498 0.019
R6989 VP.n9870 VP.n9869 0.019
R6990 VP.n9109 VP.n9108 0.019
R6991 VP.n8311 VP.n8310 0.019
R6992 VP.n7494 VP.n7493 0.019
R6993 VP.n6682 VP.n6681 0.019
R6994 VP.n5840 VP.n5839 0.019
R6995 VP.n5003 VP.n5002 0.019
R6996 VP.n10739 VP.n10727 0.019
R6997 VP.n9394 VP.n9382 0.019
R6998 VP.n8597 VP.n8587 0.019
R6999 VP.n7758 VP.n7748 0.019
R7000 VP.n6920 VP.n6909 0.019
R7001 VP.n6056 VP.n6045 0.019
R7002 VP.n5191 VP.n5181 0.019
R7003 VP.n4285 VP.n4275 0.019
R7004 VP.n3364 VP.n3354 0.019
R7005 VP.n864 VP.n863 0.019
R7006 VP.n1850 VP.n1849 0.019
R7007 VP.n2626 VP.n2616 0.019
R7008 VP.n3337 VP.n3327 0.019
R7009 VP.n4258 VP.n4248 0.019
R7010 VP.n5164 VP.n5154 0.019
R7011 VP.n6028 VP.n6018 0.019
R7012 VP.n6892 VP.n6882 0.019
R7013 VP.n7731 VP.n7721 0.019
R7014 VP.n8570 VP.n8560 0.019
R7015 VP.n9365 VP.n9354 0.019
R7016 VP.n10710 VP.n10697 0.019
R7017 VP.n1319 VP.n774 0.019
R7018 VP.n917 VP.n916 0.019
R7019 VP.n376 VP.n375 0.019
R7020 VP.n924 VP.n899 0.019
R7021 VP.n1747 VP.n1333 0.019
R7022 VP.n2295 VP.n1763 0.019
R7023 VP.n1904 VP.n1903 0.019
R7024 VP.n967 VP.n966 0.019
R7025 VP.n423 VP.n422 0.019
R7026 VP.n974 VP.n949 0.019
R7027 VP.n1480 VP.n1461 0.019
R7028 VP.n1913 VP.n1886 0.019
R7029 VP.n2708 VP.n2309 0.019
R7030 VP.n3245 VP.n2724 0.019
R7031 VP.n2885 VP.n2884 0.019
R7032 VP.n1956 VP.n1955 0.019
R7033 VP.n1017 VP.n1016 0.019
R7034 VP.n470 VP.n469 0.019
R7035 VP.n1024 VP.n999 0.019
R7036 VP.n1518 VP.n1499 0.019
R7037 VP.n1965 VP.n1938 0.019
R7038 VP.n2580 VP.n2561 0.019
R7039 VP.n2894 VP.n2867 0.019
R7040 VP.n3648 VP.n3259 0.019
R7041 VP.n4166 VP.n3664 0.019
R7042 VP.n3830 VP.n3829 0.019
R7043 VP.n2937 VP.n2936 0.019
R7044 VP.n2008 VP.n2007 0.019
R7045 VP.n1067 VP.n1066 0.019
R7046 VP.n517 VP.n516 0.019
R7047 VP.n1074 VP.n1049 0.019
R7048 VP.n1556 VP.n1537 0.019
R7049 VP.n2017 VP.n1990 0.019
R7050 VP.n2542 VP.n2523 0.019
R7051 VP.n2946 VP.n2919 0.019
R7052 VP.n3458 VP.n3439 0.019
R7053 VP.n3839 VP.n3812 0.019
R7054 VP.n4554 VP.n4180 0.019
R7055 VP.n5072 VP.n4570 0.019
R7056 VP.n4765 VP.n4764 0.019
R7057 VP.n3882 VP.n3881 0.019
R7058 VP.n2989 VP.n2988 0.019
R7059 VP.n2060 VP.n2059 0.019
R7060 VP.n1117 VP.n1116 0.019
R7061 VP.n564 VP.n563 0.019
R7062 VP.n1124 VP.n1099 0.019
R7063 VP.n1594 VP.n1575 0.019
R7064 VP.n2069 VP.n2042 0.019
R7065 VP.n2504 VP.n2485 0.019
R7066 VP.n2998 VP.n2971 0.019
R7067 VP.n3496 VP.n3477 0.019
R7068 VP.n3891 VP.n3864 0.019
R7069 VP.n4375 VP.n4356 0.019
R7070 VP.n4774 VP.n4747 0.019
R7071 VP.n5449 VP.n5086 0.019
R7072 VP.n5936 VP.n5465 0.019
R7073 VP.n1162 VP.n1149 0.019
R7074 VP.n1626 VP.n1613 0.019
R7075 VP.n2110 VP.n2094 0.019
R7076 VP.n2466 VP.n2453 0.019
R7077 VP.n3039 VP.n3023 0.019
R7078 VP.n3528 VP.n3515 0.019
R7079 VP.n3932 VP.n3916 0.019
R7080 VP.n4407 VP.n4394 0.019
R7081 VP.n4815 VP.n4799 0.019
R7082 VP.n5329 VP.n5316 0.019
R7083 VP.n5652 VP.n5636 0.019
R7084 VP.n6305 VP.n5950 0.019
R7085 VP.n6800 VP.n6321 0.019
R7086 VP.n1202 VP.n1187 0.019
R7087 VP.n1658 VP.n1645 0.019
R7088 VP.n2151 VP.n2135 0.019
R7089 VP.n2434 VP.n2421 0.019
R7090 VP.n3080 VP.n3064 0.019
R7091 VP.n3560 VP.n3547 0.019
R7092 VP.n3973 VP.n3957 0.019
R7093 VP.n4439 VP.n4426 0.019
R7094 VP.n4856 VP.n4840 0.019
R7095 VP.n5361 VP.n5348 0.019
R7096 VP.n5693 VP.n5677 0.019
R7097 VP.n6189 VP.n6176 0.019
R7098 VP.n6537 VP.n6521 0.019
R7099 VP.n7164 VP.n6814 0.019
R7100 VP.n7639 VP.n7180 0.019
R7101 VP.n1243 VP.n1227 0.019
R7102 VP.n1690 VP.n1677 0.019
R7103 VP.n2192 VP.n2176 0.019
R7104 VP.n2402 VP.n2389 0.019
R7105 VP.n3121 VP.n3105 0.019
R7106 VP.n3592 VP.n3579 0.019
R7107 VP.n4014 VP.n3998 0.019
R7108 VP.n4471 VP.n4458 0.019
R7109 VP.n4897 VP.n4881 0.019
R7110 VP.n5393 VP.n5380 0.019
R7111 VP.n5734 VP.n5718 0.019
R7112 VP.n6221 VP.n6208 0.019
R7113 VP.n6578 VP.n6562 0.019
R7114 VP.n7108 VP.n7095 0.019
R7115 VP.n7390 VP.n7374 0.019
R7116 VP.n7992 VP.n7653 0.019
R7117 VP.n8478 VP.n8008 0.019
R7118 VP.n9659 VP.n9658 0.019
R7119 VP.n8856 VP.n8855 0.019
R7120 VP.n1284 VP.n1268 0.019
R7121 VP.n1723 VP.n1709 0.019
R7122 VP.n2233 VP.n2217 0.019
R7123 VP.n2370 VP.n2357 0.019
R7124 VP.n3162 VP.n3146 0.019
R7125 VP.n3624 VP.n3611 0.019
R7126 VP.n4055 VP.n4039 0.019
R7127 VP.n4503 VP.n4490 0.019
R7128 VP.n4938 VP.n4922 0.019
R7129 VP.n5425 VP.n5412 0.019
R7130 VP.n5775 VP.n5759 0.019
R7131 VP.n6253 VP.n6240 0.019
R7132 VP.n6619 VP.n6603 0.019
R7133 VP.n7140 VP.n7127 0.019
R7134 VP.n7431 VP.n7415 0.019
R7135 VP.n7940 VP.n7927 0.019
R7136 VP.n8247 VP.n8231 0.019
R7137 VP.n8826 VP.n8492 0.019
R7138 VP.n9305 VP.n8842 0.019
R7139 VP.n8826 VP.n8825 0.019
R7140 VP.n287 VP.n286 0.019
R7141 VP.n815 VP.n814 0.019
R7142 VP.n1365 VP.n1364 0.019
R7143 VP.n1801 VP.n1800 0.019
R7144 VP.n2682 VP.n2681 0.019
R7145 VP.n2761 VP.n2760 0.019
R7146 VP.n3291 VP.n3290 0.019
R7147 VP.n3701 VP.n3700 0.019
R7148 VP.n4212 VP.n4211 0.019
R7149 VP.n4610 VP.n4609 0.019
R7150 VP.n5118 VP.n5117 0.019
R7151 VP.n5502 VP.n5501 0.019
R7152 VP.n5982 VP.n5981 0.019
R7153 VP.n6358 VP.n6357 0.019
R7154 VP.n6846 VP.n6845 0.019
R7155 VP.n7217 VP.n7216 0.019
R7156 VP.n7685 VP.n7684 0.019
R7157 VP.n8045 VP.n8044 0.019
R7158 VP.n8524 VP.n8523 0.019
R7159 VP.n8889 VP.n8888 0.019
R7160 VP.n10112 VP.n10103 0.019
R7161 VP.n10675 VP.n10123 0.019
R7162 VP.n11032 VP.n10682 0.019
R7163 VP.n9699 VP.n9698 0.019
R7164 VP.n9334 VP.n9333 0.019
R7165 VP.n8908 VP.n8907 0.019
R7166 VP.n8541 VP.n8540 0.019
R7167 VP.n8064 VP.n8063 0.019
R7168 VP.n7702 VP.n7701 0.019
R7169 VP.n7236 VP.n7235 0.019
R7170 VP.n6863 VP.n6862 0.019
R7171 VP.n6377 VP.n6376 0.019
R7172 VP.n5999 VP.n5998 0.019
R7173 VP.n5521 VP.n5520 0.019
R7174 VP.n5135 VP.n5134 0.019
R7175 VP.n4626 VP.n4625 0.019
R7176 VP.n4229 VP.n4228 0.019
R7177 VP.n3720 VP.n3719 0.019
R7178 VP.n3308 VP.n3307 0.019
R7179 VP.n2780 VP.n2779 0.019
R7180 VP.n2643 VP.n2642 0.019
R7181 VP.n1820 VP.n1819 0.019
R7182 VP.n1382 VP.n1381 0.019
R7183 VP.n836 VP.n835 0.019
R7184 VP.n9715 VP.n9712 0.019
R7185 VP.n11032 VP.n11031 0.019
R7186 VP.n10420 VP.n10419 0.019
R7187 VP.n9850 VP.n9849 0.019
R7188 VP.n9088 VP.n9087 0.019
R7189 VP.n8291 VP.n8290 0.019
R7190 VP.n7474 VP.n7473 0.019
R7191 VP.n6662 VP.n6661 0.019
R7192 VP.n5819 VP.n5818 0.019
R7193 VP.n4982 VP.n4981 0.019
R7194 VP.n4099 VP.n4098 0.019
R7195 VP.n3207 VP.n3206 0.019
R7196 VP.n3777 VP.n3776 0.019
R7197 VP.n4305 VP.n4301 0.019
R7198 VP.n5210 VP.n5206 0.019
R7199 VP.n6075 VP.n6071 0.019
R7200 VP.n6939 VP.n6935 0.019
R7201 VP.n7777 VP.n7773 0.019
R7202 VP.n8616 VP.n8612 0.019
R7203 VP.n9415 VP.n9410 0.019
R7204 VP.n8189 VP.n8188 0.018
R7205 VP.n6479 VP.n6478 0.018
R7206 VP.n4705 VP.n4704 0.018
R7207 VP.n2829 VP.n2828 0.018
R7208 VP.n8735 VP.n8734 0.018
R7209 VP.n9542 VP.n9541 0.018
R7210 VP.n7012 VP.n7011 0.018
R7211 VP.n7850 VP.n7849 0.018
R7212 VP.n8687 VP.n8686 0.018
R7213 VP.n9491 VP.n9490 0.018
R7214 VP.n5233 VP.n5232 0.018
R7215 VP.n6099 VP.n6098 0.018
R7216 VP.n6963 VP.n6962 0.018
R7217 VP.n7801 VP.n7800 0.018
R7218 VP.n8639 VP.n8638 0.018
R7219 VP.n9440 VP.n9439 0.018
R7220 VP.n10719 VP.n10718 0.018
R7221 VP.n9374 VP.n9373 0.018
R7222 VP.n8579 VP.n8578 0.018
R7223 VP.n7740 VP.n7739 0.018
R7224 VP.n6901 VP.n6900 0.018
R7225 VP.n6037 VP.n6036 0.018
R7226 VP.n5173 VP.n5172 0.018
R7227 VP.n4267 VP.n4266 0.018
R7228 VP.n3346 VP.n3345 0.018
R7229 VP.n10449 VP.n10448 0.018
R7230 VP.n9830 VP.n9829 0.018
R7231 VP.n9067 VP.n9066 0.018
R7232 VP.n8270 VP.n8269 0.018
R7233 VP.n7454 VP.n7453 0.018
R7234 VP.n6642 VP.n6641 0.018
R7235 VP.n5798 VP.n5797 0.018
R7236 VP.n4961 VP.n4960 0.018
R7237 VP.n4078 VP.n4077 0.018
R7238 VP.n3185 VP.n3184 0.018
R7239 VP.n2323 VP.n2322 0.018
R7240 VP.n9623 VP.n9622 0.018
R7241 VP.n10024 VP.n10023 0.018
R7242 VP.n7958 VP.n7957 0.018
R7243 VP.n8430 VP.n8429 0.018
R7244 VP.n9230 VP.n9229 0.018
R7245 VP.n9987 VP.n9986 0.018
R7246 VP.n6271 VP.n6270 0.018
R7247 VP.n6752 VP.n6751 0.018
R7248 VP.n7564 VP.n7563 0.018
R7249 VP.n8381 VP.n8380 0.018
R7250 VP.n9180 VP.n9179 0.018
R7251 VP.n9939 VP.n9938 0.018
R7252 VP.n4520 VP.n4519 0.018
R7253 VP.n5024 VP.n5023 0.018
R7254 VP.n5861 VP.n5860 0.018
R7255 VP.n6703 VP.n6702 0.018
R7256 VP.n7515 VP.n7514 0.018
R7257 VP.n8332 VP.n8331 0.018
R7258 VP.n9130 VP.n9129 0.018
R7259 VP.n9891 VP.n9890 0.018
R7260 VP.n8795 VP.n8794 0.017
R7261 VP.n7072 VP.n7071 0.017
R7262 VP.n5293 VP.n5292 0.017
R7263 VP.n3416 VP.n3415 0.017
R7264 VP.n922 VP.n918 0.017
R7265 VP.n1911 VP.n1905 0.017
R7266 VP.n1478 VP.n1476 0.017
R7267 VP.n972 VP.n968 0.017
R7268 VP.n2892 VP.n2886 0.017
R7269 VP.n2578 VP.n2576 0.017
R7270 VP.n1963 VP.n1957 0.017
R7271 VP.n1516 VP.n1514 0.017
R7272 VP.n1022 VP.n1018 0.017
R7273 VP.n3837 VP.n3831 0.017
R7274 VP.n3456 VP.n3454 0.017
R7275 VP.n2944 VP.n2938 0.017
R7276 VP.n2540 VP.n2538 0.017
R7277 VP.n2015 VP.n2009 0.017
R7278 VP.n1554 VP.n1552 0.017
R7279 VP.n1072 VP.n1068 0.017
R7280 VP.n4772 VP.n4766 0.017
R7281 VP.n4373 VP.n4371 0.017
R7282 VP.n3889 VP.n3883 0.017
R7283 VP.n3494 VP.n3492 0.017
R7284 VP.n2996 VP.n2990 0.017
R7285 VP.n2502 VP.n2500 0.017
R7286 VP.n2067 VP.n2061 0.017
R7287 VP.n1592 VP.n1590 0.017
R7288 VP.n1122 VP.n1118 0.017
R7289 VP.n830 VP.n829 0.017
R7290 VP.n312 VP.n311 0.017
R7291 VP.n10634 VP.n10633 0.017
R7292 VP.n10031 VP.n10026 0.017
R7293 VP.n8437 VP.n8432 0.017
R7294 VP.n6759 VP.n6754 0.017
R7295 VP.n5031 VP.n5026 0.017
R7296 VP.n3188 VP.n3187 0.017
R7297 VP.n10058 VP.n10057 0.017
R7298 VP.n10988 VP.n10987 0.017
R7299 VP.n9271 VP.n9270 0.017
R7300 VP.n9631 VP.n9630 0.017
R7301 VP.n10038 VP.n10037 0.017
R7302 VP.n10929 VP.n10928 0.017
R7303 VP.n9565 VP.n9564 0.017
R7304 VP.n7605 VP.n7604 0.017
R7305 VP.n7966 VP.n7965 0.017
R7306 VP.n8444 VP.n8443 0.017
R7307 VP.n8732 VP.n8731 0.017
R7308 VP.n9242 VP.n9241 0.017
R7309 VP.n9539 VP.n9538 0.017
R7310 VP.n9998 VP.n9997 0.017
R7311 VP.n10878 VP.n10877 0.017
R7312 VP.n7873 VP.n7872 0.017
R7313 VP.n8709 VP.n8708 0.017
R7314 VP.n9513 VP.n9512 0.017
R7315 VP.n5902 VP.n5901 0.017
R7316 VP.n6279 VP.n6278 0.017
R7317 VP.n6766 VP.n6765 0.017
R7318 VP.n7009 VP.n7008 0.017
R7319 VP.n7576 VP.n7575 0.017
R7320 VP.n7847 VP.n7846 0.017
R7321 VP.n8393 VP.n8392 0.017
R7322 VP.n8684 VP.n8683 0.017
R7323 VP.n9192 VP.n9191 0.017
R7324 VP.n9488 VP.n9487 0.017
R7325 VP.n9950 VP.n9949 0.017
R7326 VP.n10827 VP.n10826 0.017
R7327 VP.n6122 VP.n6121 0.017
R7328 VP.n6985 VP.n6984 0.017
R7329 VP.n7823 VP.n7822 0.017
R7330 VP.n8661 VP.n8660 0.017
R7331 VP.n9462 VP.n9461 0.017
R7332 VP.n4132 VP.n4131 0.017
R7333 VP.n4528 VP.n4527 0.017
R7334 VP.n5038 VP.n5037 0.017
R7335 VP.n5230 VP.n5229 0.017
R7336 VP.n5873 VP.n5872 0.017
R7337 VP.n6096 VP.n6095 0.017
R7338 VP.n6715 VP.n6714 0.017
R7339 VP.n6960 VP.n6959 0.017
R7340 VP.n7527 VP.n7526 0.017
R7341 VP.n7798 VP.n7797 0.017
R7342 VP.n8344 VP.n8343 0.017
R7343 VP.n8636 VP.n8635 0.017
R7344 VP.n9142 VP.n9141 0.017
R7345 VP.n9437 VP.n9436 0.017
R7346 VP.n9902 VP.n9901 0.017
R7347 VP.n10776 VP.n10775 0.017
R7348 VP.n10730 VP.n10729 0.017
R7349 VP.n9835 VP.n9824 0.017
R7350 VP.n9385 VP.n9384 0.017
R7351 VP.n9072 VP.n9060 0.017
R7352 VP.n8589 VP.n8588 0.017
R7353 VP.n8275 VP.n8263 0.017
R7354 VP.n7750 VP.n7749 0.017
R7355 VP.n7459 VP.n7447 0.017
R7356 VP.n6911 VP.n6910 0.017
R7357 VP.n6647 VP.n6635 0.017
R7358 VP.n6047 VP.n6046 0.017
R7359 VP.n5803 VP.n5791 0.017
R7360 VP.n5183 VP.n5182 0.017
R7361 VP.n4966 VP.n4954 0.017
R7362 VP.n4277 VP.n4276 0.017
R7363 VP.n4083 VP.n4071 0.017
R7364 VP.n3356 VP.n3355 0.017
R7365 VP.n3192 VP.n3178 0.017
R7366 VP.n2328 VP.n2321 0.017
R7367 VP.n2251 VP.n2250 0.017
R7368 VP.n2618 VP.n2617 0.017
R7369 VP.n3329 VP.n3328 0.017
R7370 VP.n4250 VP.n4249 0.017
R7371 VP.n5156 VP.n5155 0.017
R7372 VP.n6020 VP.n6019 0.017
R7373 VP.n6884 VP.n6883 0.017
R7374 VP.n7723 VP.n7722 0.017
R7375 VP.n8562 VP.n8561 0.017
R7376 VP.n9356 VP.n9355 0.017
R7377 VP.n10701 VP.n10700 0.017
R7378 VP.n264 VP.n263 0.017
R7379 VP.n1741 VP.n1740 0.017
R7380 VP.n912 VP.n911 0.017
R7381 VP.n366 VP.n365 0.017
R7382 VP.n903 VP.n902 0.017
R7383 VP.n1337 VP.n1336 0.017
R7384 VP.n2702 VP.n2701 0.017
R7385 VP.n1899 VP.n1898 0.017
R7386 VP.n1474 VP.n1473 0.017
R7387 VP.n962 VP.n961 0.017
R7388 VP.n413 VP.n412 0.017
R7389 VP.n953 VP.n952 0.017
R7390 VP.n1465 VP.n1464 0.017
R7391 VP.n1890 VP.n1889 0.017
R7392 VP.n2313 VP.n2312 0.017
R7393 VP.n3642 VP.n3641 0.017
R7394 VP.n2880 VP.n2879 0.017
R7395 VP.n2574 VP.n2573 0.017
R7396 VP.n1951 VP.n1950 0.017
R7397 VP.n1512 VP.n1511 0.017
R7398 VP.n1012 VP.n1011 0.017
R7399 VP.n460 VP.n459 0.017
R7400 VP.n1003 VP.n1002 0.017
R7401 VP.n1503 VP.n1502 0.017
R7402 VP.n1942 VP.n1941 0.017
R7403 VP.n2565 VP.n2564 0.017
R7404 VP.n2871 VP.n2870 0.017
R7405 VP.n3263 VP.n3262 0.017
R7406 VP.n4548 VP.n4547 0.017
R7407 VP.n3825 VP.n3824 0.017
R7408 VP.n3452 VP.n3451 0.017
R7409 VP.n2932 VP.n2931 0.017
R7410 VP.n2536 VP.n2535 0.017
R7411 VP.n2003 VP.n2002 0.017
R7412 VP.n1550 VP.n1549 0.017
R7413 VP.n1062 VP.n1061 0.017
R7414 VP.n507 VP.n506 0.017
R7415 VP.n1053 VP.n1052 0.017
R7416 VP.n1541 VP.n1540 0.017
R7417 VP.n1994 VP.n1993 0.017
R7418 VP.n2527 VP.n2526 0.017
R7419 VP.n2923 VP.n2922 0.017
R7420 VP.n3443 VP.n3442 0.017
R7421 VP.n3816 VP.n3815 0.017
R7422 VP.n4184 VP.n4183 0.017
R7423 VP.n5443 VP.n5442 0.017
R7424 VP.n4760 VP.n4759 0.017
R7425 VP.n4369 VP.n4368 0.017
R7426 VP.n3877 VP.n3876 0.017
R7427 VP.n3490 VP.n3489 0.017
R7428 VP.n2984 VP.n2983 0.017
R7429 VP.n2498 VP.n2497 0.017
R7430 VP.n2055 VP.n2054 0.017
R7431 VP.n1588 VP.n1587 0.017
R7432 VP.n1112 VP.n1111 0.017
R7433 VP.n554 VP.n553 0.017
R7434 VP.n1103 VP.n1102 0.017
R7435 VP.n1579 VP.n1578 0.017
R7436 VP.n2046 VP.n2045 0.017
R7437 VP.n2489 VP.n2488 0.017
R7438 VP.n2975 VP.n2974 0.017
R7439 VP.n3481 VP.n3480 0.017
R7440 VP.n3868 VP.n3867 0.017
R7441 VP.n4360 VP.n4359 0.017
R7442 VP.n4751 VP.n4750 0.017
R7443 VP.n5090 VP.n5089 0.017
R7444 VP.n6299 VP.n6298 0.017
R7445 VP.n601 VP.n600 0.017
R7446 VP.n1153 VP.n1152 0.017
R7447 VP.n1617 VP.n1616 0.017
R7448 VP.n2098 VP.n2097 0.017
R7449 VP.n2457 VP.n2456 0.017
R7450 VP.n3027 VP.n3026 0.017
R7451 VP.n3519 VP.n3518 0.017
R7452 VP.n3920 VP.n3919 0.017
R7453 VP.n4398 VP.n4397 0.017
R7454 VP.n4803 VP.n4802 0.017
R7455 VP.n5320 VP.n5319 0.017
R7456 VP.n5640 VP.n5639 0.017
R7457 VP.n5954 VP.n5953 0.017
R7458 VP.n7158 VP.n7157 0.017
R7459 VP.n641 VP.n640 0.017
R7460 VP.n1191 VP.n1190 0.017
R7461 VP.n1649 VP.n1648 0.017
R7462 VP.n2139 VP.n2138 0.017
R7463 VP.n2425 VP.n2424 0.017
R7464 VP.n3068 VP.n3067 0.017
R7465 VP.n3551 VP.n3550 0.017
R7466 VP.n3961 VP.n3960 0.017
R7467 VP.n4430 VP.n4429 0.017
R7468 VP.n4844 VP.n4843 0.017
R7469 VP.n5352 VP.n5351 0.017
R7470 VP.n5681 VP.n5680 0.017
R7471 VP.n6180 VP.n6179 0.017
R7472 VP.n6525 VP.n6524 0.017
R7473 VP.n6818 VP.n6817 0.017
R7474 VP.n7986 VP.n7985 0.017
R7475 VP.n671 VP.n670 0.017
R7476 VP.n1231 VP.n1230 0.017
R7477 VP.n1681 VP.n1680 0.017
R7478 VP.n2180 VP.n2179 0.017
R7479 VP.n2393 VP.n2392 0.017
R7480 VP.n3109 VP.n3108 0.017
R7481 VP.n3583 VP.n3582 0.017
R7482 VP.n4002 VP.n4001 0.017
R7483 VP.n4462 VP.n4461 0.017
R7484 VP.n4885 VP.n4884 0.017
R7485 VP.n5384 VP.n5383 0.017
R7486 VP.n5722 VP.n5721 0.017
R7487 VP.n6212 VP.n6211 0.017
R7488 VP.n6566 VP.n6565 0.017
R7489 VP.n7099 VP.n7098 0.017
R7490 VP.n7378 VP.n7377 0.017
R7491 VP.n7657 VP.n7656 0.017
R7492 VP.n9652 VP.n9651 0.017
R7493 VP.n703 VP.n702 0.017
R7494 VP.n1272 VP.n1271 0.017
R7495 VP.n1713 VP.n1712 0.017
R7496 VP.n2221 VP.n2220 0.017
R7497 VP.n2361 VP.n2360 0.017
R7498 VP.n3150 VP.n3149 0.017
R7499 VP.n3615 VP.n3614 0.017
R7500 VP.n4043 VP.n4042 0.017
R7501 VP.n4494 VP.n4493 0.017
R7502 VP.n4926 VP.n4925 0.017
R7503 VP.n5416 VP.n5415 0.017
R7504 VP.n5763 VP.n5762 0.017
R7505 VP.n6244 VP.n6243 0.017
R7506 VP.n6607 VP.n6606 0.017
R7507 VP.n7131 VP.n7130 0.017
R7508 VP.n7419 VP.n7418 0.017
R7509 VP.n7931 VP.n7930 0.017
R7510 VP.n8235 VP.n8234 0.017
R7511 VP.n8496 VP.n8495 0.017
R7512 VP.n8818 VP.n8817 0.017
R7513 VP.n279 VP.n278 0.017
R7514 VP.n795 VP.n794 0.017
R7515 VP.n1351 VP.n1350 0.017
R7516 VP.n1781 VP.n1780 0.017
R7517 VP.n2668 VP.n2667 0.017
R7518 VP.n2741 VP.n2740 0.017
R7519 VP.n3277 VP.n3276 0.017
R7520 VP.n3681 VP.n3680 0.017
R7521 VP.n4198 VP.n4197 0.017
R7522 VP.n4590 VP.n4589 0.017
R7523 VP.n5104 VP.n5103 0.017
R7524 VP.n5482 VP.n5481 0.017
R7525 VP.n5968 VP.n5967 0.017
R7526 VP.n6338 VP.n6337 0.017
R7527 VP.n6832 VP.n6831 0.017
R7528 VP.n7197 VP.n7196 0.017
R7529 VP.n7671 VP.n7670 0.017
R7530 VP.n8025 VP.n8024 0.017
R7531 VP.n8510 VP.n8509 0.017
R7532 VP.n8871 VP.n8870 0.017
R7533 VP.n11024 VP.n11023 0.017
R7534 VP.n4303 VP.n4302 0.017
R7535 VP.n5208 VP.n5207 0.017
R7536 VP.n6073 VP.n6072 0.017
R7537 VP.n6937 VP.n6936 0.017
R7538 VP.n7775 VP.n7774 0.017
R7539 VP.n8614 VP.n8613 0.017
R7540 VP.n9412 VP.n9411 0.017
R7541 VP.n9562 VP.n9561 0.016
R7542 VP.n7870 VP.n7869 0.016
R7543 VP.n6119 VP.n6118 0.016
R7544 VP.n2615 VP.n2614 0.016
R7545 VP.n4300 VP.n4299 0.016
R7546 VP.n9563 VP.n9562 0.016
R7547 VP.n7871 VP.n7870 0.016
R7548 VP.n8707 VP.n8706 0.016
R7549 VP.n9511 VP.n9510 0.016
R7550 VP.n6120 VP.n6119 0.016
R7551 VP.n6983 VP.n6982 0.016
R7552 VP.n7821 VP.n7820 0.016
R7553 VP.n8659 VP.n8658 0.016
R7554 VP.n9460 VP.n9459 0.016
R7555 VP.n2616 VP.n2615 0.016
R7556 VP.n3327 VP.n3326 0.016
R7557 VP.n4248 VP.n4247 0.016
R7558 VP.n5154 VP.n5153 0.016
R7559 VP.n6018 VP.n6017 0.016
R7560 VP.n6882 VP.n6881 0.016
R7561 VP.n7721 VP.n7720 0.016
R7562 VP.n8560 VP.n8559 0.016
R7563 VP.n9354 VP.n9353 0.016
R7564 VP.n10697 VP.n10696 0.016
R7565 VP.n4301 VP.n4300 0.016
R7566 VP.n5206 VP.n5205 0.016
R7567 VP.n6071 VP.n6070 0.016
R7568 VP.n6935 VP.n6934 0.016
R7569 VP.n7773 VP.n7772 0.016
R7570 VP.n8612 VP.n8611 0.016
R7571 VP.n9410 VP.n9409 0.016
R7572 VP.n10627 VP.n10626 0.016
R7573 VP.n10589 VP.n10588 0.016
R7574 VP.n10554 VP.n10553 0.016
R7575 VP.n10519 VP.n10518 0.016
R7576 VP.n10484 VP.n10483 0.016
R7577 VP.n10454 VP.n10443 0.016
R7578 VP.n10687 VP.n10686 0.016
R7579 VP.n8955 VP.n8954 0.016
R7580 VP.n8111 VP.n8110 0.016
R7581 VP.n7283 VP.n7282 0.016
R7582 VP.n6424 VP.n6423 0.016
R7583 VP.n5568 VP.n5567 0.016
R7584 VP.n4673 VP.n4672 0.016
R7585 VP.n9268 VP.n9266 0.016
R7586 VP.n9795 VP.n9794 0.016
R7587 VP.n9990 VP.n9989 0.016
R7588 VP.n9234 VP.n9233 0.016
R7589 VP.n7602 VP.n7600 0.016
R7590 VP.n9773 VP.n9772 0.016
R7591 VP.n9000 VP.n8999 0.016
R7592 VP.n8156 VP.n8155 0.016
R7593 VP.n9942 VP.n9941 0.016
R7594 VP.n9184 VP.n9183 0.016
R7595 VP.n8385 VP.n8384 0.016
R7596 VP.n7568 VP.n7567 0.016
R7597 VP.n5899 VP.n5897 0.016
R7598 VP.n9751 VP.n9750 0.016
R7599 VP.n8977 VP.n8976 0.016
R7600 VP.n8133 VP.n8132 0.016
R7601 VP.n7305 VP.n7304 0.016
R7602 VP.n6446 VP.n6445 0.016
R7603 VP.n9894 VP.n9893 0.016
R7604 VP.n9134 VP.n9133 0.016
R7605 VP.n8336 VP.n8335 0.016
R7606 VP.n7519 VP.n7518 0.016
R7607 VP.n6707 VP.n6706 0.016
R7608 VP.n5865 VP.n5864 0.016
R7609 VP.n4129 VP.n4127 0.016
R7610 VP.n10445 VP.n10444 0.016
R7611 VP.n9826 VP.n9825 0.016
R7612 VP.n9063 VP.n9062 0.016
R7613 VP.n8266 VP.n8265 0.016
R7614 VP.n7450 VP.n7449 0.016
R7615 VP.n6638 VP.n6637 0.016
R7616 VP.n5794 VP.n5793 0.016
R7617 VP.n4957 VP.n4956 0.016
R7618 VP.n4074 VP.n4073 0.016
R7619 VP.n2257 VP.n2255 0.016
R7620 VP.n9729 VP.n9728 0.016
R7621 VP.n8928 VP.n8927 0.016
R7622 VP.n8084 VP.n8083 0.016
R7623 VP.n7256 VP.n7255 0.016
R7624 VP.n6397 VP.n6396 0.016
R7625 VP.n5541 VP.n5540 0.016
R7626 VP.n4646 VP.n4645 0.016
R7627 VP.n3740 VP.n3739 0.016
R7628 VP.n2800 VP.n2799 0.016
R7629 VP.n10200 VP.n10199 0.016
R7630 VP.n10317 VP.n10316 0.016
R7631 VP.n10198 VP.n10197 0.016
R7632 VP.n10315 VP.n10314 0.016
R7633 VP.t8 VP.n10177 0.016
R7634 VP.n9836 VP.n9821 0.016
R7635 VP.n9073 VP.n9057 0.016
R7636 VP.n8276 VP.n8260 0.016
R7637 VP.n7460 VP.n7444 0.016
R7638 VP.n6648 VP.n6632 0.016
R7639 VP.n5804 VP.n5788 0.016
R7640 VP.n4967 VP.n4951 0.016
R7641 VP.n4084 VP.n4068 0.016
R7642 VP.n3193 VP.n3175 0.016
R7643 VP.n10640 VP.n10639 0.016
R7644 VP.n10039 VP.n10021 0.016
R7645 VP.n8445 VP.n8427 0.016
R7646 VP.n9243 VP.n9227 0.016
R7647 VP.n9999 VP.n9984 0.016
R7648 VP.n6767 VP.n6749 0.016
R7649 VP.n7577 VP.n7561 0.016
R7650 VP.n8394 VP.n8378 0.016
R7651 VP.n9193 VP.n9177 0.016
R7652 VP.n9951 VP.n9936 0.016
R7653 VP.n5039 VP.n5021 0.016
R7654 VP.n5874 VP.n5858 0.016
R7655 VP.n6716 VP.n6700 0.016
R7656 VP.n7528 VP.n7512 0.016
R7657 VP.n8345 VP.n8329 0.016
R7658 VP.n9143 VP.n9127 0.016
R7659 VP.n9903 VP.n9888 0.016
R7660 VP.n265 VP.n253 0.016
R7661 VP.n367 VP.n355 0.016
R7662 VP.n414 VP.n402 0.016
R7663 VP.n461 VP.n449 0.016
R7664 VP.n508 VP.n496 0.016
R7665 VP.n555 VP.n543 0.016
R7666 VP.n602 VP.n590 0.016
R7667 VP.n642 VP.n630 0.016
R7668 VP.n672 VP.n660 0.016
R7669 VP.n704 VP.n692 0.016
R7670 VP.n772 VP.n771 0.015
R7671 VP.n1761 VP.n1760 0.015
R7672 VP.n2722 VP.n2721 0.015
R7673 VP.n3662 VP.n3661 0.015
R7674 VP.n4568 VP.n4567 0.015
R7675 VP.n5463 VP.n5462 0.015
R7676 VP.n6319 VP.n6318 0.015
R7677 VP.n7178 VP.n7177 0.015
R7678 VP.n8006 VP.n8005 0.015
R7679 VP.n8840 VP.n8839 0.015
R7680 VP.n10111 VP.n10110 0.015
R7681 VP.n10121 VP.n10120 0.015
R7682 VP.n748 VP.n747 0.015
R7683 VP.t8 VP.n10288 0.015
R7684 VP.t8 VP.n10260 0.015
R7685 VP.t8 VP.n10232 0.015
R7686 VP.n8180 VP.n8179 0.015
R7687 VP.n6470 VP.n6469 0.015
R7688 VP.n4696 VP.n4695 0.015
R7689 VP.n152 VP.n151 0.015
R7690 VP.n10308 VP.n10307 0.015
R7691 VP.n10292 VP.n10291 0.015
R7692 VP.n10280 VP.n10279 0.015
R7693 VP.n10264 VP.n10263 0.015
R7694 VP.n10252 VP.n10251 0.015
R7695 VP.n10236 VP.n10235 0.015
R7696 VP.n10224 VP.n10223 0.015
R7697 VP.n10208 VP.n10207 0.015
R7698 VP.n10186 VP.n10185 0.015
R7699 VP.n380 VP.n378 0.015
R7700 VP.n427 VP.n425 0.015
R7701 VP.n474 VP.n472 0.015
R7702 VP.n521 VP.n519 0.015
R7703 VP.n568 VP.n566 0.015
R7704 VP.n10188 VP.n10187 0.015
R7705 VP.n10358 VP.n10357 0.015
R7706 VP.n10144 VP.n10135 0.015
R7707 VP.n305 VP.n304 0.014
R7708 VP.n1442 VP.n1422 0.014
R7709 VP.n10070 VP.n10069 0.014
R7710 VP.n11004 VP.n11003 0.014
R7711 VP.n10641 VP.n10640 0.014
R7712 VP.n10945 VP.n10944 0.014
R7713 VP.n9043 VP.n9031 0.014
R7714 VP.n8743 VP.n8742 0.014
R7715 VP.n9550 VP.n9549 0.014
R7716 VP.n10894 VP.n10893 0.014
R7717 VP.n9966 VP.n9964 0.014
R7718 VP.n9209 VP.n9207 0.014
R7719 VP.n8409 VP.n8407 0.014
R7720 VP.n7348 VP.n7336 0.014
R7721 VP.n7020 VP.n7019 0.014
R7722 VP.n7858 VP.n7857 0.014
R7723 VP.n8695 VP.n8694 0.014
R7724 VP.n9499 VP.n9498 0.014
R7725 VP.n10843 VP.n10842 0.014
R7726 VP.n9918 VP.n9916 0.014
R7727 VP.n9159 VP.n9157 0.014
R7728 VP.n8360 VP.n8358 0.014
R7729 VP.n7543 VP.n7541 0.014
R7730 VP.n6731 VP.n6729 0.014
R7731 VP.n5610 VP.n5598 0.014
R7732 VP.n5241 VP.n5240 0.014
R7733 VP.n6107 VP.n6106 0.014
R7734 VP.n6971 VP.n6970 0.014
R7735 VP.n7809 VP.n7808 0.014
R7736 VP.n8647 VP.n8646 0.014
R7737 VP.n9448 VP.n9447 0.014
R7738 VP.n10792 VP.n10791 0.014
R7739 VP.n9870 VP.n9868 0.014
R7740 VP.n9109 VP.n9107 0.014
R7741 VP.n8311 VP.n8309 0.014
R7742 VP.n7494 VP.n7492 0.014
R7743 VP.n6682 VP.n6680 0.014
R7744 VP.n5840 VP.n5838 0.014
R7745 VP.n5003 VP.n5001 0.014
R7746 VP.n10727 VP.n10726 0.014
R7747 VP.n9382 VP.n9381 0.014
R7748 VP.n8587 VP.n8586 0.014
R7749 VP.n7748 VP.n7747 0.014
R7750 VP.n6909 VP.n6908 0.014
R7751 VP.n6045 VP.n6044 0.014
R7752 VP.n5181 VP.n5180 0.014
R7753 VP.n4275 VP.n4274 0.014
R7754 VP.n3354 VP.n3353 0.014
R7755 VP.n873 VP.n862 0.014
R7756 VP.n1860 VP.n1848 0.014
R7757 VP.n754 VP.n753 0.014
R7758 VP.n758 VP.n752 0.014
R7759 VP.n899 VP.n898 0.014
R7760 VP.n1333 VP.n1332 0.014
R7761 VP.n949 VP.n948 0.014
R7762 VP.n1461 VP.n1460 0.014
R7763 VP.n1886 VP.n1885 0.014
R7764 VP.n2309 VP.n2308 0.014
R7765 VP.n999 VP.n998 0.014
R7766 VP.n1499 VP.n1498 0.014
R7767 VP.n1938 VP.n1937 0.014
R7768 VP.n2561 VP.n2560 0.014
R7769 VP.n2867 VP.n2866 0.014
R7770 VP.n3259 VP.n3258 0.014
R7771 VP.n1049 VP.n1048 0.014
R7772 VP.n1537 VP.n1536 0.014
R7773 VP.n1990 VP.n1989 0.014
R7774 VP.n2523 VP.n2522 0.014
R7775 VP.n2919 VP.n2918 0.014
R7776 VP.n3439 VP.n3438 0.014
R7777 VP.n3812 VP.n3811 0.014
R7778 VP.n4180 VP.n4179 0.014
R7779 VP.n1099 VP.n1098 0.014
R7780 VP.n1575 VP.n1574 0.014
R7781 VP.n2042 VP.n2041 0.014
R7782 VP.n2485 VP.n2484 0.014
R7783 VP.n2971 VP.n2970 0.014
R7784 VP.n3477 VP.n3476 0.014
R7785 VP.n3864 VP.n3863 0.014
R7786 VP.n4356 VP.n4355 0.014
R7787 VP.n4747 VP.n4746 0.014
R7788 VP.n5086 VP.n5085 0.014
R7789 VP.n1149 VP.n1148 0.014
R7790 VP.n1613 VP.n1612 0.014
R7791 VP.n2094 VP.n2093 0.014
R7792 VP.n2453 VP.n2452 0.014
R7793 VP.n3023 VP.n3022 0.014
R7794 VP.n3515 VP.n3514 0.014
R7795 VP.n3916 VP.n3915 0.014
R7796 VP.n4394 VP.n4393 0.014
R7797 VP.n4799 VP.n4798 0.014
R7798 VP.n5316 VP.n5315 0.014
R7799 VP.n5636 VP.n5635 0.014
R7800 VP.n5950 VP.n5949 0.014
R7801 VP.n1187 VP.n1186 0.014
R7802 VP.n1645 VP.n1644 0.014
R7803 VP.n2135 VP.n2134 0.014
R7804 VP.n2421 VP.n2420 0.014
R7805 VP.n3064 VP.n3063 0.014
R7806 VP.n3547 VP.n3546 0.014
R7807 VP.n3957 VP.n3956 0.014
R7808 VP.n4426 VP.n4425 0.014
R7809 VP.n4840 VP.n4839 0.014
R7810 VP.n5348 VP.n5347 0.014
R7811 VP.n5677 VP.n5676 0.014
R7812 VP.n6176 VP.n6175 0.014
R7813 VP.n6521 VP.n6520 0.014
R7814 VP.n6814 VP.n6813 0.014
R7815 VP.n1227 VP.n1226 0.014
R7816 VP.n1677 VP.n1676 0.014
R7817 VP.n2176 VP.n2175 0.014
R7818 VP.n2389 VP.n2388 0.014
R7819 VP.n3105 VP.n3104 0.014
R7820 VP.n3579 VP.n3578 0.014
R7821 VP.n3998 VP.n3997 0.014
R7822 VP.n4458 VP.n4457 0.014
R7823 VP.n4881 VP.n4880 0.014
R7824 VP.n5380 VP.n5379 0.014
R7825 VP.n5718 VP.n5717 0.014
R7826 VP.n6208 VP.n6207 0.014
R7827 VP.n6562 VP.n6561 0.014
R7828 VP.n7095 VP.n7094 0.014
R7829 VP.n7374 VP.n7373 0.014
R7830 VP.n7653 VP.n7652 0.014
R7831 VP.n8856 VP.n8854 0.014
R7832 VP.n1268 VP.n1267 0.014
R7833 VP.n1709 VP.n1708 0.014
R7834 VP.n2217 VP.n2216 0.014
R7835 VP.n2357 VP.n2356 0.014
R7836 VP.n3146 VP.n3145 0.014
R7837 VP.n3611 VP.n3610 0.014
R7838 VP.n4039 VP.n4038 0.014
R7839 VP.n4490 VP.n4489 0.014
R7840 VP.n4922 VP.n4921 0.014
R7841 VP.n5412 VP.n5411 0.014
R7842 VP.n5759 VP.n5758 0.014
R7843 VP.n6240 VP.n6239 0.014
R7844 VP.n6603 VP.n6602 0.014
R7845 VP.n7127 VP.n7126 0.014
R7846 VP.n7415 VP.n7414 0.014
R7847 VP.n7927 VP.n7926 0.014
R7848 VP.n8231 VP.n8230 0.014
R7849 VP.n8492 VP.n8491 0.014
R7850 VP.n286 VP.n285 0.014
R7851 VP.n814 VP.n813 0.014
R7852 VP.n1364 VP.n1363 0.014
R7853 VP.n1800 VP.n1799 0.014
R7854 VP.n2681 VP.n2680 0.014
R7855 VP.n2760 VP.n2759 0.014
R7856 VP.n3290 VP.n3289 0.014
R7857 VP.n3700 VP.n3699 0.014
R7858 VP.n4211 VP.n4210 0.014
R7859 VP.n4609 VP.n4608 0.014
R7860 VP.n5117 VP.n5116 0.014
R7861 VP.n5501 VP.n5500 0.014
R7862 VP.n5981 VP.n5980 0.014
R7863 VP.n6357 VP.n6356 0.014
R7864 VP.n6845 VP.n6844 0.014
R7865 VP.n7216 VP.n7215 0.014
R7866 VP.n7684 VP.n7683 0.014
R7867 VP.n8044 VP.n8043 0.014
R7868 VP.n8523 VP.n8522 0.014
R7869 VP.n8888 VP.n8887 0.014
R7870 VP.n9719 VP.n9697 0.014
R7871 VP.n9343 VP.n9332 0.014
R7872 VP.n8918 VP.n8906 0.014
R7873 VP.n8549 VP.n8539 0.014
R7874 VP.n8074 VP.n8062 0.014
R7875 VP.n7710 VP.n7700 0.014
R7876 VP.n7246 VP.n7234 0.014
R7877 VP.n6871 VP.n6861 0.014
R7878 VP.n6387 VP.n6375 0.014
R7879 VP.n6007 VP.n5997 0.014
R7880 VP.n5531 VP.n5519 0.014
R7881 VP.n5143 VP.n5133 0.014
R7882 VP.n4636 VP.n4624 0.014
R7883 VP.n4237 VP.n4227 0.014
R7884 VP.n3730 VP.n3718 0.014
R7885 VP.n3316 VP.n3306 0.014
R7886 VP.n2790 VP.n2778 0.014
R7887 VP.n2651 VP.n2641 0.014
R7888 VP.n1830 VP.n1818 0.014
R7889 VP.n1390 VP.n1380 0.014
R7890 VP.n847 VP.n834 0.014
R7891 VP.n9715 VP.n9714 0.014
R7892 VP.n10429 VP.n10418 0.014
R7893 VP.n9850 VP.n9848 0.014
R7894 VP.n9088 VP.n9086 0.014
R7895 VP.n8291 VP.n8289 0.014
R7896 VP.n7474 VP.n7472 0.014
R7897 VP.n6662 VP.n6660 0.014
R7898 VP.n5819 VP.n5817 0.014
R7899 VP.n4982 VP.n4980 0.014
R7900 VP.n4099 VP.n4097 0.014
R7901 VP.n3207 VP.n3205 0.014
R7902 VP.n3781 VP.n3775 0.014
R7903 VP.n2261 VP.n2260 0.014
R7904 VP.n1746 VP.n1745 0.014
R7905 VP.n923 VP.n922 0.014
R7906 VP.n2707 VP.n2706 0.014
R7907 VP.n1912 VP.n1911 0.014
R7908 VP.n1479 VP.n1478 0.014
R7909 VP.n973 VP.n972 0.014
R7910 VP.n3647 VP.n3646 0.014
R7911 VP.n2893 VP.n2892 0.014
R7912 VP.n2579 VP.n2578 0.014
R7913 VP.n1964 VP.n1963 0.014
R7914 VP.n1517 VP.n1516 0.014
R7915 VP.n1023 VP.n1022 0.014
R7916 VP.n4553 VP.n4552 0.014
R7917 VP.n3838 VP.n3837 0.014
R7918 VP.n3457 VP.n3456 0.014
R7919 VP.n2945 VP.n2944 0.014
R7920 VP.n2541 VP.n2540 0.014
R7921 VP.n2016 VP.n2015 0.014
R7922 VP.n1555 VP.n1554 0.014
R7923 VP.n1073 VP.n1072 0.014
R7924 VP.n5448 VP.n5447 0.014
R7925 VP.n4773 VP.n4772 0.014
R7926 VP.n4374 VP.n4373 0.014
R7927 VP.n3890 VP.n3889 0.014
R7928 VP.n3495 VP.n3494 0.014
R7929 VP.n2997 VP.n2996 0.014
R7930 VP.n2503 VP.n2502 0.014
R7931 VP.n2068 VP.n2067 0.014
R7932 VP.n1593 VP.n1592 0.014
R7933 VP.n1123 VP.n1122 0.014
R7934 VP.n6304 VP.n6303 0.014
R7935 VP.n7163 VP.n7162 0.014
R7936 VP.n7991 VP.n7990 0.014
R7937 VP.n10332 VP.n10331 0.014
R7938 VP.n9317 VP.n9311 0.014
R7939 VP.n8851 VP.n8850 0.013
R7940 VP.n9718 VP.n9717 0.013
R7941 VP.n9697 VP.n9691 0.013
R7942 VP.n9332 VP.n9328 0.013
R7943 VP.n8906 VP.n8901 0.013
R7944 VP.n8539 VP.n8535 0.013
R7945 VP.n8062 VP.n8057 0.013
R7946 VP.n7700 VP.n7696 0.013
R7947 VP.n7234 VP.n7229 0.013
R7948 VP.n6861 VP.n6857 0.013
R7949 VP.n6375 VP.n6370 0.013
R7950 VP.n5997 VP.n5993 0.013
R7951 VP.n5519 VP.n5514 0.013
R7952 VP.n5133 VP.n5129 0.013
R7953 VP.n4624 VP.n4619 0.013
R7954 VP.n4227 VP.n4223 0.013
R7955 VP.n3718 VP.n3713 0.013
R7956 VP.n3306 VP.n3302 0.013
R7957 VP.n2778 VP.n2773 0.013
R7958 VP.n2641 VP.n2637 0.013
R7959 VP.n1818 VP.n1813 0.013
R7960 VP.n1380 VP.n1376 0.013
R7961 VP.n834 VP.n827 0.013
R7962 VP.n145 VP.n144 0.013
R7963 VP.n9717 VP.n9716 0.013
R7964 VP.n10418 VP.n10417 0.013
R7965 VP.n9023 VP.n9022 0.013
R7966 VP.n7328 VP.n7327 0.013
R7967 VP.n5590 VP.n5589 0.013
R7968 VP.n9694 VP.n9693 0.013
R7969 VP.n9330 VP.n9329 0.013
R7970 VP.n8904 VP.n8903 0.013
R7971 VP.n8537 VP.n8536 0.013
R7972 VP.n8060 VP.n8059 0.013
R7973 VP.n7698 VP.n7697 0.013
R7974 VP.n7232 VP.n7231 0.013
R7975 VP.n6859 VP.n6858 0.013
R7976 VP.n6373 VP.n6372 0.013
R7977 VP.n5995 VP.n5994 0.013
R7978 VP.n5517 VP.n5516 0.013
R7979 VP.n5131 VP.n5130 0.013
R7980 VP.n4622 VP.n4621 0.013
R7981 VP.n4225 VP.n4224 0.013
R7982 VP.n3716 VP.n3715 0.013
R7983 VP.n3304 VP.n3303 0.013
R7984 VP.n2776 VP.n2775 0.013
R7985 VP.n2639 VP.n2638 0.013
R7986 VP.n1816 VP.n1815 0.013
R7987 VP.n1378 VP.n1377 0.013
R7988 VP.n742 VP.n741 0.013
R7989 VP.n385 VP.n384 0.013
R7990 VP.n432 VP.n431 0.013
R7991 VP.n479 VP.n478 0.013
R7992 VP.n526 VP.n525 0.013
R7993 VP.n573 VP.n572 0.013
R7994 VP.n613 VP.n612 0.013
R7995 VP.n715 VP.n714 0.013
R7996 VP.n9273 VP.n9272 0.012
R7997 VP.n9633 VP.n9632 0.012
R7998 VP.n10040 VP.n10039 0.012
R7999 VP.n7607 VP.n7606 0.012
R8000 VP.n7968 VP.n7967 0.012
R8001 VP.n8446 VP.n8445 0.012
R8002 VP.n9244 VP.n9243 0.012
R8003 VP.n10000 VP.n9999 0.012
R8004 VP.n5904 VP.n5903 0.012
R8005 VP.n6281 VP.n6280 0.012
R8006 VP.n6768 VP.n6767 0.012
R8007 VP.n7578 VP.n7577 0.012
R8008 VP.n8395 VP.n8394 0.012
R8009 VP.n9194 VP.n9193 0.012
R8010 VP.n9952 VP.n9951 0.012
R8011 VP.n4134 VP.n4133 0.012
R8012 VP.n4530 VP.n4529 0.012
R8013 VP.n5040 VP.n5039 0.012
R8014 VP.n5875 VP.n5874 0.012
R8015 VP.n6717 VP.n6716 0.012
R8016 VP.n7529 VP.n7528 0.012
R8017 VP.n8346 VP.n8345 0.012
R8018 VP.n9144 VP.n9143 0.012
R8019 VP.n9904 VP.n9903 0.012
R8020 VP.n758 VP.n265 0.012
R8021 VP.n392 VP.n367 0.012
R8022 VP.n439 VP.n414 0.012
R8023 VP.n486 VP.n461 0.012
R8024 VP.n533 VP.n508 0.012
R8025 VP.n580 VP.n555 0.012
R8026 VP.n620 VP.n602 0.012
R8027 VP.n650 VP.n642 0.012
R8028 VP.n682 VP.n672 0.012
R8029 VP.n722 VP.n704 0.012
R8030 VP.n7429 VP.n7427 0.012
R8031 VP.n6617 VP.n6615 0.012
R8032 VP.n5773 VP.n5771 0.012
R8033 VP.n4936 VP.n4934 0.012
R8034 VP.n4053 VP.n4051 0.012
R8035 VP.n3160 VP.n3158 0.012
R8036 VP.n2231 VP.n2229 0.012
R8037 VP.n8245 VP.n8243 0.012
R8038 VP.n1282 VP.n1280 0.012
R8039 VP.n855 VP.n854 0.012
R8040 VP.n1840 VP.n1839 0.012
R8041 VP.n3767 VP.n3766 0.012
R8042 VP.n9269 VP.n9268 0.012
R8043 VP.n9624 VP.n9623 0.012
R8044 VP.n10026 VP.n10025 0.012
R8045 VP.n10603 VP.n10602 0.012
R8046 VP.n7908 VP.n7903 0.012
R8047 VP.n7603 VP.n7602 0.012
R8048 VP.n7959 VP.n7958 0.012
R8049 VP.n8432 VP.n8431 0.012
R8050 VP.n9233 VP.n9232 0.012
R8051 VP.n9231 VP.n9230 0.012
R8052 VP.n9988 VP.n9987 0.012
R8053 VP.n10568 VP.n10567 0.012
R8054 VP.n6157 VP.n6152 0.012
R8055 VP.n5900 VP.n5899 0.012
R8056 VP.n6272 VP.n6271 0.012
R8057 VP.n6754 VP.n6753 0.012
R8058 VP.n7567 VP.n7566 0.012
R8059 VP.n7565 VP.n7564 0.012
R8060 VP.n8384 VP.n8383 0.012
R8061 VP.n8382 VP.n8381 0.012
R8062 VP.n9183 VP.n9182 0.012
R8063 VP.n9181 VP.n9180 0.012
R8064 VP.n9940 VP.n9939 0.012
R8065 VP.n10533 VP.n10532 0.012
R8066 VP.n4337 VP.n4332 0.012
R8067 VP.n4130 VP.n4129 0.012
R8068 VP.n4521 VP.n4520 0.012
R8069 VP.n5026 VP.n5025 0.012
R8070 VP.n5864 VP.n5863 0.012
R8071 VP.n5862 VP.n5861 0.012
R8072 VP.n6706 VP.n6705 0.012
R8073 VP.n6704 VP.n6703 0.012
R8074 VP.n7518 VP.n7517 0.012
R8075 VP.n7516 VP.n7515 0.012
R8076 VP.n8335 VP.n8334 0.012
R8077 VP.n8333 VP.n8332 0.012
R8078 VP.n9133 VP.n9132 0.012
R8079 VP.n9131 VP.n9130 0.012
R8080 VP.n9892 VP.n9891 0.012
R8081 VP.n10498 VP.n10497 0.012
R8082 VP.n10450 VP.n10449 0.012
R8083 VP.n9831 VP.n9830 0.012
R8084 VP.n9068 VP.n9067 0.012
R8085 VP.n9062 VP.n9061 0.012
R8086 VP.n8271 VP.n8270 0.012
R8087 VP.n8265 VP.n8264 0.012
R8088 VP.n7455 VP.n7454 0.012
R8089 VP.n7449 VP.n7448 0.012
R8090 VP.n6643 VP.n6642 0.012
R8091 VP.n6637 VP.n6636 0.012
R8092 VP.n5799 VP.n5798 0.012
R8093 VP.n5793 VP.n5792 0.012
R8094 VP.n4962 VP.n4961 0.012
R8095 VP.n4956 VP.n4955 0.012
R8096 VP.n4079 VP.n4078 0.012
R8097 VP.n4073 VP.n4072 0.012
R8098 VP.n3187 VP.n3186 0.012
R8099 VP.n2324 VP.n2323 0.012
R8100 VP.n2258 VP.n2257 0.012
R8101 VP.n380 VP.n379 0.012
R8102 VP.n392 VP.n391 0.012
R8103 VP.n427 VP.n426 0.012
R8104 VP.n439 VP.n438 0.012
R8105 VP.n474 VP.n473 0.012
R8106 VP.n486 VP.n485 0.012
R8107 VP.n521 VP.n520 0.012
R8108 VP.n533 VP.n532 0.012
R8109 VP.n568 VP.n567 0.012
R8110 VP.n580 VP.n579 0.012
R8111 VP.n10678 VP.n10677 0.012
R8112 VP.n303 VP.n301 0.012
R8113 VP.n2609 VP.n2606 0.012
R8114 VP.n9407 VP.n9406 0.012
R8115 VP.n10092 VP.n10091 0.012
R8116 VP.n9970 VP.n9969 0.012
R8117 VP.n9213 VP.n9212 0.012
R8118 VP.n8413 VP.n8412 0.012
R8119 VP.n9922 VP.n9921 0.012
R8120 VP.n9163 VP.n9162 0.012
R8121 VP.n8364 VP.n8363 0.012
R8122 VP.n7547 VP.n7546 0.012
R8123 VP.n6735 VP.n6734 0.012
R8124 VP.n9874 VP.n9873 0.012
R8125 VP.n9113 VP.n9112 0.012
R8126 VP.n8315 VP.n8314 0.012
R8127 VP.n7498 VP.n7497 0.012
R8128 VP.n6686 VP.n6685 0.012
R8129 VP.n5844 VP.n5843 0.012
R8130 VP.n5007 VP.n5006 0.012
R8131 VP.n8860 VP.n8859 0.012
R8132 VP.n9854 VP.n9853 0.012
R8133 VP.n9092 VP.n9091 0.012
R8134 VP.n8295 VP.n8294 0.012
R8135 VP.n7478 VP.n7477 0.012
R8136 VP.n6666 VP.n6665 0.012
R8137 VP.n5823 VP.n5822 0.012
R8138 VP.n4986 VP.n4985 0.012
R8139 VP.n4103 VP.n4102 0.012
R8140 VP.n3211 VP.n3210 0.012
R8141 VP.n10464 VP.n10455 0.012
R8142 VP.n9856 VP.n9836 0.012
R8143 VP.n9094 VP.n9073 0.012
R8144 VP.n8297 VP.n8276 0.012
R8145 VP.n7480 VP.n7460 0.012
R8146 VP.n6668 VP.n6648 0.012
R8147 VP.n5825 VP.n5804 0.012
R8148 VP.n4988 VP.n4967 0.012
R8149 VP.n4105 VP.n4084 0.012
R8150 VP.n3213 VP.n3193 0.012
R8151 VP.n2338 VP.n2329 0.012
R8152 VP.n8446 VP.n8414 0.012
R8153 VP.n6768 VP.n6736 0.012
R8154 VP.n5040 VP.n5008 0.012
R8155 VP.n8889 VP.n8861 0.012
R8156 VP.n3213 VP.n3212 0.012
R8157 VP.n752 VP.n751 0.011
R8158 VP.n9658 VP.n9657 0.011
R8159 VP.n8825 VP.n8823 0.011
R8160 VP.n9311 VP.n9310 0.011
R8161 VP.n10682 VP.n10678 0.011
R8162 VP.n11031 VP.n11029 0.011
R8163 VP.n1319 VP.n1318 0.011
R8164 VP.n2295 VP.n2294 0.011
R8165 VP.n3245 VP.n3244 0.011
R8166 VP.n4166 VP.n4165 0.011
R8167 VP.n5072 VP.n5071 0.011
R8168 VP.n5936 VP.n5935 0.011
R8169 VP.n6800 VP.n6799 0.011
R8170 VP.n7639 VP.n7638 0.011
R8171 VP.n8478 VP.n8477 0.011
R8172 VP.n10112 VP.n9683 0.011
R8173 VP.n9305 VP.n9304 0.011
R8174 VP.n10675 VP.n10674 0.011
R8175 VP.n10615 VP.n10613 0.011
R8176 VP.n10000 VP.n9971 0.011
R8177 VP.n9244 VP.n9214 0.011
R8178 VP.n9952 VP.n9923 0.011
R8179 VP.n9194 VP.n9164 0.011
R8180 VP.n8395 VP.n8365 0.011
R8181 VP.n7578 VP.n7548 0.011
R8182 VP.n9904 VP.n9875 0.011
R8183 VP.n9144 VP.n9114 0.011
R8184 VP.n8346 VP.n8316 0.011
R8185 VP.n7529 VP.n7499 0.011
R8186 VP.n6717 VP.n6687 0.011
R8187 VP.n5875 VP.n5845 0.011
R8188 VP.n9856 VP.n9855 0.011
R8189 VP.n9094 VP.n9093 0.011
R8190 VP.n8297 VP.n8296 0.011
R8191 VP.n7480 VP.n7479 0.011
R8192 VP.n6668 VP.n6667 0.011
R8193 VP.n5825 VP.n5824 0.011
R8194 VP.n4988 VP.n4987 0.011
R8195 VP.n4105 VP.n4104 0.011
R8196 VP.n5650 VP.n5648 0.011
R8197 VP.n4813 VP.n4811 0.011
R8198 VP.n3930 VP.n3928 0.011
R8199 VP.n3037 VP.n3035 0.011
R8200 VP.n2108 VP.n2106 0.011
R8201 VP.n6535 VP.n6533 0.011
R8202 VP.n5691 VP.n5689 0.011
R8203 VP.n4854 VP.n4852 0.011
R8204 VP.n3971 VP.n3969 0.011
R8205 VP.n3078 VP.n3076 0.011
R8206 VP.n2149 VP.n2147 0.011
R8207 VP.n7388 VP.n7386 0.011
R8208 VP.n6576 VP.n6574 0.011
R8209 VP.n5732 VP.n5730 0.011
R8210 VP.n4895 VP.n4893 0.011
R8211 VP.n4012 VP.n4010 0.011
R8212 VP.n3119 VP.n3117 0.011
R8213 VP.n2190 VP.n2188 0.011
R8214 VP.n1241 VP.n1239 0.011
R8215 VP.n9271 VP.n9264 0.011
R8216 VP.n7605 VP.n7598 0.011
R8217 VP.n5902 VP.n5895 0.011
R8218 VP.n4132 VP.n4125 0.011
R8219 VP.t8 VP.n10322 0.01
R8220 VP.t8 VP.n10304 0.01
R8221 VP.t8 VP.n10276 0.01
R8222 VP.t8 VP.n10248 0.01
R8223 VP.t8 VP.n10220 0.01
R8224 VP.n10091 VP.n10090 0.01
R8225 VP.n920 VP.n919 0.01
R8226 VP.n970 VP.n969 0.01
R8227 VP.n1020 VP.n1019 0.01
R8228 VP.n1070 VP.n1069 0.01
R8229 VP.n1120 VP.n1119 0.01
R8230 VP.t8 VP.n10202 0.01
R8231 VP.n9716 VP.n9711 0.01
R8232 VP.n37 VP.n36 0.01
R8233 VP.n27 VP.n26 0.01
R8234 VP.n138 VP.n137 0.01
R8235 VP.n9563 VP.n9560 0.01
R8236 VP.n8194 VP.n8193 0.01
R8237 VP.n7871 VP.n7868 0.01
R8238 VP.n8707 VP.n8705 0.01
R8239 VP.n9511 VP.n9509 0.01
R8240 VP.n6484 VP.n6483 0.01
R8241 VP.n6120 VP.n6117 0.01
R8242 VP.n6983 VP.n6981 0.01
R8243 VP.n7821 VP.n7819 0.01
R8244 VP.n8659 VP.n8657 0.01
R8245 VP.n9460 VP.n9458 0.01
R8246 VP.n4710 VP.n4709 0.01
R8247 VP.n2260 VP.n2259 0.01
R8248 VP.n2616 VP.n2613 0.01
R8249 VP.n3327 VP.n3325 0.01
R8250 VP.n4248 VP.n4246 0.01
R8251 VP.n5154 VP.n5152 0.01
R8252 VP.n6018 VP.n6016 0.01
R8253 VP.n6882 VP.n6880 0.01
R8254 VP.n7721 VP.n7719 0.01
R8255 VP.n8560 VP.n8558 0.01
R8256 VP.n9354 VP.n9352 0.01
R8257 VP.n312 VP.n309 0.01
R8258 VP.n4301 VP.n4298 0.01
R8259 VP.n5206 VP.n5204 0.01
R8260 VP.n6071 VP.n6069 0.01
R8261 VP.n6935 VP.n6933 0.01
R8262 VP.n7773 VP.n7771 0.01
R8263 VP.n8612 VP.n8610 0.01
R8264 VP.n9410 VP.n9408 0.01
R8265 VP.n10998 VP.n10997 0.01
R8266 VP.n10939 VP.n10938 0.01
R8267 VP.n8737 VP.n8736 0.01
R8268 VP.n9544 VP.n9543 0.01
R8269 VP.n10888 VP.n10887 0.01
R8270 VP.n7014 VP.n7013 0.01
R8271 VP.n7852 VP.n7851 0.01
R8272 VP.n8689 VP.n8688 0.01
R8273 VP.n9493 VP.n9492 0.01
R8274 VP.n10837 VP.n10836 0.01
R8275 VP.n5235 VP.n5234 0.01
R8276 VP.n6101 VP.n6100 0.01
R8277 VP.n6965 VP.n6964 0.01
R8278 VP.n7803 VP.n7802 0.01
R8279 VP.n8641 VP.n8640 0.01
R8280 VP.n9442 VP.n9441 0.01
R8281 VP.n10786 VP.n10785 0.01
R8282 VP.n10724 VP.n10723 0.01
R8283 VP.n9379 VP.n9378 0.01
R8284 VP.n8584 VP.n8583 0.01
R8285 VP.n7745 VP.n7744 0.01
R8286 VP.n6906 VP.n6905 0.01
R8287 VP.n6042 VP.n6041 0.01
R8288 VP.n5178 VP.n5177 0.01
R8289 VP.n4272 VP.n4271 0.01
R8290 VP.n3351 VP.n3350 0.01
R8291 VP.n10129 VP.n10128 0.01
R8292 VP.n1316 VP.n1315 0.01
R8293 VP.n766 VP.n765 0.01
R8294 VP.n2292 VP.n2291 0.01
R8295 VP.n893 VP.n892 0.01
R8296 VP.n1327 VP.n1326 0.01
R8297 VP.n1755 VP.n1754 0.01
R8298 VP.n3242 VP.n3241 0.01
R8299 VP.n943 VP.n942 0.01
R8300 VP.n1455 VP.n1454 0.01
R8301 VP.n1880 VP.n1879 0.01
R8302 VP.n2303 VP.n2302 0.01
R8303 VP.n2716 VP.n2715 0.01
R8304 VP.n4163 VP.n4162 0.01
R8305 VP.n993 VP.n992 0.01
R8306 VP.n1493 VP.n1492 0.01
R8307 VP.n1932 VP.n1931 0.01
R8308 VP.n2555 VP.n2554 0.01
R8309 VP.n2861 VP.n2860 0.01
R8310 VP.n3253 VP.n3252 0.01
R8311 VP.n3656 VP.n3655 0.01
R8312 VP.n5069 VP.n5068 0.01
R8313 VP.n1043 VP.n1042 0.01
R8314 VP.n1531 VP.n1530 0.01
R8315 VP.n1984 VP.n1983 0.01
R8316 VP.n2517 VP.n2516 0.01
R8317 VP.n2913 VP.n2912 0.01
R8318 VP.n3433 VP.n3432 0.01
R8319 VP.n3806 VP.n3805 0.01
R8320 VP.n4174 VP.n4173 0.01
R8321 VP.n4562 VP.n4561 0.01
R8322 VP.n5933 VP.n5932 0.01
R8323 VP.n1093 VP.n1092 0.01
R8324 VP.n1569 VP.n1568 0.01
R8325 VP.n2036 VP.n2035 0.01
R8326 VP.n2479 VP.n2478 0.01
R8327 VP.n2965 VP.n2964 0.01
R8328 VP.n3471 VP.n3470 0.01
R8329 VP.n3858 VP.n3857 0.01
R8330 VP.n4350 VP.n4349 0.01
R8331 VP.n4741 VP.n4740 0.01
R8332 VP.n5080 VP.n5079 0.01
R8333 VP.n5457 VP.n5456 0.01
R8334 VP.n6797 VP.n6796 0.01
R8335 VP.n1143 VP.n1142 0.01
R8336 VP.n1607 VP.n1606 0.01
R8337 VP.n2088 VP.n2087 0.01
R8338 VP.n2447 VP.n2446 0.01
R8339 VP.n3017 VP.n3016 0.01
R8340 VP.n3509 VP.n3508 0.01
R8341 VP.n3910 VP.n3909 0.01
R8342 VP.n4388 VP.n4387 0.01
R8343 VP.n4793 VP.n4792 0.01
R8344 VP.n5310 VP.n5309 0.01
R8345 VP.n5630 VP.n5629 0.01
R8346 VP.n5944 VP.n5943 0.01
R8347 VP.n6313 VP.n6312 0.01
R8348 VP.n7636 VP.n7635 0.01
R8349 VP.n1181 VP.n1180 0.01
R8350 VP.n1639 VP.n1638 0.01
R8351 VP.n2129 VP.n2128 0.01
R8352 VP.n2415 VP.n2414 0.01
R8353 VP.n3058 VP.n3057 0.01
R8354 VP.n3541 VP.n3540 0.01
R8355 VP.n3951 VP.n3950 0.01
R8356 VP.n4420 VP.n4419 0.01
R8357 VP.n4834 VP.n4833 0.01
R8358 VP.n5342 VP.n5341 0.01
R8359 VP.n5671 VP.n5670 0.01
R8360 VP.n6170 VP.n6169 0.01
R8361 VP.n6515 VP.n6514 0.01
R8362 VP.n6808 VP.n6807 0.01
R8363 VP.n7172 VP.n7171 0.01
R8364 VP.n8475 VP.n8474 0.01
R8365 VP.n1221 VP.n1220 0.01
R8366 VP.n1671 VP.n1670 0.01
R8367 VP.n2170 VP.n2169 0.01
R8368 VP.n2383 VP.n2382 0.01
R8369 VP.n3099 VP.n3098 0.01
R8370 VP.n3573 VP.n3572 0.01
R8371 VP.n3992 VP.n3991 0.01
R8372 VP.n4452 VP.n4451 0.01
R8373 VP.n4875 VP.n4874 0.01
R8374 VP.n5374 VP.n5373 0.01
R8375 VP.n5712 VP.n5711 0.01
R8376 VP.n6202 VP.n6201 0.01
R8377 VP.n6556 VP.n6555 0.01
R8378 VP.n7089 VP.n7088 0.01
R8379 VP.n7368 VP.n7367 0.01
R8380 VP.n7647 VP.n7646 0.01
R8381 VP.n8000 VP.n7999 0.01
R8382 VP.n9681 VP.n9680 0.01
R8383 VP.n1262 VP.n1261 0.01
R8384 VP.n1703 VP.n1702 0.01
R8385 VP.n2211 VP.n2210 0.01
R8386 VP.n2351 VP.n2350 0.01
R8387 VP.n3140 VP.n3139 0.01
R8388 VP.n3605 VP.n3604 0.01
R8389 VP.n4033 VP.n4032 0.01
R8390 VP.n4484 VP.n4483 0.01
R8391 VP.n4916 VP.n4915 0.01
R8392 VP.n5406 VP.n5405 0.01
R8393 VP.n5753 VP.n5752 0.01
R8394 VP.n6234 VP.n6233 0.01
R8395 VP.n6597 VP.n6596 0.01
R8396 VP.n7121 VP.n7120 0.01
R8397 VP.n7409 VP.n7408 0.01
R8398 VP.n7921 VP.n7920 0.01
R8399 VP.n8225 VP.n8224 0.01
R8400 VP.n8486 VP.n8485 0.01
R8401 VP.n8834 VP.n8833 0.01
R8402 VP.n9302 VP.n9301 0.01
R8403 VP.n808 VP.n807 0.01
R8404 VP.n1358 VP.n1357 0.01
R8405 VP.n1794 VP.n1793 0.01
R8406 VP.n2675 VP.n2674 0.01
R8407 VP.n2754 VP.n2753 0.01
R8408 VP.n3284 VP.n3283 0.01
R8409 VP.n3694 VP.n3693 0.01
R8410 VP.n4205 VP.n4204 0.01
R8411 VP.n4603 VP.n4602 0.01
R8412 VP.n5111 VP.n5110 0.01
R8413 VP.n5495 VP.n5494 0.01
R8414 VP.n5975 VP.n5974 0.01
R8415 VP.n6351 VP.n6350 0.01
R8416 VP.n6839 VP.n6838 0.01
R8417 VP.n7210 VP.n7209 0.01
R8418 VP.n7678 VP.n7677 0.01
R8419 VP.n8038 VP.n8037 0.01
R8420 VP.n8517 VP.n8516 0.01
R8421 VP.n8882 VP.n8881 0.01
R8422 VP.n10107 VP.n10106 0.01
R8423 VP.n10118 VP.n10117 0.01
R8424 VP.n10655 VP.n10654 0.01
R8425 VP.n10895 VP.n10868 0.01
R8426 VP.n9551 VP.n9530 0.01
R8427 VP.n10844 VP.n10817 0.01
R8428 VP.n9500 VP.n9479 0.01
R8429 VP.n7859 VP.n7839 0.01
R8430 VP.n7021 VP.n7001 0.01
R8431 VP.n10793 VP.n10766 0.01
R8432 VP.n9449 VP.n9428 0.01
R8433 VP.n7810 VP.n7790 0.01
R8434 VP.n6972 VP.n6952 0.01
R8435 VP.n6108 VP.n6088 0.01
R8436 VP.n10739 VP.n10738 0.01
R8437 VP.n9394 VP.n9393 0.01
R8438 VP.n6920 VP.n6919 0.01
R8439 VP.n6056 VP.n6055 0.01
R8440 VP.n9320 VP.n9319 0.01
R8441 VP.n9030 VP.n9029 0.009
R8442 VP.n7335 VP.n7334 0.009
R8443 VP.n5597 VP.n5596 0.009
R8444 VP.n861 VP.n860 0.009
R8445 VP.n1847 VP.n1846 0.009
R8446 VP.n3774 VP.n3773 0.009
R8447 VP.n10681 VP.n10680 0.009
R8448 VP.n9719 VP.n9718 0.009
R8449 VP.n264 VP.n260 0.009
R8450 VP.n366 VP.n362 0.009
R8451 VP.n413 VP.n409 0.009
R8452 VP.n460 VP.n456 0.009
R8453 VP.n507 VP.n503 0.009
R8454 VP.n554 VP.n550 0.009
R8455 VP.n601 VP.n597 0.009
R8456 VP.n641 VP.n637 0.009
R8457 VP.n671 VP.n667 0.009
R8458 VP.n703 VP.n699 0.009
R8459 VP.n9596 VP.n9595 0.009
R8460 VP.n10625 VP.n10624 0.009
R8461 VP.n10592 VP.n10591 0.009
R8462 VP.n10587 VP.n10586 0.009
R8463 VP.n8193 VP.n8191 0.009
R8464 VP.n10557 VP.n10556 0.009
R8465 VP.n10552 VP.n10551 0.009
R8466 VP.n6483 VP.n6481 0.009
R8467 VP.n10522 VP.n10521 0.009
R8468 VP.n10517 VP.n10516 0.009
R8469 VP.n4709 VP.n4707 0.009
R8470 VP.n10487 VP.n10486 0.009
R8471 VP.n10482 VP.n10481 0.009
R8472 VP.n10442 VP.n10441 0.009
R8473 VP.n9655 VP.n9654 0.009
R8474 VP.t116 VP.n9 0.009
R8475 VP.n8821 VP.n8820 0.009
R8476 VP.n9659 VP.n9320 0.009
R8477 VP.n10685 VP.n10684 0.009
R8478 VP.t116 VP.n150 0.009
R8479 VP.n11027 VP.n11026 0.009
R8480 VP.n11048 VP.n11047 0.009
R8481 VP.n11049 VP.n11048 0.009
R8482 VP.n11050 VP.n11049 0.009
R8483 VP.n11051 VP.n11050 0.009
R8484 VP.n11052 VP.n11051 0.009
R8485 VP.n11053 VP.n11052 0.009
R8486 VP.n11054 VP.n11053 0.009
R8487 VP.n11055 VP.n11054 0.009
R8488 VP.n11056 VP.n11055 0.009
R8489 VP.n11057 VP.n11056 0.009
R8490 VP.n11058 VP.n11057 0.009
R8491 VP.n11046 VP.n11045 0.009
R8492 VP.n11045 VP.n11044 0.009
R8493 VP.n11044 VP.n11043 0.009
R8494 VP.n11043 VP.n11042 0.009
R8495 VP.n11042 VP.n11041 0.009
R8496 VP.n11041 VP.n11040 0.009
R8497 VP.n11040 VP.n11039 0.009
R8498 VP.n11039 VP.n11038 0.009
R8499 VP.n11038 VP.n11037 0.009
R8500 VP.n11037 VP.n11036 0.009
R8501 VP.n11036 VP.n11035 0.009
R8502 VP.n722 VP.n721 0.009
R8503 VP.n9627 VP.n9625 0.009
R8504 VP.n7962 VP.n7960 0.009
R8505 VP.n9238 VP.n9236 0.009
R8506 VP.n9994 VP.n9992 0.009
R8507 VP.n6275 VP.n6273 0.009
R8508 VP.n7572 VP.n7570 0.009
R8509 VP.n8389 VP.n8387 0.009
R8510 VP.n9188 VP.n9186 0.009
R8511 VP.n9946 VP.n9944 0.009
R8512 VP.n4524 VP.n4522 0.009
R8513 VP.n5869 VP.n5867 0.009
R8514 VP.n6711 VP.n6709 0.009
R8515 VP.n7523 VP.n7521 0.009
R8516 VP.n8340 VP.n8338 0.009
R8517 VP.n9138 VP.n9136 0.009
R8518 VP.n9898 VP.n9896 0.009
R8519 VP.n10453 VP.n10451 0.009
R8520 VP.n9834 VP.n9832 0.009
R8521 VP.n9071 VP.n9069 0.009
R8522 VP.n8274 VP.n8272 0.009
R8523 VP.n7458 VP.n7456 0.009
R8524 VP.n6646 VP.n6644 0.009
R8525 VP.n5802 VP.n5800 0.009
R8526 VP.n4965 VP.n4963 0.009
R8527 VP.n4082 VP.n4080 0.009
R8528 VP.n2327 VP.n2325 0.009
R8529 VP.n1406 VP.n1404 0.009
R8530 VP.n3384 VP.n3382 0.009
R8531 VP.n8195 VP.n8194 0.009
R8532 VP.n6485 VP.n6484 0.009
R8533 VP.n4711 VP.n4710 0.009
R8534 VP.n10351 VP.n10350 0.008
R8535 VP.n2242 VP.n2241 0.008
R8536 VP.n11005 VP.n10978 0.008
R8537 VP.n9633 VP.n9613 0.008
R8538 VP.n10911 VP.n10902 0.008
R8539 VP.n10911 VP.n10910 0.008
R8540 VP.n9574 VP.n9573 0.008
R8541 VP.n7968 VP.n7948 0.008
R8542 VP.n10860 VP.n10851 0.008
R8543 VP.n10860 VP.n10859 0.008
R8544 VP.n9522 VP.n9521 0.008
R8545 VP.n6281 VP.n6261 0.008
R8546 VP.n10809 VP.n10800 0.008
R8547 VP.n10809 VP.n10808 0.008
R8548 VP.n9471 VP.n9470 0.008
R8549 VP.n10753 VP.n10751 0.008
R8550 VP.n10710 VP.n10709 0.008
R8551 VP.n9365 VP.n9364 0.008
R8552 VP.n9343 VP.n9342 0.008
R8553 VP.n2338 VP.n2337 0.008
R8554 VP.n10753 VP.n10752 0.008
R8555 VP.n9415 VP.n9414 0.008
R8556 VP.n10946 VP.n10919 0.008
R8557 VP.n5329 VP.n5328 0.008
R8558 VP.n4407 VP.n4406 0.008
R8559 VP.n3528 VP.n3527 0.008
R8560 VP.n2466 VP.n2465 0.008
R8561 VP.n1626 VP.n1625 0.008
R8562 VP.n6189 VP.n6188 0.008
R8563 VP.n5361 VP.n5360 0.008
R8564 VP.n4439 VP.n4438 0.008
R8565 VP.n3560 VP.n3559 0.008
R8566 VP.n2434 VP.n2433 0.008
R8567 VP.n1658 VP.n1657 0.008
R8568 VP.n7108 VP.n7107 0.008
R8569 VP.n6221 VP.n6220 0.008
R8570 VP.n5393 VP.n5392 0.008
R8571 VP.n4471 VP.n4470 0.008
R8572 VP.n3592 VP.n3591 0.008
R8573 VP.n2402 VP.n2401 0.008
R8574 VP.n1690 VP.n1689 0.008
R8575 VP.n682 VP.n681 0.008
R8576 VP.n10020 VP.n10016 0.008
R8577 VP.n10603 VP.n10592 0.008
R8578 VP.n8426 VP.n8422 0.008
R8579 VP.n9226 VP.n9222 0.008
R8580 VP.n9983 VP.n9979 0.008
R8581 VP.n10568 VP.n10557 0.008
R8582 VP.n6748 VP.n6744 0.008
R8583 VP.n7560 VP.n7556 0.008
R8584 VP.n8377 VP.n8373 0.008
R8585 VP.n9176 VP.n9172 0.008
R8586 VP.n9935 VP.n9931 0.008
R8587 VP.n10533 VP.n10522 0.008
R8588 VP.n5020 VP.n5016 0.008
R8589 VP.n5857 VP.n5853 0.008
R8590 VP.n6699 VP.n6695 0.008
R8591 VP.n7511 VP.n7507 0.008
R8592 VP.n8328 VP.n8324 0.008
R8593 VP.n9126 VP.n9122 0.008
R8594 VP.n9887 VP.n9883 0.008
R8595 VP.n10498 VP.n10487 0.008
R8596 VP.n9820 VP.n9819 0.008
R8597 VP.n9056 VP.n9055 0.008
R8598 VP.n8259 VP.n8258 0.008
R8599 VP.n7443 VP.n7442 0.008
R8600 VP.n6631 VP.n6630 0.008
R8601 VP.n5787 VP.n5786 0.008
R8602 VP.n4950 VP.n4949 0.008
R8603 VP.n4067 VP.n4066 0.008
R8604 VP.n3174 VP.n3173 0.008
R8605 VP.n252 VP.n251 0.008
R8606 VP.n354 VP.n353 0.008
R8607 VP.n401 VP.n400 0.008
R8608 VP.n448 VP.n447 0.008
R8609 VP.n495 VP.n494 0.008
R8610 VP.n542 VP.n541 0.008
R8611 VP.n589 VP.n588 0.008
R8612 VP.n629 VP.n628 0.008
R8613 VP.n659 VP.n658 0.008
R8614 VP.n691 VP.n690 0.008
R8615 VP VP.n11058 0.008
R8616 VP.n757 VP.n756 0.008
R8617 VP.n9969 VP.n9968 0.008
R8618 VP.n9212 VP.n9211 0.008
R8619 VP.n8412 VP.n8411 0.008
R8620 VP.n9921 VP.n9920 0.008
R8621 VP.n9162 VP.n9161 0.008
R8622 VP.n8363 VP.n8362 0.008
R8623 VP.n7546 VP.n7545 0.008
R8624 VP.n6734 VP.n6733 0.008
R8625 VP.n9873 VP.n9872 0.008
R8626 VP.n9112 VP.n9111 0.008
R8627 VP.n8314 VP.n8313 0.008
R8628 VP.n7497 VP.n7496 0.008
R8629 VP.n6685 VP.n6684 0.008
R8630 VP.n5843 VP.n5842 0.008
R8631 VP.n5006 VP.n5005 0.008
R8632 VP.n8859 VP.n8858 0.008
R8633 VP.n9853 VP.n9852 0.008
R8634 VP.n9091 VP.n9090 0.008
R8635 VP.n8294 VP.n8293 0.008
R8636 VP.n7477 VP.n7476 0.008
R8637 VP.n6665 VP.n6664 0.008
R8638 VP.n5822 VP.n5821 0.008
R8639 VP.n4985 VP.n4984 0.008
R8640 VP.n4102 VP.n4101 0.008
R8641 VP.n3210 VP.n3209 0.008
R8642 VP.n9595 VP.n9594 0.007
R8643 VP.n345 VP.n341 0.007
R8644 VP.n9971 VP.n9970 0.007
R8645 VP.n9214 VP.n9213 0.007
R8646 VP.n9923 VP.n9922 0.007
R8647 VP.n9164 VP.n9163 0.007
R8648 VP.n8365 VP.n8364 0.007
R8649 VP.n7548 VP.n7547 0.007
R8650 VP.n9875 VP.n9874 0.007
R8651 VP.n9114 VP.n9113 0.007
R8652 VP.n8316 VP.n8315 0.007
R8653 VP.n7499 VP.n7498 0.007
R8654 VP.n6687 VP.n6686 0.007
R8655 VP.n5845 VP.n5844 0.007
R8656 VP.n9855 VP.n9854 0.007
R8657 VP.n9093 VP.n9092 0.007
R8658 VP.n8296 VP.n8295 0.007
R8659 VP.n7479 VP.n7478 0.007
R8660 VP.n6667 VP.n6666 0.007
R8661 VP.n5824 VP.n5823 0.007
R8662 VP.n4987 VP.n4986 0.007
R8663 VP.n4104 VP.n4103 0.007
R8664 VP.n10034 VP.n10031 0.007
R8665 VP.n8440 VP.n8437 0.007
R8666 VP.n6762 VP.n6759 0.007
R8667 VP.n5034 VP.n5031 0.007
R8668 VP.n3191 VP.n3188 0.007
R8669 VP.n10602 VP.n10601 0.007
R8670 VP.n10567 VP.n10566 0.007
R8671 VP.n10532 VP.n10531 0.007
R8672 VP.n10497 VP.n10496 0.007
R8673 VP.n10630 VP.n10629 0.007
R8674 VP.n9601 VP.n9600 0.007
R8675 VP.n9605 VP.n9598 0.007
R8676 VP.n8799 VP.n8791 0.007
R8677 VP.n8763 VP.n8760 0.007
R8678 VP.n7076 VP.n7068 0.007
R8679 VP.n7040 VP.n7037 0.007
R8680 VP.n5297 VP.n5289 0.007
R8681 VP.n5261 VP.n5258 0.007
R8682 VP.n3420 VP.n3412 0.007
R8683 VP.n1403 VP.n1400 0.007
R8684 VP.n391 VP.n381 0.007
R8685 VP.n438 VP.n428 0.007
R8686 VP.n485 VP.n475 0.007
R8687 VP.n532 VP.n522 0.007
R8688 VP.n579 VP.n569 0.007
R8689 VP.n8825 VP.n8824 0.007
R8690 VP.n10682 VP.n10681 0.007
R8691 VP.n11031 VP.n11030 0.007
R8692 VP.n3381 VP.n3378 0.007
R8693 VP.n10121 VP.n10115 0.007
R8694 VP.n1442 VP.n1439 0.007
R8695 VP.n306 VP.n305 0.007
R8696 VP.n8414 VP.n8413 0.007
R8697 VP.n6736 VP.n6735 0.007
R8698 VP.n5008 VP.n5007 0.007
R8699 VP.n8861 VP.n8860 0.007
R8700 VP.n3212 VP.n3211 0.007
R8701 VP.n10320 VP.n10319 0.006
R8702 VP.n10302 VP.n10301 0.006
R8703 VP.n10274 VP.n10273 0.006
R8704 VP.n10246 VP.n10245 0.006
R8705 VP.n10218 VP.n10217 0.006
R8706 VP.n10195 VP.n10194 0.006
R8707 VP.n916 VP.n914 0.006
R8708 VP.n1908 VP.n1907 0.006
R8709 VP.n966 VP.n964 0.006
R8710 VP.n2884 VP.n2882 0.006
R8711 VP.n2889 VP.n2888 0.006
R8712 VP.n1960 VP.n1959 0.006
R8713 VP.n1016 VP.n1014 0.006
R8714 VP.n3834 VP.n3833 0.006
R8715 VP.n2936 VP.n2934 0.006
R8716 VP.n2941 VP.n2940 0.006
R8717 VP.n2012 VP.n2011 0.006
R8718 VP.n4764 VP.n4762 0.006
R8719 VP.n4769 VP.n4768 0.006
R8720 VP.n3881 VP.n3879 0.006
R8721 VP.n3886 VP.n3885 0.006
R8722 VP.n2988 VP.n2986 0.006
R8723 VP.n2993 VP.n2992 0.006
R8724 VP.n2064 VP.n2063 0.006
R8725 VP.n1116 VP.n1114 0.006
R8726 VP.n10071 VP.n10048 0.006
R8727 VP.n9273 VP.n9252 0.006
R8728 VP.n7607 VP.n7586 0.006
R8729 VP.n5904 VP.n5883 0.006
R8730 VP.n4134 VP.n4113 0.006
R8731 VP.n2263 VP.n2262 0.006
R8732 VP.n7889 VP.n7888 0.006
R8733 VP.n6138 VP.n6137 0.006
R8734 VP.n4318 VP.n4317 0.006
R8735 VP.n2592 VP.n2591 0.006
R8736 VP.n10070 VP.n10066 0.006
R8737 VP.n11004 VP.n10996 0.006
R8738 VP.n10641 VP.n10630 0.006
R8739 VP.n10945 VP.n10937 0.006
R8740 VP.n9031 VP.n9030 0.006
R8741 VP.n9028 VP.n9026 0.006
R8742 VP.n8770 VP.n8765 0.006
R8743 VP.n8743 VP.n8735 0.006
R8744 VP.n9550 VP.n9542 0.006
R8745 VP.n10894 VP.n10886 0.006
R8746 VP.n7336 VP.n7335 0.006
R8747 VP.n7333 VP.n7331 0.006
R8748 VP.n7047 VP.n7042 0.006
R8749 VP.n7020 VP.n7012 0.006
R8750 VP.n7858 VP.n7850 0.006
R8751 VP.n8695 VP.n8687 0.006
R8752 VP.n9499 VP.n9491 0.006
R8753 VP.n10843 VP.n10835 0.006
R8754 VP.n5598 VP.n5597 0.006
R8755 VP.n5595 VP.n5593 0.006
R8756 VP.n5268 VP.n5263 0.006
R8757 VP.n5241 VP.n5233 0.006
R8758 VP.n6107 VP.n6099 0.006
R8759 VP.n6971 VP.n6963 0.006
R8760 VP.n7809 VP.n7801 0.006
R8761 VP.n8647 VP.n8639 0.006
R8762 VP.n9448 VP.n9440 0.006
R8763 VP.n10792 VP.n10784 0.006
R8764 VP.n10727 VP.n10719 0.006
R8765 VP.n9382 VP.n9374 0.006
R8766 VP.n8587 VP.n8579 0.006
R8767 VP.n7748 VP.n7740 0.006
R8768 VP.n6909 VP.n6901 0.006
R8769 VP.n6045 VP.n6037 0.006
R8770 VP.n5181 VP.n5173 0.006
R8771 VP.n4275 VP.n4267 0.006
R8772 VP.n3354 VP.n3346 0.006
R8773 VP.n862 VP.n861 0.006
R8774 VP.n859 VP.n857 0.006
R8775 VP.n1414 VP.n1406 0.006
R8776 VP.n1848 VP.n1847 0.006
R8777 VP.n1845 VP.n1843 0.006
R8778 VP.n313 VP.n312 0.006
R8779 VP.n899 VP.n888 0.006
R8780 VP.n1333 VP.n1325 0.006
R8781 VP.n949 VP.n938 0.006
R8782 VP.n1461 VP.n1453 0.006
R8783 VP.n1886 VP.n1875 0.006
R8784 VP.n2309 VP.n2301 0.006
R8785 VP.n999 VP.n988 0.006
R8786 VP.n1499 VP.n1491 0.006
R8787 VP.n1938 VP.n1927 0.006
R8788 VP.n2561 VP.n2553 0.006
R8789 VP.n2867 VP.n2856 0.006
R8790 VP.n3259 VP.n3251 0.006
R8791 VP.n1049 VP.n1038 0.006
R8792 VP.n1537 VP.n1529 0.006
R8793 VP.n1990 VP.n1979 0.006
R8794 VP.n2523 VP.n2515 0.006
R8795 VP.n2919 VP.n2908 0.006
R8796 VP.n3439 VP.n3431 0.006
R8797 VP.n3812 VP.n3801 0.006
R8798 VP.n4180 VP.n4172 0.006
R8799 VP.n1099 VP.n1088 0.006
R8800 VP.n1575 VP.n1567 0.006
R8801 VP.n2042 VP.n2031 0.006
R8802 VP.n2485 VP.n2477 0.006
R8803 VP.n2971 VP.n2960 0.006
R8804 VP.n3477 VP.n3469 0.006
R8805 VP.n3864 VP.n3853 0.006
R8806 VP.n4356 VP.n4348 0.006
R8807 VP.n4747 VP.n4736 0.006
R8808 VP.n5086 VP.n5078 0.006
R8809 VP.n1149 VP.n1138 0.006
R8810 VP.n1613 VP.n1605 0.006
R8811 VP.n2094 VP.n2083 0.006
R8812 VP.n2453 VP.n2445 0.006
R8813 VP.n3023 VP.n3012 0.006
R8814 VP.n3515 VP.n3507 0.006
R8815 VP.n3916 VP.n3905 0.006
R8816 VP.n4394 VP.n4386 0.006
R8817 VP.n4799 VP.n4788 0.006
R8818 VP.n5316 VP.n5308 0.006
R8819 VP.n5636 VP.n5625 0.006
R8820 VP.n5950 VP.n5942 0.006
R8821 VP.n1187 VP.n1176 0.006
R8822 VP.n1645 VP.n1637 0.006
R8823 VP.n2135 VP.n2124 0.006
R8824 VP.n2421 VP.n2413 0.006
R8825 VP.n3064 VP.n3053 0.006
R8826 VP.n3547 VP.n3539 0.006
R8827 VP.n3957 VP.n3946 0.006
R8828 VP.n4426 VP.n4418 0.006
R8829 VP.n4840 VP.n4829 0.006
R8830 VP.n5348 VP.n5340 0.006
R8831 VP.n5677 VP.n5666 0.006
R8832 VP.n6176 VP.n6168 0.006
R8833 VP.n6521 VP.n6510 0.006
R8834 VP.n6814 VP.n6806 0.006
R8835 VP.n1227 VP.n1216 0.006
R8836 VP.n1677 VP.n1669 0.006
R8837 VP.n2176 VP.n2165 0.006
R8838 VP.n2389 VP.n2381 0.006
R8839 VP.n3105 VP.n3094 0.006
R8840 VP.n3579 VP.n3571 0.006
R8841 VP.n3998 VP.n3987 0.006
R8842 VP.n4458 VP.n4450 0.006
R8843 VP.n4881 VP.n4870 0.006
R8844 VP.n5380 VP.n5372 0.006
R8845 VP.n5718 VP.n5707 0.006
R8846 VP.n6208 VP.n6200 0.006
R8847 VP.n6562 VP.n6551 0.006
R8848 VP.n7095 VP.n7087 0.006
R8849 VP.n7374 VP.n7363 0.006
R8850 VP.n7653 VP.n7645 0.006
R8851 VP.n1268 VP.n1257 0.006
R8852 VP.n1709 VP.n1701 0.006
R8853 VP.n2217 VP.n2206 0.006
R8854 VP.n2357 VP.n2349 0.006
R8855 VP.n3146 VP.n3135 0.006
R8856 VP.n3611 VP.n3603 0.006
R8857 VP.n4039 VP.n4028 0.006
R8858 VP.n4490 VP.n4482 0.006
R8859 VP.n4922 VP.n4911 0.006
R8860 VP.n5412 VP.n5404 0.006
R8861 VP.n5759 VP.n5748 0.006
R8862 VP.n6240 VP.n6232 0.006
R8863 VP.n6603 VP.n6592 0.006
R8864 VP.n7127 VP.n7119 0.006
R8865 VP.n7415 VP.n7404 0.006
R8866 VP.n7927 VP.n7919 0.006
R8867 VP.n8231 VP.n8220 0.006
R8868 VP.n8492 VP.n8484 0.006
R8869 VP.n286 VP.n284 0.006
R8870 VP.n814 VP.n803 0.006
R8871 VP.n1364 VP.n1356 0.006
R8872 VP.n1800 VP.n1789 0.006
R8873 VP.n2681 VP.n2673 0.006
R8874 VP.n2760 VP.n2749 0.006
R8875 VP.n3290 VP.n3282 0.006
R8876 VP.n3700 VP.n3689 0.006
R8877 VP.n4211 VP.n4203 0.006
R8878 VP.n4609 VP.n4598 0.006
R8879 VP.n5117 VP.n5109 0.006
R8880 VP.n5501 VP.n5490 0.006
R8881 VP.n5981 VP.n5973 0.006
R8882 VP.n6357 VP.n6346 0.006
R8883 VP.n6845 VP.n6837 0.006
R8884 VP.n7216 VP.n7205 0.006
R8885 VP.n7684 VP.n7676 0.006
R8886 VP.n8044 VP.n8033 0.006
R8887 VP.n8523 VP.n8515 0.006
R8888 VP.n8888 VP.n8877 0.006
R8889 VP.n9690 VP.n9688 0.006
R8890 VP.n9327 VP.n9325 0.006
R8891 VP.n8900 VP.n8898 0.006
R8892 VP.n8534 VP.n8532 0.006
R8893 VP.n8056 VP.n8054 0.006
R8894 VP.n7695 VP.n7693 0.006
R8895 VP.n7228 VP.n7226 0.006
R8896 VP.n6856 VP.n6854 0.006
R8897 VP.n6369 VP.n6367 0.006
R8898 VP.n5992 VP.n5990 0.006
R8899 VP.n5513 VP.n5511 0.006
R8900 VP.n5128 VP.n5126 0.006
R8901 VP.n4618 VP.n4616 0.006
R8902 VP.n4222 VP.n4220 0.006
R8903 VP.n3712 VP.n3710 0.006
R8904 VP.n3301 VP.n3299 0.006
R8905 VP.n2772 VP.n2770 0.006
R8906 VP.n2636 VP.n2634 0.006
R8907 VP.n1812 VP.n1810 0.006
R8908 VP.n1375 VP.n1373 0.006
R8909 VP.n826 VP.n824 0.006
R8910 VP.n10416 VP.n10414 0.006
R8911 VP.n3386 VP.n3384 0.006
R8912 VP.n3775 VP.n3774 0.006
R8913 VP.n3772 VP.n3770 0.006
R8914 VP.n10604 VP.n10577 0.006
R8915 VP.n10040 VP.n10008 0.006
R8916 VP.n10403 VP.n10402 0.006
R8917 VP.n10403 VP.n10395 0.006
R8918 VP.n9807 VP.n9806 0.006
R8919 VP.n9043 VP.n9042 0.006
R8920 VP.n8205 VP.n8204 0.006
R8921 VP.n10569 VP.n10542 0.006
R8922 VP.n10386 VP.n10385 0.006
R8923 VP.n10386 VP.n10378 0.006
R8924 VP.n9785 VP.n9784 0.006
R8925 VP.n9013 VP.n9012 0.006
R8926 VP.n8169 VP.n8168 0.006
R8927 VP.n7348 VP.n7347 0.006
R8928 VP.n6495 VP.n6494 0.006
R8929 VP.n10534 VP.n10507 0.006
R8930 VP.n10369 VP.n10368 0.006
R8931 VP.n10369 VP.n10361 0.006
R8932 VP.n9763 VP.n9762 0.006
R8933 VP.n8990 VP.n8989 0.006
R8934 VP.n8146 VP.n8145 0.006
R8935 VP.n7318 VP.n7317 0.006
R8936 VP.n6459 VP.n6458 0.006
R8937 VP.n5610 VP.n5609 0.006
R8938 VP.n4721 VP.n4720 0.006
R8939 VP.n10499 VP.n10472 0.006
R8940 VP.n10159 VP.n10155 0.006
R8941 VP.n10144 VP.n10143 0.006
R8942 VP.n9741 VP.n9740 0.006
R8943 VP.n8941 VP.n8940 0.006
R8944 VP.n8097 VP.n8096 0.006
R8945 VP.n7269 VP.n7268 0.006
R8946 VP.n6410 VP.n6409 0.006
R8947 VP.n5554 VP.n5553 0.006
R8948 VP.n4659 VP.n4658 0.006
R8949 VP.n3753 VP.n3752 0.006
R8950 VP.n2813 VP.n2812 0.006
R8951 VP.n1860 VP.n1859 0.006
R8952 VP.n873 VP.n872 0.006
R8953 VP.n1162 VP.n1161 0.006
R8954 VP.n1202 VP.n1201 0.006
R8955 VP.n8045 VP.n8015 0.006
R8956 VP.n7217 VP.n7187 0.006
R8957 VP.n6358 VP.n6328 0.006
R8958 VP.n5502 VP.n5472 0.006
R8959 VP.n4610 VP.n4577 0.006
R8960 VP.n3701 VP.n3671 0.006
R8961 VP.n2761 VP.n2731 0.006
R8962 VP.n1801 VP.n1771 0.006
R8963 VP.n815 VP.n782 0.006
R8964 VP.n847 VP.n846 0.006
R8965 VP.n1830 VP.n1829 0.006
R8966 VP.n2790 VP.n2789 0.006
R8967 VP.n3730 VP.n3729 0.006
R8968 VP.n4636 VP.n4635 0.006
R8969 VP.n5531 VP.n5530 0.006
R8970 VP.n6387 VP.n6386 0.006
R8971 VP.n7246 VP.n7245 0.006
R8972 VP.n8074 VP.n8073 0.006
R8973 VP.n8918 VP.n8917 0.006
R8974 VP.n10429 VP.n10428 0.006
R8975 VP.n10464 VP.n10463 0.006
R8976 VP.n10159 VP.n10158 0.006
R8977 VP.n10096 VP.n10082 0.006
R8978 VP.n8962 VP.n8961 0.006
R8979 VP.n8118 VP.n8117 0.006
R8980 VP.n7290 VP.n7289 0.006
R8981 VP.n6431 VP.n6430 0.006
R8982 VP.n5575 VP.n5574 0.006
R8983 VP.n4680 VP.n4679 0.006
R8984 VP.n3781 VP.n3780 0.006
R8985 VP.n2836 VP.n2835 0.006
R8986 VP.n620 VP.n619 0.006
R8987 VP.n10970 VP.n10969 0.006
R8988 VP.n9708 VP.n9707 0.005
R8989 VP.n10064 VP.n10060 0.005
R8990 VP.n10994 VP.n10991 0.005
R8991 VP.n9605 VP.n9601 0.005
R8992 VP.n9629 VP.n9628 0.005
R8993 VP.n10935 VP.n10932 0.005
R8994 VP.n8799 VP.n8795 0.005
R8995 VP.n7964 VP.n7963 0.005
R8996 VP.n10884 VP.n10881 0.005
R8997 VP.n9969 VP.n9966 0.005
R8998 VP.n9212 VP.n9209 0.005
R8999 VP.n8412 VP.n8409 0.005
R9000 VP.n7076 VP.n7072 0.005
R9001 VP.n6277 VP.n6276 0.005
R9002 VP.n10833 VP.n10830 0.005
R9003 VP.n9921 VP.n9918 0.005
R9004 VP.n9162 VP.n9159 0.005
R9005 VP.n8363 VP.n8360 0.005
R9006 VP.n7546 VP.n7543 0.005
R9007 VP.n6734 VP.n6731 0.005
R9008 VP.n5297 VP.n5293 0.005
R9009 VP.n4526 VP.n4525 0.005
R9010 VP.n10782 VP.n10779 0.005
R9011 VP.n9873 VP.n9870 0.005
R9012 VP.n9112 VP.n9109 0.005
R9013 VP.n8314 VP.n8311 0.005
R9014 VP.n7497 VP.n7494 0.005
R9015 VP.n6685 VP.n6682 0.005
R9016 VP.n5843 VP.n5840 0.005
R9017 VP.n5006 VP.n5003 0.005
R9018 VP.n3420 VP.n3416 0.005
R9019 VP.n2320 VP.n2319 0.005
R9020 VP.n256 VP.n255 0.005
R9021 VP.n774 VP.n773 0.005
R9022 VP.n358 VP.n357 0.005
R9023 VP.n886 VP.n884 0.005
R9024 VP.n1323 VP.n1322 0.005
R9025 VP.n1763 VP.n1762 0.005
R9026 VP.n405 VP.n404 0.005
R9027 VP.n936 VP.n934 0.005
R9028 VP.n1451 VP.n1450 0.005
R9029 VP.n1873 VP.n1871 0.005
R9030 VP.n2299 VP.n2298 0.005
R9031 VP.n2724 VP.n2723 0.005
R9032 VP.n452 VP.n451 0.005
R9033 VP.n986 VP.n982 0.005
R9034 VP.n1489 VP.n1488 0.005
R9035 VP.n1925 VP.n1921 0.005
R9036 VP.n2551 VP.n2550 0.005
R9037 VP.n2854 VP.n2850 0.005
R9038 VP.n3249 VP.n3248 0.005
R9039 VP.n3664 VP.n3663 0.005
R9040 VP.n499 VP.n498 0.005
R9041 VP.n1036 VP.n1032 0.005
R9042 VP.n1527 VP.n1526 0.005
R9043 VP.n1977 VP.n1975 0.005
R9044 VP.n2513 VP.n2512 0.005
R9045 VP.n2906 VP.n2902 0.005
R9046 VP.n3429 VP.n3428 0.005
R9047 VP.n3799 VP.n3797 0.005
R9048 VP.n4170 VP.n4169 0.005
R9049 VP.n4570 VP.n4569 0.005
R9050 VP.n546 VP.n545 0.005
R9051 VP.n1086 VP.n1084 0.005
R9052 VP.n1565 VP.n1564 0.005
R9053 VP.n2029 VP.n2027 0.005
R9054 VP.n2475 VP.n2474 0.005
R9055 VP.n2958 VP.n2954 0.005
R9056 VP.n3467 VP.n3466 0.005
R9057 VP.n3851 VP.n3847 0.005
R9058 VP.n4346 VP.n4345 0.005
R9059 VP.n4734 VP.n4730 0.005
R9060 VP.n5076 VP.n5075 0.005
R9061 VP.n5465 VP.n5464 0.005
R9062 VP.n593 VP.n592 0.005
R9063 VP.n1136 VP.n1134 0.005
R9064 VP.n1603 VP.n1602 0.005
R9065 VP.n2081 VP.n2077 0.005
R9066 VP.n2443 VP.n2442 0.005
R9067 VP.n3010 VP.n3006 0.005
R9068 VP.n3505 VP.n3504 0.005
R9069 VP.n3903 VP.n3901 0.005
R9070 VP.n4384 VP.n4383 0.005
R9071 VP.n4786 VP.n4784 0.005
R9072 VP.n5306 VP.n5305 0.005
R9073 VP.n5623 VP.n5619 0.005
R9074 VP.n5940 VP.n5939 0.005
R9075 VP.n6321 VP.n6320 0.005
R9076 VP.n633 VP.n632 0.005
R9077 VP.n1174 VP.n1170 0.005
R9078 VP.n1635 VP.n1634 0.005
R9079 VP.n2122 VP.n2120 0.005
R9080 VP.n2411 VP.n2410 0.005
R9081 VP.n3051 VP.n3047 0.005
R9082 VP.n3537 VP.n3536 0.005
R9083 VP.n3944 VP.n3942 0.005
R9084 VP.n4416 VP.n4415 0.005
R9085 VP.n4827 VP.n4825 0.005
R9086 VP.n5338 VP.n5337 0.005
R9087 VP.n5664 VP.n5662 0.005
R9088 VP.n6166 VP.n6165 0.005
R9089 VP.n6508 VP.n6504 0.005
R9090 VP.n6804 VP.n6803 0.005
R9091 VP.n7180 VP.n7179 0.005
R9092 VP.n663 VP.n662 0.005
R9093 VP.n1214 VP.n1210 0.005
R9094 VP.n1667 VP.n1666 0.005
R9095 VP.n2163 VP.n2161 0.005
R9096 VP.n2379 VP.n2378 0.005
R9097 VP.n3092 VP.n3088 0.005
R9098 VP.n3569 VP.n3568 0.005
R9099 VP.n3985 VP.n3981 0.005
R9100 VP.n4448 VP.n4447 0.005
R9101 VP.n4868 VP.n4864 0.005
R9102 VP.n5370 VP.n5369 0.005
R9103 VP.n5705 VP.n5701 0.005
R9104 VP.n6198 VP.n6197 0.005
R9105 VP.n6549 VP.n6545 0.005
R9106 VP.n7085 VP.n7084 0.005
R9107 VP.n7361 VP.n7359 0.005
R9108 VP.n7643 VP.n7642 0.005
R9109 VP.n8008 VP.n8007 0.005
R9110 VP.n8859 VP.n8856 0.005
R9111 VP.n695 VP.n694 0.005
R9112 VP.n1255 VP.n1251 0.005
R9113 VP.n1699 VP.n1698 0.005
R9114 VP.n2204 VP.n2202 0.005
R9115 VP.n2347 VP.n2346 0.005
R9116 VP.n3133 VP.n3129 0.005
R9117 VP.n3601 VP.n3600 0.005
R9118 VP.n4026 VP.n4022 0.005
R9119 VP.n4480 VP.n4479 0.005
R9120 VP.n4909 VP.n4907 0.005
R9121 VP.n5402 VP.n5401 0.005
R9122 VP.n5746 VP.n5744 0.005
R9123 VP.n6230 VP.n6229 0.005
R9124 VP.n6590 VP.n6586 0.005
R9125 VP.n7117 VP.n7116 0.005
R9126 VP.n7402 VP.n7398 0.005
R9127 VP.n7917 VP.n7916 0.005
R9128 VP.n8218 VP.n8214 0.005
R9129 VP.n8482 VP.n8481 0.005
R9130 VP.n8842 VP.n8841 0.005
R9131 VP.n282 VP.n281 0.005
R9132 VP.n801 VP.n797 0.005
R9133 VP.n1354 VP.n1353 0.005
R9134 VP.n1787 VP.n1785 0.005
R9135 VP.n2671 VP.n2670 0.005
R9136 VP.n2747 VP.n2743 0.005
R9137 VP.n3280 VP.n3279 0.005
R9138 VP.n3687 VP.n3685 0.005
R9139 VP.n4201 VP.n4200 0.005
R9140 VP.n4596 VP.n4592 0.005
R9141 VP.n5107 VP.n5106 0.005
R9142 VP.n5488 VP.n5484 0.005
R9143 VP.n5971 VP.n5970 0.005
R9144 VP.n6344 VP.n6340 0.005
R9145 VP.n6835 VP.n6834 0.005
R9146 VP.n7203 VP.n7199 0.005
R9147 VP.n7674 VP.n7673 0.005
R9148 VP.n8031 VP.n8029 0.005
R9149 VP.n8513 VP.n8512 0.005
R9150 VP.n8875 VP.n8873 0.005
R9151 VP.n10103 VP.n10102 0.005
R9152 VP.n9716 VP.n9715 0.005
R9153 VP.n9853 VP.n9850 0.005
R9154 VP.n9091 VP.n9088 0.005
R9155 VP.n8294 VP.n8291 0.005
R9156 VP.n7477 VP.n7474 0.005
R9157 VP.n6665 VP.n6662 0.005
R9158 VP.n5822 VP.n5819 0.005
R9159 VP.n4985 VP.n4982 0.005
R9160 VP.n4102 VP.n4099 0.005
R9161 VP.n3210 VP.n3207 0.005
R9162 VP.n8851 VP.n8849 0.005
R9163 VP.n9272 VP.n9271 0.005
R9164 VP.n9632 VP.n9631 0.005
R9165 VP.n10039 VP.n10038 0.005
R9166 VP.n7606 VP.n7605 0.005
R9167 VP.n7967 VP.n7966 0.005
R9168 VP.n8445 VP.n8444 0.005
R9169 VP.n9243 VP.n9242 0.005
R9170 VP.n9999 VP.n9998 0.005
R9171 VP.n5903 VP.n5902 0.005
R9172 VP.n6280 VP.n6279 0.005
R9173 VP.n6767 VP.n6766 0.005
R9174 VP.n7577 VP.n7576 0.005
R9175 VP.n8394 VP.n8393 0.005
R9176 VP.n9193 VP.n9192 0.005
R9177 VP.n9951 VP.n9950 0.005
R9178 VP.n4133 VP.n4132 0.005
R9179 VP.n4529 VP.n4528 0.005
R9180 VP.n5039 VP.n5038 0.005
R9181 VP.n5874 VP.n5873 0.005
R9182 VP.n6716 VP.n6715 0.005
R9183 VP.n7528 VP.n7527 0.005
R9184 VP.n8345 VP.n8344 0.005
R9185 VP.n9143 VP.n9142 0.005
R9186 VP.n9903 VP.n9902 0.005
R9187 VP.n265 VP.n264 0.005
R9188 VP.n367 VP.n366 0.005
R9189 VP.n414 VP.n413 0.005
R9190 VP.n461 VP.n460 0.005
R9191 VP.n508 VP.n507 0.005
R9192 VP.n555 VP.n554 0.005
R9193 VP.n602 VP.n601 0.005
R9194 VP.n642 VP.n641 0.005
R9195 VP.n672 VP.n671 0.005
R9196 VP.n704 VP.n703 0.005
R9197 VP.n1722 VP.n1721 0.005
R9198 VP.n9836 VP.n9835 0.005
R9199 VP.n9073 VP.n9072 0.005
R9200 VP.n8276 VP.n8275 0.005
R9201 VP.n7460 VP.n7459 0.005
R9202 VP.n6648 VP.n6647 0.005
R9203 VP.n5804 VP.n5803 0.005
R9204 VP.n4967 VP.n4966 0.005
R9205 VP.n4084 VP.n4083 0.005
R9206 VP.n3193 VP.n3192 0.005
R9207 VP.n2329 VP.n2328 0.005
R9208 VP.n10455 VP.n10454 0.005
R9209 VP.n197 VP.n196 0.005
R9210 VP.n2839 VP.n2838 0.004
R9211 VP.n3389 VP.n3388 0.004
R9212 VP.n3784 VP.n3783 0.004
R9213 VP.n4308 VP.n4307 0.004
R9214 VP.n4683 VP.n4682 0.004
R9215 VP.n5213 VP.n5212 0.004
R9216 VP.n5578 VP.n5577 0.004
R9217 VP.n6078 VP.n6077 0.004
R9218 VP.n6434 VP.n6433 0.004
R9219 VP.n6942 VP.n6941 0.004
R9220 VP.n7293 VP.n7292 0.004
R9221 VP.n7780 VP.n7779 0.004
R9222 VP.n8121 VP.n8120 0.004
R9223 VP.n8619 VP.n8618 0.004
R9224 VP.n8965 VP.n8964 0.004
R9225 VP.n9418 VP.n9417 0.004
R9226 VP.n10756 VP.n10755 0.004
R9227 VP.n10162 VP.n10161 0.004
R9228 VP.n2249 VP.n2248 0.004
R9229 VP.n2336 VP.n2335 0.004
R9230 VP.n3200 VP.n3199 0.004
R9231 VP.n3363 VP.n3362 0.004
R9232 VP.n4091 VP.n4090 0.004
R9233 VP.n4284 VP.n4283 0.004
R9234 VP.n4974 VP.n4973 0.004
R9235 VP.n5190 VP.n5189 0.004
R9236 VP.n5811 VP.n5810 0.004
R9237 VP.n6054 VP.n6053 0.004
R9238 VP.n6655 VP.n6654 0.004
R9239 VP.n6918 VP.n6917 0.004
R9240 VP.n7467 VP.n7466 0.004
R9241 VP.n7757 VP.n7756 0.004
R9242 VP.n8283 VP.n8282 0.004
R9243 VP.n8596 VP.n8595 0.004
R9244 VP.n9080 VP.n9079 0.004
R9245 VP.n9392 VP.n9391 0.004
R9246 VP.n9843 VP.n9842 0.004
R9247 VP.n10737 VP.n10736 0.004
R9248 VP.n10462 VP.n10461 0.004
R9249 VP.n10427 VP.n10426 0.004
R9250 VP.n10955 VP.n10954 0.004
R9251 VP.n9603 VP.n9602 0.004
R9252 VP.n10051 VP.n10050 0.004
R9253 VP.n10981 VP.n10980 0.004
R9254 VP.n10618 VP.n10617 0.004
R9255 VP.n8797 VP.n8796 0.004
R9256 VP.n9255 VP.n9254 0.004
R9257 VP.n9616 VP.n9615 0.004
R9258 VP.n10011 VP.n10010 0.004
R9259 VP.n10922 VP.n10921 0.004
R9260 VP.n10580 VP.n10579 0.004
R9261 VP.n8754 VP.n8753 0.004
R9262 VP.n9040 VP.n9039 0.004
R9263 VP.n9572 VP.n9571 0.004
R9264 VP.n9805 VP.n9804 0.004
R9265 VP.n10909 VP.n10908 0.004
R9266 VP.n10398 VP.n10397 0.004
R9267 VP.n8203 VP.n8202 0.004
R9268 VP.n7906 VP.n7905 0.004
R9269 VP.n7074 VP.n7073 0.004
R9270 VP.n7589 VP.n7588 0.004
R9271 VP.n7951 VP.n7950 0.004
R9272 VP.n8417 VP.n8416 0.004
R9273 VP.n8727 VP.n8726 0.004
R9274 VP.n9217 VP.n9216 0.004
R9275 VP.n9533 VP.n9532 0.004
R9276 VP.n9974 VP.n9973 0.004
R9277 VP.n10871 VP.n10870 0.004
R9278 VP.n10545 VP.n10544 0.004
R9279 VP.n7031 VP.n7030 0.004
R9280 VP.n7345 VP.n7344 0.004
R9281 VP.n7880 VP.n7879 0.004
R9282 VP.n8166 VP.n8165 0.004
R9283 VP.n8716 VP.n8715 0.004
R9284 VP.n9010 VP.n9009 0.004
R9285 VP.n9520 VP.n9519 0.004
R9286 VP.n9783 VP.n9782 0.004
R9287 VP.n10858 VP.n10857 0.004
R9288 VP.n10381 VP.n10380 0.004
R9289 VP.n6493 VP.n6492 0.004
R9290 VP.n6155 VP.n6154 0.004
R9291 VP.n5295 VP.n5294 0.004
R9292 VP.n5886 VP.n5885 0.004
R9293 VP.n6264 VP.n6263 0.004
R9294 VP.n6739 VP.n6738 0.004
R9295 VP.n7004 VP.n7003 0.004
R9296 VP.n7551 VP.n7550 0.004
R9297 VP.n7842 VP.n7841 0.004
R9298 VP.n8368 VP.n8367 0.004
R9299 VP.n8679 VP.n8678 0.004
R9300 VP.n9167 VP.n9166 0.004
R9301 VP.n9482 VP.n9481 0.004
R9302 VP.n9926 VP.n9925 0.004
R9303 VP.n10820 VP.n10819 0.004
R9304 VP.n10510 VP.n10509 0.004
R9305 VP.n5252 VP.n5251 0.004
R9306 VP.n5607 VP.n5606 0.004
R9307 VP.n6129 VP.n6128 0.004
R9308 VP.n6456 VP.n6455 0.004
R9309 VP.n6992 VP.n6991 0.004
R9310 VP.n7315 VP.n7314 0.004
R9311 VP.n7830 VP.n7829 0.004
R9312 VP.n8143 VP.n8142 0.004
R9313 VP.n8668 VP.n8667 0.004
R9314 VP.n8987 VP.n8986 0.004
R9315 VP.n9469 VP.n9468 0.004
R9316 VP.n9761 VP.n9760 0.004
R9317 VP.n10807 VP.n10806 0.004
R9318 VP.n10364 VP.n10363 0.004
R9319 VP.n4719 VP.n4718 0.004
R9320 VP.n4335 VP.n4334 0.004
R9321 VP.n3418 VP.n3417 0.004
R9322 VP.n4116 VP.n4115 0.004
R9323 VP.n4513 VP.n4512 0.004
R9324 VP.n5011 VP.n5010 0.004
R9325 VP.n5225 VP.n5224 0.004
R9326 VP.n5848 VP.n5847 0.004
R9327 VP.n6091 VP.n6090 0.004
R9328 VP.n6690 VP.n6689 0.004
R9329 VP.n6955 VP.n6954 0.004
R9330 VP.n7502 VP.n7501 0.004
R9331 VP.n7793 VP.n7792 0.004
R9332 VP.n8319 VP.n8318 0.004
R9333 VP.n8631 VP.n8630 0.004
R9334 VP.n9117 VP.n9116 0.004
R9335 VP.n9431 VP.n9430 0.004
R9336 VP.n9878 VP.n9877 0.004
R9337 VP.n10769 VP.n10768 0.004
R9338 VP.n10475 VP.n10474 0.004
R9339 VP.n343 VP.n342 0.004
R9340 VP.n871 VP.n870 0.004
R9341 VP.n1413 VP.n1412 0.004
R9342 VP.n1857 VP.n1856 0.004
R9343 VP.n2625 VP.n2624 0.004
R9344 VP.n2810 VP.n2809 0.004
R9345 VP.n3336 VP.n3335 0.004
R9346 VP.n3750 VP.n3749 0.004
R9347 VP.n4257 VP.n4256 0.004
R9348 VP.n4656 VP.n4655 0.004
R9349 VP.n5163 VP.n5162 0.004
R9350 VP.n5551 VP.n5550 0.004
R9351 VP.n6027 VP.n6026 0.004
R9352 VP.n6407 VP.n6406 0.004
R9353 VP.n6891 VP.n6890 0.004
R9354 VP.n7266 VP.n7265 0.004
R9355 VP.n7730 VP.n7729 0.004
R9356 VP.n8094 VP.n8093 0.004
R9357 VP.n8569 VP.n8568 0.004
R9358 VP.n8938 VP.n8937 0.004
R9359 VP.n9363 VP.n9362 0.004
R9360 VP.n9739 VP.n9738 0.004
R9361 VP.n10708 VP.n10707 0.004
R9362 VP.n10142 VP.n10141 0.004
R9363 VP.n11020 VP.n11019 0.004
R9364 VP.n9706 VP.n9705 0.004
R9365 VP.n9341 VP.n9340 0.004
R9366 VP.n8915 VP.n8914 0.004
R9367 VP.n8548 VP.n8547 0.004
R9368 VP.n8071 VP.n8070 0.004
R9369 VP.n7709 VP.n7708 0.004
R9370 VP.n7243 VP.n7242 0.004
R9371 VP.n6870 VP.n6869 0.004
R9372 VP.n6384 VP.n6383 0.004
R9373 VP.n6006 VP.n6005 0.004
R9374 VP.n5528 VP.n5527 0.004
R9375 VP.n5142 VP.n5141 0.004
R9376 VP.n4633 VP.n4632 0.004
R9377 VP.n4236 VP.n4235 0.004
R9378 VP.n3727 VP.n3726 0.004
R9379 VP.n3315 VP.n3314 0.004
R9380 VP.n2787 VP.n2786 0.004
R9381 VP.n2650 VP.n2649 0.004
R9382 VP.n1827 VP.n1826 0.004
R9383 VP.n1389 VP.n1388 0.004
R9384 VP.n843 VP.n842 0.004
R9385 VP.n300 VP.n299 0.004
R9386 VP.n737 VP.n736 0.004
R9387 VP.n374 VP.n373 0.004
R9388 VP.n910 VP.n909 0.004
R9389 VP.n1738 VP.n1737 0.004
R9390 VP.n421 VP.n420 0.004
R9391 VP.n960 VP.n959 0.004
R9392 VP.n1472 VP.n1471 0.004
R9393 VP.n1897 VP.n1896 0.004
R9394 VP.n2699 VP.n2698 0.004
R9395 VP.n468 VP.n467 0.004
R9396 VP.n1010 VP.n1009 0.004
R9397 VP.n1510 VP.n1509 0.004
R9398 VP.n1949 VP.n1948 0.004
R9399 VP.n2572 VP.n2571 0.004
R9400 VP.n2878 VP.n2877 0.004
R9401 VP.n3639 VP.n3638 0.004
R9402 VP.n515 VP.n514 0.004
R9403 VP.n1060 VP.n1059 0.004
R9404 VP.n1548 VP.n1547 0.004
R9405 VP.n2001 VP.n2000 0.004
R9406 VP.n2534 VP.n2533 0.004
R9407 VP.n2930 VP.n2929 0.004
R9408 VP.n3450 VP.n3449 0.004
R9409 VP.n3823 VP.n3822 0.004
R9410 VP.n4545 VP.n4544 0.004
R9411 VP.n562 VP.n561 0.004
R9412 VP.n1110 VP.n1109 0.004
R9413 VP.n1586 VP.n1585 0.004
R9414 VP.n2053 VP.n2052 0.004
R9415 VP.n2496 VP.n2495 0.004
R9416 VP.n2982 VP.n2981 0.004
R9417 VP.n3488 VP.n3487 0.004
R9418 VP.n3875 VP.n3874 0.004
R9419 VP.n4367 VP.n4366 0.004
R9420 VP.n4758 VP.n4757 0.004
R9421 VP.n5440 VP.n5439 0.004
R9422 VP.n609 VP.n608 0.004
R9423 VP.n1160 VP.n1159 0.004
R9424 VP.n1624 VP.n1623 0.004
R9425 VP.n2105 VP.n2104 0.004
R9426 VP.n2464 VP.n2463 0.004
R9427 VP.n3034 VP.n3033 0.004
R9428 VP.n3526 VP.n3525 0.004
R9429 VP.n3927 VP.n3926 0.004
R9430 VP.n4405 VP.n4404 0.004
R9431 VP.n4810 VP.n4809 0.004
R9432 VP.n5327 VP.n5326 0.004
R9433 VP.n5647 VP.n5646 0.004
R9434 VP.n6296 VP.n6295 0.004
R9435 VP.n649 VP.n648 0.004
R9436 VP.n1198 VP.n1197 0.004
R9437 VP.n1656 VP.n1655 0.004
R9438 VP.n2146 VP.n2145 0.004
R9439 VP.n2432 VP.n2431 0.004
R9440 VP.n3075 VP.n3074 0.004
R9441 VP.n3558 VP.n3557 0.004
R9442 VP.n3968 VP.n3967 0.004
R9443 VP.n4437 VP.n4436 0.004
R9444 VP.n4851 VP.n4850 0.004
R9445 VP.n5359 VP.n5358 0.004
R9446 VP.n5688 VP.n5687 0.004
R9447 VP.n6187 VP.n6186 0.004
R9448 VP.n6532 VP.n6531 0.004
R9449 VP.n7155 VP.n7154 0.004
R9450 VP.n679 VP.n678 0.004
R9451 VP.n1238 VP.n1237 0.004
R9452 VP.n1688 VP.n1687 0.004
R9453 VP.n2187 VP.n2186 0.004
R9454 VP.n2400 VP.n2399 0.004
R9455 VP.n3116 VP.n3115 0.004
R9456 VP.n3590 VP.n3589 0.004
R9457 VP.n4009 VP.n4008 0.004
R9458 VP.n4469 VP.n4468 0.004
R9459 VP.n4892 VP.n4891 0.004
R9460 VP.n5391 VP.n5390 0.004
R9461 VP.n5729 VP.n5728 0.004
R9462 VP.n6219 VP.n6218 0.004
R9463 VP.n6573 VP.n6572 0.004
R9464 VP.n7106 VP.n7105 0.004
R9465 VP.n7385 VP.n7384 0.004
R9466 VP.n7983 VP.n7982 0.004
R9467 VP.n272 VP.n271 0.004
R9468 VP.n785 VP.n784 0.004
R9469 VP.n1344 VP.n1343 0.004
R9470 VP.n1774 VP.n1773 0.004
R9471 VP.n2661 VP.n2660 0.004
R9472 VP.n2734 VP.n2733 0.004
R9473 VP.n3270 VP.n3269 0.004
R9474 VP.n3674 VP.n3673 0.004
R9475 VP.n4191 VP.n4190 0.004
R9476 VP.n4580 VP.n4579 0.004
R9477 VP.n5097 VP.n5096 0.004
R9478 VP.n5475 VP.n5474 0.004
R9479 VP.n5961 VP.n5960 0.004
R9480 VP.n6331 VP.n6330 0.004
R9481 VP.n6825 VP.n6824 0.004
R9482 VP.n7190 VP.n7189 0.004
R9483 VP.n7664 VP.n7663 0.004
R9484 VP.n8018 VP.n8017 0.004
R9485 VP.n8503 VP.n8502 0.004
R9486 VP.n8864 VP.n8863 0.004
R9487 VP.n9648 VP.n9647 0.004
R9488 VP.n2228 VP.n2227 0.004
R9489 VP.n2368 VP.n2367 0.004
R9490 VP.n3157 VP.n3156 0.004
R9491 VP.n3622 VP.n3621 0.004
R9492 VP.n4050 VP.n4049 0.004
R9493 VP.n4501 VP.n4500 0.004
R9494 VP.n4933 VP.n4932 0.004
R9495 VP.n5423 VP.n5422 0.004
R9496 VP.n5770 VP.n5769 0.004
R9497 VP.n6251 VP.n6250 0.004
R9498 VP.n6614 VP.n6613 0.004
R9499 VP.n7138 VP.n7137 0.004
R9500 VP.n7426 VP.n7425 0.004
R9501 VP.n7938 VP.n7937 0.004
R9502 VP.n8242 VP.n8241 0.004
R9503 VP.n8814 VP.n8813 0.004
R9504 VP.n711 VP.n710 0.004
R9505 VP.n1279 VP.n1278 0.004
R9506 VP.n1720 VP.n1719 0.004
R9507 VP.n1441 VP.n1440 0.004
R9508 VP.n10095 VP.n10094 0.004
R9509 VP.n9961 VP.n9960 0.004
R9510 VP.n9204 VP.n9203 0.004
R9511 VP.n8404 VP.n8403 0.004
R9512 VP.n9913 VP.n9912 0.004
R9513 VP.n9154 VP.n9153 0.004
R9514 VP.n8355 VP.n8354 0.004
R9515 VP.n7538 VP.n7537 0.004
R9516 VP.n6726 VP.n6725 0.004
R9517 VP.n9865 VP.n9864 0.004
R9518 VP.n9104 VP.n9103 0.004
R9519 VP.n8306 VP.n8305 0.004
R9520 VP.n7489 VP.n7488 0.004
R9521 VP.n6677 VP.n6676 0.004
R9522 VP.n5835 VP.n5834 0.004
R9523 VP.n4998 VP.n4997 0.004
R9524 VP.n9845 VP.n9844 0.004
R9525 VP.n9083 VP.n9082 0.004
R9526 VP.n8286 VP.n8285 0.004
R9527 VP.n7469 VP.n7468 0.004
R9528 VP.n6657 VP.n6656 0.004
R9529 VP.n5814 VP.n5813 0.004
R9530 VP.n4977 VP.n4976 0.004
R9531 VP.n4094 VP.n4093 0.004
R9532 VP.n3202 VP.n3201 0.004
R9533 VP.n2822 VP.n2821 0.004
R9534 VP.n3373 VP.n3372 0.004
R9535 VP.n3762 VP.n3761 0.004
R9536 VP.n4294 VP.n4293 0.004
R9537 VP.n4668 VP.n4667 0.004
R9538 VP.n5200 VP.n5199 0.004
R9539 VP.n5563 VP.n5562 0.004
R9540 VP.n6065 VP.n6064 0.004
R9541 VP.n6419 VP.n6418 0.004
R9542 VP.n6929 VP.n6928 0.004
R9543 VP.n7278 VP.n7277 0.004
R9544 VP.n7767 VP.n7766 0.004
R9545 VP.n8106 VP.n8105 0.004
R9546 VP.n8606 VP.n8605 0.004
R9547 VP.n8950 VP.n8949 0.004
R9548 VP.n9403 VP.n9402 0.004
R9549 VP.n10748 VP.n10747 0.004
R9550 VP.n10153 VP.n10152 0.004
R9551 VP.n2263 VP.n2261 0.004
R9552 VP.n1747 VP.n1746 0.004
R9553 VP.n924 VP.n923 0.004
R9554 VP.n2708 VP.n2707 0.004
R9555 VP.n1913 VP.n1912 0.004
R9556 VP.n1480 VP.n1479 0.004
R9557 VP.n974 VP.n973 0.004
R9558 VP.n3648 VP.n3647 0.004
R9559 VP.n2894 VP.n2893 0.004
R9560 VP.n2580 VP.n2579 0.004
R9561 VP.n1965 VP.n1964 0.004
R9562 VP.n1518 VP.n1517 0.004
R9563 VP.n1024 VP.n1023 0.004
R9564 VP.n4554 VP.n4553 0.004
R9565 VP.n3839 VP.n3838 0.004
R9566 VP.n3458 VP.n3457 0.004
R9567 VP.n2946 VP.n2945 0.004
R9568 VP.n2542 VP.n2541 0.004
R9569 VP.n2017 VP.n2016 0.004
R9570 VP.n1556 VP.n1555 0.004
R9571 VP.n1074 VP.n1073 0.004
R9572 VP.n5449 VP.n5448 0.004
R9573 VP.n4774 VP.n4773 0.004
R9574 VP.n4375 VP.n4374 0.004
R9575 VP.n3891 VP.n3890 0.004
R9576 VP.n3496 VP.n3495 0.004
R9577 VP.n2998 VP.n2997 0.004
R9578 VP.n2504 VP.n2503 0.004
R9579 VP.n2069 VP.n2068 0.004
R9580 VP.n1594 VP.n1593 0.004
R9581 VP.n1124 VP.n1123 0.004
R9582 VP.n6305 VP.n6304 0.004
R9583 VP.n7164 VP.n7163 0.004
R9584 VP.n7992 VP.n7991 0.004
R9585 VP.n832 VP.n831 0.004
R9586 VP.n10021 VP.n10020 0.004
R9587 VP.n8770 VP.n8769 0.004
R9588 VP.n8183 VP.n8180 0.004
R9589 VP.n8427 VP.n8426 0.004
R9590 VP.n9227 VP.n9226 0.004
R9591 VP.n9984 VP.n9983 0.004
R9592 VP.n7047 VP.n7046 0.004
R9593 VP.n6473 VP.n6470 0.004
R9594 VP.n6749 VP.n6748 0.004
R9595 VP.n7561 VP.n7560 0.004
R9596 VP.n8378 VP.n8377 0.004
R9597 VP.n9177 VP.n9176 0.004
R9598 VP.n9936 VP.n9935 0.004
R9599 VP.n5268 VP.n5267 0.004
R9600 VP.n4699 VP.n4696 0.004
R9601 VP.n5021 VP.n5020 0.004
R9602 VP.n5858 VP.n5857 0.004
R9603 VP.n6700 VP.n6699 0.004
R9604 VP.n7512 VP.n7511 0.004
R9605 VP.n8329 VP.n8328 0.004
R9606 VP.n9127 VP.n9126 0.004
R9607 VP.n9888 VP.n9887 0.004
R9608 VP.n9821 VP.n9820 0.004
R9609 VP.n9057 VP.n9056 0.004
R9610 VP.n8260 VP.n8259 0.004
R9611 VP.n7444 VP.n7443 0.004
R9612 VP.n6632 VP.n6631 0.004
R9613 VP.n5788 VP.n5787 0.004
R9614 VP.n4951 VP.n4950 0.004
R9615 VP.n4068 VP.n4067 0.004
R9616 VP.n3175 VP.n3174 0.004
R9617 VP.n1442 VP.n1426 0.004
R9618 VP.n313 VP.n303 0.004
R9619 VP.n253 VP.n252 0.004
R9620 VP.n355 VP.n354 0.004
R9621 VP.n402 VP.n401 0.004
R9622 VP.n449 VP.n448 0.004
R9623 VP.n496 VP.n495 0.004
R9624 VP.n543 VP.n542 0.004
R9625 VP.n590 VP.n589 0.004
R9626 VP.n630 VP.n629 0.004
R9627 VP.n660 VP.n659 0.004
R9628 VP.n9656 VP.n9655 0.004
R9629 VP.n692 VP.n691 0.004
R9630 VP.n8822 VP.n8821 0.004
R9631 VP.n156 VP.n152 0.004
R9632 VP.n11028 VP.n11027 0.004
R9633 VP.n2844 VP.n2843 0.004
R9634 VP.n3394 VP.n3393 0.004
R9635 VP.n3789 VP.n3788 0.004
R9636 VP.n4313 VP.n4312 0.004
R9637 VP.n4688 VP.n4687 0.004
R9638 VP.n5218 VP.n5217 0.004
R9639 VP.n5583 VP.n5582 0.004
R9640 VP.n6083 VP.n6082 0.004
R9641 VP.n6439 VP.n6438 0.004
R9642 VP.n6947 VP.n6946 0.004
R9643 VP.n7298 VP.n7297 0.004
R9644 VP.n7785 VP.n7784 0.004
R9645 VP.n8126 VP.n8125 0.004
R9646 VP.n8624 VP.n8623 0.004
R9647 VP.n8970 VP.n8969 0.004
R9648 VP.n9423 VP.n9422 0.004
R9649 VP.n10761 VP.n10760 0.004
R9650 VP.n10167 VP.n10166 0.004
R9651 VP.t8 VP.n10204 0.004
R9652 VP.t8 VP.n10336 0.004
R9653 VP.t8 VP.n10324 0.004
R9654 VP.t8 VP.n10306 0.004
R9655 VP.t8 VP.n10290 0.004
R9656 VP.t8 VP.n10278 0.004
R9657 VP.t8 VP.n10262 0.004
R9658 VP.t8 VP.n10250 0.004
R9659 VP.t8 VP.n10234 0.004
R9660 VP.t8 VP.n10222 0.004
R9661 VP.t8 VP.n10339 0.004
R9662 VP.t116 VP.n129 0.004
R9663 VP.t6 VP.n10125 0.004
R9664 VP.t49 VP.n776 0.004
R9665 VP.t53 VP.n1765 0.004
R9666 VP.t108 VP.n2726 0.004
R9667 VP.t76 VP.n3666 0.004
R9668 VP.t169 VP.n4572 0.004
R9669 VP.t26 VP.n5467 0.004
R9670 VP.t159 VP.n6323 0.004
R9671 VP.t134 VP.n7182 0.004
R9672 VP.t18 VP.n8010 0.004
R9673 VP.t126 VP.n9685 0.004
R9674 VP.t207 VP.n8844 0.004
R9675 VP.t8 VP.n10341 0.004
R9676 VP.t116 VP.n201 0.004
R9677 VP.t116 VP.n205 0.004
R9678 VP.t116 VP.n209 0.004
R9679 VP.t116 VP.n213 0.004
R9680 VP.t116 VP.n217 0.004
R9681 VP.t116 VP.n221 0.004
R9682 VP.t116 VP.n225 0.004
R9683 VP.t116 VP.n229 0.004
R9684 VP.t116 VP.n233 0.004
R9685 VP.t116 VP.n237 0.004
R9686 VP.t116 VP.n142 0.004
R9687 VP.t116 VP.n241 0.004
R9688 VP.t8 VP.n10206 0.004
R9689 VP.t91 VP.n2690 0.004
R9690 VP.n2847 VP.n2846 0.003
R9691 VP.n3397 VP.n3396 0.003
R9692 VP.n3792 VP.n3791 0.003
R9693 VP.n4316 VP.n4315 0.003
R9694 VP.n4691 VP.n4690 0.003
R9695 VP.n5221 VP.n5220 0.003
R9696 VP.n5586 VP.n5585 0.003
R9697 VP.n6086 VP.n6085 0.003
R9698 VP.n6442 VP.n6441 0.003
R9699 VP.n6950 VP.n6949 0.003
R9700 VP.n7301 VP.n7300 0.003
R9701 VP.n7788 VP.n7787 0.003
R9702 VP.n8129 VP.n8128 0.003
R9703 VP.n8627 VP.n8626 0.003
R9704 VP.n8973 VP.n8972 0.003
R9705 VP.n9426 VP.n9425 0.003
R9706 VP.n10764 VP.n10763 0.003
R9707 VP.n10170 VP.n10169 0.003
R9708 VP.n1447 VP.n1446 0.003
R9709 VP.n2266 VP.n2265 0.003
R9710 VP.n2344 VP.n2343 0.003
R9711 VP.n3216 VP.n3215 0.003
R9712 VP.n3370 VP.n3369 0.003
R9713 VP.n4108 VP.n4107 0.003
R9714 VP.n4291 VP.n4290 0.003
R9715 VP.n4991 VP.n4990 0.003
R9716 VP.n5197 VP.n5196 0.003
R9717 VP.n5828 VP.n5827 0.003
R9718 VP.n6062 VP.n6061 0.003
R9719 VP.n6671 VP.n6670 0.003
R9720 VP.n6926 VP.n6925 0.003
R9721 VP.n7483 VP.n7482 0.003
R9722 VP.n7764 VP.n7763 0.003
R9723 VP.n8300 VP.n8299 0.003
R9724 VP.n8603 VP.n8602 0.003
R9725 VP.n9097 VP.n9096 0.003
R9726 VP.n9400 VP.n9399 0.003
R9727 VP.n9859 VP.n9858 0.003
R9728 VP.n10745 VP.n10744 0.003
R9729 VP.n10467 VP.n10466 0.003
R9730 VP.n10435 VP.n10434 0.003
R9731 VP.n10975 VP.n10974 0.003
R9732 VP.n9610 VP.n9609 0.003
R9733 VP.n10074 VP.n10073 0.003
R9734 VP.n11008 VP.n11007 0.003
R9735 VP.n10645 VP.n10644 0.003
R9736 VP.n8804 VP.n8803 0.003
R9737 VP.n9276 VP.n9275 0.003
R9738 VP.n9636 VP.n9635 0.003
R9739 VP.n10043 VP.n10042 0.003
R9740 VP.n10952 VP.n10951 0.003
R9741 VP.n10607 VP.n10606 0.003
R9742 VP.n8776 VP.n8775 0.003
R9743 VP.n9049 VP.n9048 0.003
R9744 VP.n9580 VP.n9579 0.003
R9745 VP.n9813 VP.n9812 0.003
R9746 VP.n10917 VP.n10916 0.003
R9747 VP.n10409 VP.n10408 0.003
R9748 VP.n8211 VP.n8210 0.003
R9749 VP.n7913 VP.n7912 0.003
R9750 VP.n7081 VP.n7080 0.003
R9751 VP.n7610 VP.n7609 0.003
R9752 VP.n7971 VP.n7970 0.003
R9753 VP.n8449 VP.n8448 0.003
R9754 VP.n8750 VP.n8749 0.003
R9755 VP.n9247 VP.n9246 0.003
R9756 VP.n9557 VP.n9556 0.003
R9757 VP.n10003 VP.n10002 0.003
R9758 VP.n10901 VP.n10900 0.003
R9759 VP.n10572 VP.n10571 0.003
R9760 VP.n7053 VP.n7052 0.003
R9761 VP.n7354 VP.n7353 0.003
R9762 VP.n7887 VP.n7886 0.003
R9763 VP.n8175 VP.n8174 0.003
R9764 VP.n8723 VP.n8722 0.003
R9765 VP.n9019 VP.n9018 0.003
R9766 VP.n9528 VP.n9527 0.003
R9767 VP.n9791 VP.n9790 0.003
R9768 VP.n10866 VP.n10865 0.003
R9769 VP.n10392 VP.n10391 0.003
R9770 VP.n6501 VP.n6500 0.003
R9771 VP.n6162 VP.n6161 0.003
R9772 VP.n5302 VP.n5301 0.003
R9773 VP.n5907 VP.n5906 0.003
R9774 VP.n6284 VP.n6283 0.003
R9775 VP.n6771 VP.n6770 0.003
R9776 VP.n7027 VP.n7026 0.003
R9777 VP.n7581 VP.n7580 0.003
R9778 VP.n7865 VP.n7864 0.003
R9779 VP.n8398 VP.n8397 0.003
R9780 VP.n8702 VP.n8701 0.003
R9781 VP.n9197 VP.n9196 0.003
R9782 VP.n9506 VP.n9505 0.003
R9783 VP.n9955 VP.n9954 0.003
R9784 VP.n10850 VP.n10849 0.003
R9785 VP.n10537 VP.n10536 0.003
R9786 VP.n5274 VP.n5273 0.003
R9787 VP.n5616 VP.n5615 0.003
R9788 VP.n6136 VP.n6135 0.003
R9789 VP.n6465 VP.n6464 0.003
R9790 VP.n6999 VP.n6998 0.003
R9791 VP.n7324 VP.n7323 0.003
R9792 VP.n7837 VP.n7836 0.003
R9793 VP.n8152 VP.n8151 0.003
R9794 VP.n8675 VP.n8674 0.003
R9795 VP.n8996 VP.n8995 0.003
R9796 VP.n9477 VP.n9476 0.003
R9797 VP.n9769 VP.n9768 0.003
R9798 VP.n10815 VP.n10814 0.003
R9799 VP.n10375 VP.n10374 0.003
R9800 VP.n4727 VP.n4726 0.003
R9801 VP.n4342 VP.n4341 0.003
R9802 VP.n3425 VP.n3424 0.003
R9803 VP.n4137 VP.n4136 0.003
R9804 VP.n4533 VP.n4532 0.003
R9805 VP.n5043 VP.n5042 0.003
R9806 VP.n5248 VP.n5247 0.003
R9807 VP.n5878 VP.n5877 0.003
R9808 VP.n6114 VP.n6113 0.003
R9809 VP.n6720 VP.n6719 0.003
R9810 VP.n6978 VP.n6977 0.003
R9811 VP.n7532 VP.n7531 0.003
R9812 VP.n7816 VP.n7815 0.003
R9813 VP.n8349 VP.n8348 0.003
R9814 VP.n8654 VP.n8653 0.003
R9815 VP.n9147 VP.n9146 0.003
R9816 VP.n9455 VP.n9454 0.003
R9817 VP.n9907 VP.n9906 0.003
R9818 VP.n10799 VP.n10798 0.003
R9819 VP.n10502 VP.n10501 0.003
R9820 VP.n350 VP.n349 0.003
R9821 VP.n879 VP.n878 0.003
R9822 VP.n1420 VP.n1419 0.003
R9823 VP.n1866 VP.n1865 0.003
R9824 VP.n2629 VP.n2628 0.003
R9825 VP.n2819 VP.n2818 0.003
R9826 VP.n3343 VP.n3342 0.003
R9827 VP.n3759 VP.n3758 0.003
R9828 VP.n4264 VP.n4263 0.003
R9829 VP.n4665 VP.n4664 0.003
R9830 VP.n5170 VP.n5169 0.003
R9831 VP.n5560 VP.n5559 0.003
R9832 VP.n6034 VP.n6033 0.003
R9833 VP.n6416 VP.n6415 0.003
R9834 VP.n6898 VP.n6897 0.003
R9835 VP.n7275 VP.n7274 0.003
R9836 VP.n7737 VP.n7736 0.003
R9837 VP.n8103 VP.n8102 0.003
R9838 VP.n8576 VP.n8575 0.003
R9839 VP.n8947 VP.n8946 0.003
R9840 VP.n9371 VP.n9370 0.003
R9841 VP.n9747 VP.n9746 0.003
R9842 VP.n10716 VP.n10715 0.003
R9843 VP.n10150 VP.n10149 0.003
R9844 VP.n11014 VP.n11013 0.003
R9845 VP.n9725 VP.n9724 0.003
R9846 VP.n9349 VP.n9348 0.003
R9847 VP.n8924 VP.n8923 0.003
R9848 VP.n8555 VP.n8554 0.003
R9849 VP.n8080 VP.n8079 0.003
R9850 VP.n7716 VP.n7715 0.003
R9851 VP.n7252 VP.n7251 0.003
R9852 VP.n6877 VP.n6876 0.003
R9853 VP.n6393 VP.n6392 0.003
R9854 VP.n6013 VP.n6012 0.003
R9855 VP.n5537 VP.n5536 0.003
R9856 VP.n5149 VP.n5148 0.003
R9857 VP.n4642 VP.n4641 0.003
R9858 VP.n4243 VP.n4242 0.003
R9859 VP.n3736 VP.n3735 0.003
R9860 VP.n3322 VP.n3321 0.003
R9861 VP.n2796 VP.n2795 0.003
R9862 VP.n2654 VP.n2653 0.003
R9863 VP.n1836 VP.n1835 0.003
R9864 VP.n1396 VP.n1395 0.003
R9865 VP.n850 VP.n849 0.003
R9866 VP.n319 VP.n318 0.003
R9867 VP.n731 VP.n730 0.003
R9868 VP.n395 VP.n394 0.003
R9869 VP.n927 VP.n926 0.003
R9870 VP.n1732 VP.n1731 0.003
R9871 VP.n442 VP.n441 0.003
R9872 VP.n977 VP.n976 0.003
R9873 VP.n1483 VP.n1482 0.003
R9874 VP.n1916 VP.n1915 0.003
R9875 VP.n2693 VP.n2692 0.003
R9876 VP.n489 VP.n488 0.003
R9877 VP.n1027 VP.n1026 0.003
R9878 VP.n1521 VP.n1520 0.003
R9879 VP.n1968 VP.n1967 0.003
R9880 VP.n2586 VP.n2585 0.003
R9881 VP.n2897 VP.n2896 0.003
R9882 VP.n3633 VP.n3632 0.003
R9883 VP.n536 VP.n535 0.003
R9884 VP.n1077 VP.n1076 0.003
R9885 VP.n1559 VP.n1558 0.003
R9886 VP.n2020 VP.n2019 0.003
R9887 VP.n2548 VP.n2547 0.003
R9888 VP.n2949 VP.n2948 0.003
R9889 VP.n3461 VP.n3460 0.003
R9890 VP.n3842 VP.n3841 0.003
R9891 VP.n4539 VP.n4538 0.003
R9892 VP.n583 VP.n582 0.003
R9893 VP.n1127 VP.n1126 0.003
R9894 VP.n1597 VP.n1596 0.003
R9895 VP.n2072 VP.n2071 0.003
R9896 VP.n2510 VP.n2509 0.003
R9897 VP.n3001 VP.n3000 0.003
R9898 VP.n3499 VP.n3498 0.003
R9899 VP.n3894 VP.n3893 0.003
R9900 VP.n4378 VP.n4377 0.003
R9901 VP.n4777 VP.n4776 0.003
R9902 VP.n5434 VP.n5433 0.003
R9903 VP.n623 VP.n622 0.003
R9904 VP.n1165 VP.n1164 0.003
R9905 VP.n1629 VP.n1628 0.003
R9906 VP.n2113 VP.n2112 0.003
R9907 VP.n2472 VP.n2471 0.003
R9908 VP.n3042 VP.n3041 0.003
R9909 VP.n3531 VP.n3530 0.003
R9910 VP.n3935 VP.n3934 0.003
R9911 VP.n4410 VP.n4409 0.003
R9912 VP.n4818 VP.n4817 0.003
R9913 VP.n5332 VP.n5331 0.003
R9914 VP.n5655 VP.n5654 0.003
R9915 VP.n6290 VP.n6289 0.003
R9916 VP.n653 VP.n652 0.003
R9917 VP.n1205 VP.n1204 0.003
R9918 VP.n1661 VP.n1660 0.003
R9919 VP.n2154 VP.n2153 0.003
R9920 VP.n2440 VP.n2439 0.003
R9921 VP.n3083 VP.n3082 0.003
R9922 VP.n3563 VP.n3562 0.003
R9923 VP.n3976 VP.n3975 0.003
R9924 VP.n4442 VP.n4441 0.003
R9925 VP.n4859 VP.n4858 0.003
R9926 VP.n5364 VP.n5363 0.003
R9927 VP.n5696 VP.n5695 0.003
R9928 VP.n6192 VP.n6191 0.003
R9929 VP.n6540 VP.n6539 0.003
R9930 VP.n7149 VP.n7148 0.003
R9931 VP.n685 VP.n684 0.003
R9932 VP.n1246 VP.n1245 0.003
R9933 VP.n1693 VP.n1692 0.003
R9934 VP.n2195 VP.n2194 0.003
R9935 VP.n2408 VP.n2407 0.003
R9936 VP.n3124 VP.n3123 0.003
R9937 VP.n3595 VP.n3594 0.003
R9938 VP.n4017 VP.n4016 0.003
R9939 VP.n4474 VP.n4473 0.003
R9940 VP.n4900 VP.n4899 0.003
R9941 VP.n5396 VP.n5395 0.003
R9942 VP.n5737 VP.n5736 0.003
R9943 VP.n6224 VP.n6223 0.003
R9944 VP.n6581 VP.n6580 0.003
R9945 VP.n7111 VP.n7110 0.003
R9946 VP.n7393 VP.n7392 0.003
R9947 VP.n7977 VP.n7976 0.003
R9948 VP.n293 VP.n292 0.003
R9949 VP.n788 VP.n787 0.003
R9950 VP.n1371 VP.n1370 0.003
R9951 VP.n1807 VP.n1806 0.003
R9952 VP.n2685 VP.n2684 0.003
R9953 VP.n2767 VP.n2766 0.003
R9954 VP.n3297 VP.n3296 0.003
R9955 VP.n3707 VP.n3706 0.003
R9956 VP.n4218 VP.n4217 0.003
R9957 VP.n4583 VP.n4582 0.003
R9958 VP.n5124 VP.n5123 0.003
R9959 VP.n5508 VP.n5507 0.003
R9960 VP.n5988 VP.n5987 0.003
R9961 VP.n6364 VP.n6363 0.003
R9962 VP.n6852 VP.n6851 0.003
R9963 VP.n7223 VP.n7222 0.003
R9964 VP.n7691 VP.n7690 0.003
R9965 VP.n8051 VP.n8050 0.003
R9966 VP.n8530 VP.n8529 0.003
R9967 VP.n8895 VP.n8894 0.003
R9968 VP.n9642 VP.n9641 0.003
R9969 VP.n2236 VP.n2235 0.003
R9970 VP.n2376 VP.n2375 0.003
R9971 VP.n3165 VP.n3164 0.003
R9972 VP.n3627 VP.n3626 0.003
R9973 VP.n4058 VP.n4057 0.003
R9974 VP.n4506 VP.n4505 0.003
R9975 VP.n4941 VP.n4940 0.003
R9976 VP.n5428 VP.n5427 0.003
R9977 VP.n5778 VP.n5777 0.003
R9978 VP.n6256 VP.n6255 0.003
R9979 VP.n6622 VP.n6621 0.003
R9980 VP.n7143 VP.n7142 0.003
R9981 VP.n7434 VP.n7433 0.003
R9982 VP.n7943 VP.n7942 0.003
R9983 VP.n8250 VP.n8249 0.003
R9984 VP.n8808 VP.n8807 0.003
R9985 VP.n725 VP.n724 0.003
R9986 VP.n1287 VP.n1286 0.003
R9987 VP.n1726 VP.n1725 0.003
R9988 VP.n2263 VP.n2246 0.003
R9989 VP.n2338 VP.n2333 0.003
R9990 VP.n3213 VP.n3197 0.003
R9991 VP.n3364 VP.n3360 0.003
R9992 VP.n4105 VP.n4088 0.003
R9993 VP.n4285 VP.n4281 0.003
R9994 VP.n4988 VP.n4971 0.003
R9995 VP.n5191 VP.n5187 0.003
R9996 VP.n5825 VP.n5808 0.003
R9997 VP.n6056 VP.n6051 0.003
R9998 VP.n6668 VP.n6652 0.003
R9999 VP.n6920 VP.n6915 0.003
R10000 VP.n7480 VP.n7464 0.003
R10001 VP.n7758 VP.n7754 0.003
R10002 VP.n8297 VP.n8280 0.003
R10003 VP.n8597 VP.n8593 0.003
R10004 VP.n9094 VP.n9077 0.003
R10005 VP.n9394 VP.n9389 0.003
R10006 VP.n9856 VP.n9840 0.003
R10007 VP.n10739 VP.n10734 0.003
R10008 VP.n10464 VP.n10459 0.003
R10009 VP.n10429 VP.n10424 0.003
R10010 VP.n10071 VP.n10054 0.003
R10011 VP.n11005 VP.n10984 0.003
R10012 VP.n10642 VP.n10621 0.003
R10013 VP.n9273 VP.n9258 0.003
R10014 VP.n9633 VP.n9619 0.003
R10015 VP.n10040 VP.n10014 0.003
R10016 VP.n10946 VP.n10925 0.003
R10017 VP.n10604 VP.n10583 0.003
R10018 VP.n8770 VP.n8757 0.003
R10019 VP.n9043 VP.n9037 0.003
R10020 VP.n9574 VP.n9569 0.003
R10021 VP.n9807 VP.n9802 0.003
R10022 VP.n10911 VP.n10906 0.003
R10023 VP.n10403 VP.n10401 0.003
R10024 VP.n8205 VP.n8200 0.003
R10025 VP.n7607 VP.n7592 0.003
R10026 VP.n7968 VP.n7954 0.003
R10027 VP.n8446 VP.n8420 0.003
R10028 VP.n8744 VP.n8730 0.003
R10029 VP.n9244 VP.n9220 0.003
R10030 VP.n9551 VP.n9536 0.003
R10031 VP.n10000 VP.n9977 0.003
R10032 VP.n10895 VP.n10874 0.003
R10033 VP.n10569 VP.n10548 0.003
R10034 VP.n7047 VP.n7034 0.003
R10035 VP.n7348 VP.n7342 0.003
R10036 VP.n7881 VP.n7877 0.003
R10037 VP.n8169 VP.n8163 0.003
R10038 VP.n8717 VP.n8713 0.003
R10039 VP.n9013 VP.n9007 0.003
R10040 VP.n9522 VP.n9517 0.003
R10041 VP.n9785 VP.n9780 0.003
R10042 VP.n10860 VP.n10855 0.003
R10043 VP.n10386 VP.n10384 0.003
R10044 VP.n6495 VP.n6490 0.003
R10045 VP.n5904 VP.n5889 0.003
R10046 VP.n6281 VP.n6267 0.003
R10047 VP.n6768 VP.n6742 0.003
R10048 VP.n7021 VP.n7007 0.003
R10049 VP.n7578 VP.n7554 0.003
R10050 VP.n7859 VP.n7845 0.003
R10051 VP.n8395 VP.n8371 0.003
R10052 VP.n8696 VP.n8682 0.003
R10053 VP.n9194 VP.n9170 0.003
R10054 VP.n9500 VP.n9485 0.003
R10055 VP.n9952 VP.n9929 0.003
R10056 VP.n10844 VP.n10823 0.003
R10057 VP.n10534 VP.n10513 0.003
R10058 VP.n5268 VP.n5255 0.003
R10059 VP.n5610 VP.n5604 0.003
R10060 VP.n6130 VP.n6126 0.003
R10061 VP.n6459 VP.n6453 0.003
R10062 VP.n6993 VP.n6989 0.003
R10063 VP.n7318 VP.n7312 0.003
R10064 VP.n7831 VP.n7827 0.003
R10065 VP.n8146 VP.n8140 0.003
R10066 VP.n8669 VP.n8665 0.003
R10067 VP.n8990 VP.n8984 0.003
R10068 VP.n9471 VP.n9466 0.003
R10069 VP.n9763 VP.n9758 0.003
R10070 VP.n10809 VP.n10804 0.003
R10071 VP.n10369 VP.n10367 0.003
R10072 VP.n4721 VP.n4716 0.003
R10073 VP.n4134 VP.n4119 0.003
R10074 VP.n4530 VP.n4516 0.003
R10075 VP.n5040 VP.n5014 0.003
R10076 VP.n5242 VP.n5228 0.003
R10077 VP.n5875 VP.n5851 0.003
R10078 VP.n6108 VP.n6094 0.003
R10079 VP.n6717 VP.n6693 0.003
R10080 VP.n6972 VP.n6958 0.003
R10081 VP.n7529 VP.n7505 0.003
R10082 VP.n7810 VP.n7796 0.003
R10083 VP.n8346 VP.n8322 0.003
R10084 VP.n8648 VP.n8634 0.003
R10085 VP.n9144 VP.n9120 0.003
R10086 VP.n9449 VP.n9434 0.003
R10087 VP.n9904 VP.n9881 0.003
R10088 VP.n10793 VP.n10772 0.003
R10089 VP.n10499 VP.n10478 0.003
R10090 VP.n873 VP.n868 0.003
R10091 VP.n1414 VP.n1410 0.003
R10092 VP.n1860 VP.n1854 0.003
R10093 VP.n2626 VP.n2622 0.003
R10094 VP.n2813 VP.n2807 0.003
R10095 VP.n3337 VP.n3333 0.003
R10096 VP.n3753 VP.n3747 0.003
R10097 VP.n4258 VP.n4254 0.003
R10098 VP.n4659 VP.n4653 0.003
R10099 VP.n5164 VP.n5160 0.003
R10100 VP.n5554 VP.n5548 0.003
R10101 VP.n6028 VP.n6024 0.003
R10102 VP.n6410 VP.n6404 0.003
R10103 VP.n6892 VP.n6888 0.003
R10104 VP.n7269 VP.n7263 0.003
R10105 VP.n7731 VP.n7727 0.003
R10106 VP.n8097 VP.n8091 0.003
R10107 VP.n8570 VP.n8566 0.003
R10108 VP.n8941 VP.n8935 0.003
R10109 VP.n9365 VP.n9360 0.003
R10110 VP.n9741 VP.n9736 0.003
R10111 VP.n10710 VP.n10705 0.003
R10112 VP.n10144 VP.n10139 0.003
R10113 VP.n11032 VP.n10690 0.003
R10114 VP.n9719 VP.n9703 0.003
R10115 VP.n9343 VP.n9338 0.003
R10116 VP.n8918 VP.n8912 0.003
R10117 VP.n8549 VP.n8545 0.003
R10118 VP.n8074 VP.n8068 0.003
R10119 VP.n7710 VP.n7706 0.003
R10120 VP.n7246 VP.n7240 0.003
R10121 VP.n6871 VP.n6867 0.003
R10122 VP.n6387 VP.n6381 0.003
R10123 VP.n6007 VP.n6003 0.003
R10124 VP.n5531 VP.n5525 0.003
R10125 VP.n5143 VP.n5139 0.003
R10126 VP.n4636 VP.n4630 0.003
R10127 VP.n4237 VP.n4233 0.003
R10128 VP.n3730 VP.n3724 0.003
R10129 VP.n3316 VP.n3312 0.003
R10130 VP.n2790 VP.n2784 0.003
R10131 VP.n2651 VP.n2647 0.003
R10132 VP.n1830 VP.n1824 0.003
R10133 VP.n1390 VP.n1386 0.003
R10134 VP.n847 VP.n840 0.003
R10135 VP.n313 VP.n297 0.003
R10136 VP.n758 VP.n268 0.003
R10137 VP.n392 VP.n371 0.003
R10138 VP.n924 VP.n907 0.003
R10139 VP.n1747 VP.n1340 0.003
R10140 VP.n439 VP.n418 0.003
R10141 VP.n974 VP.n957 0.003
R10142 VP.n1480 VP.n1469 0.003
R10143 VP.n1913 VP.n1894 0.003
R10144 VP.n2708 VP.n2316 0.003
R10145 VP.n486 VP.n465 0.003
R10146 VP.n1024 VP.n1007 0.003
R10147 VP.n1518 VP.n1507 0.003
R10148 VP.n1965 VP.n1946 0.003
R10149 VP.n2580 VP.n2569 0.003
R10150 VP.n2894 VP.n2875 0.003
R10151 VP.n3648 VP.n3266 0.003
R10152 VP.n533 VP.n512 0.003
R10153 VP.n1074 VP.n1057 0.003
R10154 VP.n1556 VP.n1545 0.003
R10155 VP.n2017 VP.n1998 0.003
R10156 VP.n2542 VP.n2531 0.003
R10157 VP.n2946 VP.n2927 0.003
R10158 VP.n3458 VP.n3447 0.003
R10159 VP.n3839 VP.n3820 0.003
R10160 VP.n4554 VP.n4187 0.003
R10161 VP.n580 VP.n559 0.003
R10162 VP.n1124 VP.n1107 0.003
R10163 VP.n1594 VP.n1583 0.003
R10164 VP.n2069 VP.n2050 0.003
R10165 VP.n2504 VP.n2493 0.003
R10166 VP.n2998 VP.n2979 0.003
R10167 VP.n3496 VP.n3485 0.003
R10168 VP.n3891 VP.n3872 0.003
R10169 VP.n4375 VP.n4364 0.003
R10170 VP.n4774 VP.n4755 0.003
R10171 VP.n5449 VP.n5093 0.003
R10172 VP.n620 VP.n606 0.003
R10173 VP.n1162 VP.n1157 0.003
R10174 VP.n1626 VP.n1621 0.003
R10175 VP.n2110 VP.n2102 0.003
R10176 VP.n2466 VP.n2461 0.003
R10177 VP.n3039 VP.n3031 0.003
R10178 VP.n3528 VP.n3523 0.003
R10179 VP.n3932 VP.n3924 0.003
R10180 VP.n4407 VP.n4402 0.003
R10181 VP.n4815 VP.n4807 0.003
R10182 VP.n5329 VP.n5324 0.003
R10183 VP.n5652 VP.n5644 0.003
R10184 VP.n6305 VP.n5957 0.003
R10185 VP.n650 VP.n646 0.003
R10186 VP.n1202 VP.n1195 0.003
R10187 VP.n1658 VP.n1653 0.003
R10188 VP.n2151 VP.n2143 0.003
R10189 VP.n2434 VP.n2429 0.003
R10190 VP.n3080 VP.n3072 0.003
R10191 VP.n3560 VP.n3555 0.003
R10192 VP.n3973 VP.n3965 0.003
R10193 VP.n4439 VP.n4434 0.003
R10194 VP.n4856 VP.n4848 0.003
R10195 VP.n5361 VP.n5356 0.003
R10196 VP.n5693 VP.n5685 0.003
R10197 VP.n6189 VP.n6184 0.003
R10198 VP.n6537 VP.n6529 0.003
R10199 VP.n7164 VP.n6821 0.003
R10200 VP.n682 VP.n676 0.003
R10201 VP.n1243 VP.n1235 0.003
R10202 VP.n1690 VP.n1685 0.003
R10203 VP.n2192 VP.n2184 0.003
R10204 VP.n2402 VP.n2397 0.003
R10205 VP.n3121 VP.n3113 0.003
R10206 VP.n3592 VP.n3587 0.003
R10207 VP.n4014 VP.n4006 0.003
R10208 VP.n4471 VP.n4466 0.003
R10209 VP.n4897 VP.n4889 0.003
R10210 VP.n5393 VP.n5388 0.003
R10211 VP.n5734 VP.n5726 0.003
R10212 VP.n6221 VP.n6216 0.003
R10213 VP.n6578 VP.n6570 0.003
R10214 VP.n7108 VP.n7103 0.003
R10215 VP.n7390 VP.n7382 0.003
R10216 VP.n7992 VP.n7660 0.003
R10217 VP.n287 VP.n275 0.003
R10218 VP.n815 VP.n791 0.003
R10219 VP.n1365 VP.n1347 0.003
R10220 VP.n1801 VP.n1777 0.003
R10221 VP.n2682 VP.n2664 0.003
R10222 VP.n2761 VP.n2737 0.003
R10223 VP.n3291 VP.n3273 0.003
R10224 VP.n3701 VP.n3677 0.003
R10225 VP.n4212 VP.n4194 0.003
R10226 VP.n4610 VP.n4586 0.003
R10227 VP.n5118 VP.n5100 0.003
R10228 VP.n5502 VP.n5478 0.003
R10229 VP.n5982 VP.n5964 0.003
R10230 VP.n6358 VP.n6334 0.003
R10231 VP.n6846 VP.n6828 0.003
R10232 VP.n7217 VP.n7193 0.003
R10233 VP.n7685 VP.n7667 0.003
R10234 VP.n8045 VP.n8021 0.003
R10235 VP.n8524 VP.n8506 0.003
R10236 VP.n8889 VP.n8867 0.003
R10237 VP.n9659 VP.n9323 0.003
R10238 VP.n2233 VP.n2225 0.003
R10239 VP.n2370 VP.n2365 0.003
R10240 VP.n3162 VP.n3154 0.003
R10241 VP.n3624 VP.n3619 0.003
R10242 VP.n4055 VP.n4047 0.003
R10243 VP.n4503 VP.n4498 0.003
R10244 VP.n4938 VP.n4930 0.003
R10245 VP.n5425 VP.n5420 0.003
R10246 VP.n5775 VP.n5767 0.003
R10247 VP.n6253 VP.n6248 0.003
R10248 VP.n6619 VP.n6611 0.003
R10249 VP.n7140 VP.n7135 0.003
R10250 VP.n7431 VP.n7423 0.003
R10251 VP.n7940 VP.n7935 0.003
R10252 VP.n8247 VP.n8239 0.003
R10253 VP.n8826 VP.n8499 0.003
R10254 VP.n722 VP.n708 0.003
R10255 VP.n1284 VP.n1276 0.003
R10256 VP.n1723 VP.n1717 0.003
R10257 VP.n10123 VP.n10122 0.003
R10258 VP.n10096 VP.n10079 0.003
R10259 VP.n10096 VP.n10081 0.003
R10260 VP.n9657 VP.n9656 0.003
R10261 VP.n8823 VP.n8822 0.003
R10262 VP.n11029 VP.n11028 0.003
R10263 VP.n196 VP.n192 0.003
R10264 VP.n196 VP.n189 0.003
R10265 VP.n196 VP.n186 0.003
R10266 VP.n196 VP.n183 0.003
R10267 VP.n196 VP.n180 0.003
R10268 VP.n196 VP.n177 0.003
R10269 VP.n196 VP.n174 0.003
R10270 VP.n196 VP.n171 0.003
R10271 VP.n196 VP.n168 0.003
R10272 VP.n196 VP.n165 0.003
R10273 VP.n2832 VP.n2830 0.003
R10274 VP.n196 VP.n162 0.002
R10275 VP.n164 VP.n163 0.002
R10276 VP.n167 VP.n166 0.002
R10277 VP.n170 VP.n169 0.002
R10278 VP.n173 VP.n172 0.002
R10279 VP.n176 VP.n175 0.002
R10280 VP.n179 VP.n178 0.002
R10281 VP.n182 VP.n181 0.002
R10282 VP.n185 VP.n184 0.002
R10283 VP.n188 VP.n187 0.002
R10284 VP.n191 VP.n190 0.002
R10285 VP.n194 VP.n193 0.002
R10286 VP.n161 VP.n160 0.002
R10287 VP.n10454 VP.n10453 0.002
R10288 VP.n9835 VP.n9834 0.002
R10289 VP.n9072 VP.n9071 0.002
R10290 VP.n8275 VP.n8274 0.002
R10291 VP.n7459 VP.n7458 0.002
R10292 VP.n6647 VP.n6646 0.002
R10293 VP.n5803 VP.n5802 0.002
R10294 VP.n4966 VP.n4965 0.002
R10295 VP.n4083 VP.n4082 0.002
R10296 VP.n2328 VP.n2327 0.002
R10297 VP.n9631 VP.n9627 0.002
R10298 VP.n7966 VP.n7962 0.002
R10299 VP.n9242 VP.n9238 0.002
R10300 VP.n9998 VP.n9994 0.002
R10301 VP.n6279 VP.n6275 0.002
R10302 VP.n7576 VP.n7572 0.002
R10303 VP.n8393 VP.n8389 0.002
R10304 VP.n9192 VP.n9188 0.002
R10305 VP.n9950 VP.n9946 0.002
R10306 VP.n4528 VP.n4524 0.002
R10307 VP.n5873 VP.n5869 0.002
R10308 VP.n6715 VP.n6711 0.002
R10309 VP.n7527 VP.n7523 0.002
R10310 VP.n8344 VP.n8340 0.002
R10311 VP.n9142 VP.n9138 0.002
R10312 VP.n9902 VP.n9898 0.002
R10313 VP.n2241 VP.n2240 0.002
R10314 VP.n8196 VP.n8185 0.002
R10315 VP.n6486 VP.n6475 0.002
R10316 VP.n4712 VP.n4701 0.002
R10317 VP.n10065 VP.n10064 0.002
R10318 VP.n10066 VP.n10065 0.002
R10319 VP.n10995 VP.n10994 0.002
R10320 VP.n10996 VP.n10995 0.002
R10321 VP.n10936 VP.n10935 0.002
R10322 VP.n10937 VP.n10936 0.002
R10323 VP.n10885 VP.n10884 0.002
R10324 VP.n10886 VP.n10885 0.002
R10325 VP.n10834 VP.n10833 0.002
R10326 VP.n10835 VP.n10834 0.002
R10327 VP.n10783 VP.n10782 0.002
R10328 VP.n10784 VP.n10783 0.002
R10329 VP.n1426 VP.n1424 0.002
R10330 VP.n756 VP.n755 0.002
R10331 VP.n887 VP.n886 0.002
R10332 VP.n888 VP.n887 0.002
R10333 VP.n1324 VP.n1323 0.002
R10334 VP.n1325 VP.n1324 0.002
R10335 VP.n937 VP.n936 0.002
R10336 VP.n938 VP.n937 0.002
R10337 VP.n1452 VP.n1451 0.002
R10338 VP.n1453 VP.n1452 0.002
R10339 VP.n1874 VP.n1873 0.002
R10340 VP.n1875 VP.n1874 0.002
R10341 VP.n2300 VP.n2299 0.002
R10342 VP.n2301 VP.n2300 0.002
R10343 VP.n987 VP.n986 0.002
R10344 VP.n988 VP.n987 0.002
R10345 VP.n1490 VP.n1489 0.002
R10346 VP.n1491 VP.n1490 0.002
R10347 VP.n1926 VP.n1925 0.002
R10348 VP.n1927 VP.n1926 0.002
R10349 VP.n2552 VP.n2551 0.002
R10350 VP.n2553 VP.n2552 0.002
R10351 VP.n2855 VP.n2854 0.002
R10352 VP.n2856 VP.n2855 0.002
R10353 VP.n3250 VP.n3249 0.002
R10354 VP.n3251 VP.n3250 0.002
R10355 VP.n1037 VP.n1036 0.002
R10356 VP.n1038 VP.n1037 0.002
R10357 VP.n1528 VP.n1527 0.002
R10358 VP.n1529 VP.n1528 0.002
R10359 VP.n1978 VP.n1977 0.002
R10360 VP.n1979 VP.n1978 0.002
R10361 VP.n2514 VP.n2513 0.002
R10362 VP.n2515 VP.n2514 0.002
R10363 VP.n2907 VP.n2906 0.002
R10364 VP.n2908 VP.n2907 0.002
R10365 VP.n3430 VP.n3429 0.002
R10366 VP.n3431 VP.n3430 0.002
R10367 VP.n3800 VP.n3799 0.002
R10368 VP.n3801 VP.n3800 0.002
R10369 VP.n4171 VP.n4170 0.002
R10370 VP.n4172 VP.n4171 0.002
R10371 VP.n1087 VP.n1086 0.002
R10372 VP.n1088 VP.n1087 0.002
R10373 VP.n1566 VP.n1565 0.002
R10374 VP.n1567 VP.n1566 0.002
R10375 VP.n2030 VP.n2029 0.002
R10376 VP.n2031 VP.n2030 0.002
R10377 VP.n2476 VP.n2475 0.002
R10378 VP.n2477 VP.n2476 0.002
R10379 VP.n2959 VP.n2958 0.002
R10380 VP.n2960 VP.n2959 0.002
R10381 VP.n3468 VP.n3467 0.002
R10382 VP.n3469 VP.n3468 0.002
R10383 VP.n3852 VP.n3851 0.002
R10384 VP.n3853 VP.n3852 0.002
R10385 VP.n4347 VP.n4346 0.002
R10386 VP.n4348 VP.n4347 0.002
R10387 VP.n4735 VP.n4734 0.002
R10388 VP.n4736 VP.n4735 0.002
R10389 VP.n5077 VP.n5076 0.002
R10390 VP.n5078 VP.n5077 0.002
R10391 VP.n1137 VP.n1136 0.002
R10392 VP.n1138 VP.n1137 0.002
R10393 VP.n1604 VP.n1603 0.002
R10394 VP.n1605 VP.n1604 0.002
R10395 VP.n2082 VP.n2081 0.002
R10396 VP.n2083 VP.n2082 0.002
R10397 VP.n2444 VP.n2443 0.002
R10398 VP.n2445 VP.n2444 0.002
R10399 VP.n3011 VP.n3010 0.002
R10400 VP.n3012 VP.n3011 0.002
R10401 VP.n3506 VP.n3505 0.002
R10402 VP.n3507 VP.n3506 0.002
R10403 VP.n3904 VP.n3903 0.002
R10404 VP.n3905 VP.n3904 0.002
R10405 VP.n4385 VP.n4384 0.002
R10406 VP.n4386 VP.n4385 0.002
R10407 VP.n4787 VP.n4786 0.002
R10408 VP.n4788 VP.n4787 0.002
R10409 VP.n5307 VP.n5306 0.002
R10410 VP.n5308 VP.n5307 0.002
R10411 VP.n5624 VP.n5623 0.002
R10412 VP.n5625 VP.n5624 0.002
R10413 VP.n5941 VP.n5940 0.002
R10414 VP.n5942 VP.n5941 0.002
R10415 VP.n1175 VP.n1174 0.002
R10416 VP.n1176 VP.n1175 0.002
R10417 VP.n1636 VP.n1635 0.002
R10418 VP.n1637 VP.n1636 0.002
R10419 VP.n2123 VP.n2122 0.002
R10420 VP.n2124 VP.n2123 0.002
R10421 VP.n2412 VP.n2411 0.002
R10422 VP.n2413 VP.n2412 0.002
R10423 VP.n3052 VP.n3051 0.002
R10424 VP.n3053 VP.n3052 0.002
R10425 VP.n3538 VP.n3537 0.002
R10426 VP.n3539 VP.n3538 0.002
R10427 VP.n3945 VP.n3944 0.002
R10428 VP.n3946 VP.n3945 0.002
R10429 VP.n4417 VP.n4416 0.002
R10430 VP.n4418 VP.n4417 0.002
R10431 VP.n4828 VP.n4827 0.002
R10432 VP.n4829 VP.n4828 0.002
R10433 VP.n5339 VP.n5338 0.002
R10434 VP.n5340 VP.n5339 0.002
R10435 VP.n5665 VP.n5664 0.002
R10436 VP.n5666 VP.n5665 0.002
R10437 VP.n6167 VP.n6166 0.002
R10438 VP.n6168 VP.n6167 0.002
R10439 VP.n6509 VP.n6508 0.002
R10440 VP.n6510 VP.n6509 0.002
R10441 VP.n6805 VP.n6804 0.002
R10442 VP.n6806 VP.n6805 0.002
R10443 VP.n1215 VP.n1214 0.002
R10444 VP.n1216 VP.n1215 0.002
R10445 VP.n1668 VP.n1667 0.002
R10446 VP.n1669 VP.n1668 0.002
R10447 VP.n2164 VP.n2163 0.002
R10448 VP.n2165 VP.n2164 0.002
R10449 VP.n2380 VP.n2379 0.002
R10450 VP.n2381 VP.n2380 0.002
R10451 VP.n3093 VP.n3092 0.002
R10452 VP.n3094 VP.n3093 0.002
R10453 VP.n3570 VP.n3569 0.002
R10454 VP.n3571 VP.n3570 0.002
R10455 VP.n3986 VP.n3985 0.002
R10456 VP.n3987 VP.n3986 0.002
R10457 VP.n4449 VP.n4448 0.002
R10458 VP.n4450 VP.n4449 0.002
R10459 VP.n4869 VP.n4868 0.002
R10460 VP.n4870 VP.n4869 0.002
R10461 VP.n5371 VP.n5370 0.002
R10462 VP.n5372 VP.n5371 0.002
R10463 VP.n5706 VP.n5705 0.002
R10464 VP.n5707 VP.n5706 0.002
R10465 VP.n6199 VP.n6198 0.002
R10466 VP.n6200 VP.n6199 0.002
R10467 VP.n6550 VP.n6549 0.002
R10468 VP.n6551 VP.n6550 0.002
R10469 VP.n7086 VP.n7085 0.002
R10470 VP.n7087 VP.n7086 0.002
R10471 VP.n7362 VP.n7361 0.002
R10472 VP.n7363 VP.n7362 0.002
R10473 VP.n7644 VP.n7643 0.002
R10474 VP.n7645 VP.n7644 0.002
R10475 VP.n1256 VP.n1255 0.002
R10476 VP.n1257 VP.n1256 0.002
R10477 VP.n1700 VP.n1699 0.002
R10478 VP.n1701 VP.n1700 0.002
R10479 VP.n2205 VP.n2204 0.002
R10480 VP.n2206 VP.n2205 0.002
R10481 VP.n2348 VP.n2347 0.002
R10482 VP.n2349 VP.n2348 0.002
R10483 VP.n3134 VP.n3133 0.002
R10484 VP.n3135 VP.n3134 0.002
R10485 VP.n3602 VP.n3601 0.002
R10486 VP.n3603 VP.n3602 0.002
R10487 VP.n4027 VP.n4026 0.002
R10488 VP.n4028 VP.n4027 0.002
R10489 VP.n4481 VP.n4480 0.002
R10490 VP.n4482 VP.n4481 0.002
R10491 VP.n4910 VP.n4909 0.002
R10492 VP.n4911 VP.n4910 0.002
R10493 VP.n5403 VP.n5402 0.002
R10494 VP.n5404 VP.n5403 0.002
R10495 VP.n5747 VP.n5746 0.002
R10496 VP.n5748 VP.n5747 0.002
R10497 VP.n6231 VP.n6230 0.002
R10498 VP.n6232 VP.n6231 0.002
R10499 VP.n6591 VP.n6590 0.002
R10500 VP.n6592 VP.n6591 0.002
R10501 VP.n7118 VP.n7117 0.002
R10502 VP.n7119 VP.n7118 0.002
R10503 VP.n7403 VP.n7402 0.002
R10504 VP.n7404 VP.n7403 0.002
R10505 VP.n7918 VP.n7917 0.002
R10506 VP.n7919 VP.n7918 0.002
R10507 VP.n8219 VP.n8218 0.002
R10508 VP.n8220 VP.n8219 0.002
R10509 VP.n8483 VP.n8482 0.002
R10510 VP.n8484 VP.n8483 0.002
R10511 VP.n283 VP.n282 0.002
R10512 VP.n284 VP.n283 0.002
R10513 VP.n802 VP.n801 0.002
R10514 VP.n803 VP.n802 0.002
R10515 VP.n1355 VP.n1354 0.002
R10516 VP.n1356 VP.n1355 0.002
R10517 VP.n1788 VP.n1787 0.002
R10518 VP.n1789 VP.n1788 0.002
R10519 VP.n2672 VP.n2671 0.002
R10520 VP.n2673 VP.n2672 0.002
R10521 VP.n2748 VP.n2747 0.002
R10522 VP.n2749 VP.n2748 0.002
R10523 VP.n3281 VP.n3280 0.002
R10524 VP.n3282 VP.n3281 0.002
R10525 VP.n3688 VP.n3687 0.002
R10526 VP.n3689 VP.n3688 0.002
R10527 VP.n4202 VP.n4201 0.002
R10528 VP.n4203 VP.n4202 0.002
R10529 VP.n4597 VP.n4596 0.002
R10530 VP.n4598 VP.n4597 0.002
R10531 VP.n5108 VP.n5107 0.002
R10532 VP.n5109 VP.n5108 0.002
R10533 VP.n5489 VP.n5488 0.002
R10534 VP.n5490 VP.n5489 0.002
R10535 VP.n5972 VP.n5971 0.002
R10536 VP.n5973 VP.n5972 0.002
R10537 VP.n6345 VP.n6344 0.002
R10538 VP.n6346 VP.n6345 0.002
R10539 VP.n6836 VP.n6835 0.002
R10540 VP.n6837 VP.n6836 0.002
R10541 VP.n7204 VP.n7203 0.002
R10542 VP.n7205 VP.n7204 0.002
R10543 VP.n7675 VP.n7674 0.002
R10544 VP.n7676 VP.n7675 0.002
R10545 VP.n8032 VP.n8031 0.002
R10546 VP.n8033 VP.n8032 0.002
R10547 VP.n8514 VP.n8513 0.002
R10548 VP.n8515 VP.n8514 0.002
R10549 VP.n8876 VP.n8875 0.002
R10550 VP.n8877 VP.n8876 0.002
R10551 VP.n157 VP.n156 0.002
R10552 VP.n10350 VP.n10349 0.002
R10553 VP.n3192 VP.n3191 0.002
R10554 VP.n10038 VP.n10034 0.002
R10555 VP.n8444 VP.n8440 0.002
R10556 VP.n6766 VP.n6762 0.002
R10557 VP.n5038 VP.n5034 0.002
R10558 VP.t8 VP.n10182 0.002
R10559 VP.n1771 VP.n1769 0.002
R10560 VP.n196 VP.n195 0.002
R10561 VP.n10352 VP.n10351 0.001
R10562 VP.t8 VP.n10352 0.001
R10563 VP.n10174 VP.n10172 0.001
R10564 VP.n8205 VP.n8197 0.001
R10565 VP.n8770 VP.n8751 0.001
R10566 VP.n9043 VP.n9034 0.001
R10567 VP.n9574 VP.n9566 0.001
R10568 VP.n9807 VP.n9799 0.001
R10569 VP.n10911 VP.n10903 0.001
R10570 VP.n6495 VP.n6487 0.001
R10571 VP.n7047 VP.n7028 0.001
R10572 VP.n7348 VP.n7339 0.001
R10573 VP.n7881 VP.n7874 0.001
R10574 VP.n8169 VP.n8160 0.001
R10575 VP.n8717 VP.n8710 0.001
R10576 VP.n9013 VP.n9004 0.001
R10577 VP.n9522 VP.n9514 0.001
R10578 VP.n9785 VP.n9777 0.001
R10579 VP.n10860 VP.n10852 0.001
R10580 VP.n4721 VP.n4713 0.001
R10581 VP.n5268 VP.n5249 0.001
R10582 VP.n5610 VP.n5601 0.001
R10583 VP.n6130 VP.n6123 0.001
R10584 VP.n6459 VP.n6450 0.001
R10585 VP.n6993 VP.n6986 0.001
R10586 VP.n7318 VP.n7309 0.001
R10587 VP.n7831 VP.n7824 0.001
R10588 VP.n8146 VP.n8137 0.001
R10589 VP.n8669 VP.n8662 0.001
R10590 VP.n8990 VP.n8981 0.001
R10591 VP.n9471 VP.n9463 0.001
R10592 VP.n9763 VP.n9755 0.001
R10593 VP.n10809 VP.n10801 0.001
R10594 VP.n2836 VP.n2834 0.001
R10595 VP.n3386 VP.n3385 0.001
R10596 VP.n3781 VP.n3778 0.001
R10597 VP.n4305 VP.n4304 0.001
R10598 VP.n4680 VP.n4677 0.001
R10599 VP.n5210 VP.n5209 0.001
R10600 VP.n5575 VP.n5572 0.001
R10601 VP.n6075 VP.n6074 0.001
R10602 VP.n6431 VP.n6428 0.001
R10603 VP.n6939 VP.n6938 0.001
R10604 VP.n7290 VP.n7287 0.001
R10605 VP.n7777 VP.n7776 0.001
R10606 VP.n8118 VP.n8115 0.001
R10607 VP.n8616 VP.n8615 0.001
R10608 VP.n8962 VP.n8959 0.001
R10609 VP.n9415 VP.n9413 0.001
R10610 VP.n10096 VP.n10083 0.001
R10611 VP.n10753 VP.n10750 0.001
R10612 VP.n873 VP.n865 0.001
R10613 VP.n1414 VP.n1407 0.001
R10614 VP.n1860 VP.n1851 0.001
R10615 VP.n2626 VP.n2619 0.001
R10616 VP.n2813 VP.n2804 0.001
R10617 VP.n3337 VP.n3330 0.001
R10618 VP.n3753 VP.n3744 0.001
R10619 VP.n4258 VP.n4251 0.001
R10620 VP.n4659 VP.n4650 0.001
R10621 VP.n5164 VP.n5157 0.001
R10622 VP.n5554 VP.n5545 0.001
R10623 VP.n6028 VP.n6021 0.001
R10624 VP.n6410 VP.n6401 0.001
R10625 VP.n6892 VP.n6885 0.001
R10626 VP.n7269 VP.n7260 0.001
R10627 VP.n7731 VP.n7724 0.001
R10628 VP.n8097 VP.n8088 0.001
R10629 VP.n8570 VP.n8563 0.001
R10630 VP.n8941 VP.n8932 0.001
R10631 VP.n9365 VP.n9357 0.001
R10632 VP.n9741 VP.n9733 0.001
R10633 VP.n10710 VP.n10702 0.001
R10634 VP.n10144 VP.n10136 0.001
R10635 VP.n313 VP.n294 0.001
R10636 VP.n847 VP.n837 0.001
R10637 VP.n1390 VP.n1383 0.001
R10638 VP.n1830 VP.n1821 0.001
R10639 VP.n2651 VP.n2644 0.001
R10640 VP.n2790 VP.n2781 0.001
R10641 VP.n3316 VP.n3309 0.001
R10642 VP.n3730 VP.n3721 0.001
R10643 VP.n4237 VP.n4230 0.001
R10644 VP.n4636 VP.n4627 0.001
R10645 VP.n5143 VP.n5136 0.001
R10646 VP.n5531 VP.n5522 0.001
R10647 VP.n6007 VP.n6000 0.001
R10648 VP.n6387 VP.n6378 0.001
R10649 VP.n6871 VP.n6864 0.001
R10650 VP.n7246 VP.n7237 0.001
R10651 VP.n7710 VP.n7703 0.001
R10652 VP.n8074 VP.n8065 0.001
R10653 VP.n8549 VP.n8542 0.001
R10654 VP.n8918 VP.n8909 0.001
R10655 VP.n9343 VP.n9335 0.001
R10656 VP.n9719 VP.n9700 0.001
R10657 VP.n10671 VP.n10670 0.001
R10658 VP.n9671 VP.n9670 0.001
R10659 VP.n9292 VP.n9291 0.001
R10660 VP.n8465 VP.n8464 0.001
R10661 VP.n7626 VP.n7625 0.001
R10662 VP.n6787 VP.n6786 0.001
R10663 VP.n5923 VP.n5922 0.001
R10664 VP.n5059 VP.n5058 0.001
R10665 VP.n4153 VP.n4152 0.001
R10666 VP.n3232 VP.n3231 0.001
R10667 VP.n2282 VP.n2281 0.001
R10668 VP.n1305 VP.n1304 0.001
R10669 VP.n325 VP.n324 0.001
R10670 VP.n10966 VP.n10965 0.001
R10671 VP.n9591 VP.n9590 0.001
R10672 VP.n8787 VP.n8786 0.001
R10673 VP.n7900 VP.n7899 0.001
R10674 VP.n7064 VP.n7063 0.001
R10675 VP.n6149 VP.n6148 0.001
R10676 VP.n5285 VP.n5284 0.001
R10677 VP.n4329 VP.n4328 0.001
R10678 VP.n3408 VP.n3407 0.001
R10679 VP.n2603 VP.n2602 0.001
R10680 VP.n1437 VP.n1436 0.001
R10681 VP.n339 VP.n338 0.001
R10682 VP.n10695 VP.n10694 0.001
R10683 VP.n249 VP.n244 0.001
R10684 VP.n1319 VP.n1292 0.001
R10685 VP.n2295 VP.n2271 0.001
R10686 VP.n3245 VP.n3221 0.001
R10687 VP.n4166 VP.n4142 0.001
R10688 VP.n5072 VP.n5048 0.001
R10689 VP.n5936 VP.n5912 0.001
R10690 VP.n6800 VP.n6776 0.001
R10691 VP.n7639 VP.n7615 0.001
R10692 VP.n8478 VP.n8454 0.001
R10693 VP.n10112 VP.n10101 0.001
R10694 VP.n9305 VP.n9281 0.001
R10695 VP.n10675 VP.n10650 0.001
R10696 VP.n2610 VP.n2609 0.001
R10697 VP.n10063 VP.n10062 0.001
R10698 VP.n10993 VP.n10992 0.001
R10699 VP.n10019 VP.n10018 0.001
R10700 VP.n10934 VP.n10933 0.001
R10701 VP.n8425 VP.n8424 0.001
R10702 VP.n9225 VP.n9224 0.001
R10703 VP.n9982 VP.n9981 0.001
R10704 VP.n10883 VP.n10882 0.001
R10705 VP.n6747 VP.n6746 0.001
R10706 VP.n7559 VP.n7558 0.001
R10707 VP.n8376 VP.n8375 0.001
R10708 VP.n9175 VP.n9174 0.001
R10709 VP.n9934 VP.n9933 0.001
R10710 VP.n10832 VP.n10831 0.001
R10711 VP.n5019 VP.n5018 0.001
R10712 VP.n5856 VP.n5855 0.001
R10713 VP.n6698 VP.n6697 0.001
R10714 VP.n7510 VP.n7509 0.001
R10715 VP.n8327 VP.n8326 0.001
R10716 VP.n9125 VP.n9124 0.001
R10717 VP.n9886 VP.n9885 0.001
R10718 VP.n10781 VP.n10780 0.001
R10719 VP.n9817 VP.n9816 0.001
R10720 VP.n9053 VP.n9052 0.001
R10721 VP.n8256 VP.n8255 0.001
R10722 VP.n7440 VP.n7439 0.001
R10723 VP.n6628 VP.n6627 0.001
R10724 VP.n5784 VP.n5783 0.001
R10725 VP.n4947 VP.n4946 0.001
R10726 VP.n4064 VP.n4063 0.001
R10727 VP.n3171 VP.n3170 0.001
R10728 VP.n1414 VP.n1397 0.001
R10729 VP.n744 VP.n743 0.001
R10730 VP.t116 VP.n128 0.001
R10731 VP.t116 VP.n120 0.001
R10732 VP.n763 VP.n762 0.001
R10733 VP.n2289 VP.n2288 0.001
R10734 VP.n387 VP.n386 0.001
R10735 VP.t116 VP.n115 0.001
R10736 VP.t116 VP.n107 0.001
R10737 VP.n890 VP.n889 0.001
R10738 VP.n1752 VP.n1751 0.001
R10739 VP.n3239 VP.n3238 0.001
R10740 VP.n434 VP.n433 0.001
R10741 VP.t116 VP.n102 0.001
R10742 VP.t116 VP.n96 0.001
R10743 VP.n940 VP.n939 0.001
R10744 VP.n1877 VP.n1876 0.001
R10745 VP.n2713 VP.n2712 0.001
R10746 VP.n4160 VP.n4159 0.001
R10747 VP.n481 VP.n480 0.001
R10748 VP.t116 VP.n89 0.001
R10749 VP.t116 VP.n81 0.001
R10750 VP.n990 VP.n989 0.001
R10751 VP.n985 VP.n984 0.001
R10752 VP.n1929 VP.n1928 0.001
R10753 VP.n1924 VP.n1923 0.001
R10754 VP.n2858 VP.n2857 0.001
R10755 VP.n2853 VP.n2852 0.001
R10756 VP.n3653 VP.n3652 0.001
R10757 VP.n5066 VP.n5065 0.001
R10758 VP.n528 VP.n527 0.001
R10759 VP.t116 VP.n76 0.001
R10760 VP.t116 VP.n70 0.001
R10761 VP.n1040 VP.n1039 0.001
R10762 VP.n1035 VP.n1034 0.001
R10763 VP.n1981 VP.n1980 0.001
R10764 VP.n2910 VP.n2909 0.001
R10765 VP.n2905 VP.n2904 0.001
R10766 VP.n3803 VP.n3802 0.001
R10767 VP.n4559 VP.n4558 0.001
R10768 VP.n5930 VP.n5929 0.001
R10769 VP.n575 VP.n574 0.001
R10770 VP.t116 VP.n63 0.001
R10771 VP.t116 VP.n55 0.001
R10772 VP.n1090 VP.n1089 0.001
R10773 VP.n2033 VP.n2032 0.001
R10774 VP.n2962 VP.n2961 0.001
R10775 VP.n2957 VP.n2956 0.001
R10776 VP.n3855 VP.n3854 0.001
R10777 VP.n3850 VP.n3849 0.001
R10778 VP.n4738 VP.n4737 0.001
R10779 VP.n4733 VP.n4732 0.001
R10780 VP.n5454 VP.n5453 0.001
R10781 VP.n6794 VP.n6793 0.001
R10782 VP.n615 VP.n614 0.001
R10783 VP.t116 VP.n50 0.001
R10784 VP.t116 VP.n44 0.001
R10785 VP.n1140 VP.n1139 0.001
R10786 VP.n2085 VP.n2084 0.001
R10787 VP.n2080 VP.n2079 0.001
R10788 VP.n3014 VP.n3013 0.001
R10789 VP.n3009 VP.n3008 0.001
R10790 VP.n3907 VP.n3906 0.001
R10791 VP.n4790 VP.n4789 0.001
R10792 VP.n5627 VP.n5626 0.001
R10793 VP.n5622 VP.n5621 0.001
R10794 VP.n6310 VP.n6309 0.001
R10795 VP.n7633 VP.n7632 0.001
R10796 VP.t116 VP.n34 0.001
R10797 VP.n1178 VP.n1177 0.001
R10798 VP.n1173 VP.n1172 0.001
R10799 VP.n2126 VP.n2125 0.001
R10800 VP.n3055 VP.n3054 0.001
R10801 VP.n3050 VP.n3049 0.001
R10802 VP.n3948 VP.n3947 0.001
R10803 VP.n4831 VP.n4830 0.001
R10804 VP.n5668 VP.n5667 0.001
R10805 VP.n6512 VP.n6511 0.001
R10806 VP.n6507 VP.n6506 0.001
R10807 VP.n7169 VP.n7168 0.001
R10808 VP.n8472 VP.n8471 0.001
R10809 VP.t116 VP.n24 0.001
R10810 VP.n1218 VP.n1217 0.001
R10811 VP.n1213 VP.n1212 0.001
R10812 VP.n2167 VP.n2166 0.001
R10813 VP.n3096 VP.n3095 0.001
R10814 VP.n3091 VP.n3090 0.001
R10815 VP.n3989 VP.n3988 0.001
R10816 VP.n3984 VP.n3983 0.001
R10817 VP.n4872 VP.n4871 0.001
R10818 VP.n4867 VP.n4866 0.001
R10819 VP.n5709 VP.n5708 0.001
R10820 VP.n5704 VP.n5703 0.001
R10821 VP.n6553 VP.n6552 0.001
R10822 VP.n6548 VP.n6547 0.001
R10823 VP.n7365 VP.n7364 0.001
R10824 VP.n7997 VP.n7996 0.001
R10825 VP.n9678 VP.n9677 0.001
R10826 VP.n717 VP.n716 0.001
R10827 VP.t116 VP.n17 0.001
R10828 VP.n1259 VP.n1258 0.001
R10829 VP.n1254 VP.n1253 0.001
R10830 VP.n2208 VP.n2207 0.001
R10831 VP.n3137 VP.n3136 0.001
R10832 VP.n3132 VP.n3131 0.001
R10833 VP.n4030 VP.n4029 0.001
R10834 VP.n4025 VP.n4024 0.001
R10835 VP.n4913 VP.n4912 0.001
R10836 VP.n5750 VP.n5749 0.001
R10837 VP.n6594 VP.n6593 0.001
R10838 VP.n6589 VP.n6588 0.001
R10839 VP.n7406 VP.n7405 0.001
R10840 VP.n7401 VP.n7400 0.001
R10841 VP.n8222 VP.n8221 0.001
R10842 VP.n8217 VP.n8216 0.001
R10843 VP.n8831 VP.n8830 0.001
R10844 VP.n9299 VP.n9298 0.001
R10845 VP.t116 VP.n135 0.001
R10846 VP.n805 VP.n804 0.001
R10847 VP.n800 VP.n799 0.001
R10848 VP.n1791 VP.n1790 0.001
R10849 VP.n2751 VP.n2750 0.001
R10850 VP.n2746 VP.n2745 0.001
R10851 VP.n3691 VP.n3690 0.001
R10852 VP.n4600 VP.n4599 0.001
R10853 VP.n4595 VP.n4594 0.001
R10854 VP.n5492 VP.n5491 0.001
R10855 VP.n5487 VP.n5486 0.001
R10856 VP.n6348 VP.n6347 0.001
R10857 VP.n6343 VP.n6342 0.001
R10858 VP.n7207 VP.n7206 0.001
R10859 VP.n7202 VP.n7201 0.001
R10860 VP.n8035 VP.n8034 0.001
R10861 VP.n8879 VP.n8878 0.001
R10862 VP.n10652 VP.n10651 0.001
R10863 VP.n249 VP.n248 0.001
R10864 VP.n249 VP.n4 0.001
R10865 VP.n3386 VP.n3375 0.001
R10866 VP.n2844 VP.n2841 0.001
R10867 VP.t108 VP.n2844 0.001
R10868 VP.n3394 VP.n3391 0.001
R10869 VP.t72 VP.n3394 0.001
R10870 VP.n3789 VP.n3786 0.001
R10871 VP.t76 VP.n3789 0.001
R10872 VP.n4313 VP.n4310 0.001
R10873 VP.t140 VP.n4313 0.001
R10874 VP.n4688 VP.n4685 0.001
R10875 VP.t169 VP.n4688 0.001
R10876 VP.n5218 VP.n5215 0.001
R10877 VP.t119 VP.n5218 0.001
R10878 VP.n5583 VP.n5580 0.001
R10879 VP.t26 VP.n5583 0.001
R10880 VP.n6083 VP.n6080 0.001
R10881 VP.t24 VP.n6083 0.001
R10882 VP.n6439 VP.n6436 0.001
R10883 VP.t159 VP.n6439 0.001
R10884 VP.n6947 VP.n6944 0.001
R10885 VP.t195 VP.n6947 0.001
R10886 VP.n7298 VP.n7295 0.001
R10887 VP.t134 VP.n7298 0.001
R10888 VP.n7785 VP.n7782 0.001
R10889 VP.t111 VP.n7785 0.001
R10890 VP.n8126 VP.n8123 0.001
R10891 VP.t18 VP.n8126 0.001
R10892 VP.n8624 VP.n8621 0.001
R10893 VP.t28 VP.n8624 0.001
R10894 VP.n8970 VP.n8967 0.001
R10895 VP.t207 VP.n8970 0.001
R10896 VP.n9423 VP.n9420 0.001
R10897 VP.t143 VP.n9423 0.001
R10898 VP.n10761 VP.n10758 0.001
R10899 VP.t16 VP.n10761 0.001
R10900 VP.n10167 VP.n10164 0.001
R10901 VP.t6 VP.n10167 0.001
R10902 VP.n10964 VP.n10963 0.001
R10903 VP.n9589 VP.n9588 0.001
R10904 VP.n8785 VP.n8784 0.001
R10905 VP.n7898 VP.n7897 0.001
R10906 VP.n7062 VP.n7061 0.001
R10907 VP.n6147 VP.n6146 0.001
R10908 VP.n5283 VP.n5282 0.001
R10909 VP.n4327 VP.n4326 0.001
R10910 VP.n3406 VP.n3405 0.001
R10911 VP.n2601 VP.n2600 0.001
R10912 VP.n1435 VP.n1434 0.001
R10913 VP.n337 VP.n336 0.001
R10914 VP.t91 VP.n2610 0.001
R10915 VP.n10650 VP.t6 0.001
R10916 VP.n1292 VP.t49 0.001
R10917 VP.n2271 VP.t53 0.001
R10918 VP.n3221 VP.t108 0.001
R10919 VP.n4142 VP.t76 0.001
R10920 VP.n5048 VP.t169 0.001
R10921 VP.n5912 VP.t26 0.001
R10922 VP.n6776 VP.t159 0.001
R10923 VP.n7615 VP.t134 0.001
R10924 VP.n8454 VP.t18 0.001
R10925 VP.n10101 VP.t126 0.001
R10926 VP.n9281 VP.t207 0.001
R10927 VP.n244 VP.t116 0.001
R10928 VP.n10695 VP.n10693 0.001
R10929 VP.n196 VP.n194 0.001
R10930 VP.n196 VP.n191 0.001
R10931 VP.n196 VP.n188 0.001
R10932 VP.n196 VP.n185 0.001
R10933 VP.n196 VP.n182 0.001
R10934 VP.n196 VP.n179 0.001
R10935 VP.n196 VP.n176 0.001
R10936 VP.n196 VP.n173 0.001
R10937 VP.n196 VP.n170 0.001
R10938 VP.n196 VP.n167 0.001
R10939 VP.n196 VP.n164 0.001
R10940 VP.n11034 VP.n10675 0.001
R10941 VP.n1320 VP.n1319 0.001
R10942 VP.n2296 VP.n2295 0.001
R10943 VP.n3246 VP.n3245 0.001
R10944 VP.n4167 VP.n4166 0.001
R10945 VP.n5073 VP.n5072 0.001
R10946 VP.n5937 VP.n5936 0.001
R10947 VP.n6801 VP.n6800 0.001
R10948 VP.n7640 VP.n7639 0.001
R10949 VP.n8479 VP.n8478 0.001
R10950 VP.n10113 VP.n10112 0.001
R10951 VP.n10965 VP.n10964 0.001
R10952 VP.n9590 VP.n9589 0.001
R10953 VP.n8786 VP.n8785 0.001
R10954 VP.n7899 VP.n7898 0.001
R10955 VP.n7063 VP.n7062 0.001
R10956 VP.n6148 VP.n6147 0.001
R10957 VP.n5284 VP.n5283 0.001
R10958 VP.n4328 VP.n4327 0.001
R10959 VP.n3407 VP.n3406 0.001
R10960 VP.n2602 VP.n2601 0.001
R10961 VP.n1436 VP.n1435 0.001
R10962 VP.n338 VP.n337 0.001
R10963 VP.n10174 VP.n10173 0.001
R10964 VP.n10672 VP.n10671 0.001
R10965 VP.n9672 VP.n9671 0.001
R10966 VP.n9293 VP.n9292 0.001
R10967 VP.n8466 VP.n8465 0.001
R10968 VP.n7627 VP.n7626 0.001
R10969 VP.n6788 VP.n6787 0.001
R10970 VP.n5924 VP.n5923 0.001
R10971 VP.n5060 VP.n5059 0.001
R10972 VP.n4154 VP.n4153 0.001
R10973 VP.n3233 VP.n3232 0.001
R10974 VP.n2283 VP.n2282 0.001
R10975 VP.n1306 VP.n1305 0.001
R10976 VP.n324 VP.n323 0.001
R10977 VP.n10403 VP.n10394 0.001
R10978 VP.n10386 VP.n10377 0.001
R10979 VP.n10369 VP.n10360 0.001
R10980 VP.n10159 VP.n10157 0.001
R10981 VP.n11033 VP.n11032 0.001
R10982 VP.n9660 VP.n9659 0.001
R10983 VP.n10429 VP.n10421 0.001
R10984 VP.n10351 VP.n10343 0.001
R10985 VP.n10970 VP.n10953 0.001
R10986 VP.n9605 VP.n9604 0.001
R10987 VP.n8799 VP.n8798 0.001
R10988 VP.n7908 VP.n7907 0.001
R10989 VP.n7076 VP.n7075 0.001
R10990 VP.n6157 VP.n6156 0.001
R10991 VP.n5297 VP.n5296 0.001
R10992 VP.n4337 VP.n4336 0.001
R10993 VP.n3420 VP.n3419 0.001
R10994 VP.n345 VP.n344 0.001
R10995 VP.n1442 VP.n1421 0.001
R10996 VP.n2609 VP.n2608 0.001
R10997 VP.n9306 VP.n9305 0.001
R10998 VP.n2246 VP.n2245 0.001
R10999 VP.n2333 VP.n2332 0.001
R11000 VP.n3197 VP.n3196 0.001
R11001 VP.n3360 VP.n3359 0.001
R11002 VP.n4088 VP.n4087 0.001
R11003 VP.n4281 VP.n4280 0.001
R11004 VP.n4971 VP.n4970 0.001
R11005 VP.n5187 VP.n5186 0.001
R11006 VP.n5808 VP.n5807 0.001
R11007 VP.n6051 VP.n6050 0.001
R11008 VP.n6652 VP.n6651 0.001
R11009 VP.n6915 VP.n6914 0.001
R11010 VP.n7464 VP.n7463 0.001
R11011 VP.n7754 VP.n7753 0.001
R11012 VP.n8280 VP.n8279 0.001
R11013 VP.n8593 VP.n8592 0.001
R11014 VP.n9077 VP.n9076 0.001
R11015 VP.n9389 VP.n9388 0.001
R11016 VP.n9840 VP.n9839 0.001
R11017 VP.n10734 VP.n10733 0.001
R11018 VP.n10459 VP.n10458 0.001
R11019 VP.n10424 VP.n10423 0.001
R11020 VP.n10054 VP.n10053 0.001
R11021 VP.n10984 VP.n10983 0.001
R11022 VP.n10621 VP.n10620 0.001
R11023 VP.n9258 VP.n9257 0.001
R11024 VP.n9619 VP.n9618 0.001
R11025 VP.n10014 VP.n10013 0.001
R11026 VP.n10925 VP.n10924 0.001
R11027 VP.n10583 VP.n10582 0.001
R11028 VP.n8757 VP.n8756 0.001
R11029 VP.n9037 VP.n9036 0.001
R11030 VP.n9569 VP.n9568 0.001
R11031 VP.n9802 VP.n9801 0.001
R11032 VP.n10906 VP.n10905 0.001
R11033 VP.n10401 VP.n10400 0.001
R11034 VP.n8200 VP.n8199 0.001
R11035 VP.n7592 VP.n7591 0.001
R11036 VP.n7954 VP.n7953 0.001
R11037 VP.n8420 VP.n8419 0.001
R11038 VP.n8730 VP.n8729 0.001
R11039 VP.n9220 VP.n9219 0.001
R11040 VP.n9536 VP.n9535 0.001
R11041 VP.n9977 VP.n9976 0.001
R11042 VP.n10874 VP.n10873 0.001
R11043 VP.n10548 VP.n10547 0.001
R11044 VP.n7034 VP.n7033 0.001
R11045 VP.n7342 VP.n7341 0.001
R11046 VP.n7877 VP.n7876 0.001
R11047 VP.n8163 VP.n8162 0.001
R11048 VP.n8713 VP.n8712 0.001
R11049 VP.n9007 VP.n9006 0.001
R11050 VP.n9517 VP.n9516 0.001
R11051 VP.n9780 VP.n9779 0.001
R11052 VP.n10855 VP.n10854 0.001
R11053 VP.n10384 VP.n10383 0.001
R11054 VP.n6490 VP.n6489 0.001
R11055 VP.n5889 VP.n5888 0.001
R11056 VP.n6267 VP.n6266 0.001
R11057 VP.n6742 VP.n6741 0.001
R11058 VP.n7007 VP.n7006 0.001
R11059 VP.n7554 VP.n7553 0.001
R11060 VP.n7845 VP.n7844 0.001
R11061 VP.n8371 VP.n8370 0.001
R11062 VP.n8682 VP.n8681 0.001
R11063 VP.n9170 VP.n9169 0.001
R11064 VP.n9485 VP.n9484 0.001
R11065 VP.n9929 VP.n9928 0.001
R11066 VP.n10823 VP.n10822 0.001
R11067 VP.n10513 VP.n10512 0.001
R11068 VP.n5255 VP.n5254 0.001
R11069 VP.n5604 VP.n5603 0.001
R11070 VP.n6126 VP.n6125 0.001
R11071 VP.n6453 VP.n6452 0.001
R11072 VP.n6989 VP.n6988 0.001
R11073 VP.n7312 VP.n7311 0.001
R11074 VP.n7827 VP.n7826 0.001
R11075 VP.n8140 VP.n8139 0.001
R11076 VP.n8665 VP.n8664 0.001
R11077 VP.n8984 VP.n8983 0.001
R11078 VP.n9466 VP.n9465 0.001
R11079 VP.n9758 VP.n9757 0.001
R11080 VP.n10804 VP.n10803 0.001
R11081 VP.n10367 VP.n10366 0.001
R11082 VP.n4716 VP.n4715 0.001
R11083 VP.n4119 VP.n4118 0.001
R11084 VP.n4516 VP.n4515 0.001
R11085 VP.n5014 VP.n5013 0.001
R11086 VP.n5228 VP.n5227 0.001
R11087 VP.n5851 VP.n5850 0.001
R11088 VP.n6094 VP.n6093 0.001
R11089 VP.n6693 VP.n6692 0.001
R11090 VP.n6958 VP.n6957 0.001
R11091 VP.n7505 VP.n7504 0.001
R11092 VP.n7796 VP.n7795 0.001
R11093 VP.n8322 VP.n8321 0.001
R11094 VP.n8634 VP.n8633 0.001
R11095 VP.n9120 VP.n9119 0.001
R11096 VP.n9434 VP.n9433 0.001
R11097 VP.n9881 VP.n9880 0.001
R11098 VP.n10772 VP.n10771 0.001
R11099 VP.n10478 VP.n10477 0.001
R11100 VP.n868 VP.n867 0.001
R11101 VP.n1410 VP.n1409 0.001
R11102 VP.n1854 VP.n1853 0.001
R11103 VP.n2622 VP.n2621 0.001
R11104 VP.n2807 VP.n2806 0.001
R11105 VP.n3333 VP.n3332 0.001
R11106 VP.n3747 VP.n3746 0.001
R11107 VP.n4254 VP.n4253 0.001
R11108 VP.n4653 VP.n4652 0.001
R11109 VP.n5160 VP.n5159 0.001
R11110 VP.n5548 VP.n5547 0.001
R11111 VP.n6024 VP.n6023 0.001
R11112 VP.n6404 VP.n6403 0.001
R11113 VP.n6888 VP.n6887 0.001
R11114 VP.n7263 VP.n7262 0.001
R11115 VP.n7727 VP.n7726 0.001
R11116 VP.n8091 VP.n8090 0.001
R11117 VP.n8566 VP.n8565 0.001
R11118 VP.n8935 VP.n8934 0.001
R11119 VP.n9360 VP.n9359 0.001
R11120 VP.n9736 VP.n9735 0.001
R11121 VP.n10705 VP.n10704 0.001
R11122 VP.n10139 VP.n10138 0.001
R11123 VP.n10690 VP.n10689 0.001
R11124 VP.n9703 VP.n9702 0.001
R11125 VP.n9338 VP.n9337 0.001
R11126 VP.n8912 VP.n8911 0.001
R11127 VP.n8545 VP.n8544 0.001
R11128 VP.n8068 VP.n8067 0.001
R11129 VP.n7706 VP.n7705 0.001
R11130 VP.n7240 VP.n7239 0.001
R11131 VP.n6867 VP.n6866 0.001
R11132 VP.n6381 VP.n6380 0.001
R11133 VP.n6003 VP.n6002 0.001
R11134 VP.n5525 VP.n5524 0.001
R11135 VP.n5139 VP.n5138 0.001
R11136 VP.n4630 VP.n4629 0.001
R11137 VP.n4233 VP.n4232 0.001
R11138 VP.n3724 VP.n3723 0.001
R11139 VP.n3312 VP.n3311 0.001
R11140 VP.n2784 VP.n2783 0.001
R11141 VP.n2647 VP.n2646 0.001
R11142 VP.n1824 VP.n1823 0.001
R11143 VP.n1386 VP.n1385 0.001
R11144 VP.n840 VP.n839 0.001
R11145 VP.n297 VP.n296 0.001
R11146 VP.n268 VP.n267 0.001
R11147 VP.n371 VP.n370 0.001
R11148 VP.n907 VP.n906 0.001
R11149 VP.n1340 VP.n1339 0.001
R11150 VP.n418 VP.n417 0.001
R11151 VP.n957 VP.n956 0.001
R11152 VP.n1469 VP.n1468 0.001
R11153 VP.n1894 VP.n1893 0.001
R11154 VP.n2316 VP.n2315 0.001
R11155 VP.n465 VP.n464 0.001
R11156 VP.n1007 VP.n1006 0.001
R11157 VP.n1507 VP.n1506 0.001
R11158 VP.n1946 VP.n1945 0.001
R11159 VP.n2569 VP.n2568 0.001
R11160 VP.n2875 VP.n2874 0.001
R11161 VP.n3266 VP.n3265 0.001
R11162 VP.n512 VP.n511 0.001
R11163 VP.n1057 VP.n1056 0.001
R11164 VP.n1545 VP.n1544 0.001
R11165 VP.n1998 VP.n1997 0.001
R11166 VP.n2531 VP.n2530 0.001
R11167 VP.n2927 VP.n2926 0.001
R11168 VP.n3447 VP.n3446 0.001
R11169 VP.n3820 VP.n3819 0.001
R11170 VP.n4187 VP.n4186 0.001
R11171 VP.n559 VP.n558 0.001
R11172 VP.n1107 VP.n1106 0.001
R11173 VP.n1583 VP.n1582 0.001
R11174 VP.n2050 VP.n2049 0.001
R11175 VP.n2493 VP.n2492 0.001
R11176 VP.n2979 VP.n2978 0.001
R11177 VP.n3485 VP.n3484 0.001
R11178 VP.n3872 VP.n3871 0.001
R11179 VP.n4364 VP.n4363 0.001
R11180 VP.n4755 VP.n4754 0.001
R11181 VP.n5093 VP.n5092 0.001
R11182 VP.n606 VP.n605 0.001
R11183 VP.n1157 VP.n1156 0.001
R11184 VP.n1621 VP.n1620 0.001
R11185 VP.n2102 VP.n2101 0.001
R11186 VP.n2461 VP.n2460 0.001
R11187 VP.n3031 VP.n3030 0.001
R11188 VP.n3523 VP.n3522 0.001
R11189 VP.n3924 VP.n3923 0.001
R11190 VP.n4402 VP.n4401 0.001
R11191 VP.n4807 VP.n4806 0.001
R11192 VP.n5324 VP.n5323 0.001
R11193 VP.n5644 VP.n5643 0.001
R11194 VP.n5957 VP.n5956 0.001
R11195 VP.n646 VP.n645 0.001
R11196 VP.n1195 VP.n1194 0.001
R11197 VP.n1653 VP.n1652 0.001
R11198 VP.n2143 VP.n2142 0.001
R11199 VP.n2429 VP.n2428 0.001
R11200 VP.n3072 VP.n3071 0.001
R11201 VP.n3555 VP.n3554 0.001
R11202 VP.n3965 VP.n3964 0.001
R11203 VP.n4434 VP.n4433 0.001
R11204 VP.n4848 VP.n4847 0.001
R11205 VP.n5356 VP.n5355 0.001
R11206 VP.n5685 VP.n5684 0.001
R11207 VP.n6184 VP.n6183 0.001
R11208 VP.n6529 VP.n6528 0.001
R11209 VP.n6821 VP.n6820 0.001
R11210 VP.n676 VP.n675 0.001
R11211 VP.n1235 VP.n1234 0.001
R11212 VP.n1685 VP.n1684 0.001
R11213 VP.n2184 VP.n2183 0.001
R11214 VP.n2397 VP.n2396 0.001
R11215 VP.n3113 VP.n3112 0.001
R11216 VP.n3587 VP.n3586 0.001
R11217 VP.n4006 VP.n4005 0.001
R11218 VP.n4466 VP.n4465 0.001
R11219 VP.n4889 VP.n4888 0.001
R11220 VP.n5388 VP.n5387 0.001
R11221 VP.n5726 VP.n5725 0.001
R11222 VP.n6216 VP.n6215 0.001
R11223 VP.n6570 VP.n6569 0.001
R11224 VP.n7103 VP.n7102 0.001
R11225 VP.n7382 VP.n7381 0.001
R11226 VP.n7660 VP.n7659 0.001
R11227 VP.n275 VP.n274 0.001
R11228 VP.n791 VP.n790 0.001
R11229 VP.n1347 VP.n1346 0.001
R11230 VP.n1777 VP.n1776 0.001
R11231 VP.n2664 VP.n2663 0.001
R11232 VP.n2737 VP.n2736 0.001
R11233 VP.n3273 VP.n3272 0.001
R11234 VP.n3677 VP.n3676 0.001
R11235 VP.n4194 VP.n4193 0.001
R11236 VP.n4586 VP.n4585 0.001
R11237 VP.n5100 VP.n5099 0.001
R11238 VP.n5478 VP.n5477 0.001
R11239 VP.n5964 VP.n5963 0.001
R11240 VP.n6334 VP.n6333 0.001
R11241 VP.n6828 VP.n6827 0.001
R11242 VP.n7193 VP.n7192 0.001
R11243 VP.n7667 VP.n7666 0.001
R11244 VP.n8021 VP.n8020 0.001
R11245 VP.n8506 VP.n8505 0.001
R11246 VP.n8867 VP.n8866 0.001
R11247 VP.n9323 VP.n9322 0.001
R11248 VP.n2225 VP.n2224 0.001
R11249 VP.n2365 VP.n2364 0.001
R11250 VP.n3154 VP.n3153 0.001
R11251 VP.n3619 VP.n3618 0.001
R11252 VP.n4047 VP.n4046 0.001
R11253 VP.n4498 VP.n4497 0.001
R11254 VP.n4930 VP.n4929 0.001
R11255 VP.n5420 VP.n5419 0.001
R11256 VP.n5767 VP.n5766 0.001
R11257 VP.n6248 VP.n6247 0.001
R11258 VP.n6611 VP.n6610 0.001
R11259 VP.n7135 VP.n7134 0.001
R11260 VP.n7423 VP.n7422 0.001
R11261 VP.n7935 VP.n7934 0.001
R11262 VP.n8239 VP.n8238 0.001
R11263 VP.n8499 VP.n8498 0.001
R11264 VP.n708 VP.n707 0.001
R11265 VP.n1276 VP.n1275 0.001
R11266 VP.n1717 VP.n1716 0.001
R11267 VP.n162 VP.n161 0.001
R11268 VP.n10071 VP.n10047 0.001
R11269 VP.n9273 VP.n9251 0.001
R11270 VP.n7607 VP.n7585 0.001
R11271 VP.n5904 VP.n5882 0.001
R11272 VP.n4134 VP.n4112 0.001
R11273 VP.n2263 VP.n2243 0.001
R11274 VP.t8 VP.n10313 0.001
R11275 VP.t8 VP.n10297 0.001
R11276 VP.t8 VP.n10269 0.001
R11277 VP.t8 VP.n10241 0.001
R11278 VP.n10359 VP.t8 0.001
R11279 VP.t8 VP.n10213 0.001
R11280 VP.t8 VP.n10193 0.001
R11281 VP.t8 VP.n10329 0.001
R11282 VP.n8889 VP.n8847 0.001
R11283 VP.n11005 VP.n10977 0.001
R11284 VP.n10642 VP.n10611 0.001
R11285 VP.n9633 VP.n9612 0.001
R11286 VP.n10040 VP.n10007 0.001
R11287 VP.n10946 VP.n10918 0.001
R11288 VP.n10604 VP.n10576 0.001
R11289 VP.n7968 VP.n7947 0.001
R11290 VP.n8446 VP.n8402 0.001
R11291 VP.n8744 VP.n8724 0.001
R11292 VP.n9244 VP.n9201 0.001
R11293 VP.n9551 VP.n9529 0.001
R11294 VP.n10000 VP.n9959 0.001
R11295 VP.n10895 VP.n10867 0.001
R11296 VP.n10569 VP.n10541 0.001
R11297 VP.n6281 VP.n6260 0.001
R11298 VP.n6768 VP.n6724 0.001
R11299 VP.n7021 VP.n7000 0.001
R11300 VP.n7578 VP.n7536 0.001
R11301 VP.n7859 VP.n7838 0.001
R11302 VP.n8395 VP.n8353 0.001
R11303 VP.n8696 VP.n8676 0.001
R11304 VP.n9194 VP.n9151 0.001
R11305 VP.n9500 VP.n9478 0.001
R11306 VP.n9952 VP.n9911 0.001
R11307 VP.n10844 VP.n10816 0.001
R11308 VP.n10534 VP.n10506 0.001
R11309 VP.n4530 VP.n4510 0.001
R11310 VP.n5040 VP.n4995 0.001
R11311 VP.n5242 VP.n5222 0.001
R11312 VP.n5875 VP.n5832 0.001
R11313 VP.n6108 VP.n6087 0.001
R11314 VP.n6717 VP.n6675 0.001
R11315 VP.n6972 VP.n6951 0.001
R11316 VP.n7529 VP.n7487 0.001
R11317 VP.n7810 VP.n7789 0.001
R11318 VP.n8346 VP.n8304 0.001
R11319 VP.n8648 VP.n8628 0.001
R11320 VP.n9144 VP.n9101 0.001
R11321 VP.n9449 VP.n9427 0.001
R11322 VP.n9904 VP.n9863 0.001
R11323 VP.n10793 VP.n10765 0.001
R11324 VP.n10499 VP.n10471 0.001
R11325 VP.n2338 VP.n2330 0.001
R11326 VP.n3213 VP.n3194 0.001
R11327 VP.n3364 VP.n3357 0.001
R11328 VP.n4105 VP.n4085 0.001
R11329 VP.n4285 VP.n4278 0.001
R11330 VP.n4988 VP.n4968 0.001
R11331 VP.n5191 VP.n5184 0.001
R11332 VP.n5825 VP.n5805 0.001
R11333 VP.n6056 VP.n6048 0.001
R11334 VP.n6668 VP.n6649 0.001
R11335 VP.n6920 VP.n6912 0.001
R11336 VP.n7480 VP.n7461 0.001
R11337 VP.n7758 VP.n7751 0.001
R11338 VP.n8297 VP.n8277 0.001
R11339 VP.n8597 VP.n8590 0.001
R11340 VP.n9094 VP.n9074 0.001
R11341 VP.n9394 VP.n9386 0.001
R11342 VP.n9856 VP.n9837 0.001
R11343 VP.n10739 VP.n10731 0.001
R11344 VP.n10464 VP.n10456 0.001
R11345 VP.n759 VP.n758 0.001
R11346 VP.n1748 VP.n1747 0.001
R11347 VP.n924 VP.n904 0.001
R11348 VP.n392 VP.n368 0.001
R11349 VP.n2709 VP.n2708 0.001
R11350 VP.n1913 VP.n1891 0.001
R11351 VP.n1480 VP.n1466 0.001
R11352 VP.n974 VP.n954 0.001
R11353 VP.n439 VP.n415 0.001
R11354 VP.n3649 VP.n3648 0.001
R11355 VP.n2894 VP.n2872 0.001
R11356 VP.n2580 VP.n2566 0.001
R11357 VP.n1965 VP.n1943 0.001
R11358 VP.n1518 VP.n1504 0.001
R11359 VP.n1024 VP.n1004 0.001
R11360 VP.n486 VP.n462 0.001
R11361 VP.n4555 VP.n4554 0.001
R11362 VP.n3839 VP.n3817 0.001
R11363 VP.n3458 VP.n3444 0.001
R11364 VP.n2946 VP.n2924 0.001
R11365 VP.n2542 VP.n2528 0.001
R11366 VP.n2017 VP.n1995 0.001
R11367 VP.n1556 VP.n1542 0.001
R11368 VP.n1074 VP.n1054 0.001
R11369 VP.n533 VP.n509 0.001
R11370 VP.n5450 VP.n5449 0.001
R11371 VP.n4774 VP.n4752 0.001
R11372 VP.n4375 VP.n4361 0.001
R11373 VP.n3891 VP.n3869 0.001
R11374 VP.n3496 VP.n3482 0.001
R11375 VP.n2998 VP.n2976 0.001
R11376 VP.n2504 VP.n2490 0.001
R11377 VP.n2069 VP.n2047 0.001
R11378 VP.n1594 VP.n1580 0.001
R11379 VP.n1124 VP.n1104 0.001
R11380 VP.n580 VP.n556 0.001
R11381 VP.n6306 VP.n6305 0.001
R11382 VP.n5652 VP.n5641 0.001
R11383 VP.n5329 VP.n5321 0.001
R11384 VP.n4815 VP.n4804 0.001
R11385 VP.n4407 VP.n4399 0.001
R11386 VP.n3932 VP.n3921 0.001
R11387 VP.n3528 VP.n3520 0.001
R11388 VP.n3039 VP.n3028 0.001
R11389 VP.n2466 VP.n2458 0.001
R11390 VP.n2110 VP.n2099 0.001
R11391 VP.n1626 VP.n1618 0.001
R11392 VP.n1162 VP.n1154 0.001
R11393 VP.n620 VP.n603 0.001
R11394 VP.n7165 VP.n7164 0.001
R11395 VP.n6537 VP.n6526 0.001
R11396 VP.n6189 VP.n6181 0.001
R11397 VP.n5693 VP.n5682 0.001
R11398 VP.n5361 VP.n5353 0.001
R11399 VP.n4856 VP.n4845 0.001
R11400 VP.n4439 VP.n4431 0.001
R11401 VP.n3973 VP.n3962 0.001
R11402 VP.n3560 VP.n3552 0.001
R11403 VP.n3080 VP.n3069 0.001
R11404 VP.n2434 VP.n2426 0.001
R11405 VP.n2151 VP.n2140 0.001
R11406 VP.n1658 VP.n1650 0.001
R11407 VP.n1202 VP.n1192 0.001
R11408 VP.n650 VP.n643 0.001
R11409 VP.n7993 VP.n7992 0.001
R11410 VP.n7390 VP.n7379 0.001
R11411 VP.n7108 VP.n7100 0.001
R11412 VP.n6578 VP.n6567 0.001
R11413 VP.n6221 VP.n6213 0.001
R11414 VP.n5734 VP.n5723 0.001
R11415 VP.n5393 VP.n5385 0.001
R11416 VP.n4897 VP.n4886 0.001
R11417 VP.n4471 VP.n4463 0.001
R11418 VP.n4014 VP.n4003 0.001
R11419 VP.n3592 VP.n3584 0.001
R11420 VP.n3121 VP.n3110 0.001
R11421 VP.n2402 VP.n2394 0.001
R11422 VP.n2192 VP.n2181 0.001
R11423 VP.n1690 VP.n1682 0.001
R11424 VP.n1243 VP.n1232 0.001
R11425 VP.n682 VP.n673 0.001
R11426 VP.n8524 VP.n8500 0.001
R11427 VP.n8045 VP.n8013 0.001
R11428 VP.n7685 VP.n7661 0.001
R11429 VP.n7217 VP.n7185 0.001
R11430 VP.n6846 VP.n6822 0.001
R11431 VP.n6358 VP.n6326 0.001
R11432 VP.n5982 VP.n5958 0.001
R11433 VP.n5502 VP.n5470 0.001
R11434 VP.n5118 VP.n5094 0.001
R11435 VP.n4610 VP.n4575 0.001
R11436 VP.n4212 VP.n4188 0.001
R11437 VP.n3701 VP.n3669 0.001
R11438 VP.n3291 VP.n3267 0.001
R11439 VP.n2761 VP.n2729 0.001
R11440 VP.n2682 VP.n2658 0.001
R11441 VP.n1801 VP.n1768 0.001
R11442 VP.n1365 VP.n1341 0.001
R11443 VP.n815 VP.n779 0.001
R11444 VP.n287 VP.n269 0.001
R11445 VP.n8827 VP.n8826 0.001
R11446 VP.n8247 VP.n8236 0.001
R11447 VP.n7940 VP.n7932 0.001
R11448 VP.n7431 VP.n7420 0.001
R11449 VP.n7140 VP.n7132 0.001
R11450 VP.n6619 VP.n6608 0.001
R11451 VP.n6253 VP.n6245 0.001
R11452 VP.n5775 VP.n5764 0.001
R11453 VP.n5425 VP.n5417 0.001
R11454 VP.n4938 VP.n4927 0.001
R11455 VP.n4503 VP.n4495 0.001
R11456 VP.n4055 VP.n4044 0.001
R11457 VP.n3624 VP.n3616 0.001
R11458 VP.n3162 VP.n3151 0.001
R11459 VP.n2370 VP.n2362 0.001
R11460 VP.n2233 VP.n2222 0.001
R11461 VP.n1723 VP.n1714 0.001
R11462 VP.n1284 VP.n1273 0.001
R11463 VP.n722 VP.n705 0.001
R11464 VP.n10348 VP.n10347 0.001
R11465 VP.n10968 VP.n10967 0.001
R11466 VP.n9593 VP.n9592 0.001
R11467 VP.n8789 VP.n8788 0.001
R11468 VP.n7902 VP.n7901 0.001
R11469 VP.n7066 VP.n7065 0.001
R11470 VP.n6151 VP.n6150 0.001
R11471 VP.n5287 VP.n5286 0.001
R11472 VP.n4331 VP.n4330 0.001
R11473 VP.n3410 VP.n3409 0.001
R11474 VP.n2605 VP.n2604 0.001
R11475 VP.t108 VP.n2847 0.001
R11476 VP.n2841 VP.n2840 0.001
R11477 VP.t72 VP.n3397 0.001
R11478 VP.n3391 VP.n3390 0.001
R11479 VP.t76 VP.n3792 0.001
R11480 VP.n3786 VP.n3785 0.001
R11481 VP.t140 VP.n4316 0.001
R11482 VP.n4310 VP.n4309 0.001
R11483 VP.t169 VP.n4691 0.001
R11484 VP.n4685 VP.n4684 0.001
R11485 VP.t119 VP.n5221 0.001
R11486 VP.n5215 VP.n5214 0.001
R11487 VP.t26 VP.n5586 0.001
R11488 VP.n5580 VP.n5579 0.001
R11489 VP.t24 VP.n6086 0.001
R11490 VP.n6080 VP.n6079 0.001
R11491 VP.t159 VP.n6442 0.001
R11492 VP.n6436 VP.n6435 0.001
R11493 VP.t195 VP.n6950 0.001
R11494 VP.n6944 VP.n6943 0.001
R11495 VP.t134 VP.n7301 0.001
R11496 VP.n7295 VP.n7294 0.001
R11497 VP.t111 VP.n7788 0.001
R11498 VP.n7782 VP.n7781 0.001
R11499 VP.t18 VP.n8129 0.001
R11500 VP.n8123 VP.n8122 0.001
R11501 VP.t28 VP.n8627 0.001
R11502 VP.n8621 VP.n8620 0.001
R11503 VP.t207 VP.n8973 0.001
R11504 VP.n8967 VP.n8966 0.001
R11505 VP.t143 VP.n9426 0.001
R11506 VP.n9420 VP.n9419 0.001
R11507 VP.t16 VP.n10764 0.001
R11508 VP.n10758 VP.n10757 0.001
R11509 VP.t6 VP.n10170 0.001
R11510 VP.n10164 VP.n10163 0.001
R11511 VP.t34 VP.n1447 0.001
R11512 VP.t53 VP.n2266 0.001
R11513 VP.t53 VP.n2269 0.001
R11514 VP.t91 VP.n2344 0.001
R11515 VP.t91 VP.n2341 0.001
R11516 VP.n2341 VP.n2338 0.001
R11517 VP.t108 VP.n3216 0.001
R11518 VP.t108 VP.n3219 0.001
R11519 VP.t72 VP.n3370 0.001
R11520 VP.t72 VP.n3367 0.001
R11521 VP.n3367 VP.n3364 0.001
R11522 VP.t76 VP.n4108 0.001
R11523 VP.t76 VP.n4111 0.001
R11524 VP.t140 VP.n4291 0.001
R11525 VP.t140 VP.n4288 0.001
R11526 VP.n4288 VP.n4285 0.001
R11527 VP.t169 VP.n4991 0.001
R11528 VP.t169 VP.n4994 0.001
R11529 VP.t119 VP.n5197 0.001
R11530 VP.t119 VP.n5194 0.001
R11531 VP.n5194 VP.n5191 0.001
R11532 VP.t26 VP.n5828 0.001
R11533 VP.t26 VP.n5831 0.001
R11534 VP.t24 VP.n6062 0.001
R11535 VP.t24 VP.n6059 0.001
R11536 VP.n6059 VP.n6056 0.001
R11537 VP.t159 VP.n6671 0.001
R11538 VP.t159 VP.n6674 0.001
R11539 VP.t195 VP.n6926 0.001
R11540 VP.t195 VP.n6923 0.001
R11541 VP.n6923 VP.n6920 0.001
R11542 VP.t134 VP.n7483 0.001
R11543 VP.t134 VP.n7486 0.001
R11544 VP.t111 VP.n7764 0.001
R11545 VP.t111 VP.n7761 0.001
R11546 VP.n7761 VP.n7758 0.001
R11547 VP.t18 VP.n8300 0.001
R11548 VP.t18 VP.n8303 0.001
R11549 VP.t28 VP.n8603 0.001
R11550 VP.t28 VP.n8600 0.001
R11551 VP.n8600 VP.n8597 0.001
R11552 VP.t207 VP.n9097 0.001
R11553 VP.t207 VP.n9100 0.001
R11554 VP.t143 VP.n9400 0.001
R11555 VP.t143 VP.n9397 0.001
R11556 VP.n9397 VP.n9394 0.001
R11557 VP.t126 VP.n9859 0.001
R11558 VP.t126 VP.n9862 0.001
R11559 VP.t16 VP.n10745 0.001
R11560 VP.t16 VP.n10742 0.001
R11561 VP.n10742 VP.n10739 0.001
R11562 VP.t6 VP.n10467 0.001
R11563 VP.t6 VP.n10470 0.001
R11564 VP.t6 VP.n10435 0.001
R11565 VP.t6 VP.n10432 0.001
R11566 VP.n10432 VP.n10429 0.001
R11567 VP.t16 VP.n10975 0.001
R11568 VP.t16 VP.n10972 0.001
R11569 VP.n10972 VP.n10970 0.001
R11570 VP.t143 VP.n9610 0.001
R11571 VP.t143 VP.n9607 0.001
R11572 VP.n9607 VP.n9605 0.001
R11573 VP.t126 VP.n10074 0.001
R11574 VP.t126 VP.n10077 0.001
R11575 VP.t16 VP.n11008 0.001
R11576 VP.t16 VP.n11011 0.001
R11577 VP.t6 VP.n10645 0.001
R11578 VP.t6 VP.n10648 0.001
R11579 VP.t28 VP.n8804 0.001
R11580 VP.t28 VP.n8801 0.001
R11581 VP.n8801 VP.n8799 0.001
R11582 VP.t207 VP.n9276 0.001
R11583 VP.t207 VP.n9279 0.001
R11584 VP.t143 VP.n9636 0.001
R11585 VP.t143 VP.n9639 0.001
R11586 VP.t126 VP.n10043 0.001
R11587 VP.t126 VP.n10046 0.001
R11588 VP.t16 VP.n10952 0.001
R11589 VP.t16 VP.n10949 0.001
R11590 VP.n10949 VP.n10946 0.001
R11591 VP.t6 VP.n10607 0.001
R11592 VP.t6 VP.n10610 0.001
R11593 VP.t28 VP.n8776 0.001
R11594 VP.t28 VP.n8773 0.001
R11595 VP.n8773 VP.n8770 0.001
R11596 VP.t207 VP.n9049 0.001
R11597 VP.t207 VP.n9046 0.001
R11598 VP.n9046 VP.n9043 0.001
R11599 VP.t143 VP.n9580 0.001
R11600 VP.t143 VP.n9577 0.001
R11601 VP.n9577 VP.n9574 0.001
R11602 VP.t126 VP.n9813 0.001
R11603 VP.t126 VP.n9810 0.001
R11604 VP.n9810 VP.n9807 0.001
R11605 VP.t16 VP.n10917 0.001
R11606 VP.t16 VP.n10914 0.001
R11607 VP.n10914 VP.n10911 0.001
R11608 VP.t6 VP.n10409 0.001
R11609 VP.t6 VP.n10406 0.001
R11610 VP.n10406 VP.n10403 0.001
R11611 VP.t18 VP.n8211 0.001
R11612 VP.t18 VP.n8208 0.001
R11613 VP.n8208 VP.n8205 0.001
R11614 VP.t111 VP.n7913 0.001
R11615 VP.t111 VP.n7910 0.001
R11616 VP.n7910 VP.n7908 0.001
R11617 VP.t195 VP.n7081 0.001
R11618 VP.t195 VP.n7078 0.001
R11619 VP.n7078 VP.n7076 0.001
R11620 VP.t134 VP.n7610 0.001
R11621 VP.t134 VP.n7613 0.001
R11622 VP.t111 VP.n7971 0.001
R11623 VP.t111 VP.n7974 0.001
R11624 VP.t18 VP.n8449 0.001
R11625 VP.t18 VP.n8452 0.001
R11626 VP.t28 VP.n8750 0.001
R11627 VP.t28 VP.n8747 0.001
R11628 VP.n8747 VP.n8744 0.001
R11629 VP.t207 VP.n9247 0.001
R11630 VP.t207 VP.n9250 0.001
R11631 VP.t143 VP.n9557 0.001
R11632 VP.t143 VP.n9554 0.001
R11633 VP.n9554 VP.n9551 0.001
R11634 VP.t126 VP.n10003 0.001
R11635 VP.t126 VP.n10006 0.001
R11636 VP.t16 VP.n10901 0.001
R11637 VP.t16 VP.n10898 0.001
R11638 VP.n10898 VP.n10895 0.001
R11639 VP.t6 VP.n10572 0.001
R11640 VP.t6 VP.n10575 0.001
R11641 VP.t195 VP.n7053 0.001
R11642 VP.t195 VP.n7050 0.001
R11643 VP.n7050 VP.n7047 0.001
R11644 VP.t134 VP.n7354 0.001
R11645 VP.t134 VP.n7351 0.001
R11646 VP.n7351 VP.n7348 0.001
R11647 VP.t111 VP.n7887 0.001
R11648 VP.t111 VP.n7884 0.001
R11649 VP.n7884 VP.n7881 0.001
R11650 VP.t18 VP.n8175 0.001
R11651 VP.t18 VP.n8172 0.001
R11652 VP.n8172 VP.n8169 0.001
R11653 VP.t28 VP.n8723 0.001
R11654 VP.t28 VP.n8720 0.001
R11655 VP.n8720 VP.n8717 0.001
R11656 VP.t207 VP.n9019 0.001
R11657 VP.t207 VP.n9016 0.001
R11658 VP.n9016 VP.n9013 0.001
R11659 VP.t143 VP.n9528 0.001
R11660 VP.t143 VP.n9525 0.001
R11661 VP.n9525 VP.n9522 0.001
R11662 VP.t126 VP.n9791 0.001
R11663 VP.t126 VP.n9788 0.001
R11664 VP.n9788 VP.n9785 0.001
R11665 VP.t16 VP.n10866 0.001
R11666 VP.t16 VP.n10863 0.001
R11667 VP.n10863 VP.n10860 0.001
R11668 VP.t6 VP.n10392 0.001
R11669 VP.t6 VP.n10389 0.001
R11670 VP.n10389 VP.n10386 0.001
R11671 VP.t159 VP.n6501 0.001
R11672 VP.t159 VP.n6498 0.001
R11673 VP.n6498 VP.n6495 0.001
R11674 VP.t24 VP.n6162 0.001
R11675 VP.t24 VP.n6159 0.001
R11676 VP.n6159 VP.n6157 0.001
R11677 VP.t119 VP.n5302 0.001
R11678 VP.t119 VP.n5299 0.001
R11679 VP.n5299 VP.n5297 0.001
R11680 VP.t26 VP.n5907 0.001
R11681 VP.t26 VP.n5910 0.001
R11682 VP.t24 VP.n6284 0.001
R11683 VP.t24 VP.n6287 0.001
R11684 VP.t159 VP.n6771 0.001
R11685 VP.t159 VP.n6774 0.001
R11686 VP.t195 VP.n7027 0.001
R11687 VP.t195 VP.n7024 0.001
R11688 VP.n7024 VP.n7021 0.001
R11689 VP.t134 VP.n7581 0.001
R11690 VP.t134 VP.n7584 0.001
R11691 VP.t111 VP.n7865 0.001
R11692 VP.t111 VP.n7862 0.001
R11693 VP.n7862 VP.n7859 0.001
R11694 VP.t18 VP.n8398 0.001
R11695 VP.t18 VP.n8401 0.001
R11696 VP.t28 VP.n8702 0.001
R11697 VP.t28 VP.n8699 0.001
R11698 VP.n8699 VP.n8696 0.001
R11699 VP.t207 VP.n9197 0.001
R11700 VP.t207 VP.n9200 0.001
R11701 VP.t143 VP.n9506 0.001
R11702 VP.t143 VP.n9503 0.001
R11703 VP.n9503 VP.n9500 0.001
R11704 VP.t126 VP.n9955 0.001
R11705 VP.t126 VP.n9958 0.001
R11706 VP.t16 VP.n10850 0.001
R11707 VP.t16 VP.n10847 0.001
R11708 VP.n10847 VP.n10844 0.001
R11709 VP.t6 VP.n10537 0.001
R11710 VP.t6 VP.n10540 0.001
R11711 VP.t119 VP.n5274 0.001
R11712 VP.t119 VP.n5271 0.001
R11713 VP.n5271 VP.n5268 0.001
R11714 VP.t26 VP.n5616 0.001
R11715 VP.t26 VP.n5613 0.001
R11716 VP.n5613 VP.n5610 0.001
R11717 VP.t24 VP.n6136 0.001
R11718 VP.t24 VP.n6133 0.001
R11719 VP.n6133 VP.n6130 0.001
R11720 VP.t159 VP.n6465 0.001
R11721 VP.t159 VP.n6462 0.001
R11722 VP.n6462 VP.n6459 0.001
R11723 VP.t195 VP.n6999 0.001
R11724 VP.t195 VP.n6996 0.001
R11725 VP.n6996 VP.n6993 0.001
R11726 VP.t134 VP.n7324 0.001
R11727 VP.t134 VP.n7321 0.001
R11728 VP.n7321 VP.n7318 0.001
R11729 VP.t111 VP.n7837 0.001
R11730 VP.t111 VP.n7834 0.001
R11731 VP.n7834 VP.n7831 0.001
R11732 VP.t18 VP.n8152 0.001
R11733 VP.t18 VP.n8149 0.001
R11734 VP.n8149 VP.n8146 0.001
R11735 VP.t28 VP.n8675 0.001
R11736 VP.t28 VP.n8672 0.001
R11737 VP.n8672 VP.n8669 0.001
R11738 VP.t207 VP.n8996 0.001
R11739 VP.t207 VP.n8993 0.001
R11740 VP.n8993 VP.n8990 0.001
R11741 VP.t143 VP.n9477 0.001
R11742 VP.t143 VP.n9474 0.001
R11743 VP.n9474 VP.n9471 0.001
R11744 VP.t126 VP.n9769 0.001
R11745 VP.t126 VP.n9766 0.001
R11746 VP.n9766 VP.n9763 0.001
R11747 VP.t16 VP.n10815 0.001
R11748 VP.t16 VP.n10812 0.001
R11749 VP.n10812 VP.n10809 0.001
R11750 VP.t6 VP.n10375 0.001
R11751 VP.t6 VP.n10372 0.001
R11752 VP.n10372 VP.n10369 0.001
R11753 VP.t169 VP.n4727 0.001
R11754 VP.t169 VP.n4724 0.001
R11755 VP.n4724 VP.n4721 0.001
R11756 VP.t140 VP.n4342 0.001
R11757 VP.t140 VP.n4339 0.001
R11758 VP.n4339 VP.n4337 0.001
R11759 VP.t72 VP.n3425 0.001
R11760 VP.t72 VP.n3422 0.001
R11761 VP.n3422 VP.n3420 0.001
R11762 VP.t76 VP.n4137 0.001
R11763 VP.t76 VP.n4140 0.001
R11764 VP.t140 VP.n4533 0.001
R11765 VP.t140 VP.n4536 0.001
R11766 VP.t169 VP.n5043 0.001
R11767 VP.t169 VP.n5046 0.001
R11768 VP.t119 VP.n5248 0.001
R11769 VP.t119 VP.n5245 0.001
R11770 VP.n5245 VP.n5242 0.001
R11771 VP.t26 VP.n5878 0.001
R11772 VP.t26 VP.n5881 0.001
R11773 VP.t24 VP.n6114 0.001
R11774 VP.t24 VP.n6111 0.001
R11775 VP.n6111 VP.n6108 0.001
R11776 VP.t159 VP.n6720 0.001
R11777 VP.t159 VP.n6723 0.001
R11778 VP.t195 VP.n6978 0.001
R11779 VP.t195 VP.n6975 0.001
R11780 VP.n6975 VP.n6972 0.001
R11781 VP.t134 VP.n7532 0.001
R11782 VP.t134 VP.n7535 0.001
R11783 VP.t111 VP.n7816 0.001
R11784 VP.t111 VP.n7813 0.001
R11785 VP.n7813 VP.n7810 0.001
R11786 VP.t18 VP.n8349 0.001
R11787 VP.t18 VP.n8352 0.001
R11788 VP.t28 VP.n8654 0.001
R11789 VP.t28 VP.n8651 0.001
R11790 VP.n8651 VP.n8648 0.001
R11791 VP.t207 VP.n9147 0.001
R11792 VP.t207 VP.n9150 0.001
R11793 VP.t143 VP.n9455 0.001
R11794 VP.t143 VP.n9452 0.001
R11795 VP.n9452 VP.n9449 0.001
R11796 VP.t126 VP.n9907 0.001
R11797 VP.t126 VP.n9910 0.001
R11798 VP.t16 VP.n10799 0.001
R11799 VP.t16 VP.n10796 0.001
R11800 VP.n10796 VP.n10793 0.001
R11801 VP.t6 VP.n10502 0.001
R11802 VP.t6 VP.n10505 0.001
R11803 VP.t57 VP.n350 0.001
R11804 VP.t57 VP.n347 0.001
R11805 VP.n347 VP.n345 0.001
R11806 VP.t49 VP.n879 0.001
R11807 VP.t49 VP.n876 0.001
R11808 VP.n876 VP.n873 0.001
R11809 VP.t34 VP.n1420 0.001
R11810 VP.t34 VP.n1417 0.001
R11811 VP.n1417 VP.n1414 0.001
R11812 VP.t53 VP.n1866 0.001
R11813 VP.t53 VP.n1863 0.001
R11814 VP.n1863 VP.n1860 0.001
R11815 VP.t91 VP.n2629 0.001
R11816 VP.t91 VP.n2632 0.001
R11817 VP.t108 VP.n2819 0.001
R11818 VP.t108 VP.n2816 0.001
R11819 VP.n2816 VP.n2813 0.001
R11820 VP.t72 VP.n3343 0.001
R11821 VP.t72 VP.n3340 0.001
R11822 VP.n3340 VP.n3337 0.001
R11823 VP.t76 VP.n3759 0.001
R11824 VP.t76 VP.n3756 0.001
R11825 VP.n3756 VP.n3753 0.001
R11826 VP.t140 VP.n4264 0.001
R11827 VP.t140 VP.n4261 0.001
R11828 VP.n4261 VP.n4258 0.001
R11829 VP.t169 VP.n4665 0.001
R11830 VP.t169 VP.n4662 0.001
R11831 VP.n4662 VP.n4659 0.001
R11832 VP.t119 VP.n5170 0.001
R11833 VP.t119 VP.n5167 0.001
R11834 VP.n5167 VP.n5164 0.001
R11835 VP.t26 VP.n5560 0.001
R11836 VP.t26 VP.n5557 0.001
R11837 VP.n5557 VP.n5554 0.001
R11838 VP.t24 VP.n6034 0.001
R11839 VP.t24 VP.n6031 0.001
R11840 VP.n6031 VP.n6028 0.001
R11841 VP.t159 VP.n6416 0.001
R11842 VP.t159 VP.n6413 0.001
R11843 VP.n6413 VP.n6410 0.001
R11844 VP.t195 VP.n6898 0.001
R11845 VP.t195 VP.n6895 0.001
R11846 VP.n6895 VP.n6892 0.001
R11847 VP.t134 VP.n7275 0.001
R11848 VP.t134 VP.n7272 0.001
R11849 VP.n7272 VP.n7269 0.001
R11850 VP.t111 VP.n7737 0.001
R11851 VP.t111 VP.n7734 0.001
R11852 VP.n7734 VP.n7731 0.001
R11853 VP.t18 VP.n8103 0.001
R11854 VP.t18 VP.n8100 0.001
R11855 VP.n8100 VP.n8097 0.001
R11856 VP.t28 VP.n8576 0.001
R11857 VP.t28 VP.n8573 0.001
R11858 VP.n8573 VP.n8570 0.001
R11859 VP.t207 VP.n8947 0.001
R11860 VP.t207 VP.n8944 0.001
R11861 VP.n8944 VP.n8941 0.001
R11862 VP.t143 VP.n9371 0.001
R11863 VP.t143 VP.n9368 0.001
R11864 VP.n9368 VP.n9365 0.001
R11865 VP.t126 VP.n9747 0.001
R11866 VP.t126 VP.n9744 0.001
R11867 VP.n9744 VP.n9741 0.001
R11868 VP.t16 VP.n10716 0.001
R11869 VP.t16 VP.n10713 0.001
R11870 VP.n10713 VP.n10710 0.001
R11871 VP.t6 VP.n10150 0.001
R11872 VP.t6 VP.n10147 0.001
R11873 VP.n10147 VP.n10144 0.001
R11874 VP.n11014 VP.t16 0.001
R11875 VP.n11032 VP.n11017 0.001
R11876 VP.t126 VP.n9725 0.001
R11877 VP.t126 VP.n9722 0.001
R11878 VP.n9722 VP.n9719 0.001
R11879 VP.t143 VP.n9349 0.001
R11880 VP.t143 VP.n9346 0.001
R11881 VP.n9346 VP.n9343 0.001
R11882 VP.t207 VP.n8924 0.001
R11883 VP.t207 VP.n8921 0.001
R11884 VP.n8921 VP.n8918 0.001
R11885 VP.t28 VP.n8555 0.001
R11886 VP.t28 VP.n8552 0.001
R11887 VP.n8552 VP.n8549 0.001
R11888 VP.t18 VP.n8080 0.001
R11889 VP.t18 VP.n8077 0.001
R11890 VP.n8077 VP.n8074 0.001
R11891 VP.t111 VP.n7716 0.001
R11892 VP.t111 VP.n7713 0.001
R11893 VP.n7713 VP.n7710 0.001
R11894 VP.t134 VP.n7252 0.001
R11895 VP.t134 VP.n7249 0.001
R11896 VP.n7249 VP.n7246 0.001
R11897 VP.t195 VP.n6877 0.001
R11898 VP.t195 VP.n6874 0.001
R11899 VP.n6874 VP.n6871 0.001
R11900 VP.t159 VP.n6393 0.001
R11901 VP.t159 VP.n6390 0.001
R11902 VP.n6390 VP.n6387 0.001
R11903 VP.t24 VP.n6013 0.001
R11904 VP.t24 VP.n6010 0.001
R11905 VP.n6010 VP.n6007 0.001
R11906 VP.t26 VP.n5537 0.001
R11907 VP.t26 VP.n5534 0.001
R11908 VP.n5534 VP.n5531 0.001
R11909 VP.t119 VP.n5149 0.001
R11910 VP.t119 VP.n5146 0.001
R11911 VP.n5146 VP.n5143 0.001
R11912 VP.t169 VP.n4642 0.001
R11913 VP.t169 VP.n4639 0.001
R11914 VP.n4639 VP.n4636 0.001
R11915 VP.t140 VP.n4243 0.001
R11916 VP.t140 VP.n4240 0.001
R11917 VP.n4240 VP.n4237 0.001
R11918 VP.t76 VP.n3736 0.001
R11919 VP.t76 VP.n3733 0.001
R11920 VP.n3733 VP.n3730 0.001
R11921 VP.t72 VP.n3322 0.001
R11922 VP.t72 VP.n3319 0.001
R11923 VP.n3319 VP.n3316 0.001
R11924 VP.t108 VP.n2796 0.001
R11925 VP.t108 VP.n2793 0.001
R11926 VP.n2793 VP.n2790 0.001
R11927 VP.t91 VP.n2654 0.001
R11928 VP.t91 VP.n2657 0.001
R11929 VP.t53 VP.n1836 0.001
R11930 VP.t53 VP.n1833 0.001
R11931 VP.n1833 VP.n1830 0.001
R11932 VP.t34 VP.n1396 0.001
R11933 VP.t34 VP.n1393 0.001
R11934 VP.n1393 VP.n1390 0.001
R11935 VP.t49 VP.n850 0.001
R11936 VP.t49 VP.n821 0.001
R11937 VP.t57 VP.n319 0.001
R11938 VP.t57 VP.n316 0.001
R11939 VP.n316 VP.n313 0.001
R11940 VP.n731 VP.t57 0.001
R11941 VP.n758 VP.n734 0.001
R11942 VP.t57 VP.n395 0.001
R11943 VP.t57 VP.n398 0.001
R11944 VP.t49 VP.n927 0.001
R11945 VP.t49 VP.n930 0.001
R11946 VP.n1732 VP.t34 0.001
R11947 VP.n1747 VP.n1735 0.001
R11948 VP.t57 VP.n442 0.001
R11949 VP.t57 VP.n445 0.001
R11950 VP.t49 VP.n977 0.001
R11951 VP.t49 VP.n980 0.001
R11952 VP.t34 VP.n1483 0.001
R11953 VP.t34 VP.n1486 0.001
R11954 VP.t53 VP.n1916 0.001
R11955 VP.t53 VP.n1919 0.001
R11956 VP.n2693 VP.t91 0.001
R11957 VP.n2708 VP.n2696 0.001
R11958 VP.t57 VP.n489 0.001
R11959 VP.t57 VP.n492 0.001
R11960 VP.t49 VP.n1027 0.001
R11961 VP.t49 VP.n1030 0.001
R11962 VP.t34 VP.n1521 0.001
R11963 VP.t34 VP.n1524 0.001
R11964 VP.t53 VP.n1968 0.001
R11965 VP.t53 VP.n1971 0.001
R11966 VP.t91 VP.n2586 0.001
R11967 VP.t91 VP.n2583 0.001
R11968 VP.n2583 VP.n2580 0.001
R11969 VP.t108 VP.n2897 0.001
R11970 VP.t108 VP.n2900 0.001
R11971 VP.n3633 VP.t72 0.001
R11972 VP.n3648 VP.n3636 0.001
R11973 VP.t57 VP.n536 0.001
R11974 VP.t57 VP.n539 0.001
R11975 VP.t49 VP.n1077 0.001
R11976 VP.t49 VP.n1080 0.001
R11977 VP.t34 VP.n1559 0.001
R11978 VP.t34 VP.n1562 0.001
R11979 VP.t53 VP.n2020 0.001
R11980 VP.t53 VP.n2023 0.001
R11981 VP.t91 VP.n2548 0.001
R11982 VP.t91 VP.n2545 0.001
R11983 VP.n2545 VP.n2542 0.001
R11984 VP.t108 VP.n2949 0.001
R11985 VP.t108 VP.n2952 0.001
R11986 VP.t72 VP.n3461 0.001
R11987 VP.t72 VP.n3464 0.001
R11988 VP.t76 VP.n3842 0.001
R11989 VP.t76 VP.n3845 0.001
R11990 VP.n4539 VP.t140 0.001
R11991 VP.n4554 VP.n4542 0.001
R11992 VP.t57 VP.n583 0.001
R11993 VP.t57 VP.n586 0.001
R11994 VP.t49 VP.n1127 0.001
R11995 VP.t49 VP.n1130 0.001
R11996 VP.t34 VP.n1597 0.001
R11997 VP.t34 VP.n1600 0.001
R11998 VP.t53 VP.n2072 0.001
R11999 VP.t53 VP.n2075 0.001
R12000 VP.t91 VP.n2510 0.001
R12001 VP.t91 VP.n2507 0.001
R12002 VP.n2507 VP.n2504 0.001
R12003 VP.t108 VP.n3001 0.001
R12004 VP.t108 VP.n3004 0.001
R12005 VP.t72 VP.n3499 0.001
R12006 VP.t72 VP.n3502 0.001
R12007 VP.t76 VP.n3894 0.001
R12008 VP.t76 VP.n3897 0.001
R12009 VP.t140 VP.n4378 0.001
R12010 VP.t140 VP.n4381 0.001
R12011 VP.t169 VP.n4777 0.001
R12012 VP.t169 VP.n4780 0.001
R12013 VP.n5434 VP.t119 0.001
R12014 VP.n5449 VP.n5437 0.001
R12015 VP.t57 VP.n623 0.001
R12016 VP.t57 VP.n626 0.001
R12017 VP.t49 VP.n1165 0.001
R12018 VP.t49 VP.n1168 0.001
R12019 VP.t34 VP.n1629 0.001
R12020 VP.t34 VP.n1632 0.001
R12021 VP.t53 VP.n2113 0.001
R12022 VP.t53 VP.n2116 0.001
R12023 VP.t91 VP.n2472 0.001
R12024 VP.t91 VP.n2469 0.001
R12025 VP.n2469 VP.n2466 0.001
R12026 VP.t108 VP.n3042 0.001
R12027 VP.t108 VP.n3045 0.001
R12028 VP.t72 VP.n3531 0.001
R12029 VP.t72 VP.n3534 0.001
R12030 VP.t76 VP.n3935 0.001
R12031 VP.t76 VP.n3938 0.001
R12032 VP.t140 VP.n4410 0.001
R12033 VP.t140 VP.n4413 0.001
R12034 VP.t169 VP.n4818 0.001
R12035 VP.t169 VP.n4821 0.001
R12036 VP.t119 VP.n5332 0.001
R12037 VP.t119 VP.n5335 0.001
R12038 VP.t26 VP.n5655 0.001
R12039 VP.t26 VP.n5658 0.001
R12040 VP.n6290 VP.t24 0.001
R12041 VP.n6305 VP.n6293 0.001
R12042 VP.t57 VP.n653 0.001
R12043 VP.t57 VP.n656 0.001
R12044 VP.t49 VP.n1205 0.001
R12045 VP.t49 VP.n1208 0.001
R12046 VP.t34 VP.n1661 0.001
R12047 VP.t34 VP.n1664 0.001
R12048 VP.t53 VP.n2154 0.001
R12049 VP.t53 VP.n2157 0.001
R12050 VP.t91 VP.n2440 0.001
R12051 VP.t91 VP.n2437 0.001
R12052 VP.n2437 VP.n2434 0.001
R12053 VP.t108 VP.n3083 0.001
R12054 VP.t108 VP.n3086 0.001
R12055 VP.t72 VP.n3563 0.001
R12056 VP.t72 VP.n3566 0.001
R12057 VP.t76 VP.n3976 0.001
R12058 VP.t76 VP.n3979 0.001
R12059 VP.t140 VP.n4442 0.001
R12060 VP.t140 VP.n4445 0.001
R12061 VP.t169 VP.n4859 0.001
R12062 VP.t169 VP.n4862 0.001
R12063 VP.t119 VP.n5364 0.001
R12064 VP.t119 VP.n5367 0.001
R12065 VP.t26 VP.n5696 0.001
R12066 VP.t26 VP.n5699 0.001
R12067 VP.t24 VP.n6192 0.001
R12068 VP.t24 VP.n6195 0.001
R12069 VP.t159 VP.n6540 0.001
R12070 VP.t159 VP.n6543 0.001
R12071 VP.n7149 VP.t195 0.001
R12072 VP.n7164 VP.n7152 0.001
R12073 VP.t57 VP.n685 0.001
R12074 VP.t57 VP.n688 0.001
R12075 VP.t49 VP.n1246 0.001
R12076 VP.t49 VP.n1249 0.001
R12077 VP.t34 VP.n1693 0.001
R12078 VP.t34 VP.n1696 0.001
R12079 VP.t53 VP.n2195 0.001
R12080 VP.t53 VP.n2198 0.001
R12081 VP.t91 VP.n2408 0.001
R12082 VP.t91 VP.n2405 0.001
R12083 VP.n2405 VP.n2402 0.001
R12084 VP.t108 VP.n3124 0.001
R12085 VP.t108 VP.n3127 0.001
R12086 VP.t72 VP.n3595 0.001
R12087 VP.t72 VP.n3598 0.001
R12088 VP.t76 VP.n4017 0.001
R12089 VP.t76 VP.n4020 0.001
R12090 VP.t140 VP.n4474 0.001
R12091 VP.t140 VP.n4477 0.001
R12092 VP.t169 VP.n4900 0.001
R12093 VP.t169 VP.n4903 0.001
R12094 VP.t119 VP.n5396 0.001
R12095 VP.t119 VP.n5399 0.001
R12096 VP.t26 VP.n5737 0.001
R12097 VP.t26 VP.n5740 0.001
R12098 VP.t24 VP.n6224 0.001
R12099 VP.t24 VP.n6227 0.001
R12100 VP.t159 VP.n6581 0.001
R12101 VP.t159 VP.n6584 0.001
R12102 VP.t195 VP.n7111 0.001
R12103 VP.t195 VP.n7114 0.001
R12104 VP.t134 VP.n7393 0.001
R12105 VP.t134 VP.n7396 0.001
R12106 VP.n7977 VP.t111 0.001
R12107 VP.n7992 VP.n7980 0.001
R12108 VP.t57 VP.n293 0.001
R12109 VP.t57 VP.n290 0.001
R12110 VP.n290 VP.n287 0.001
R12111 VP.t49 VP.n818 0.001
R12112 VP.n818 VP.n815 0.001
R12113 VP.t34 VP.n1371 0.001
R12114 VP.t34 VP.n1368 0.001
R12115 VP.n1368 VP.n1365 0.001
R12116 VP.t53 VP.n1807 0.001
R12117 VP.t53 VP.n1804 0.001
R12118 VP.n1804 VP.n1801 0.001
R12119 VP.t91 VP.n2685 0.001
R12120 VP.t91 VP.n2688 0.001
R12121 VP.t108 VP.n2767 0.001
R12122 VP.t108 VP.n2764 0.001
R12123 VP.n2764 VP.n2761 0.001
R12124 VP.t72 VP.n3297 0.001
R12125 VP.t72 VP.n3294 0.001
R12126 VP.n3294 VP.n3291 0.001
R12127 VP.t76 VP.n3707 0.001
R12128 VP.t76 VP.n3704 0.001
R12129 VP.n3704 VP.n3701 0.001
R12130 VP.t140 VP.n4218 0.001
R12131 VP.t140 VP.n4215 0.001
R12132 VP.n4215 VP.n4212 0.001
R12133 VP.t169 VP.n4613 0.001
R12134 VP.n4613 VP.n4610 0.001
R12135 VP.t119 VP.n5124 0.001
R12136 VP.t119 VP.n5121 0.001
R12137 VP.n5121 VP.n5118 0.001
R12138 VP.t26 VP.n5508 0.001
R12139 VP.t26 VP.n5505 0.001
R12140 VP.n5505 VP.n5502 0.001
R12141 VP.t24 VP.n5988 0.001
R12142 VP.t24 VP.n5985 0.001
R12143 VP.n5985 VP.n5982 0.001
R12144 VP.t159 VP.n6364 0.001
R12145 VP.t159 VP.n6361 0.001
R12146 VP.n6361 VP.n6358 0.001
R12147 VP.t195 VP.n6852 0.001
R12148 VP.t195 VP.n6849 0.001
R12149 VP.n6849 VP.n6846 0.001
R12150 VP.t134 VP.n7223 0.001
R12151 VP.t134 VP.n7220 0.001
R12152 VP.n7220 VP.n7217 0.001
R12153 VP.t111 VP.n7691 0.001
R12154 VP.t111 VP.n7688 0.001
R12155 VP.n7688 VP.n7685 0.001
R12156 VP.t18 VP.n8051 0.001
R12157 VP.t18 VP.n8048 0.001
R12158 VP.n8048 VP.n8045 0.001
R12159 VP.t28 VP.n8530 0.001
R12160 VP.t28 VP.n8527 0.001
R12161 VP.n8527 VP.n8524 0.001
R12162 VP.t207 VP.n8895 0.001
R12163 VP.t207 VP.n8892 0.001
R12164 VP.n8892 VP.n8889 0.001
R12165 VP.n9642 VP.t143 0.001
R12166 VP.n9659 VP.n9645 0.001
R12167 VP.t53 VP.n2236 0.001
R12168 VP.t53 VP.n2239 0.001
R12169 VP.t91 VP.n2376 0.001
R12170 VP.t91 VP.n2373 0.001
R12171 VP.n2373 VP.n2370 0.001
R12172 VP.t108 VP.n3165 0.001
R12173 VP.t108 VP.n3168 0.001
R12174 VP.t72 VP.n3627 0.001
R12175 VP.t72 VP.n3630 0.001
R12176 VP.t76 VP.n4058 0.001
R12177 VP.t76 VP.n4061 0.001
R12178 VP.t140 VP.n4506 0.001
R12179 VP.t140 VP.n4509 0.001
R12180 VP.t169 VP.n4941 0.001
R12181 VP.t169 VP.n4944 0.001
R12182 VP.t119 VP.n5428 0.001
R12183 VP.t119 VP.n5431 0.001
R12184 VP.t26 VP.n5778 0.001
R12185 VP.t26 VP.n5781 0.001
R12186 VP.t24 VP.n6256 0.001
R12187 VP.t24 VP.n6259 0.001
R12188 VP.t159 VP.n6622 0.001
R12189 VP.t159 VP.n6625 0.001
R12190 VP.t195 VP.n7143 0.001
R12191 VP.t195 VP.n7146 0.001
R12192 VP.t134 VP.n7434 0.001
R12193 VP.t134 VP.n7437 0.001
R12194 VP.t111 VP.n7943 0.001
R12195 VP.t111 VP.n7946 0.001
R12196 VP.t18 VP.n8250 0.001
R12197 VP.t18 VP.n8253 0.001
R12198 VP.n8808 VP.t28 0.001
R12199 VP.n8826 VP.n8811 0.001
R12200 VP.t57 VP.n725 0.001
R12201 VP.t57 VP.n728 0.001
R12202 VP.t49 VP.n1287 0.001
R12203 VP.t49 VP.n1290 0.001
R12204 VP.t34 VP.n1726 0.001
R12205 VP.t34 VP.n1729 0.001
R12206 VP.t34 VP.n1444 0.001
R12207 VP.n1444 VP.n1442 0.001
R12208 VP.n2629 VP.n2626 0.001
R12209 VP.n11032 VP.n11014 0.001
R12210 VP.n2654 VP.n2651 0.001
R12211 VP.n850 VP.n847 0.001
R12212 VP.n9659 VP.n9642 0.001
R12213 VP.n4610 VP.n4583 0.001
R12214 VP.n2685 VP.n2682 0.001
R12215 VP.n815 VP.n788 0.001
R12216 VP.n758 VP.n731 0.001
R12217 VP.n927 VP.n924 0.001
R12218 VP.n1747 VP.n1732 0.001
R12219 VP.n395 VP.n392 0.001
R12220 VP.n977 VP.n974 0.001
R12221 VP.n1483 VP.n1480 0.001
R12222 VP.n1916 VP.n1913 0.001
R12223 VP.n2708 VP.n2693 0.001
R12224 VP.n442 VP.n439 0.001
R12225 VP.n1027 VP.n1024 0.001
R12226 VP.n1521 VP.n1518 0.001
R12227 VP.n1968 VP.n1965 0.001
R12228 VP.n2897 VP.n2894 0.001
R12229 VP.n3648 VP.n3633 0.001
R12230 VP.n489 VP.n486 0.001
R12231 VP.n1077 VP.n1074 0.001
R12232 VP.n1559 VP.n1556 0.001
R12233 VP.n2020 VP.n2017 0.001
R12234 VP.n2949 VP.n2946 0.001
R12235 VP.n3461 VP.n3458 0.001
R12236 VP.n3842 VP.n3839 0.001
R12237 VP.n4554 VP.n4539 0.001
R12238 VP.n536 VP.n533 0.001
R12239 VP.n1127 VP.n1124 0.001
R12240 VP.n1597 VP.n1594 0.001
R12241 VP.n2072 VP.n2069 0.001
R12242 VP.n3001 VP.n2998 0.001
R12243 VP.n3499 VP.n3496 0.001
R12244 VP.n3894 VP.n3891 0.001
R12245 VP.n4378 VP.n4375 0.001
R12246 VP.n4777 VP.n4774 0.001
R12247 VP.n5449 VP.n5434 0.001
R12248 VP.n583 VP.n580 0.001
R12249 VP.n1165 VP.n1162 0.001
R12250 VP.n1629 VP.n1626 0.001
R12251 VP.n2113 VP.n2110 0.001
R12252 VP.n3042 VP.n3039 0.001
R12253 VP.n3531 VP.n3528 0.001
R12254 VP.n3935 VP.n3932 0.001
R12255 VP.n4410 VP.n4407 0.001
R12256 VP.n4818 VP.n4815 0.001
R12257 VP.n5332 VP.n5329 0.001
R12258 VP.n5655 VP.n5652 0.001
R12259 VP.n6305 VP.n6290 0.001
R12260 VP.n623 VP.n620 0.001
R12261 VP.n653 VP.n650 0.001
R12262 VP.n1661 VP.n1658 0.001
R12263 VP.n3563 VP.n3560 0.001
R12264 VP.n4442 VP.n4439 0.001
R12265 VP.n5364 VP.n5361 0.001
R12266 VP.n6192 VP.n6189 0.001
R12267 VP.n7164 VP.n7149 0.001
R12268 VP.n6540 VP.n6537 0.001
R12269 VP.n5696 VP.n5693 0.001
R12270 VP.n4859 VP.n4856 0.001
R12271 VP.n3976 VP.n3973 0.001
R12272 VP.n3083 VP.n3080 0.001
R12273 VP.n2154 VP.n2151 0.001
R12274 VP.n1205 VP.n1202 0.001
R12275 VP.n685 VP.n682 0.001
R12276 VP.n1693 VP.n1690 0.001
R12277 VP.n3595 VP.n3592 0.001
R12278 VP.n4474 VP.n4471 0.001
R12279 VP.n5396 VP.n5393 0.001
R12280 VP.n6224 VP.n6221 0.001
R12281 VP.n7111 VP.n7108 0.001
R12282 VP.n7992 VP.n7977 0.001
R12283 VP.n7393 VP.n7390 0.001
R12284 VP.n6581 VP.n6578 0.001
R12285 VP.n5737 VP.n5734 0.001
R12286 VP.n4900 VP.n4897 0.001
R12287 VP.n4017 VP.n4014 0.001
R12288 VP.n3124 VP.n3121 0.001
R12289 VP.n2195 VP.n2192 0.001
R12290 VP.n1246 VP.n1243 0.001
R12291 VP.n1287 VP.n1284 0.001
R12292 VP.n1726 VP.n1723 0.001
R12293 VP.n2236 VP.n2233 0.001
R12294 VP.n3165 VP.n3162 0.001
R12295 VP.n3627 VP.n3624 0.001
R12296 VP.n4058 VP.n4055 0.001
R12297 VP.n4506 VP.n4503 0.001
R12298 VP.n4941 VP.n4938 0.001
R12299 VP.n5428 VP.n5425 0.001
R12300 VP.n5778 VP.n5775 0.001
R12301 VP.n6256 VP.n6253 0.001
R12302 VP.n6622 VP.n6619 0.001
R12303 VP.n7143 VP.n7140 0.001
R12304 VP.n7434 VP.n7431 0.001
R12305 VP.n7943 VP.n7940 0.001
R12306 VP.n8250 VP.n8247 0.001
R12307 VP.n8826 VP.n8808 0.001
R12308 VP.n725 VP.n722 0.001
R12309 VP.n10467 VP.n10464 0.001
R12310 VP.n9859 VP.n9856 0.001
R12311 VP.n9097 VP.n9094 0.001
R12312 VP.n8300 VP.n8297 0.001
R12313 VP.n7483 VP.n7480 0.001
R12314 VP.n6671 VP.n6668 0.001
R12315 VP.n5828 VP.n5825 0.001
R12316 VP.n4991 VP.n4988 0.001
R12317 VP.n4108 VP.n4105 0.001
R12318 VP.n3216 VP.n3213 0.001
R12319 VP.n2266 VP.n2263 0.001
R12320 VP.n10502 VP.n10499 0.001
R12321 VP.n9907 VP.n9904 0.001
R12322 VP.n9147 VP.n9144 0.001
R12323 VP.n8349 VP.n8346 0.001
R12324 VP.n7532 VP.n7529 0.001
R12325 VP.n6720 VP.n6717 0.001
R12326 VP.n5878 VP.n5875 0.001
R12327 VP.n5043 VP.n5040 0.001
R12328 VP.n4533 VP.n4530 0.001
R12329 VP.n4137 VP.n4134 0.001
R12330 VP.n10537 VP.n10534 0.001
R12331 VP.n9955 VP.n9952 0.001
R12332 VP.n9197 VP.n9194 0.001
R12333 VP.n8398 VP.n8395 0.001
R12334 VP.n7581 VP.n7578 0.001
R12335 VP.n6771 VP.n6768 0.001
R12336 VP.n6284 VP.n6281 0.001
R12337 VP.n5907 VP.n5904 0.001
R12338 VP.n10572 VP.n10569 0.001
R12339 VP.n10003 VP.n10000 0.001
R12340 VP.n9247 VP.n9244 0.001
R12341 VP.n8449 VP.n8446 0.001
R12342 VP.n7971 VP.n7968 0.001
R12343 VP.n7610 VP.n7607 0.001
R12344 VP.n10607 VP.n10604 0.001
R12345 VP.n10043 VP.n10040 0.001
R12346 VP.n9636 VP.n9633 0.001
R12347 VP.n9276 VP.n9273 0.001
R12348 VP.n10645 VP.n10642 0.001
R12349 VP.n11008 VP.n11005 0.001
R12350 VP.n10074 VP.n10071 0.001
R12351 VP.n10670 VP.n10669 0.001
R12352 VP.n9670 VP.n9669 0.001
R12353 VP.n9291 VP.n9290 0.001
R12354 VP.n8464 VP.n8463 0.001
R12355 VP.n7625 VP.n7624 0.001
R12356 VP.n6786 VP.n6785 0.001
R12357 VP.n5922 VP.n5921 0.001
R12358 VP.n5058 VP.n5057 0.001
R12359 VP.n4152 VP.n4151 0.001
R12360 VP.n3231 VP.n3230 0.001
R12361 VP.n2281 VP.n2280 0.001
R12362 VP.n1304 VP.n1303 0.001
R12363 VP.n326 VP.n325 0.001
R12364 VP.n1294 VP.n1293 0.001
R12365 VP.n1307 VP.n1298 0.001
R12366 VP.n2284 VP.n2275 0.001
R12367 VP.n3234 VP.n3225 0.001
R12368 VP.n4155 VP.n4146 0.001
R12369 VP.n5061 VP.n5052 0.001
R12370 VP.n5925 VP.n5916 0.001
R12371 VP.n6789 VP.n6780 0.001
R12372 VP.n7628 VP.n7619 0.001
R12373 VP.n8467 VP.n8458 0.001
R12374 VP.n9294 VP.n9285 0.001
R12375 VP.n9673 VP.n9664 0.001
R12376 VP.n10673 VP.n10664 0.001
R12377 VP.n327 VP.n326 0.001
R12378 VP.n10669 VP.n10668 0.001
R12379 VP.n9669 VP.n9668 0.001
R12380 VP.n9290 VP.n9289 0.001
R12381 VP.n8463 VP.n8462 0.001
R12382 VP.n7624 VP.n7623 0.001
R12383 VP.n6785 VP.n6784 0.001
R12384 VP.n5921 VP.n5920 0.001
R12385 VP.n5057 VP.n5056 0.001
R12386 VP.n4151 VP.n4150 0.001
R12387 VP.n3230 VP.n3229 0.001
R12388 VP.n2280 VP.n2279 0.001
R12389 VP.n1303 VP.n1302 0.001
R12390 VP.n10163 VP.n10159 0.001
R12391 VP.n10757 VP.n10753 0.001
R12392 VP.n9419 VP.n9415 0.001
R12393 VP.n8966 VP.n8962 0.001
R12394 VP.n8620 VP.n8616 0.001
R12395 VP.n8122 VP.n8118 0.001
R12396 VP.n7781 VP.n7777 0.001
R12397 VP.n7294 VP.n7290 0.001
R12398 VP.n6943 VP.n6939 0.001
R12399 VP.n6435 VP.n6431 0.001
R12400 VP.n6079 VP.n6075 0.001
R12401 VP.n5579 VP.n5575 0.001
R12402 VP.n5214 VP.n5210 0.001
R12403 VP.n4684 VP.n4680 0.001
R12404 VP.n4309 VP.n4305 0.001
R12405 VP.n3785 VP.n3781 0.001
R12406 VP.n3390 VP.n3386 0.001
R12407 VP.n2840 VP.n2836 0.001
R12408 VP.t126 VP.n10099 0.001
R12409 VP.n10099 VP.n10096 0.001
R12410 fc2.n2640 fc2.n2639 180.813
R12411 fc2.n1515 fc2.n1514 168.716
R12412 fc2.n2798 fc2.n2797 138.352
R12413 fc2.n551 fc2.n550 138.352
R12414 fc2.n2436 fc2.n2435 138.352
R12415 fc2.n1009 fc2.n1008 138.352
R12416 fc2.n1538 fc2.n1537 138.352
R12417 fc2.n1520 fc2.n1519 138.352
R12418 fc2.n84 fc2.n83 138.125
R12419 fc2.n2792 fc2.n2791 138.125
R12420 fc2.n545 fc2.n544 138.125
R12421 fc2.n2430 fc2.n2429 138.125
R12422 fc2.n1003 fc2.n1002 138.125
R12423 fc2.n1533 fc2.n1532 138.125
R12424 fc2.n2795 fc2.n2794 129.015
R12425 fc2.n548 fc2.n547 129.015
R12426 fc2.n2433 fc2.n2432 129.015
R12427 fc2.n1006 fc2.n1005 129.015
R12428 fc2.n1535 fc2.n1534 129.015
R12429 fc2.n1513 fc2.n1512 129.015
R12430 fc2.n2640 fc2.t69 119.146
R12431 fc2.n2801 fc2.t19 119.146
R12432 fc2.n131 fc2.t8 119.146
R12433 fc2.n554 fc2.t43 119.146
R12434 fc2.n2001 fc2.t34 119.146
R12435 fc2.n2439 fc2.t0 119.146
R12436 fc2.n628 fc2.t2 119.146
R12437 fc2.n1012 fc2.t26 119.146
R12438 fc2.n1685 fc2.t16 119.146
R12439 fc2.n1541 fc2.t50 119.146
R12440 fc2.n1087 fc2.t41 119.146
R12441 fc2.n1523 fc2.t6 119.146
R12442 fc2.t14 fc2.n8 114.696
R12443 fc2.t4 fc2.n2658 114.696
R12444 fc2.t38 fc2.n2454 114.696
R12445 fc2.t66 fc2.n173 114.696
R12446 fc2.t62 fc2.n504 114.696
R12447 fc2.t98 fc2.n2074 114.696
R12448 fc2.t23 fc2.n2265 114.696
R12449 fc2.t52 fc2.n702 114.696
R12450 fc2.t47 fc2.n883 114.696
R12451 fc2.t12 fc2.n1759 114.696
R12452 fc2.t28 fc2.n1906 114.696
R12453 fc2.t10 fc2.n1132 114.696
R12454 fc2.t94 fc2.n1445 114.696
R12455 fc2.n2655 fc2.n2654 91.65
R12456 fc2.n1108 fc2.n1107 91.65
R12457 fc2.n1701 fc2.n1700 91.65
R12458 fc2.n644 fc2.n643 91.65
R12459 fc2.n2017 fc2.n2016 91.65
R12460 fc2.n147 fc2.n146 91.65
R12461 fc2.n541 fc2.n540 91.389
R12462 fc2.n2785 fc2.n2784 91.389
R12463 fc2.n2423 fc2.n2422 91.389
R12464 fc2.n1976 fc2.n1975 91.389
R12465 fc2.n1504 fc2.n1503 91.389
R12466 fc2.n996 fc2.n995 91.389
R12467 fc2.n7 fc2.n6 87.222
R12468 fc2.n47 fc2.n46 87.222
R12469 fc2.n41 fc2.n40 87.222
R12470 fc2.n27 fc2.n26 87.222
R12471 fc2.n20 fc2.n19 87.222
R12472 fc2.n34 fc2.n33 87.222
R12473 fc2.n3425 fc2.n3424 86.961
R12474 fc2.n3408 fc2.n3407 86.961
R12475 fc2.n3391 fc2.n3390 86.961
R12476 fc2.n3379 fc2.n3378 86.961
R12477 fc2.n3364 fc2.n3363 86.961
R12478 fc2.n3442 fc2.n3441 86.961
R12479 fc2.n1445 fc2.t21 21.258
R12480 fc2.n77 fc2.n76 7.273
R12481 fc2.n3292 fc2.t565 4.535
R12482 fc2.n3282 fc2.t725 4.535
R12483 fc2.n3272 fc2.t477 4.535
R12484 fc2.n3262 fc2.t436 4.535
R12485 fc2.n3252 fc2.t691 4.535
R12486 fc2.n3242 fc2.t545 4.535
R12487 fc2.n3232 fc2.t644 4.535
R12488 fc2.n3222 fc2.t713 4.535
R12489 fc2.n3212 fc2.t675 4.535
R12490 fc2.n3202 fc2.t699 4.535
R12491 fc2.n3191 fc2.t416 4.535
R12492 fc2.n3182 fc2.t568 4.535
R12493 fc2.n3084 fc2.t621 4.535
R12494 fc2.n3094 fc2.t503 4.535
R12495 fc2.n3114 fc2.t701 4.535
R12496 fc2.n3134 fc2.t752 4.535
R12497 fc2.n3154 fc2.t607 4.535
R12498 fc2.n3072 fc2.t423 4.535
R12499 fc2.n3162 fc2.t554 4.535
R12500 fc2.n3142 fc2.t459 4.535
R12501 fc2.n3122 fc2.t747 4.535
R12502 fc2.n3102 fc2.t659 4.535
R12503 fc2.n3013 fc2.t522 4.535
R12504 fc2.n3023 fc2.t695 4.535
R12505 fc2.n3043 fc2.t507 4.535
R12506 fc2.n3001 fc2.t419 4.535
R12507 fc2.n3051 fc2.t573 4.535
R12508 fc2.n3031 fc2.t438 4.535
R12509 fc2.n2979 fc2.t722 4.535
R12510 fc2.n2970 fc2.t418 4.535
R12511 fc2.n2919 fc2.t527 4.535
R12512 fc2.n2929 fc2.t724 4.535
R12513 fc2.n2907 fc2.t512 4.535
R12514 fc2.n2937 fc2.t618 4.535
R12515 fc2.n2828 fc2.t455 4.535
R12516 fc2.n2838 fc2.t581 4.535
R12517 fc2.n2858 fc2.t634 4.535
R12518 fc2.n2878 fc2.t622 4.535
R12519 fc2.n2816 fc2.t457 4.535
R12520 fc2.n2886 fc2.t739 4.535
R12521 fc2.n2866 fc2.t705 4.535
R12522 fc2.n2846 fc2.t600 4.535
R12523 fc2.n3689 fc2.t602 4.535
R12524 fc2.n3460 fc2.t587 4.535
R12525 fc2.n3561 fc2.t617 4.535
R12526 fc2.n3550 fc2.t543 4.535
R12527 fc2.n3540 fc2.t466 4.535
R12528 fc2.n3530 fc2.t413 4.535
R12529 fc2.n3520 fc2.t469 4.535
R12530 fc2.n3510 fc2.t401 4.535
R12531 fc2.n3500 fc2.t470 4.535
R12532 fc2.n3490 fc2.t681 4.535
R12533 fc2.n3480 fc2.t474 4.535
R12534 fc2.n3469 fc2.t537 4.535
R12535 fc2.n3870 fc2.t393 4.535
R12536 fc2.n3951 fc2.t670 4.535
R12537 fc2.n3941 fc2.t696 4.535
R12538 fc2.n3931 fc2.t519 4.535
R12539 fc2.n3921 fc2.t710 4.535
R12540 fc2.n3911 fc2.t505 4.535
R12541 fc2.n3901 fc2.t484 4.535
R12542 fc2.n3891 fc2.t569 4.535
R12543 fc2.n3878 fc2.t513 4.535
R12544 fc2.n3600 fc2.t683 4.535
R12545 fc2.n3661 fc2.t433 4.535
R12546 fc2.n3650 fc2.t561 4.535
R12547 fc2.n3640 fc2.t638 4.535
R12548 fc2.n3630 fc2.t479 4.535
R12549 fc2.n3620 fc2.t396 4.535
R12550 fc2.n3609 fc2.t597 4.535
R12551 fc2.n3787 fc2.t541 4.535
R12552 fc2.n3828 fc2.t407 4.535
R12553 fc2.n3818 fc2.t591 4.535
R12554 fc2.n3808 fc2.t735 4.535
R12555 fc2.n3795 fc2.t726 4.535
R12556 fc2.n3701 fc2.t652 4.535
R12557 fc2.n3711 fc2.t431 4.535
R12558 fc2.n3748 fc2.t446 4.535
R12559 fc2.n3296 fc2.t481 4.472
R12560 fc2.n3286 fc2.t440 4.472
R12561 fc2.n3276 fc2.t676 4.472
R12562 fc2.n3266 fc2.t647 4.472
R12563 fc2.n3256 fc2.t449 4.472
R12564 fc2.n3246 fc2.t627 4.472
R12565 fc2.n3236 fc2.t511 4.472
R12566 fc2.n3226 fc2.t640 4.472
R12567 fc2.n3216 fc2.t628 4.472
R12568 fc2.n3206 fc2.t542 4.472
R12569 fc2.n3195 fc2.t590 4.472
R12570 fc2.n3186 fc2.t506 4.472
R12571 fc2.n3766 fc2.t490 4.472
R12572 fc2.n3087 fc2.t398 4.472
R12573 fc2.n3097 fc2.t662 4.472
R12574 fc2.n3117 fc2.t692 4.472
R12575 fc2.n3137 fc2.t744 4.472
R12576 fc2.n3157 fc2.t698 4.472
R12577 fc2.n3075 fc2.t672 4.472
R12578 fc2.n3166 fc2.t635 4.472
R12579 fc2.n3146 fc2.t584 4.472
R12580 fc2.n3126 fc2.t564 4.472
R12581 fc2.n3106 fc2.t454 4.472
R12582 fc2.n3016 fc2.t482 4.472
R12583 fc2.n3026 fc2.t421 4.472
R12584 fc2.n3046 fc2.t478 4.472
R12585 fc2.n3004 fc2.t492 4.472
R12586 fc2.n3055 fc2.t500 4.472
R12587 fc2.n3035 fc2.t552 4.472
R12588 fc2.n2982 fc2.t468 4.472
R12589 fc2.n2973 fc2.t444 4.472
R12590 fc2.n2922 fc2.t462 4.472
R12591 fc2.n2932 fc2.t430 4.472
R12592 fc2.n2910 fc2.t605 4.472
R12593 fc2.n2941 fc2.t624 4.472
R12594 fc2.n2831 fc2.t677 4.472
R12595 fc2.n2841 fc2.t595 4.472
R12596 fc2.n2861 fc2.t749 4.472
R12597 fc2.n2881 fc2.t667 4.472
R12598 fc2.n2819 fc2.t708 4.472
R12599 fc2.n2890 fc2.t671 4.472
R12600 fc2.n2870 fc2.t690 4.472
R12601 fc2.n2850 fc2.t737 4.472
R12602 fc2.n3692 fc2.t653 4.472
R12603 fc2.n3571 fc2.t633 4.472
R12604 fc2.n3565 fc2.t405 4.472
R12605 fc2.n3554 fc2.t495 4.472
R12606 fc2.n3544 fc2.t411 4.472
R12607 fc2.n3534 fc2.t452 4.472
R12608 fc2.n3524 fc2.t571 4.472
R12609 fc2.n3514 fc2.t551 4.472
R12610 fc2.n3504 fc2.t585 4.472
R12611 fc2.n3494 fc2.t504 4.472
R12612 fc2.n3484 fc2.t528 4.472
R12613 fc2.n3473 fc2.t656 4.472
R12614 fc2.n3970 fc2.t738 4.472
R12615 fc2.n3955 fc2.t576 4.472
R12616 fc2.n3945 fc2.t753 4.472
R12617 fc2.n3935 fc2.t494 4.472
R12618 fc2.n3925 fc2.t697 4.472
R12619 fc2.n3915 fc2.t533 4.472
R12620 fc2.n3905 fc2.t711 4.472
R12621 fc2.n3895 fc2.t535 4.472
R12622 fc2.n3882 fc2.t465 4.472
R12623 fc2.n3671 fc2.t748 4.472
R12624 fc2.n3665 fc2.t451 4.472
R12625 fc2.n3654 fc2.t733 4.472
R12626 fc2.n3644 fc2.t435 4.472
R12627 fc2.n3634 fc2.t403 4.472
R12628 fc2.n3624 fc2.t460 4.472
R12629 fc2.n3613 fc2.t402 4.472
R12630 fc2.n3847 fc2.t577 4.472
R12631 fc2.n3832 fc2.t650 4.472
R12632 fc2.n3822 fc2.t408 4.472
R12633 fc2.n3812 fc2.t530 4.472
R12634 fc2.n3799 fc2.t728 4.472
R12635 fc2.n3731 fc2.t593 4.472
R12636 fc2.n3705 fc2.t463 4.472
R12637 fc2.n3295 fc2.t502 4.237
R12638 fc2.n3285 fc2.t727 4.237
R12639 fc2.n3275 fc2.t532 4.237
R12640 fc2.n3265 fc2.t499 4.237
R12641 fc2.n3255 fc2.t694 4.237
R12642 fc2.n3245 fc2.t615 4.237
R12643 fc2.n3235 fc2.t574 4.237
R12644 fc2.n3225 fc2.t736 4.237
R12645 fc2.n3215 fc2.t442 4.237
R12646 fc2.n3205 fc2.t501 4.237
R12647 fc2.n3194 fc2.t458 4.237
R12648 fc2.n3185 fc2.t529 4.237
R12649 fc2.n3086 fc2.t680 4.237
R12650 fc2.n3096 fc2.t559 4.237
R12651 fc2.n3116 fc2.t734 4.237
R12652 fc2.n3136 fc2.t417 4.237
R12653 fc2.n3156 fc2.t723 4.237
R12654 fc2.n3074 fc2.t439 4.237
R12655 fc2.n3066 fc2.t611 4.237
R12656 fc2.n3165 fc2.t580 4.237
R12657 fc2.n3145 fc2.t447 4.237
R12658 fc2.n3125 fc2.t480 4.237
R12659 fc2.n3105 fc2.t473 4.237
R12660 fc2.n3015 fc2.t626 4.237
R12661 fc2.n3025 fc2.t497 4.237
R12662 fc2.n3045 fc2.t707 4.237
R12663 fc2.n3003 fc2.t437 4.237
R12664 fc2.n2995 fc2.t601 4.237
R12665 fc2.n3054 fc2.t623 4.237
R12666 fc2.n3034 fc2.t685 4.237
R12667 fc2.n2981 fc2.t714 4.237
R12668 fc2.n2972 fc2.t488 4.237
R12669 fc2.n2963 fc2.t472 4.237
R12670 fc2.n2953 fc2.t415 4.237
R12671 fc2.n2921 fc2.t406 4.237
R12672 fc2.n2931 fc2.t646 4.237
R12673 fc2.n2909 fc2.t718 4.237
R12674 fc2.n2901 fc2.t630 4.237
R12675 fc2.n2940 fc2.t538 4.237
R12676 fc2.n2830 fc2.t750 4.237
R12677 fc2.n2840 fc2.t556 4.237
R12678 fc2.n2860 fc2.t616 4.237
R12679 fc2.n2880 fc2.t654 4.237
R12680 fc2.n2818 fc2.t570 4.237
R12681 fc2.n2810 fc2.t562 4.237
R12682 fc2.n2889 fc2.t575 4.237
R12683 fc2.n2869 fc2.t660 4.237
R12684 fc2.n2849 fc2.t663 4.237
R12685 fc2.n3691 fc2.t510 4.237
R12686 fc2.n3564 fc2.t703 4.237
R12687 fc2.n3553 fc2.t521 4.237
R12688 fc2.n3543 fc2.t429 4.237
R12689 fc2.n3533 fc2.t746 4.237
R12690 fc2.n3523 fc2.t567 4.237
R12691 fc2.n3513 fc2.t489 4.237
R12692 fc2.n3503 fc2.t606 4.237
R12693 fc2.n3493 fc2.t400 4.237
R12694 fc2.n3483 fc2.t731 4.237
R12695 fc2.n3472 fc2.t609 4.237
R12696 fc2.n3954 fc2.t594 4.237
R12697 fc2.n3944 fc2.t516 4.237
R12698 fc2.n3934 fc2.t420 4.237
R12699 fc2.n3924 fc2.t674 4.237
R12700 fc2.n3914 fc2.t448 4.237
R12701 fc2.n3904 fc2.t534 4.237
R12702 fc2.n3894 fc2.t592 4.237
R12703 fc2.n3881 fc2.t441 4.237
R12704 fc2.n3664 fc2.t456 4.237
R12705 fc2.n3653 fc2.t404 4.237
R12706 fc2.n3643 fc2.t544 4.237
R12707 fc2.n3633 fc2.t673 4.237
R12708 fc2.n3623 fc2.t550 4.237
R12709 fc2.n3612 fc2.t655 4.237
R12710 fc2.n3831 fc2.t651 4.237
R12711 fc2.n3821 fc2.t665 4.237
R12712 fc2.n3811 fc2.t612 4.237
R12713 fc2.n3798 fc2.t399 4.237
R12714 fc2.n3704 fc2.t599 4.237
R12715 fc2.n3079 fc2.t547 4.231
R12716 fc2.n3008 fc2.t471 4.231
R12717 fc2.n2957 fc2.t719 4.231
R12718 fc2.n2914 fc2.t524 4.231
R12719 fc2.n2823 fc2.t432 4.231
R12720 fc2.n3179 fc2.t555 4.231
R12721 fc2.n3767 fc2.t648 4.231
R12722 fc2.n3572 fc2.t686 4.231
R12723 fc2.n3971 fc2.t525 4.231
R12724 fc2.n3672 fc2.t625 4.231
R12725 fc2.n3848 fc2.t709 4.231
R12726 fc2.n3732 fc2.t588 4.231
R12727 fc2.n3177 fc2.t682 4.221
R12728 fc2.n3067 fc2.t526 4.221
R12729 fc2.n2996 fc2.t572 4.221
R12730 fc2.n2964 fc2.t642 4.221
R12731 fc2.n2954 fc2.t740 4.221
R12732 fc2.n2902 fc2.t476 4.221
R12733 fc2.n2811 fc2.t428 4.221
R12734 fc2.n3461 fc2.t742 4.221
R12735 fc2.n3871 fc2.t536 4.221
R12736 fc2.n3601 fc2.t464 4.221
R12737 fc2.n3788 fc2.t409 4.221
R12738 fc2.n3712 fc2.t730 4.221
R12739 fc2.n3749 fc2.t422 4.221
R12740 fc2.n2988 fc2.t467 4.196
R12741 fc2.n3293 fc2.t517 4.182
R12742 fc2.n3283 fc2.t632 4.182
R12743 fc2.n3273 fc2.t729 4.182
R12744 fc2.n3263 fc2.t687 4.182
R12745 fc2.n3253 fc2.t598 4.182
R12746 fc2.n3243 fc2.t397 4.182
R12747 fc2.n3233 fc2.t391 4.182
R12748 fc2.n3223 fc2.t434 4.182
R12749 fc2.n3213 fc2.t596 4.182
R12750 fc2.n3203 fc2.t486 4.182
R12751 fc2.n3192 fc2.t485 4.182
R12752 fc2.n3183 fc2.t716 4.182
R12753 fc2.n3083 fc2.t540 4.182
R12754 fc2.n3093 fc2.t548 4.182
R12755 fc2.n3113 fc2.t549 4.182
R12756 fc2.n3133 fc2.t520 4.182
R12757 fc2.n3153 fc2.t491 4.182
R12758 fc2.n3071 fc2.t583 4.182
R12759 fc2.n3163 fc2.t610 4.182
R12760 fc2.n3143 fc2.t712 4.182
R12761 fc2.n3123 fc2.t743 4.182
R12762 fc2.n3103 fc2.t678 4.182
R12763 fc2.n3078 fc2.t410 4.182
R12764 fc2.n3012 fc2.t483 4.182
R12765 fc2.n3022 fc2.t426 4.182
R12766 fc2.n3042 fc2.t498 4.182
R12767 fc2.n3000 fc2.t563 4.182
R12768 fc2.n3052 fc2.t717 4.182
R12769 fc2.n3032 fc2.t578 4.182
R12770 fc2.n3007 fc2.t531 4.182
R12771 fc2.n2978 fc2.t445 4.182
R12772 fc2.n2969 fc2.t720 4.182
R12773 fc2.n2986 fc2.t450 4.182
R12774 fc2.n2956 fc2.t523 4.182
R12775 fc2.n2918 fc2.t629 4.182
R12776 fc2.n2928 fc2.t496 4.182
R12777 fc2.n2906 fc2.t639 4.182
R12778 fc2.n2938 fc2.t664 4.182
R12779 fc2.n2913 fc2.t741 4.182
R12780 fc2.n2827 fc2.t509 4.182
R12781 fc2.n2837 fc2.t461 4.182
R12782 fc2.n2857 fc2.t636 4.182
R12783 fc2.n2877 fc2.t508 4.182
R12784 fc2.n2815 fc2.t589 4.182
R12785 fc2.n2887 fc2.t631 4.182
R12786 fc2.n2867 fc2.t700 4.182
R12787 fc2.n2847 fc2.t425 4.182
R12788 fc2.n2822 fc2.t643 4.182
R12789 fc2.n3688 fc2.t751 4.182
R12790 fc2.n3562 fc2.t518 4.182
R12791 fc2.n3551 fc2.t553 4.182
R12792 fc2.n3541 fc2.t453 4.182
R12793 fc2.n3531 fc2.t688 4.182
R12794 fc2.n3521 fc2.t414 4.182
R12795 fc2.n3511 fc2.t539 4.182
R12796 fc2.n3501 fc2.t582 4.182
R12797 fc2.n3491 fc2.t604 4.182
R12798 fc2.n3481 fc2.t637 4.182
R12799 fc2.n3470 fc2.t721 4.182
R12800 fc2.n3952 fc2.t669 4.182
R12801 fc2.n3942 fc2.t560 4.182
R12802 fc2.n3932 fc2.t754 4.182
R12803 fc2.n3922 fc2.t392 4.182
R12804 fc2.n3912 fc2.t608 4.182
R12805 fc2.n3902 fc2.t658 4.182
R12806 fc2.n3892 fc2.t546 4.182
R12807 fc2.n3879 fc2.t475 4.182
R12808 fc2.n3662 fc2.t649 4.182
R12809 fc2.n3651 fc2.t586 4.182
R12810 fc2.n3641 fc2.t412 4.182
R12811 fc2.n3631 fc2.t566 4.182
R12812 fc2.n3621 fc2.t702 4.182
R12813 fc2.n3610 fc2.t666 4.182
R12814 fc2.n3829 fc2.t645 4.182
R12815 fc2.n3819 fc2.t614 4.182
R12816 fc2.n3809 fc2.t684 4.182
R12817 fc2.n3796 fc2.t732 4.182
R12818 fc2.n3702 fc2.t668 4.182
R12819 fc2.n2987 fc2.t693 3.951
R12820 fc2.n3177 fc2.t745 3.921
R12821 fc2.n3768 fc2.t493 3.917
R12822 fc2.n3080 fc2.t619 3.917
R12823 fc2.n3009 fc2.t443 3.917
R12824 fc2.n2958 fc2.t715 3.917
R12825 fc2.n2915 fc2.t613 3.917
R12826 fc2.n2824 fc2.t706 3.917
R12827 fc2.n3573 fc2.t487 3.917
R12828 fc2.n3972 fc2.t679 3.917
R12829 fc2.n3673 fc2.t603 3.917
R12830 fc2.n3849 fc2.t395 3.917
R12831 fc2.n3733 fc2.t689 3.917
R12832 fc2.n2632 fc2.t295 3.904
R12833 fc2.n2634 fc2.n2633 3.904
R12834 fc2.n289 fc2.n288 3.904
R12835 fc2.n296 fc2.t82 3.904
R12836 fc2.n300 fc2.n299 3.904
R12837 fc2.n292 fc2.t25 3.904
R12838 fc2.n50 fc2.t146 3.904
R12839 fc2.n2616 fc2.n2615 3.904
R12840 fc2.n2583 fc2.t367 3.904
R12841 fc2.n2610 fc2.n2609 3.904
R12842 fc2.n2585 fc2.t292 3.904
R12843 fc2.n541 fc2.t193 3.904
R12844 fc2.n339 fc2.t125 3.904
R12845 fc2.n9 fc2.t278 3.904
R12846 fc2.n2656 fc2.t255 3.904
R12847 fc2.n2463 fc2.n2462 3.904
R12848 fc2.n2474 fc2.t39 3.904
R12849 fc2.n2477 fc2.t359 3.904
R12850 fc2.n2460 fc2.n2459 3.904
R12851 fc2.n159 fc2.n158 3.904
R12852 fc2.n171 fc2.t152 3.904
R12853 fc2.n168 fc2.t84 3.904
R12854 fc2.n156 fc2.n155 3.904
R12855 fc2.n521 fc2.n520 3.904
R12856 fc2.n535 fc2.t245 3.904
R12857 fc2.n538 fc2.t388 3.904
R12858 fc2.n518 fc2.n517 3.904
R12859 fc2.n2061 fc2.n2060 3.904
R12860 fc2.n2072 fc2.t253 3.904
R12861 fc2.n2069 fc2.t116 3.904
R12862 fc2.n2058 fc2.n2057 3.904
R12863 fc2.n2255 fc2.n2254 3.904
R12864 fc2.n2263 fc2.t345 3.904
R12865 fc2.n2237 fc2.t293 3.904
R12866 fc2.n2252 fc2.n2251 3.904
R12867 fc2.n689 fc2.n688 3.904
R12868 fc2.n700 fc2.t83 3.904
R12869 fc2.n697 fc2.t385 3.904
R12870 fc2.n686 fc2.n685 3.904
R12871 fc2.n870 fc2.n869 3.904
R12872 fc2.n881 fc2.t176 3.904
R12873 fc2.n878 fc2.t126 3.904
R12874 fc2.n867 fc2.n866 3.904
R12875 fc2.n1746 fc2.n1745 3.904
R12876 fc2.n1757 fc2.t285 3.904
R12877 fc2.n1754 fc2.t211 3.904
R12878 fc2.n1743 fc2.n1742 3.904
R12879 fc2.n1893 fc2.n1892 3.904
R12880 fc2.n1904 fc2.t379 3.904
R12881 fc2.n1901 fc2.t324 3.904
R12882 fc2.n1890 fc2.n1889 3.904
R12883 fc2.n1119 fc2.n1118 3.904
R12884 fc2.n1130 fc2.t119 3.904
R12885 fc2.n1127 fc2.t42 3.904
R12886 fc2.n1116 fc2.n1115 3.904
R12887 fc2.n1430 fc2.n1429 3.904
R12888 fc2.n1443 fc2.t224 3.904
R12889 fc2.n1440 fc2.t155 3.904
R12890 fc2.n1427 fc2.n1426 3.904
R12891 fc2.n45 fc2.t30 3.904
R12892 fc2.n2730 fc2.n2729 3.904
R12893 fc2.n2742 fc2.t167 3.904
R12894 fc2.n2745 fc2.t77 3.904
R12895 fc2.n2727 fc2.n2726 3.904
R12896 fc2.n2785 fc2.t237 3.904
R12897 fc2.n2787 fc2.t164 3.904
R12898 fc2.n38 fc2.t269 3.904
R12899 fc2.n2713 fc2.n2712 3.904
R12900 fc2.n2720 fc2.t49 3.904
R12901 fc2.n2723 fc2.t313 3.904
R12902 fc2.n2716 fc2.n2715 3.904
R12903 fc2.n2552 fc2.n2551 3.904
R12904 fc2.n2577 fc2.t107 3.904
R12905 fc2.n2580 fc2.t45 3.904
R12906 fc2.n2549 fc2.n2548 3.904
R12907 fc2.n247 fc2.n246 3.904
R12908 fc2.n267 fc2.t206 3.904
R12909 fc2.n270 fc2.t143 3.904
R12910 fc2.n244 fc2.n243 3.904
R12911 fc2.n357 fc2.n356 3.904
R12912 fc2.n383 fc2.t323 3.904
R12913 fc2.n380 fc2.t250 3.904
R12914 fc2.n354 fc2.n353 3.904
R12915 fc2.n2165 fc2.n2164 3.904
R12916 fc2.n2162 fc2.t118 3.904
R12917 fc2.n2159 fc2.t362 3.904
R12918 fc2.n1990 fc2.n1989 3.904
R12919 fc2.n2423 fc2.t223 3.904
R12920 fc2.n2425 fc2.t153 3.904
R12921 fc2.n1976 fc2.t142 3.904
R12922 fc2.n1973 fc2.t68 3.904
R12923 fc2.n1765 fc2.n1764 3.904
R12924 fc2.n1784 fc2.t13 3.904
R12925 fc2.n1787 fc2.t350 3.904
R12926 fc2.n1762 fc2.n1761 3.904
R12927 fc2.n937 fc2.n936 3.904
R12928 fc2.n960 fc2.t312 3.904
R12929 fc2.n963 fc2.t238 3.904
R12930 fc2.n934 fc2.n933 3.904
R12931 fc2.n712 fc2.n711 3.904
R12932 fc2.n731 fc2.t197 3.904
R12933 fc2.n734 fc2.t133 3.904
R12934 fc2.n709 fc2.n708 3.904
R12935 fc2.n2320 fc2.n2319 3.904
R12936 fc2.n2343 fc2.t93 3.904
R12937 fc2.n2346 fc2.t31 3.904
R12938 fc2.n2317 fc2.n2316 3.904
R12939 fc2.n2084 fc2.n2083 3.904
R12940 fc2.n2103 fc2.t369 3.904
R12941 fc2.n2106 fc2.t225 3.904
R12942 fc2.n2081 fc2.n2080 3.904
R12943 fc2.n433 fc2.n432 3.904
R12944 fc2.n459 fc2.t186 3.904
R12945 fc2.n456 fc2.t135 3.904
R12946 fc2.n430 fc2.n429 3.904
R12947 fc2.n183 fc2.n182 3.904
R12948 fc2.n203 fc2.t97 3.904
R12949 fc2.n206 fc2.t9 3.904
R12950 fc2.n180 fc2.n179 3.904
R12951 fc2.n2485 fc2.n2484 3.904
R12952 fc2.n2509 fc2.t356 3.904
R12953 fc2.n2512 fc2.t303 3.904
R12954 fc2.n2482 fc2.n2481 3.904
R12955 fc2.n2664 fc2.n2663 3.904
R12956 fc2.n2675 fc2.t307 3.904
R12957 fc2.n2678 fc2.t195 3.904
R12958 fc2.n2661 fc2.n2660 3.904
R12959 fc2.n23 fc2.t328 3.904
R12960 fc2.n17 fc2.t87 3.904
R12961 fc2.n2756 fc2.n2755 3.904
R12962 fc2.n2753 fc2.t233 3.904
R12963 fc2.n2750 fc2.t129 3.904
R12964 fc2.n2619 fc2.n2618 3.904
R12965 fc2.n2772 fc2.n2771 3.904
R12966 fc2.n2779 fc2.t288 3.904
R12967 fc2.n2782 fc2.t61 3.904
R12968 fc2.n2769 fc2.n2768 3.904
R12969 fc2.n275 fc2.n274 3.904
R12970 fc2.n283 fc2.t218 3.904
R12971 fc2.n286 fc2.t157 3.904
R12972 fc2.n278 fc2.n277 3.904
R12973 fc2.n324 fc2.n323 3.904
R12974 fc2.n337 fc2.t316 3.904
R12975 fc2.n327 fc2.t260 3.904
R12976 fc2.n330 fc2.n329 3.904
R12977 fc2.n2144 fc2.n2143 3.904
R12978 fc2.n2153 fc2.t128 3.904
R12979 fc2.n2156 fc2.t352 3.904
R12980 fc2.n2147 fc2.n2146 3.904
R12981 fc2.n2399 fc2.n2398 3.904
R12982 fc2.n2417 fc2.t214 3.904
R12983 fc2.n2420 fc2.t165 3.904
R12984 fc2.n2402 fc2.n2401 3.904
R12985 fc2.n769 fc2.n768 3.904
R12986 fc2.n780 fc2.t325 3.904
R12987 fc2.n783 fc2.t258 3.904
R12988 fc2.n772 fc2.n771 3.904
R12989 fc2.n972 fc2.n971 3.904
R12990 fc2.n990 fc2.t48 3.904
R12991 fc2.n993 fc2.t368 3.904
R12992 fc2.n975 fc2.n974 3.904
R12993 fc2.n1792 fc2.n1791 3.904
R12994 fc2.n1803 fc2.t160 3.904
R12995 fc2.n1806 fc2.t89 3.904
R12996 fc2.n1795 fc2.n1794 3.904
R12997 fc2.n1952 fc2.n1951 3.904
R12998 fc2.n1968 fc2.t266 3.904
R12999 fc2.n1971 fc2.t194 3.904
R13000 fc2.n1955 fc2.n1954 3.904
R13001 fc2.n1167 fc2.n1166 3.904
R13002 fc2.n1181 fc2.t354 3.904
R13003 fc2.n1184 fc2.t310 3.904
R13004 fc2.n1170 fc2.n1169 3.904
R13005 fc2.n1504 fc2.t103 3.904
R13006 fc2.n1501 fc2.t7 3.904
R13007 fc2.n31 fc2.t15 3.904
R13008 fc2.n2689 fc2.n2688 3.904
R13009 fc2.n2696 fc2.t178 3.904
R13010 fc2.n2699 fc2.t70 3.904
R13011 fc2.n2692 fc2.n2691 3.904
R13012 fc2.n2534 fc2.n2533 3.904
R13013 fc2.n2542 fc2.t227 3.904
R13014 fc2.n2545 fc2.t175 3.904
R13015 fc2.n2537 fc2.n2536 3.904
R13016 fc2.n213 fc2.n212 3.904
R13017 fc2.n233 fc2.t338 3.904
R13018 fc2.n236 fc2.t267 3.904
R13019 fc2.n210 fc2.n209 3.904
R13020 fc2.n391 fc2.n390 3.904
R13021 fc2.n417 fc2.t63 3.904
R13022 fc2.n414 fc2.t377 3.904
R13023 fc2.n388 fc2.n387 3.904
R13024 fc2.n2117 fc2.n2116 3.904
R13025 fc2.n2136 fc2.t241 3.904
R13026 fc2.n2139 fc2.t104 3.904
R13027 fc2.n2114 fc2.n2113 3.904
R13028 fc2.n2364 fc2.n2363 3.904
R13029 fc2.n2387 fc2.t351 3.904
R13030 fc2.n2390 fc2.t280 3.904
R13031 fc2.n2361 fc2.n2360 3.904
R13032 fc2.n742 fc2.n741 3.904
R13033 fc2.n761 fc2.t73 3.904
R13034 fc2.n764 fc2.t3 3.904
R13035 fc2.n739 fc2.n738 3.904
R13036 fc2.n996 fc2.t183 3.904
R13037 fc2.n998 fc2.t113 3.904
R13038 fc2.n3314 fc2.t22 3.904
R13039 fc2.n1109 fc2.t120 3.904
R13040 fc2.n1472 fc2.n1471 3.904
R13041 fc2.n1496 fc2.t276 3.904
R13042 fc2.n1499 fc2.t219 3.904
R13043 fc2.n1469 fc2.n1468 3.904
R13044 fc2.n3425 fc2.t273 3.904
R13045 fc2.n3419 fc2.t384 3.904
R13046 fc2.n1702 fc2.t161 3.904
R13047 fc2.n1919 fc2.n1918 3.904
R13048 fc2.n1940 fc2.t319 3.904
R13049 fc2.n1943 fc2.t264 3.904
R13050 fc2.n1916 fc2.n1915 3.904
R13051 fc2.n1139 fc2.n1138 3.904
R13052 fc2.n1159 fc2.t55 3.904
R13053 fc2.n1162 fc2.t357 3.904
R13054 fc2.n1136 fc2.n1135 3.904
R13055 fc2.n1039 fc2.n1038 3.904
R13056 fc2.n1068 fc2.t150 3.904
R13057 fc2.n1065 fc2.t294 3.904
R13058 fc2.n1036 fc2.n1035 3.904
R13059 fc2.n3408 fc2.t344 3.904
R13060 fc2.n3396 fc2.t85 3.904
R13061 fc2.n645 fc2.t199 3.904
R13062 fc2.n896 fc2.n895 3.904
R13063 fc2.n918 fc2.t361 3.904
R13064 fc2.n921 fc2.t308 3.904
R13065 fc2.n893 fc2.n892 3.904
R13066 fc2.n1714 fc2.n1713 3.904
R13067 fc2.n1736 fc2.t101 3.904
R13068 fc2.n1733 fc2.t17 3.904
R13069 fc2.n1711 fc2.n1710 3.904
R13070 fc2.n1563 fc2.n1562 3.904
R13071 fc2.n1589 fc2.t189 3.904
R13072 fc2.n1586 fc2.t335 3.904
R13073 fc2.n1560 fc2.n1559 3.904
R13074 fc2.n1193 fc2.n1192 3.904
R13075 fc2.n1190 fc2.t130 3.904
R13076 fc2.n1187 fc2.t59 3.904
R13077 fc2.n1074 fc2.n1073 3.904
R13078 fc2.n1227 fc2.n1226 3.904
R13079 fc2.n1256 fc2.t215 3.904
R13080 fc2.n1253 fc2.t166 3.904
R13081 fc2.n1224 fc2.n1223 3.904
R13082 fc2.n3391 fc2.t213 3.904
R13083 fc2.n3382 fc2.t326 3.904
R13084 fc2.n2018 fc2.t169 3.904
R13085 fc2.n2281 fc2.n2280 3.904
R13086 fc2.n2304 fc2.t24 3.904
R13087 fc2.n2278 fc2.t349 3.904
R13088 fc2.n2275 fc2.n2274 3.904
R13089 fc2.n657 fc2.n656 3.904
R13090 fc2.n679 fc2.t140 3.904
R13091 fc2.n676 fc2.t74 3.904
R13092 fc2.n654 fc2.n653 3.904
R13093 fc2.n583 fc2.n582 3.904
R13094 fc2.n609 fc2.t231 3.904
R13095 fc2.n606 fc2.t378 3.904
R13096 fc2.n580 fc2.n579 3.904
R13097 fc2.n1606 fc2.n1605 3.904
R13098 fc2.n1603 fc2.t168 3.904
R13099 fc2.n1600 fc2.t106 3.904
R13100 fc2.n1597 fc2.n1596 3.904
R13101 fc2.n1639 fc2.n1638 3.904
R13102 fc2.n1665 fc2.t261 3.904
R13103 fc2.n1662 fc2.t205 3.904
R13104 fc2.n1636 fc2.n1635 3.904
R13105 fc2.n1271 fc2.n1270 3.904
R13106 fc2.n1268 fc2.t370 3.904
R13107 fc2.n1265 fc2.t301 3.904
R13108 fc2.n1262 fc2.n1261 3.904
R13109 fc2.n1305 fc2.n1304 3.904
R13110 fc2.n1334 fc2.t95 3.904
R13111 fc2.n1331 fc2.t32 3.904
R13112 fc2.n1302 fc2.n1301 3.904
R13113 fc2.n3379 fc2.t92 3.904
R13114 fc2.n3367 fc2.t200 3.904
R13115 fc2.n148 fc2.t208 3.904
R13116 fc2.n476 fc2.n475 3.904
R13117 fc2.n502 fc2.t373 3.904
R13118 fc2.n499 fc2.t318 3.904
R13119 fc2.n473 fc2.n472 3.904
R13120 fc2.n2029 fc2.n2028 3.904
R13121 fc2.n2051 fc2.t181 3.904
R13122 fc2.n2048 fc2.t35 3.904
R13123 fc2.n2026 fc2.n2025 3.904
R13124 fc2.n2208 fc2.n2207 3.904
R13125 fc2.n2234 fc2.t274 3.904
R13126 fc2.n2231 fc2.t46 3.904
R13127 fc2.n2205 fc2.n2204 3.904
R13128 fc2.n792 fc2.n791 3.904
R13129 fc2.n789 fc2.t207 3.904
R13130 fc2.n786 fc2.t144 3.904
R13131 fc2.n616 fc2.n615 3.904
R13132 fc2.n826 fc2.n825 3.904
R13133 fc2.n852 fc2.t305 3.904
R13134 fc2.n849 fc2.t251 3.904
R13135 fc2.n823 fc2.n822 3.904
R13136 fc2.n1815 fc2.n1814 3.904
R13137 fc2.n1812 fc2.t33 3.904
R13138 fc2.n1809 fc2.t342 3.904
R13139 fc2.n1672 fc2.n1671 3.904
R13140 fc2.n1849 fc2.n1848 3.904
R13141 fc2.n1875 fc2.t136 3.904
R13142 fc2.n1872 fc2.t81 3.904
R13143 fc2.n1846 fc2.n1845 3.904
R13144 fc2.n1349 fc2.n1348 3.904
R13145 fc2.n1346 fc2.t242 3.904
R13146 fc2.n1343 fc2.t174 3.904
R13147 fc2.n1340 fc2.n1339 3.904
R13148 fc2.n1383 fc2.n1382 3.904
R13149 fc2.n1412 fc2.t336 3.904
R13150 fc2.n1409 fc2.t282 3.904
R13151 fc2.n1380 fc2.n1379 3.904
R13152 fc2.n3364 fc2.t333 3.904
R13153 fc2.n3351 fc2.t75 3.904
R13154 fc2.n3440 fc2.t314 3.904
R13155 fc2.n3442 fc2.t221 3.904
R13156 fc2.n2622 fc2.t184 3.904
R13157 fc2.n2748 fc2.n2747 3.904
R13158 fc2.n3179 fc2.t558 3.897
R13159 fc2.n3065 fc2.t394 3.894
R13160 fc2.n2994 fc2.t704 3.894
R13161 fc2.n2965 fc2.t514 3.894
R13162 fc2.n2952 fc2.t557 3.894
R13163 fc2.n2900 fc2.t620 3.894
R13164 fc2.n2809 fc2.t579 3.894
R13165 fc2.n3459 fc2.t661 3.894
R13166 fc2.n3869 fc2.t427 3.894
R13167 fc2.n3599 fc2.t424 3.894
R13168 fc2.n3786 fc2.t641 3.894
R13169 fc2.n3713 fc2.t657 3.894
R13170 fc2.n3750 fc2.t515 3.894
R13171 fc2.n2632 fc2.n2631 3.643
R13172 fc2.n2634 fc2.t284 3.643
R13173 fc2.n289 fc2.t76 3.643
R13174 fc2.n296 fc2.n295 3.643
R13175 fc2.n300 fc2.t240 3.643
R13176 fc2.n292 fc2.n291 3.643
R13177 fc2.n7 fc2.t209 3.643
R13178 fc2.n49 fc2.t40 3.643
R13179 fc2.n2616 fc2.t247 3.643
R13180 fc2.n2583 fc2.n2582 3.643
R13181 fc2.n2610 fc2.t36 3.643
R13182 fc2.n2585 fc2.n2584 3.643
R13183 fc2.n316 fc2.t243 3.643
R13184 fc2.n4 fc2.t327 3.643
R13185 fc2.n2655 fc2.t334 3.643
R13186 fc2.n2635 fc2.t90 3.643
R13187 fc2.n2463 fc2.t315 3.643
R13188 fc2.n2474 fc2.n2473 3.643
R13189 fc2.n2477 fc2.n2476 3.643
R13190 fc2.n2460 fc2.t115 3.643
R13191 fc2.n159 fc2.t127 3.643
R13192 fc2.n171 fc2.n170 3.643
R13193 fc2.n168 fc2.n167 3.643
R13194 fc2.n156 fc2.t290 3.643
R13195 fc2.n521 fc2.t343 3.643
R13196 fc2.n535 fc2.n534 3.643
R13197 fc2.n538 fc2.n537 3.643
R13198 fc2.n518 fc2.t141 3.643
R13199 fc2.n2061 fc2.t220 3.643
R13200 fc2.n2072 fc2.n2071 3.643
R13201 fc2.n2069 fc2.n2068 3.643
R13202 fc2.n2058 fc2.t1 3.643
R13203 fc2.n2255 fc2.t248 3.643
R13204 fc2.n2263 fc2.n2262 3.643
R13205 fc2.n2237 fc2.n2236 3.643
R13206 fc2.n2252 fc2.t37 3.643
R13207 fc2.n689 fc2.t53 3.643
R13208 fc2.n700 fc2.n699 3.643
R13209 fc2.n697 fc2.n696 3.643
R13210 fc2.n686 fc2.t217 3.643
R13211 fc2.n870 fc2.t80 3.643
R13212 fc2.n881 fc2.n880 3.643
R13213 fc2.n878 fc2.n877 3.643
R13214 fc2.n867 fc2.t244 3.643
R13215 fc2.n1746 fc2.t256 3.643
R13216 fc2.n1757 fc2.n1756 3.643
R13217 fc2.n1754 fc2.n1753 3.643
R13218 fc2.n1743 fc2.t51 3.643
R13219 fc2.n1893 fc2.t279 3.643
R13220 fc2.n1904 fc2.n1903 3.643
R13221 fc2.n1901 fc2.n1900 3.643
R13222 fc2.n1890 fc2.t78 3.643
R13223 fc2.n1119 fc2.t109 3.643
R13224 fc2.n1130 fc2.n1129 3.643
R13225 fc2.n1127 fc2.n1126 3.643
R13226 fc2.n1116 fc2.t254 3.643
R13227 fc2.n1430 fc2.t112 3.643
R13228 fc2.n1443 fc2.n1442 3.643
R13229 fc2.n1440 fc2.n1439 3.643
R13230 fc2.n1427 fc2.t232 3.643
R13231 fc2.n47 fc2.t86 3.643
R13232 fc2.n48 fc2.t289 3.643
R13233 fc2.n2730 fc2.t159 3.643
R13234 fc2.n2742 fc2.n2741 3.643
R13235 fc2.n2745 fc2.n2744 3.643
R13236 fc2.n2727 fc2.t283 3.643
R13237 fc2.n2789 fc2.t286 3.643
R13238 fc2.n41 fc2.t340 3.643
R13239 fc2.n37 fc2.t173 3.643
R13240 fc2.n2713 fc2.t5 3.643
R13241 fc2.n2720 fc2.n2719 3.643
R13242 fc2.n2723 fc2.n2722 3.643
R13243 fc2.n2716 fc2.t148 3.643
R13244 fc2.n2552 fc2.t375 3.643
R13245 fc2.n2577 fc2.n2576 3.643
R13246 fc2.n2580 fc2.n2579 3.643
R13247 fc2.n2549 fc2.t170 3.643
R13248 fc2.n247 fc2.t198 3.643
R13249 fc2.n267 fc2.n266 3.643
R13250 fc2.n270 fc2.n269 3.643
R13251 fc2.n244 fc2.t347 3.643
R13252 fc2.n357 fc2.t202 3.643
R13253 fc2.n383 fc2.n382 3.643
R13254 fc2.n380 fc2.n379 3.643
R13255 fc2.n354 fc2.t371 3.643
R13256 fc2.n2165 fc2.t108 3.643
R13257 fc2.n2162 fc2.n2161 3.643
R13258 fc2.n2159 fc2.n2158 3.643
R13259 fc2.n1990 fc2.t268 3.643
R13260 fc2.n2427 fc2.t271 3.643
R13261 fc2.n1546 fc2.t188 3.643
R13262 fc2.n1765 fc2.t389 3.643
R13263 fc2.n1784 fc2.n1783 3.643
R13264 fc2.n1787 fc2.n1786 3.643
R13265 fc2.n1762 fc2.t185 3.643
R13266 fc2.n937 fc2.t190 3.643
R13267 fc2.n960 fc2.n959 3.643
R13268 fc2.n963 fc2.n962 3.643
R13269 fc2.n934 fc2.t358 3.643
R13270 fc2.n712 fc2.t187 3.643
R13271 fc2.n731 fc2.n730 3.643
R13272 fc2.n734 fc2.n733 3.643
R13273 fc2.n709 fc2.t337 3.643
R13274 fc2.n2320 fc2.t364 3.643
R13275 fc2.n2343 fc2.n2342 3.643
R13276 fc2.n2346 fc2.n2345 3.643
R13277 fc2.n2317 fc2.t162 3.643
R13278 fc2.n2084 fc2.t339 3.643
R13279 fc2.n2103 fc2.n2102 3.643
R13280 fc2.n2106 fc2.n2105 3.643
R13281 fc2.n2081 fc2.t137 3.643
R13282 fc2.n433 fc2.t91 3.643
R13283 fc2.n459 fc2.n458 3.643
R13284 fc2.n456 fc2.n455 3.643
R13285 fc2.n430 fc2.t257 3.643
R13286 fc2.n183 fc2.t67 3.643
R13287 fc2.n203 fc2.n202 3.643
R13288 fc2.n206 fc2.n205 3.643
R13289 fc2.n180 fc2.t230 3.643
R13290 fc2.n2485 fc2.t259 3.643
R13291 fc2.n2509 fc2.n2508 3.643
R13292 fc2.n2512 fc2.n2511 3.643
R13293 fc2.n2482 fc2.t54 3.643
R13294 fc2.n2664 fc2.t275 3.643
R13295 fc2.n2675 fc2.n2674 3.643
R13296 fc2.n2678 fc2.n2677 3.643
R13297 fc2.n2661 fc2.t20 3.643
R13298 fc2.n27 fc2.t222 3.643
R13299 fc2.n24 fc2.t58 3.643
R13300 fc2.n20 fc2.t156 3.643
R13301 fc2.n18 fc2.t355 3.643
R13302 fc2.n2756 fc2.t204 3.643
R13303 fc2.n2753 fc2.n2752 3.643
R13304 fc2.n2750 fc2.n2749 3.643
R13305 fc2.n2619 fc2.t330 3.643
R13306 fc2.n2772 fc2.t386 3.643
R13307 fc2.n2779 fc2.n2778 3.643
R13308 fc2.n2782 fc2.n2781 3.643
R13309 fc2.n2769 fc2.t182 3.643
R13310 fc2.n275 fc2.t191 3.643
R13311 fc2.n283 fc2.n282 3.643
R13312 fc2.n286 fc2.n285 3.643
R13313 fc2.n278 fc2.t360 3.643
R13314 fc2.n324 fc2.t212 3.643
R13315 fc2.n337 fc2.n336 3.643
R13316 fc2.n327 fc2.n326 3.643
R13317 fc2.n330 fc2.t383 3.643
R13318 fc2.n2144 fc2.t99 3.643
R13319 fc2.n2153 fc2.n2152 3.643
R13320 fc2.n2156 fc2.n2155 3.643
R13321 fc2.n2147 fc2.t263 3.643
R13322 fc2.n2399 fc2.t123 3.643
R13323 fc2.n2417 fc2.n2416 3.643
R13324 fc2.n2420 fc2.n2419 3.643
R13325 fc2.n2402 fc2.t287 3.643
R13326 fc2.n769 fc2.t297 3.643
R13327 fc2.n780 fc2.n779 3.643
R13328 fc2.n783 fc2.n782 3.643
R13329 fc2.n772 fc2.t96 3.643
R13330 fc2.n972 fc2.t321 3.643
R13331 fc2.n990 fc2.n989 3.643
R13332 fc2.n993 fc2.n992 3.643
R13333 fc2.n975 fc2.t121 3.643
R13334 fc2.n1792 fc2.t147 3.643
R13335 fc2.n1803 fc2.n1802 3.643
R13336 fc2.n1806 fc2.n1805 3.643
R13337 fc2.n1795 fc2.t296 3.643
R13338 fc2.n1952 fc2.t151 3.643
R13339 fc2.n1968 fc2.n1967 3.643
R13340 fc2.n1971 fc2.n1970 3.643
R13341 fc2.n1955 fc2.t317 3.643
R13342 fc2.n1167 fc2.t346 3.643
R13343 fc2.n1181 fc2.n1180 3.643
R13344 fc2.n1184 fc2.n1183 3.643
R13345 fc2.n1170 fc2.t145 3.643
R13346 fc2.n1019 fc2.t111 3.643
R13347 fc2.n34 fc2.t100 3.643
R13348 fc2.n30 fc2.t300 3.643
R13349 fc2.n2689 fc2.t149 3.643
R13350 fc2.n2696 fc2.n2695 3.643
R13351 fc2.n2699 fc2.n2698 3.643
R13352 fc2.n2692 fc2.t272 3.643
R13353 fc2.n2534 fc2.t134 3.643
R13354 fc2.n2542 fc2.n2541 3.643
R13355 fc2.n2545 fc2.n2544 3.643
R13356 fc2.n2537 fc2.t298 3.643
R13357 fc2.n213 fc2.t311 3.643
R13358 fc2.n233 fc2.n232 3.643
R13359 fc2.n236 fc2.n235 3.643
R13360 fc2.n210 fc2.t110 3.643
R13361 fc2.n391 fc2.t331 3.643
R13362 fc2.n417 fc2.n416 3.643
R13363 fc2.n414 fc2.n413 3.643
R13364 fc2.n388 fc2.t131 3.643
R13365 fc2.n2117 fc2.t228 3.643
R13366 fc2.n2136 fc2.n2135 3.643
R13367 fc2.n2139 fc2.n2138 3.643
R13368 fc2.n2114 fc2.t380 3.643
R13369 fc2.n2364 fc2.t234 3.643
R13370 fc2.n2387 fc2.n2386 3.643
R13371 fc2.n2390 fc2.n2389 3.643
R13372 fc2.n2361 fc2.t18 3.643
R13373 fc2.n742 fc2.t64 3.643
R13374 fc2.n761 fc2.n760 3.643
R13375 fc2.n764 fc2.n763 3.643
R13376 fc2.n739 fc2.t226 3.643
R13377 fc2.n1000 fc2.t229 3.643
R13378 fc2.n3341 fc2.t117 3.643
R13379 fc2.n1108 fc2.t158 3.643
R13380 fc2.n1076 fc2.t322 3.643
R13381 fc2.n1472 fc2.t177 3.643
R13382 fc2.n1496 fc2.n1495 3.643
R13383 fc2.n1499 fc2.n1498 3.643
R13384 fc2.n1469 fc2.t302 3.643
R13385 fc2.n3418 fc2.t353 3.643
R13386 fc2.n1701 fc2.t196 3.643
R13387 fc2.n1674 fc2.t365 3.643
R13388 fc2.n1919 fc2.t216 3.643
R13389 fc2.n1940 fc2.n1939 3.643
R13390 fc2.n1943 fc2.n1942 3.643
R13391 fc2.n1916 fc2.t387 3.643
R13392 fc2.n1139 fc2.t11 3.643
R13393 fc2.n1159 fc2.n1158 3.643
R13394 fc2.n1162 fc2.n1161 3.643
R13395 fc2.n1136 fc2.t192 3.643
R13396 fc2.n1039 fc2.t249 3.643
R13397 fc2.n1068 fc2.n1067 3.643
R13398 fc2.n1065 fc2.n1064 3.643
R13399 fc2.n1036 fc2.t374 3.643
R13400 fc2.n3395 fc2.t57 3.643
R13401 fc2.n644 fc2.t239 3.643
R13402 fc2.n618 fc2.t27 3.643
R13403 fc2.n896 fc2.t262 3.643
R13404 fc2.n918 fc2.n917 3.643
R13405 fc2.n921 fc2.n920 3.643
R13406 fc2.n893 fc2.t60 3.643
R13407 fc2.n1714 fc2.t71 3.643
R13408 fc2.n1736 fc2.n1735 3.643
R13409 fc2.n1733 fc2.n1732 3.643
R13410 fc2.n1711 fc2.t235 3.643
R13411 fc2.n1563 fc2.t291 3.643
R13412 fc2.n1589 fc2.n1588 3.643
R13413 fc2.n1586 fc2.n1585 3.643
R13414 fc2.n1560 fc2.t88 3.643
R13415 fc2.n1193 fc2.t102 3.643
R13416 fc2.n1190 fc2.n1189 3.643
R13417 fc2.n1187 fc2.n1186 3.643
R13418 fc2.n1074 fc2.t265 3.643
R13419 fc2.n1227 fc2.t124 3.643
R13420 fc2.n1256 fc2.n1255 3.643
R13421 fc2.n1253 fc2.n1252 3.643
R13422 fc2.n1224 fc2.t246 3.643
R13423 fc2.n3381 fc2.t299 3.643
R13424 fc2.n2017 fc2.t281 3.643
R13425 fc2.n1992 fc2.t79 3.643
R13426 fc2.n2281 fc2.t304 3.643
R13427 fc2.n2304 fc2.n2303 3.643
R13428 fc2.n2278 fc2.n2277 3.643
R13429 fc2.n2275 fc2.t105 3.643
R13430 fc2.n657 fc2.t114 3.643
R13431 fc2.n679 fc2.n678 3.643
R13432 fc2.n676 fc2.n675 3.643
R13433 fc2.n654 fc2.t277 3.643
R13434 fc2.n583 fc2.t332 3.643
R13435 fc2.n609 fc2.n608 3.643
R13436 fc2.n606 fc2.n605 3.643
R13437 fc2.n580 fc2.t132 3.643
R13438 fc2.n1606 fc2.t139 3.643
R13439 fc2.n1603 fc2.n1602 3.643
R13440 fc2.n1600 fc2.n1599 3.643
R13441 fc2.n1597 fc2.t309 3.643
R13442 fc2.n1639 fc2.t163 3.643
R13443 fc2.n1665 fc2.n1664 3.643
R13444 fc2.n1662 fc2.n1661 3.643
R13445 fc2.n1636 fc2.t329 3.643
R13446 fc2.n1271 fc2.t341 3.643
R13447 fc2.n1268 fc2.n1267 3.643
R13448 fc2.n1265 fc2.n1264 3.643
R13449 fc2.n1262 fc2.t138 3.643
R13450 fc2.n1305 fc2.t366 3.643
R13451 fc2.n1334 fc2.n1333 3.643
R13452 fc2.n1331 fc2.n1330 3.643
R13453 fc2.n1302 fc2.t122 3.643
R13454 fc2.n3366 fc2.t172 3.643
R13455 fc2.n147 fc2.t252 3.643
R13456 fc2.n122 fc2.t44 3.643
R13457 fc2.n476 fc2.t270 3.643
R13458 fc2.n502 fc2.n501 3.643
R13459 fc2.n499 fc2.n498 3.643
R13460 fc2.n473 fc2.t72 3.643
R13461 fc2.n2029 fc2.t154 3.643
R13462 fc2.n2051 fc2.n2050 3.643
R13463 fc2.n2048 fc2.n2047 3.643
R13464 fc2.n2026 fc2.t320 3.643
R13465 fc2.n2208 fc2.t376 3.643
R13466 fc2.n2234 fc2.n2233 3.643
R13467 fc2.n2231 fc2.n2230 3.643
R13468 fc2.n2205 fc2.t171 3.643
R13469 fc2.n792 fc2.t180 3.643
R13470 fc2.n789 fc2.n788 3.643
R13471 fc2.n786 fc2.n785 3.643
R13472 fc2.n616 fc2.t348 3.643
R13473 fc2.n826 fc2.t203 3.643
R13474 fc2.n852 fc2.n851 3.643
R13475 fc2.n849 fc2.n848 3.643
R13476 fc2.n823 fc2.t372 3.643
R13477 fc2.n1815 fc2.t382 3.643
R13478 fc2.n1812 fc2.n1811 3.643
R13479 fc2.n1809 fc2.n1808 3.643
R13480 fc2.n1672 fc2.t179 3.643
R13481 fc2.n1849 fc2.t29 3.643
R13482 fc2.n1875 fc2.n1874 3.643
R13483 fc2.n1872 fc2.n1871 3.643
R13484 fc2.n1846 fc2.t201 3.643
R13485 fc2.n1349 fc2.t210 3.643
R13486 fc2.n1346 fc2.n1345 3.643
R13487 fc2.n1343 fc2.n1342 3.643
R13488 fc2.n1340 fc2.t381 3.643
R13489 fc2.n1383 fc2.t236 3.643
R13490 fc2.n1412 fc2.n1411 3.643
R13491 fc2.n1409 fc2.n1408 3.643
R13492 fc2.n1380 fc2.t363 3.643
R13493 fc2.n3350 fc2.t65 3.643
R13494 fc2.n3439 fc2.t306 3.643
R13495 fc2.n2622 fc2.n2621 3.643
R13496 fc2.n2748 fc2.t390 3.643
R13497 fc2.n2796 fc2.n2795 2.494
R13498 fc2.n549 fc2.n548 2.494
R13499 fc2.n2434 fc2.n2433 2.494
R13500 fc2.n1007 fc2.n1006 2.494
R13501 fc2.n1536 fc2.n1535 2.494
R13502 fc2.n1515 fc2.n1513 2.494
R13503 fc2.n3476 fc2.n3475 0.21
R13504 fc2.n3887 fc2.n3886 0.21
R13505 fc2.n3616 fc2.n3615 0.21
R13506 fc2.n3804 fc2.n3803 0.21
R13507 fc2.n3394 fc2.n3393 0.2
R13508 fc2.n106 fc2.n82 0.178
R13509 fc2.n2451 fc2.n2448 0.176
R13510 fc2.n1979 fc2.n1978 0.176
R13511 fc2.n118 fc2.n115 0.176
R13512 fc2.n3773 fc2.n3772 0.174
R13513 fc2.n1527 fc2.n1526 0.171
R13514 fc2.n3335 fc2.n3329 0.157
R13515 fc2.n3401 fc2.n3400 0.154
R13516 fc2.n1984 fc2.n1983 0.153
R13517 fc2.n3189 fc2.n3180 0.147
R13518 fc2.n366 fc2.n364 0.145
R13519 fc2.n2561 fc2.n2560 0.145
R13520 fc2.n946 fc2.n945 0.145
R13521 fc2.n2329 fc2.n2328 0.145
R13522 fc2.n442 fc2.n441 0.145
R13523 fc2.n2494 fc2.n2493 0.145
R13524 fc2.n400 fc2.n398 0.145
R13525 fc2.n2373 fc2.n2371 0.145
R13526 fc2.n2519 fc2.n2516 0.145
R13527 fc2.n2593 fc2.n2590 0.145
R13528 fc2.n1449 fc2.n1448 0.145
R13529 fc2.n1060 fc2.n1058 0.145
R13530 fc2.n904 fc2.n902 0.145
R13531 fc2.n1572 fc2.n1570 0.145
R13532 fc2.n1248 fc2.n1246 0.145
R13533 fc2.n2290 fc2.n2288 0.145
R13534 fc2.n592 fc2.n590 0.145
R13535 fc2.n1648 fc2.n1646 0.145
R13536 fc2.n1326 fc2.n1324 0.145
R13537 fc2.n485 fc2.n483 0.145
R13538 fc2.n2217 fc2.n2215 0.145
R13539 fc2.n835 fc2.n833 0.145
R13540 fc2.n1858 fc2.n1856 0.145
R13541 fc2.n1404 fc2.n1402 0.145
R13542 fc2.n251 fc2.n250 0.144
R13543 fc2.n361 fc2.n360 0.144
R13544 fc2.n2169 fc2.n2168 0.144
R13545 fc2.n1769 fc2.n1767 0.144
R13546 fc2.n941 fc2.n939 0.144
R13547 fc2.n716 fc2.n714 0.144
R13548 fc2.n2324 fc2.n2322 0.144
R13549 fc2.n2088 fc2.n2086 0.144
R13550 fc2.n437 fc2.n435 0.144
R13551 fc2.n187 fc2.n185 0.144
R13552 fc2.n395 fc2.n394 0.144
R13553 fc2.n2121 fc2.n2120 0.144
R13554 fc2.n2368 fc2.n2367 0.144
R13555 fc2.n746 fc2.n745 0.144
R13556 fc2.n217 fc2.n216 0.144
R13557 fc2.n1923 fc2.n1922 0.144
R13558 fc2.n1143 fc2.n1142 0.144
R13559 fc2.n1043 fc2.n1042 0.144
R13560 fc2.n900 fc2.n899 0.144
R13561 fc2.n1718 fc2.n1717 0.144
R13562 fc2.n1567 fc2.n1566 0.144
R13563 fc2.n1197 fc2.n1196 0.144
R13564 fc2.n1231 fc2.n1230 0.144
R13565 fc2.n2285 fc2.n2284 0.144
R13566 fc2.n661 fc2.n660 0.144
R13567 fc2.n587 fc2.n586 0.144
R13568 fc2.n1610 fc2.n1609 0.144
R13569 fc2.n1643 fc2.n1642 0.144
R13570 fc2.n1275 fc2.n1274 0.144
R13571 fc2.n1309 fc2.n1308 0.144
R13572 fc2.n470 fc2.n468 0.144
R13573 fc2.n480 fc2.n479 0.144
R13574 fc2.n2033 fc2.n2032 0.144
R13575 fc2.n2212 fc2.n2211 0.144
R13576 fc2.n796 fc2.n795 0.144
R13577 fc2.n830 fc2.n829 0.144
R13578 fc2.n1819 fc2.n1818 0.144
R13579 fc2.n1853 fc2.n1852 0.144
R13580 fc2.n1353 fc2.n1352 0.144
R13581 fc2.n1387 fc2.n1386 0.144
R13582 fc2.n3581 fc2.n3580 0.143
R13583 fc2.n3581 fc2.n3447 0.143
R13584 fc2.n3982 fc2.n3981 0.143
R13585 fc2.n3982 fc2.n3865 0.143
R13586 fc2.n3681 fc2.n3680 0.143
R13587 fc2.n3681 fc2.n3587 0.143
R13588 fc2.n3859 fc2.n3858 0.143
R13589 fc2.n3859 fc2.n3782 0.143
R13590 fc2.n3777 fc2.n3746 0.143
R13591 fc2.n3741 fc2.n3723 0.143
R13592 fc2.n3741 fc2.n3740 0.143
R13593 fc2.n3777 fc2.n3776 0.143
R13594 fc2.n3779 fc2.n3778 0.142
R13595 fc2.n2962 fc2.n2961 0.141
R13596 fc2.n3876 fc2.n3866 0.14
R13597 fc2.n3793 fc2.n3783 0.14
R13598 fc2.n1521 fc2.n1518 0.136
R13599 fc2.n3775 fc2.n3773 0.133
R13600 fc2.n3765 fc2.n3763 0.126
R13601 fc2.n3305 fc2.n3304 0.125
R13602 fc2.n3984 fc2.n3983 0.123
R13603 fc2.n3861 fc2.n3860 0.123
R13604 fc2.n1482 fc2.n1478 0.122
R13605 fc2.n1029 fc2.n1028 0.122
R13606 fc2.n3444 fc2.n3443 0.119
R13607 fc2.n85 fc2.n84 0.119
R13608 fc2.n2793 fc2.n2792 0.119
R13609 fc2.n546 fc2.n545 0.119
R13610 fc2.n2431 fc2.n2430 0.119
R13611 fc2.n1004 fc2.n1003 0.119
R13612 fc2.n1544 fc2.n1533 0.119
R13613 fc2.n2807 fc2.n109 0.117
R13614 fc2.n3464 fc2.n3456 0.115
R13615 fc2.n3874 fc2.n3873 0.115
R13616 fc2.n3604 fc2.n3596 0.115
R13617 fc2.n3791 fc2.n3790 0.115
R13618 fc2.n3719 fc2.n3718 0.115
R13619 fc2.n2807 fc2.n1531 0.115
R13620 fc2.n2807 fc2.n1987 0.115
R13621 fc2.n1461 fc2.n1460 0.115
R13622 fc2.n3308 fc2.n3174 0.113
R13623 fc2.n3308 fc2.n3063 0.113
R13624 fc2.n3308 fc2.n2949 0.113
R13625 fc2.n3308 fc2.n2898 0.113
R13626 fc2.n3969 fc2.n3960 0.113
R13627 fc2.n3846 fc2.n3837 0.113
R13628 fc2.n3308 fc2.n2992 0.113
R13629 fc2.n3308 fc2.n2960 0.113
R13630 fc2.n2807 fc2.n1017 0.111
R13631 fc2.n2807 fc2.n2444 0.111
R13632 fc2.n2807 fc2.n2806 0.111
R13633 fc2.n2807 fc2.n559 0.11
R13634 fc2.n3759 fc2.n3758 0.109
R13635 fc2.n3585 fc2.n3584 0.108
R13636 fc2.n3685 fc2.n3684 0.108
R13637 fc2.n3745 fc2.n3744 0.108
R13638 fc2.n1912 fc2.n1907 0.108
R13639 fc2.n889 fc2.n884 0.108
R13640 fc2.n2271 fc2.n2266 0.108
R13641 fc2.n467 fc2.n461 0.108
R13642 fc2.n1486 fc2.n1485 0.107
R13643 fc2.n3422 fc2.n3421 0.107
R13644 fc2.n3781 fc2.n3780 0.105
R13645 fc2.n3987 fc2.n3986 0.105
R13646 fc2.n3864 fc2.n3863 0.105
R13647 fc2.n3417 fc2.n3416 0.105
R13648 fc2.n3423 fc2.n3422 0.105
R13649 fc2.n3406 fc2.n3405 0.105
R13650 fc2.n3389 fc2.n3388 0.105
R13651 fc2.n3377 fc2.n3376 0.105
R13652 fc2.n3362 fc2.n3361 0.105
R13653 fc2.n3985 fc2.n3585 0.105
R13654 fc2.n3862 fc2.n3685 0.105
R13655 fc2.n3779 fc2.n3745 0.105
R13656 fc2.n3752 fc2.n3751 0.102
R13657 fc2.n1083 fc2.n1078 0.101
R13658 fc2.n1681 fc2.n1676 0.101
R13659 fc2.n624 fc2.n620 0.101
R13660 fc2.n1997 fc2.n1994 0.101
R13661 fc2.n127 fc2.n124 0.101
R13662 fc2.n2650 fc2.n2647 0.101
R13663 fc2.n1032 fc2.n1031 0.101
R13664 fc2.n1693 fc2.n1692 0.101
R13665 fc2.n636 fc2.n635 0.101
R13666 fc2.n2009 fc2.n2008 0.101
R13667 fc2.n139 fc2.n138 0.101
R13668 fc2.n3583 fc2.n3582 0.1
R13669 fc2.n3683 fc2.n3682 0.1
R13670 fc2.n3743 fc2.n3742 0.1
R13671 fc2.n262 fc2.n259 0.096
R13672 fc2.n375 fc2.n370 0.096
R13673 fc2.n2179 fc2.n2176 0.096
R13674 fc2.n1779 fc2.n1778 0.096
R13675 fc2.n955 fc2.n954 0.096
R13676 fc2.n726 fc2.n725 0.096
R13677 fc2.n2338 fc2.n2337 0.096
R13678 fc2.n2098 fc2.n2097 0.096
R13679 fc2.n451 fc2.n450 0.096
R13680 fc2.n198 fc2.n197 0.096
R13681 fc2.n227 fc2.n224 0.096
R13682 fc2.n409 fc2.n404 0.096
R13683 fc2.n2131 fc2.n2128 0.096
R13684 fc2.n2382 fc2.n2377 0.096
R13685 fc2.n756 fc2.n753 0.096
R13686 fc2.n2527 fc2.n2522 0.096
R13687 fc2.n2601 fc2.n2596 0.096
R13688 fc2.n1935 fc2.n1930 0.096
R13689 fc2.n1154 fc2.n1150 0.096
R13690 fc2.n913 fc2.n908 0.096
R13691 fc2.n1728 fc2.n1725 0.096
R13692 fc2.n1581 fc2.n1576 0.096
R13693 fc2.n1208 fc2.n1204 0.096
R13694 fc2.n2299 fc2.n2294 0.096
R13695 fc2.n671 fc2.n668 0.096
R13696 fc2.n601 fc2.n596 0.096
R13697 fc2.n1620 fc2.n1617 0.096
R13698 fc2.n1657 fc2.n1652 0.096
R13699 fc2.n1286 fc2.n1282 0.096
R13700 fc2.n494 fc2.n489 0.096
R13701 fc2.n2043 fc2.n2040 0.096
R13702 fc2.n2226 fc2.n2221 0.096
R13703 fc2.n806 fc2.n803 0.096
R13704 fc2.n844 fc2.n839 0.096
R13705 fc2.n1829 fc2.n1826 0.096
R13706 fc2.n1867 fc2.n1862 0.096
R13707 fc2.n1364 fc2.n1360 0.096
R13708 fc2.n2737 fc2.n2734 0.096
R13709 fc2.n307 fc2.n306 0.096
R13710 fc2.n2571 fc2.n2565 0.095
R13711 fc2.n2707 fc2.n2704 0.095
R13712 fc2.n2504 fc2.n2503 0.095
R13713 fc2.n1483 fc2.n1476 0.095
R13714 fc2.n1100 fc2.n1095 0.093
R13715 fc2.n1053 fc2.n1051 0.092
R13716 fc2.n1241 fc2.n1239 0.092
R13717 fc2.n1319 fc2.n1317 0.092
R13718 fc2.n1397 fc2.n1395 0.092
R13719 fc2.n2671 fc2.n2670 0.091
R13720 fc2.n2685 fc2.n2682 0.091
R13721 fc2.n2628 fc2.n2625 0.091
R13722 fc2.n3417 fc2.n3415 0.089
R13723 fc2.n3406 fc2.n3404 0.089
R13724 fc2.n3389 fc2.n3387 0.089
R13725 fc2.n3377 fc2.n3375 0.089
R13726 fc2.n3362 fc2.n3360 0.089
R13727 fc2.n1462 fc2.n1453 0.087
R13728 fc2.n1507 fc2.n1506 0.086
R13729 fc2.n2569 fc2.n2568 0.085
R13730 fc2.n2499 fc2.n2498 0.085
R13731 fc2.n3308 fc2.n3307 0.085
R13732 fc2.n1098 fc2.n1097 0.085
R13733 fc2.n1488 fc2.n1474 0.084
R13734 fc2.n3438 fc2.n3437 0.084
R13735 fc2.n2471 fc2.n2469 0.083
R13736 fc2.n3414 fc2.n3413 0.082
R13737 fc2.n3412 fc2.n3411 0.082
R13738 fc2.n3399 fc2.n3398 0.082
R13739 fc2.n3385 fc2.n3384 0.082
R13740 fc2.n3372 fc2.n3369 0.082
R13741 fc2.n3356 fc2.n3353 0.082
R13742 fc2.n1023 fc2.n1022 0.082
R13743 fc2.n2804 fc2.n2803 0.081
R13744 fc2.n557 fc2.n556 0.081
R13745 fc2.n2442 fc2.n2441 0.081
R13746 fc2.n1015 fc2.n1014 0.081
R13747 fc2.n1544 fc2.n1543 0.081
R13748 fc2.n1527 fc2.n1525 0.081
R13749 fc2.n1447 fc2.n1446 0.08
R13750 fc2.n1487 fc2.n1486 0.08
R13751 fc2.n15 fc2.n13 0.08
R13752 fc2.n2990 fc2.n2989 0.079
R13753 fc2.n3082 fc2.n3081 0.079
R13754 fc2.n3011 fc2.n3010 0.079
R13755 fc2.n2917 fc2.n2916 0.079
R13756 fc2.n2826 fc2.n2825 0.079
R13757 fc2.n74 fc2.n73 0.078
R13758 fc2.n104 fc2.n102 0.078
R13759 fc2.n3700 fc2.n3699 0.078
R13760 fc2.n3468 fc2.n3467 0.078
R13761 fc2.n3889 fc2.n3876 0.078
R13762 fc2.n3608 fc2.n3607 0.078
R13763 fc2.n3806 fc2.n3793 0.078
R13764 fc2.n2960 fc2.n2959 0.077
R13765 fc2.n3458 fc2.n3457 0.077
R13766 fc2.n3463 fc2.n3462 0.077
R13767 fc2.n3868 fc2.n3867 0.077
R13768 fc2.n3598 fc2.n3597 0.077
R13769 fc2.n3603 fc2.n3602 0.077
R13770 fc2.n3785 fc2.n3784 0.077
R13771 fc2.n3715 fc2.n3714 0.077
R13772 fc2.n3710 fc2.n3709 0.077
R13773 fc2.n1104 fc2.n1103 0.075
R13774 fc2.n349 fc2.n346 0.075
R13775 fc2.n425 fc2.n424 0.075
R13776 fc2.n2312 fc2.n2311 0.075
R13777 fc2.n929 fc2.n928 0.075
R13778 fc2.n980 fc2.n977 0.075
R13779 fc2.n2407 fc2.n2404 0.075
R13780 fc2.n2356 fc2.n2353 0.075
R13781 fc2.n1555 fc2.n1553 0.075
R13782 fc2.n1631 fc2.n1629 0.075
R13783 fc2.n575 fc2.n573 0.075
R13784 fc2.n1841 fc2.n1838 0.075
R13785 fc2.n818 fc2.n815 0.075
R13786 fc2.n2200 fc2.n2197 0.075
R13787 fc2.n1422 fc2.n1419 0.075
R13788 fc2.n1885 fc2.n1882 0.075
R13789 fc2.n862 fc2.n859 0.075
R13790 fc2.n2247 fc2.n2244 0.075
R13791 fc2.n513 fc2.n510 0.075
R13792 fc2.n1912 fc2.n1910 0.075
R13793 fc2.n889 fc2.n887 0.075
R13794 fc2.n2271 fc2.n2269 0.075
R13795 fc2.n467 fc2.n465 0.075
R13796 fc2.n1697 fc2.n1696 0.074
R13797 fc2.n640 fc2.n639 0.074
R13798 fc2.n2013 fc2.n2012 0.074
R13799 fc2.n143 fc2.n142 0.074
R13800 fc2.n1092 fc2.n1091 0.074
R13801 fc2.n1690 fc2.n1689 0.074
R13802 fc2.n633 fc2.n632 0.074
R13803 fc2.n2006 fc2.n2005 0.074
R13804 fc2.n136 fc2.n135 0.074
R13805 fc2.n1982 fc2.n1981 0.074
R13806 fc2.n3171 fc2.n3170 0.074
R13807 fc2.n3160 fc2.n3150 0.074
R13808 fc2.n3140 fc2.n3130 0.074
R13809 fc2.n3120 fc2.n3110 0.074
R13810 fc2.n3060 fc2.n3059 0.074
R13811 fc2.n3049 fc2.n3039 0.074
R13812 fc2.n2946 fc2.n2945 0.074
R13813 fc2.n2895 fc2.n2894 0.074
R13814 fc2.n2884 fc2.n2874 0.074
R13815 fc2.n2864 fc2.n2854 0.074
R13816 fc2.n2645 fc2.n2644 0.073
R13817 fc2.n3410 fc2.n3409 0.073
R13818 fc2.n100 fc2.n87 0.073
R13819 fc2.n71 fc2.n58 0.073
R13820 fc2.n3977 fc2.n3976 0.073
R13821 fc2.n3965 fc2.n3964 0.073
R13822 fc2.n96 fc2.n89 0.073
R13823 fc2.n67 fc2.n60 0.073
R13824 fc2.n3854 fc2.n3853 0.073
R13825 fc2.n3842 fc2.n3841 0.073
R13826 fc2.n63 fc2.n62 0.073
R13827 fc2.n92 fc2.n91 0.073
R13828 fc2.n3198 fc2.n3197 0.072
R13829 fc2.n3899 fc2.n3889 0.072
R13830 fc2.n3816 fc2.n3806 0.072
R13831 fc2.n3100 fc2.n3090 0.072
R13832 fc2.n3029 fc2.n3019 0.072
R13833 fc2.n2935 fc2.n2925 0.072
R13834 fc2.n2844 fc2.n2834 0.072
R13835 fc2.n3909 fc2.n3899 0.072
R13836 fc2.n3919 fc2.n3909 0.072
R13837 fc2.n3929 fc2.n3919 0.072
R13838 fc2.n3939 fc2.n3929 0.072
R13839 fc2.n3949 fc2.n3939 0.072
R13840 fc2.n3959 fc2.n3949 0.072
R13841 fc2.n3826 fc2.n3816 0.072
R13842 fc2.n3836 fc2.n3826 0.072
R13843 fc2.n3210 fc2.n3200 0.072
R13844 fc2.n3220 fc2.n3210 0.072
R13845 fc2.n3230 fc2.n3220 0.072
R13846 fc2.n3240 fc2.n3230 0.072
R13847 fc2.n3250 fc2.n3240 0.072
R13848 fc2.n3260 fc2.n3250 0.072
R13849 fc2.n3270 fc2.n3260 0.072
R13850 fc2.n3280 fc2.n3270 0.072
R13851 fc2.n3290 fc2.n3280 0.072
R13852 fc2.n3300 fc2.n3290 0.072
R13853 fc2.n3200 fc2.n3189 0.072
R13854 fc2.n3130 fc2.n3120 0.072
R13855 fc2.n3150 fc2.n3140 0.072
R13856 fc2.n3170 fc2.n3160 0.072
R13857 fc2.n3110 fc2.n3100 0.072
R13858 fc2.n3059 fc2.n3049 0.072
R13859 fc2.n3039 fc2.n3029 0.072
R13860 fc2.n2945 fc2.n2935 0.072
R13861 fc2.n2874 fc2.n2864 0.072
R13862 fc2.n2894 fc2.n2884 0.072
R13863 fc2.n2854 fc2.n2844 0.072
R13864 fc2.n3328 fc2.n3327 0.07
R13865 fc2.n3321 fc2.n3320 0.07
R13866 fc2.n3374 fc2.n3373 0.068
R13867 fc2.n2451 fc2.n2450 0.068
R13868 fc2.n2189 fc2.n2188 0.068
R13869 fc2.n565 fc2.n564 0.068
R13870 fc2.n118 fc2.n117 0.068
R13871 fc2.n106 fc2.n105 0.067
R13872 fc2.n106 fc2.n75 0.067
R13873 fc2.n3337 fc2.n3336 0.067
R13874 fc2.n43 fc2.n42 0.067
R13875 fc2.n36 fc2.n35 0.067
R13876 fc2.n3359 fc2.n3358 0.066
R13877 fc2.n3437 fc2.n3436 0.066
R13878 fc2.n558 fc2.n557 0.065
R13879 fc2.n2805 fc2.n2804 0.065
R13880 fc2.n2443 fc2.n2442 0.065
R13881 fc2.n1016 fc2.n1015 0.065
R13882 fc2.n22 fc2.n21 0.064
R13883 fc2.n112 fc2.n111 0.063
R13884 fc2.n1545 fc2.n1544 0.063
R13885 fc2.n1457 fc2.n1456 0.062
R13886 fc2.n3372 fc2.n3371 0.062
R13887 fc2.n3356 fc2.n3355 0.062
R13888 fc2.n2557 fc2.n2556 0.061
R13889 fc2.n254 fc2.n253 0.061
R13890 fc2.n190 fc2.n189 0.061
R13891 fc2.n2490 fc2.n2489 0.061
R13892 fc2.n2518 fc2.n2517 0.061
R13893 fc2.n2592 fc2.n2591 0.061
R13894 fc2.n3991 fc2.n3990 0.061
R13895 fc2.n3301 fc2.n3300 0.061
R13896 fc2.n2466 fc2.n2465 0.06
R13897 fc2.n1466 fc2.n1465 0.06
R13898 fc2.n3174 fc2.n3173 0.06
R13899 fc2.n3063 fc2.n3062 0.06
R13900 fc2.n2949 fc2.n2948 0.06
R13901 fc2.n2898 fc2.n2897 0.06
R13902 fc2.n1528 fc2.n1527 0.058
R13903 fc2.n3306 fc2.n3305 0.056
R13904 fc2.n3340 fc2.n3314 0.056
R13905 fc2.n53 fc2.n4 0.055
R13906 fc2.n2788 fc2.n2787 0.055
R13907 fc2.n2426 fc2.n2425 0.055
R13908 fc2.n1974 fc2.n1973 0.055
R13909 fc2.n1502 fc2.n1501 0.055
R13910 fc2.n999 fc2.n998 0.055
R13911 fc2.n542 fc2.n316 0.054
R13912 fc2.n2653 fc2.n2635 0.054
R13913 fc2.n1106 fc2.n1076 0.054
R13914 fc2.n1699 fc2.n1674 0.054
R13915 fc2.n642 fc2.n618 0.054
R13916 fc2.n2015 fc2.n1992 0.054
R13917 fc2.n145 fc2.n122 0.054
R13918 fc2.n2776 fc2.n2775 0.054
R13919 fc2.n1177 fc2.n1176 0.054
R13920 fc2.n1494 fc2.n1493 0.054
R13921 fc2.n3763 fc2.n3762 0.054
R13922 fc2.n2478 fc2.n2477 0.054
R13923 fc2.n169 fc2.n168 0.054
R13924 fc2.n539 fc2.n538 0.054
R13925 fc2.n2070 fc2.n2069 0.054
R13926 fc2.n2238 fc2.n2237 0.054
R13927 fc2.n698 fc2.n697 0.054
R13928 fc2.n879 fc2.n878 0.054
R13929 fc2.n1755 fc2.n1754 0.054
R13930 fc2.n1902 fc2.n1901 0.054
R13931 fc2.n1128 fc2.n1127 0.054
R13932 fc2.n1441 fc2.n1440 0.054
R13933 fc2.n2746 fc2.n2745 0.054
R13934 fc2.n2724 fc2.n2723 0.054
R13935 fc2.n2581 fc2.n2580 0.054
R13936 fc2.n271 fc2.n270 0.054
R13937 fc2.n381 fc2.n380 0.054
R13938 fc2.n2160 fc2.n2159 0.054
R13939 fc2.n1788 fc2.n1787 0.054
R13940 fc2.n964 fc2.n963 0.054
R13941 fc2.n735 fc2.n734 0.054
R13942 fc2.n2347 fc2.n2346 0.054
R13943 fc2.n2107 fc2.n2106 0.054
R13944 fc2.n457 fc2.n456 0.054
R13945 fc2.n207 fc2.n206 0.054
R13946 fc2.n2513 fc2.n2512 0.054
R13947 fc2.n2679 fc2.n2678 0.054
R13948 fc2.n2751 fc2.n2750 0.054
R13949 fc2.n2783 fc2.n2782 0.054
R13950 fc2.n287 fc2.n286 0.054
R13951 fc2.n328 fc2.n327 0.054
R13952 fc2.n2157 fc2.n2156 0.054
R13953 fc2.n2421 fc2.n2420 0.054
R13954 fc2.n784 fc2.n783 0.054
R13955 fc2.n994 fc2.n993 0.054
R13956 fc2.n1807 fc2.n1806 0.054
R13957 fc2.n1972 fc2.n1971 0.054
R13958 fc2.n1185 fc2.n1184 0.054
R13959 fc2.n2700 fc2.n2699 0.054
R13960 fc2.n2546 fc2.n2545 0.054
R13961 fc2.n237 fc2.n236 0.054
R13962 fc2.n415 fc2.n414 0.054
R13963 fc2.n2140 fc2.n2139 0.054
R13964 fc2.n2391 fc2.n2390 0.054
R13965 fc2.n765 fc2.n764 0.054
R13966 fc2.n1500 fc2.n1499 0.054
R13967 fc2.n1944 fc2.n1943 0.054
R13968 fc2.n1163 fc2.n1162 0.054
R13969 fc2.n1066 fc2.n1065 0.054
R13970 fc2.n922 fc2.n921 0.054
R13971 fc2.n1734 fc2.n1733 0.054
R13972 fc2.n1587 fc2.n1586 0.054
R13973 fc2.n1188 fc2.n1187 0.054
R13974 fc2.n1254 fc2.n1253 0.054
R13975 fc2.n2279 fc2.n2278 0.054
R13976 fc2.n677 fc2.n676 0.054
R13977 fc2.n607 fc2.n606 0.054
R13978 fc2.n1601 fc2.n1600 0.054
R13979 fc2.n1663 fc2.n1662 0.054
R13980 fc2.n1266 fc2.n1265 0.054
R13981 fc2.n1332 fc2.n1331 0.054
R13982 fc2.n500 fc2.n499 0.054
R13983 fc2.n2049 fc2.n2048 0.054
R13984 fc2.n2232 fc2.n2231 0.054
R13985 fc2.n787 fc2.n786 0.054
R13986 fc2.n850 fc2.n849 0.054
R13987 fc2.n1810 fc2.n1809 0.054
R13988 fc2.n1873 fc2.n1872 0.054
R13989 fc2.n1344 fc2.n1343 0.054
R13990 fc2.n1410 fc2.n1409 0.054
R13991 fc2.n1435 fc2.n1434 0.054
R13992 fc2.n3765 fc2.n3764 0.053
R13993 fc2.n3775 fc2.n3774 0.053
R13994 fc2.n2643 fc2.n2642 0.053
R13995 fc2.n134 fc2.n133 0.053
R13996 fc2.n2004 fc2.n2003 0.053
R13997 fc2.n631 fc2.n630 0.053
R13998 fc2.n1688 fc2.n1687 0.053
R13999 fc2.n1090 fc2.n1089 0.053
R14000 fc2.n15 fc2.n14 0.053
R14001 fc2.n12 fc2.n11 0.053
R14002 fc2.n3445 fc2.n3444 0.053
R14003 fc2.n3560 fc2.n3559 0.053
R14004 fc2.n3960 fc2.n3959 0.053
R14005 fc2.n3660 fc2.n3659 0.053
R14006 fc2.n3837 fc2.n3836 0.053
R14007 fc2.n3695 fc2.n3694 0.053
R14008 fc2.n2469 fc2.n2468 0.052
R14009 fc2.t4 fc2.n2622 0.052
R14010 fc2.n3297 fc2.n3296 0.052
R14011 fc2.n3287 fc2.n3286 0.052
R14012 fc2.n3277 fc2.n3276 0.052
R14013 fc2.n3267 fc2.n3266 0.052
R14014 fc2.n3257 fc2.n3256 0.052
R14015 fc2.n3247 fc2.n3246 0.052
R14016 fc2.n3237 fc2.n3236 0.052
R14017 fc2.n3227 fc2.n3226 0.052
R14018 fc2.n3217 fc2.n3216 0.052
R14019 fc2.n3207 fc2.n3206 0.052
R14020 fc2.n3196 fc2.n3195 0.052
R14021 fc2.n3187 fc2.n3186 0.052
R14022 fc2.n3088 fc2.n3087 0.052
R14023 fc2.n3098 fc2.n3097 0.052
R14024 fc2.n3118 fc2.n3117 0.052
R14025 fc2.n3138 fc2.n3137 0.052
R14026 fc2.n3158 fc2.n3157 0.052
R14027 fc2.n3076 fc2.n3075 0.052
R14028 fc2.n3167 fc2.n3166 0.052
R14029 fc2.n3147 fc2.n3146 0.052
R14030 fc2.n3127 fc2.n3126 0.052
R14031 fc2.n3107 fc2.n3106 0.052
R14032 fc2.n3017 fc2.n3016 0.052
R14033 fc2.n3027 fc2.n3026 0.052
R14034 fc2.n3047 fc2.n3046 0.052
R14035 fc2.n3005 fc2.n3004 0.052
R14036 fc2.n3056 fc2.n3055 0.052
R14037 fc2.n3036 fc2.n3035 0.052
R14038 fc2.n2983 fc2.n2982 0.052
R14039 fc2.n2974 fc2.n2973 0.052
R14040 fc2.n2923 fc2.n2922 0.052
R14041 fc2.n2933 fc2.n2932 0.052
R14042 fc2.n2911 fc2.n2910 0.052
R14043 fc2.n2942 fc2.n2941 0.052
R14044 fc2.n2832 fc2.n2831 0.052
R14045 fc2.n2842 fc2.n2841 0.052
R14046 fc2.n2862 fc2.n2861 0.052
R14047 fc2.n2882 fc2.n2881 0.052
R14048 fc2.n2820 fc2.n2819 0.052
R14049 fc2.n2891 fc2.n2890 0.052
R14050 fc2.n2871 fc2.n2870 0.052
R14051 fc2.n2851 fc2.n2850 0.052
R14052 fc2.n3693 fc2.n3692 0.052
R14053 fc2.n3566 fc2.n3565 0.052
R14054 fc2.n3555 fc2.n3554 0.052
R14055 fc2.n3545 fc2.n3544 0.052
R14056 fc2.n3535 fc2.n3534 0.052
R14057 fc2.n3525 fc2.n3524 0.052
R14058 fc2.n3515 fc2.n3514 0.052
R14059 fc2.n3505 fc2.n3504 0.052
R14060 fc2.n3495 fc2.n3494 0.052
R14061 fc2.n3485 fc2.n3484 0.052
R14062 fc2.n3474 fc2.n3473 0.052
R14063 fc2.n3956 fc2.n3955 0.052
R14064 fc2.n3946 fc2.n3945 0.052
R14065 fc2.n3936 fc2.n3935 0.052
R14066 fc2.n3926 fc2.n3925 0.052
R14067 fc2.n3916 fc2.n3915 0.052
R14068 fc2.n3906 fc2.n3905 0.052
R14069 fc2.n3896 fc2.n3895 0.052
R14070 fc2.n3883 fc2.n3882 0.052
R14071 fc2.n3666 fc2.n3665 0.052
R14072 fc2.n3655 fc2.n3654 0.052
R14073 fc2.n3645 fc2.n3644 0.052
R14074 fc2.n3635 fc2.n3634 0.052
R14075 fc2.n3625 fc2.n3624 0.052
R14076 fc2.n3614 fc2.n3613 0.052
R14077 fc2.n3833 fc2.n3832 0.052
R14078 fc2.n3823 fc2.n3822 0.052
R14079 fc2.n3813 fc2.n3812 0.052
R14080 fc2.n3800 fc2.n3799 0.052
R14081 fc2.n3706 fc2.n3705 0.052
R14082 fc2.n29 fc2.n28 0.052
R14083 fc2.n52 fc2.n51 0.052
R14084 fc2.n108 fc2.n56 0.052
R14085 fc2.t4 fc2.n2748 0.051
R14086 fc2.n3294 fc2.n3293 0.051
R14087 fc2.n3284 fc2.n3283 0.051
R14088 fc2.n3274 fc2.n3273 0.051
R14089 fc2.n3264 fc2.n3263 0.051
R14090 fc2.n3254 fc2.n3253 0.051
R14091 fc2.n3244 fc2.n3243 0.051
R14092 fc2.n3234 fc2.n3233 0.051
R14093 fc2.n3224 fc2.n3223 0.051
R14094 fc2.n3214 fc2.n3213 0.051
R14095 fc2.n3204 fc2.n3203 0.051
R14096 fc2.n3193 fc2.n3192 0.051
R14097 fc2.n3184 fc2.n3183 0.051
R14098 fc2.n3085 fc2.n3083 0.051
R14099 fc2.n3095 fc2.n3093 0.051
R14100 fc2.n3115 fc2.n3113 0.051
R14101 fc2.n3135 fc2.n3133 0.051
R14102 fc2.n3155 fc2.n3153 0.051
R14103 fc2.n3073 fc2.n3071 0.051
R14104 fc2.n3164 fc2.n3163 0.051
R14105 fc2.n3144 fc2.n3143 0.051
R14106 fc2.n3124 fc2.n3123 0.051
R14107 fc2.n3104 fc2.n3103 0.051
R14108 fc2.n3014 fc2.n3012 0.051
R14109 fc2.n3024 fc2.n3022 0.051
R14110 fc2.n3044 fc2.n3042 0.051
R14111 fc2.n3002 fc2.n3000 0.051
R14112 fc2.n3053 fc2.n3052 0.051
R14113 fc2.n3033 fc2.n3032 0.051
R14114 fc2.n2980 fc2.n2978 0.051
R14115 fc2.n2971 fc2.n2969 0.051
R14116 fc2.n2920 fc2.n2918 0.051
R14117 fc2.n2930 fc2.n2928 0.051
R14118 fc2.n2908 fc2.n2906 0.051
R14119 fc2.n2939 fc2.n2938 0.051
R14120 fc2.n2829 fc2.n2827 0.051
R14121 fc2.n2839 fc2.n2837 0.051
R14122 fc2.n2859 fc2.n2857 0.051
R14123 fc2.n2879 fc2.n2877 0.051
R14124 fc2.n2817 fc2.n2815 0.051
R14125 fc2.n2888 fc2.n2887 0.051
R14126 fc2.n2868 fc2.n2867 0.051
R14127 fc2.n2848 fc2.n2847 0.051
R14128 fc2.n3690 fc2.n3688 0.051
R14129 fc2.n3563 fc2.n3562 0.051
R14130 fc2.n3552 fc2.n3551 0.051
R14131 fc2.n3542 fc2.n3541 0.051
R14132 fc2.n3532 fc2.n3531 0.051
R14133 fc2.n3522 fc2.n3521 0.051
R14134 fc2.n3512 fc2.n3511 0.051
R14135 fc2.n3502 fc2.n3501 0.051
R14136 fc2.n3492 fc2.n3491 0.051
R14137 fc2.n3482 fc2.n3481 0.051
R14138 fc2.n3471 fc2.n3470 0.051
R14139 fc2.n3953 fc2.n3952 0.051
R14140 fc2.n3943 fc2.n3942 0.051
R14141 fc2.n3933 fc2.n3932 0.051
R14142 fc2.n3923 fc2.n3922 0.051
R14143 fc2.n3913 fc2.n3912 0.051
R14144 fc2.n3903 fc2.n3902 0.051
R14145 fc2.n3893 fc2.n3892 0.051
R14146 fc2.n3880 fc2.n3879 0.051
R14147 fc2.n3663 fc2.n3662 0.051
R14148 fc2.n3652 fc2.n3651 0.051
R14149 fc2.n3642 fc2.n3641 0.051
R14150 fc2.n3632 fc2.n3631 0.051
R14151 fc2.n3622 fc2.n3621 0.051
R14152 fc2.n3611 fc2.n3610 0.051
R14153 fc2.n3830 fc2.n3829 0.051
R14154 fc2.n3820 fc2.n3819 0.051
R14155 fc2.n3810 fc2.n3809 0.051
R14156 fc2.n3797 fc2.n3796 0.051
R14157 fc2.n3703 fc2.n3702 0.051
R14158 fc2.n3762 fc2.n3761 0.051
R14159 fc2.n3069 fc2.n3065 0.05
R14160 fc2.n2998 fc2.n2994 0.05
R14161 fc2.n2967 fc2.n2965 0.05
R14162 fc2.n2955 fc2.n2952 0.05
R14163 fc2.n2904 fc2.n2900 0.05
R14164 fc2.n2813 fc2.n2809 0.05
R14165 fc2.n3464 fc2.n3459 0.05
R14166 fc2.n3873 fc2.n3869 0.05
R14167 fc2.n3604 fc2.n3599 0.05
R14168 fc2.n3790 fc2.n3786 0.05
R14169 fc2.n3719 fc2.n3713 0.05
R14170 fc2.n3755 fc2.n3750 0.05
R14171 fc2.n302 fc2.n301 0.05
R14172 fc2.n2612 fc2.n2611 0.05
R14173 fc2.n3569 fc2.n3558 0.049
R14174 fc2.n3558 fc2.n3548 0.049
R14175 fc2.n3548 fc2.n3538 0.049
R14176 fc2.n3538 fc2.n3528 0.049
R14177 fc2.n3528 fc2.n3518 0.049
R14178 fc2.n3518 fc2.n3508 0.049
R14179 fc2.n3508 fc2.n3498 0.049
R14180 fc2.n3498 fc2.n3488 0.049
R14181 fc2.n3488 fc2.n3478 0.049
R14182 fc2.n3669 fc2.n3658 0.049
R14183 fc2.n3658 fc2.n3648 0.049
R14184 fc2.n3648 fc2.n3638 0.049
R14185 fc2.n3638 fc2.n3628 0.049
R14186 fc2.n3628 fc2.n3618 0.049
R14187 fc2.n2991 fc2.n2990 0.049
R14188 fc2.n3721 fc2.n3720 0.049
R14189 fc2.n1460 fc2.n1459 0.048
R14190 fc2.n56 fc2.n55 0.048
R14191 fc2.n107 fc2.n106 0.048
R14192 fc2.n2992 fc2.n2991 0.047
R14193 fc2.n2565 fc2.n2564 0.047
R14194 fc2.n2704 fc2.n2703 0.047
R14195 fc2.n2503 fc2.n2502 0.047
R14196 fc2.n2670 fc2.n2669 0.047
R14197 fc2.n2682 fc2.n2681 0.047
R14198 fc2.n2625 fc2.n2624 0.047
R14199 fc2.n1453 fc2.n1452 0.047
R14200 fc2.n1095 fc2.n1094 0.047
R14201 fc2.n2472 fc2.n2461 0.047
R14202 fc2.n166 fc2.n157 0.047
R14203 fc2.n533 fc2.n519 0.047
R14204 fc2.n2067 fc2.n2059 0.047
R14205 fc2.n2261 fc2.n2253 0.047
R14206 fc2.n695 fc2.n687 0.047
R14207 fc2.n876 fc2.n868 0.047
R14208 fc2.n1752 fc2.n1744 0.047
R14209 fc2.n1899 fc2.n1891 0.047
R14210 fc2.n1125 fc2.n1117 0.047
R14211 fc2.n1438 fc2.n1428 0.047
R14212 fc2.n2740 fc2.n2728 0.047
R14213 fc2.n2806 fc2.n2790 0.047
R14214 fc2.n2718 fc2.n2717 0.047
R14215 fc2.n2575 fc2.n2550 0.047
R14216 fc2.n265 fc2.n245 0.047
R14217 fc2.n378 fc2.n355 0.047
R14218 fc2.n2182 fc2.n1991 0.047
R14219 fc2.n2444 fc2.n2428 0.047
R14220 fc2.n1986 fc2.n1547 0.047
R14221 fc2.n1782 fc2.n1763 0.047
R14222 fc2.n958 fc2.n935 0.047
R14223 fc2.n729 fc2.n710 0.047
R14224 fc2.n2341 fc2.n2318 0.047
R14225 fc2.n2101 fc2.n2082 0.047
R14226 fc2.n454 fc2.n431 0.047
R14227 fc2.n201 fc2.n181 0.047
R14228 fc2.n2507 fc2.n2483 0.047
R14229 fc2.n2673 fc2.n2662 0.047
R14230 fc2.n2766 fc2.n2620 0.047
R14231 fc2.n2777 fc2.n2770 0.047
R14232 fc2.n281 fc2.n279 0.047
R14233 fc2.n335 fc2.n331 0.047
R14234 fc2.n2151 fc2.n2148 0.047
R14235 fc2.n2415 fc2.n2403 0.047
R14236 fc2.n778 fc2.n773 0.047
R14237 fc2.n988 fc2.n976 0.047
R14238 fc2.n1801 fc2.n1796 0.047
R14239 fc2.n1966 fc2.n1956 0.047
R14240 fc2.n1179 fc2.n1171 0.047
R14241 fc2.n1530 fc2.n1020 0.047
R14242 fc2.n2694 fc2.n2693 0.047
R14243 fc2.n2540 fc2.n2538 0.047
R14244 fc2.n231 fc2.n211 0.047
R14245 fc2.n412 fc2.n389 0.047
R14246 fc2.n2134 fc2.n2115 0.047
R14247 fc2.n2385 fc2.n2362 0.047
R14248 fc2.n759 fc2.n740 0.047
R14249 fc2.n1017 fc2.n1001 0.047
R14250 fc2.n1494 fc2.n1470 0.047
R14251 fc2.n1938 fc2.n1917 0.047
R14252 fc2.n1157 fc2.n1137 0.047
R14253 fc2.n1063 fc2.n1037 0.047
R14254 fc2.n916 fc2.n894 0.047
R14255 fc2.n1731 fc2.n1712 0.047
R14256 fc2.n1584 fc2.n1561 0.047
R14257 fc2.n1211 fc2.n1075 0.047
R14258 fc2.n1251 fc2.n1225 0.047
R14259 fc2.n2302 fc2.n2276 0.047
R14260 fc2.n674 fc2.n655 0.047
R14261 fc2.n604 fc2.n581 0.047
R14262 fc2.n1623 fc2.n1598 0.047
R14263 fc2.n1660 fc2.n1637 0.047
R14264 fc2.n1289 fc2.n1263 0.047
R14265 fc2.n1329 fc2.n1303 0.047
R14266 fc2.n497 fc2.n474 0.047
R14267 fc2.n2046 fc2.n2027 0.047
R14268 fc2.n2229 fc2.n2206 0.047
R14269 fc2.n809 fc2.n617 0.047
R14270 fc2.n847 fc2.n824 0.047
R14271 fc2.n1832 fc2.n1673 0.047
R14272 fc2.n1870 fc2.n1847 0.047
R14273 fc2.n1367 fc2.n1341 0.047
R14274 fc2.n1407 fc2.n1381 0.047
R14275 fc2.n1157 fc2.n1134 0.047
R14276 fc2.n2457 fc2.n2455 0.047
R14277 fc2.n3570 fc2.n3569 0.047
R14278 fc2.n3670 fc2.n3669 0.047
R14279 fc2.n3722 fc2.n3721 0.047
R14280 fc2.n1964 fc2.n1958 0.046
R14281 fc2.n3478 fc2.n3464 0.046
R14282 fc2.n3618 fc2.n3604 0.046
R14283 fc2.n2739 fc2.n2733 0.046
R14284 fc2.n2709 fc2.n2701 0.046
R14285 fc2 fc2.n3991 0.046
R14286 fc2.n3772 fc2.n3771 0.045
R14287 fc2.n334 fc2.n333 0.045
R14288 fc2.n3339 fc2.n3337 0.045
R14289 fc2.n3720 fc2.n3719 0.045
R14290 fc2.n2737 fc2.n2736 0.045
R14291 fc2.n3575 fc2.n3574 0.045
R14292 fc2.n3449 fc2.n3448 0.045
R14293 fc2.n3974 fc2.n3973 0.045
R14294 fc2.n3962 fc2.n3961 0.045
R14295 fc2.n3675 fc2.n3674 0.045
R14296 fc2.n3589 fc2.n3588 0.045
R14297 fc2.n3851 fc2.n3850 0.045
R14298 fc2.n3839 fc2.n3838 0.045
R14299 fc2.n3725 fc2.n3724 0.045
R14300 fc2.n3735 fc2.n3734 0.045
R14301 fc2.n251 fc2.n249 0.045
R14302 fc2.n361 fc2.n359 0.045
R14303 fc2.n2169 fc2.n2167 0.045
R14304 fc2.n1769 fc2.n1768 0.045
R14305 fc2.n941 fc2.n940 0.045
R14306 fc2.n716 fc2.n715 0.045
R14307 fc2.n2324 fc2.n2323 0.045
R14308 fc2.n2088 fc2.n2087 0.045
R14309 fc2.n437 fc2.n436 0.045
R14310 fc2.n187 fc2.n186 0.045
R14311 fc2.n395 fc2.n393 0.045
R14312 fc2.n2121 fc2.n2119 0.045
R14313 fc2.n2368 fc2.n2366 0.045
R14314 fc2.n746 fc2.n744 0.045
R14315 fc2.n217 fc2.n215 0.045
R14316 fc2.n1923 fc2.n1921 0.045
R14317 fc2.n1143 fc2.n1141 0.045
R14318 fc2.n1043 fc2.n1041 0.045
R14319 fc2.n900 fc2.n898 0.045
R14320 fc2.n1718 fc2.n1716 0.045
R14321 fc2.n1567 fc2.n1565 0.045
R14322 fc2.n1197 fc2.n1195 0.045
R14323 fc2.n1231 fc2.n1229 0.045
R14324 fc2.n2285 fc2.n2283 0.045
R14325 fc2.n661 fc2.n659 0.045
R14326 fc2.n587 fc2.n585 0.045
R14327 fc2.n1610 fc2.n1608 0.045
R14328 fc2.n1643 fc2.n1641 0.045
R14329 fc2.n1275 fc2.n1273 0.045
R14330 fc2.n1309 fc2.n1307 0.045
R14331 fc2.n470 fc2.n469 0.045
R14332 fc2.n480 fc2.n478 0.045
R14333 fc2.n2033 fc2.n2031 0.045
R14334 fc2.n2212 fc2.n2210 0.045
R14335 fc2.n796 fc2.n794 0.045
R14336 fc2.n830 fc2.n828 0.045
R14337 fc2.n1819 fc2.n1817 0.045
R14338 fc2.n1853 fc2.n1851 0.045
R14339 fc2.n1353 fc2.n1351 0.045
R14340 fc2.n1387 fc2.n1385 0.045
R14341 fc2.n3772 fc2.n3769 0.044
R14342 fc2.n3762 fc2.n3759 0.044
R14343 fc2.n2 fc2.n1 0.044
R14344 fc2.n1178 fc2.n1174 0.044
R14345 fc2.n1450 fc2.n1449 0.044
R14346 fc2.n1491 fc2.n1490 0.044
R14347 fc2.n313 fc2.n312 0.044
R14348 fc2.n558 fc2.n543 0.043
R14349 fc2.n3886 fc2.n3885 0.043
R14350 fc2.n3803 fc2.n3802 0.043
R14351 fc2.n3717 fc2.n3716 0.043
R14352 fc2.n1080 fc2.n1079 0.043
R14353 fc2.n3467 fc2.n3466 0.043
R14354 fc2.n3876 fc2.n3875 0.043
R14355 fc2.n3607 fc2.n3606 0.043
R14356 fc2.n3793 fc2.n3792 0.043
R14357 fc2.n3699 fc2.n3698 0.043
R14358 fc2.n320 fc2.n319 0.043
R14359 fc2.n2395 fc2.n2394 0.043
R14360 fc2.n968 fc2.n967 0.043
R14361 fc2.n1949 fc2.n1948 0.043
R14362 fc2.n11 fc2.n10 0.042
R14363 fc2.n2444 fc2.n2183 0.042
R14364 fc2.n559 fc2.n315 0.042
R14365 fc2.n3990 fc2.n3989 0.041
R14366 fc2.n2480 fc2.n2479 0.041
R14367 fc2.n1518 fc2.n1517 0.04
R14368 fc2.n2643 fc2.n2636 0.04
R14369 fc2.n134 fc2.n128 0.04
R14370 fc2.n2004 fc2.n1998 0.04
R14371 fc2.n631 fc2.n625 0.04
R14372 fc2.n1688 fc2.n1682 0.04
R14373 fc2.n1090 fc2.n1084 0.04
R14374 fc2.n261 fc2.n260 0.04
R14375 fc2.n374 fc2.n373 0.04
R14376 fc2.n2178 fc2.n2177 0.04
R14377 fc2.n1777 fc2.n1776 0.04
R14378 fc2.n952 fc2.n951 0.04
R14379 fc2.n723 fc2.n722 0.04
R14380 fc2.n2335 fc2.n2334 0.04
R14381 fc2.n2095 fc2.n2094 0.04
R14382 fc2.n448 fc2.n447 0.04
R14383 fc2.n195 fc2.n194 0.04
R14384 fc2.n226 fc2.n225 0.04
R14385 fc2.n408 fc2.n407 0.04
R14386 fc2.n2130 fc2.n2129 0.04
R14387 fc2.n2381 fc2.n2380 0.04
R14388 fc2.n755 fc2.n754 0.04
R14389 fc2.n2526 fc2.n2525 0.04
R14390 fc2.n2600 fc2.n2599 0.04
R14391 fc2.n1934 fc2.n1933 0.04
R14392 fc2.n1153 fc2.n1152 0.04
R14393 fc2.n912 fc2.n911 0.04
R14394 fc2.n1727 fc2.n1726 0.04
R14395 fc2.n1580 fc2.n1579 0.04
R14396 fc2.n1207 fc2.n1206 0.04
R14397 fc2.n2298 fc2.n2297 0.04
R14398 fc2.n670 fc2.n669 0.04
R14399 fc2.n600 fc2.n599 0.04
R14400 fc2.n1619 fc2.n1618 0.04
R14401 fc2.n1656 fc2.n1655 0.04
R14402 fc2.n1285 fc2.n1284 0.04
R14403 fc2.n493 fc2.n492 0.04
R14404 fc2.n2042 fc2.n2041 0.04
R14405 fc2.n2225 fc2.n2224 0.04
R14406 fc2.n805 fc2.n804 0.04
R14407 fc2.n843 fc2.n842 0.04
R14408 fc2.n1828 fc2.n1827 0.04
R14409 fc2.n1866 fc2.n1865 0.04
R14410 fc2.n1363 fc2.n1362 0.04
R14411 fc2.n507 fc2.n506 0.039
R14412 fc2.n2241 fc2.n2240 0.039
R14413 fc2.n856 fc2.n855 0.039
R14414 fc2.n1879 fc2.n1878 0.039
R14415 fc2.n1416 fc2.n1415 0.039
R14416 fc2.n343 fc2.n342 0.039
R14417 fc2.n420 fc2.n419 0.039
R14418 fc2.n2307 fc2.n2306 0.039
R14419 fc2.n924 fc2.n923 0.039
R14420 fc2.n2412 fc2.n2411 0.039
R14421 fc2.n985 fc2.n984 0.039
R14422 fc2.n2763 fc2.n2762 0.039
R14423 fc2.n2350 fc2.n2349 0.039
R14424 fc2.n1550 fc2.n1549 0.039
R14425 fc2.n570 fc2.n569 0.039
R14426 fc2.n1626 fc2.n1625 0.039
R14427 fc2.n2194 fc2.n2193 0.039
R14428 fc2.n812 fc2.n811 0.039
R14429 fc2.n1835 fc2.n1834 0.039
R14430 fc2.n3579 fc2.n3578 0.039
R14431 fc2.n3581 fc2.n3579 0.039
R14432 fc2.n3453 fc2.n3452 0.039
R14433 fc2.n3980 fc2.n3979 0.039
R14434 fc2.n3982 fc2.n3980 0.039
R14435 fc2.n3968 fc2.n3967 0.039
R14436 fc2.n3679 fc2.n3678 0.039
R14437 fc2.n3681 fc2.n3679 0.039
R14438 fc2.n3593 fc2.n3592 0.039
R14439 fc2.n3857 fc2.n3856 0.039
R14440 fc2.n3859 fc2.n3857 0.039
R14441 fc2.n3845 fc2.n3844 0.039
R14442 fc2.n3761 fc2.n3760 0.039
R14443 fc2.n3757 fc2.n3756 0.039
R14444 fc2.n3729 fc2.n3728 0.039
R14445 fc2.n3739 fc2.n3738 0.039
R14446 fc2.n3741 fc2.n3739 0.039
R14447 fc2.n3771 fc2.n3770 0.039
R14448 fc2.n3754 fc2.n3753 0.039
R14449 fc2.n2642 fc2.n2637 0.039
R14450 fc2.n133 fc2.n129 0.039
R14451 fc2.n2003 fc2.n1999 0.039
R14452 fc2.n630 fc2.n626 0.039
R14453 fc2.n1687 fc2.n1683 0.039
R14454 fc2.n1089 fc2.n1085 0.039
R14455 fc2.n1212 fc2.n1211 0.039
R14456 fc2.n1290 fc2.n1289 0.039
R14457 fc2.n1624 fc2.n1623 0.039
R14458 fc2.n1368 fc2.n1367 0.039
R14459 fc2.n1833 fc2.n1832 0.039
R14460 fc2.n810 fc2.n809 0.039
R14461 fc2.t56 fc2.n3394 0.038
R14462 fc2.n1047 fc2.n1046 0.038
R14463 fc2.n1235 fc2.n1234 0.038
R14464 fc2.n1313 fc2.n1312 0.038
R14465 fc2.n1391 fc2.n1390 0.038
R14466 fc2.t56 fc2.n3428 0.038
R14467 fc2.n2641 fc2.n2638 0.037
R14468 fc2.n132 fc2.n130 0.037
R14469 fc2.n2002 fc2.n2000 0.037
R14470 fc2.n629 fc2.n627 0.037
R14471 fc2.n1686 fc2.n1684 0.037
R14472 fc2.n1088 fc2.n1086 0.037
R14473 fc2.n1483 fc2.n1482 0.037
R14474 fc2.n2176 fc2.n2175 0.037
R14475 fc2.n753 fc2.n752 0.037
R14476 fc2.n1452 fc2.n1451 0.037
R14477 fc2.n79 fc2.n77 0.037
R14478 fc2.n2800 fc2.n2796 0.037
R14479 fc2.n553 fc2.n549 0.037
R14480 fc2.n2438 fc2.n2434 0.037
R14481 fc2.n1011 fc2.n1007 0.037
R14482 fc2.n1540 fc2.n1536 0.037
R14483 fc2.n1522 fc2.n1515 0.037
R14484 fc2.n1083 fc2.n1082 0.037
R14485 fc2.n1032 fc2.n1029 0.037
R14486 fc2.n1681 fc2.n1680 0.037
R14487 fc2.n624 fc2.n623 0.037
R14488 fc2.n1997 fc2.n1996 0.037
R14489 fc2.n127 fc2.n126 0.037
R14490 fc2.n2650 fc2.n2649 0.037
R14491 fc2.n1494 fc2.n1464 0.036
R14492 fc2.n1965 fc2.n1964 0.036
R14493 fc2.n2671 fc2.n2667 0.036
R14494 fc2.n2685 fc2.n2684 0.036
R14495 fc2.n2628 fc2.n2627 0.036
R14496 fc2.t56 fc2.n3440 0.036
R14497 fc2.n340 fc2.n339 0.035
R14498 fc2.n2657 fc2.n2656 0.035
R14499 fc2.n1110 fc2.n1109 0.035
R14500 fc2.n1703 fc2.n1702 0.035
R14501 fc2.n646 fc2.n645 0.035
R14502 fc2.n2019 fc2.n2018 0.035
R14503 fc2.n149 fc2.n148 0.035
R14504 fc2.n265 fc2.n252 0.035
R14505 fc2.n378 fc2.n362 0.035
R14506 fc2.n2182 fc2.n2170 0.035
R14507 fc2.n378 fc2.n352 0.035
R14508 fc2.n265 fc2.n242 0.035
R14509 fc2.n201 fc2.n178 0.035
R14510 fc2.n454 fc2.n428 0.035
R14511 fc2.n2101 fc2.n2079 0.035
R14512 fc2.n2341 fc2.n2315 0.035
R14513 fc2.n729 fc2.n707 0.035
R14514 fc2.n958 fc2.n932 0.035
R14515 fc2.n1782 fc2.n1770 0.035
R14516 fc2.n958 fc2.n942 0.035
R14517 fc2.n729 fc2.n717 0.035
R14518 fc2.n2341 fc2.n2325 0.035
R14519 fc2.n2101 fc2.n2089 0.035
R14520 fc2.n454 fc2.n438 0.035
R14521 fc2.n201 fc2.n188 0.035
R14522 fc2.n335 fc2.n322 0.035
R14523 fc2.n2415 fc2.n2397 0.035
R14524 fc2.n988 fc2.n970 0.035
R14525 fc2.n1801 fc2.n1797 0.035
R14526 fc2.n988 fc2.n983 0.035
R14527 fc2.n778 fc2.n774 0.035
R14528 fc2.n2415 fc2.n2410 0.035
R14529 fc2.n412 fc2.n396 0.035
R14530 fc2.n2134 fc2.n2122 0.035
R14531 fc2.n2385 fc2.n2369 0.035
R14532 fc2.n759 fc2.n747 0.035
R14533 fc2.n2385 fc2.n2359 0.035
R14534 fc2.n2134 fc2.n2112 0.035
R14535 fc2.n231 fc2.n218 0.035
R14536 fc2.n1938 fc2.n1924 0.035
R14537 fc2.n1157 fc2.n1144 0.035
R14538 fc2.n916 fc2.n901 0.035
R14539 fc2.n1731 fc2.n1719 0.035
R14540 fc2.n1584 fc2.n1568 0.035
R14541 fc2.n1211 fc2.n1198 0.035
R14542 fc2.n2302 fc2.n2286 0.035
R14543 fc2.n674 fc2.n662 0.035
R14544 fc2.n604 fc2.n588 0.035
R14545 fc2.n1623 fc2.n1611 0.035
R14546 fc2.n1660 fc2.n1644 0.035
R14547 fc2.n1289 fc2.n1276 0.035
R14548 fc2.n1407 fc2.n1378 0.035
R14549 fc2.n1870 fc2.n1844 0.035
R14550 fc2.n1832 fc2.n1670 0.035
R14551 fc2.n847 fc2.n821 0.035
R14552 fc2.n809 fc2.n614 0.035
R14553 fc2.n2229 fc2.n2203 0.035
R14554 fc2.n2046 fc2.n2024 0.035
R14555 fc2.n497 fc2.n471 0.035
R14556 fc2.n497 fc2.n481 0.035
R14557 fc2.n2046 fc2.n2034 0.035
R14558 fc2.n2229 fc2.n2213 0.035
R14559 fc2.n809 fc2.n797 0.035
R14560 fc2.n847 fc2.n831 0.035
R14561 fc2.n1832 fc2.n1820 0.035
R14562 fc2.n1870 fc2.n1854 0.035
R14563 fc2.n1367 fc2.n1354 0.035
R14564 fc2.n1438 fc2.n1425 0.035
R14565 fc2.n1125 fc2.n1114 0.035
R14566 fc2.n1899 fc2.n1888 0.035
R14567 fc2.n1752 fc2.n1741 0.035
R14568 fc2.n876 fc2.n865 0.035
R14569 fc2.n695 fc2.n684 0.035
R14570 fc2.n2261 fc2.n2250 0.035
R14571 fc2.n2067 fc2.n2056 0.035
R14572 fc2.n533 fc2.n516 0.035
R14573 fc2.n166 fc2.n154 0.035
R14574 fc2.n166 fc2.n161 0.035
R14575 fc2.n533 fc2.n529 0.035
R14576 fc2.n2067 fc2.n2063 0.035
R14577 fc2.n2261 fc2.n2257 0.035
R14578 fc2.n695 fc2.n691 0.035
R14579 fc2.n876 fc2.n872 0.035
R14580 fc2.n1125 fc2.n1121 0.035
R14581 fc2.t14 fc2.n50 0.035
R14582 fc2.t14 fc2.n45 0.035
R14583 fc2.t14 fc2.n38 0.035
R14584 fc2.t14 fc2.n23 0.035
R14585 fc2.t14 fc2.n17 0.035
R14586 fc2.t14 fc2.n31 0.035
R14587 fc2.t56 fc2.n3419 0.035
R14588 fc2.t56 fc2.n3396 0.035
R14589 fc2.t56 fc2.n3382 0.035
R14590 fc2.t56 fc2.n3367 0.035
R14591 fc2.t56 fc2.n3351 0.035
R14592 fc2.n1174 fc2.n1173 0.034
R14593 fc2.n2989 fc2.n2988 0.034
R14594 fc2.n2806 fc2.n2452 0.034
R14595 fc2.n2444 fc2.n2190 0.034
R14596 fc2.n1017 fc2.n566 0.034
R14597 fc2.n559 fc2.n119 0.034
R14598 fc2.t14 fc2.n49 0.034
R14599 fc2.t14 fc2.n48 0.034
R14600 fc2.t14 fc2.n37 0.034
R14601 fc2.t14 fc2.n24 0.034
R14602 fc2.t14 fc2.n18 0.034
R14603 fc2.t14 fc2.n30 0.034
R14604 fc2.t56 fc2.n3418 0.034
R14605 fc2.t56 fc2.n3395 0.034
R14606 fc2.t56 fc2.n3381 0.034
R14607 fc2.t56 fc2.n3366 0.034
R14608 fc2.t56 fc2.n3350 0.034
R14609 fc2.t56 fc2.n3439 0.034
R14610 fc2.n1055 fc2.n1054 0.033
R14611 fc2.n1243 fc2.n1242 0.033
R14612 fc2.n1321 fc2.n1320 0.033
R14613 fc2.n1399 fc2.n1398 0.033
R14614 fc2.n3777 fc2.n3768 0.033
R14615 fc2.n3081 fc2.n3080 0.033
R14616 fc2.n3010 fc2.n3009 0.033
R14617 fc2.n2959 fc2.n2958 0.033
R14618 fc2.n2916 fc2.n2915 0.033
R14619 fc2.n2825 fc2.n2824 0.033
R14620 fc2.n1963 fc2.n1962 0.033
R14621 fc2.n3581 fc2.n3573 0.033
R14622 fc2.n3982 fc2.n3972 0.033
R14623 fc2.n3681 fc2.n3673 0.033
R14624 fc2.n3859 fc2.n3849 0.033
R14625 fc2.n3741 fc2.n3733 0.033
R14626 fc2.n109 fc2.n3 0.033
R14627 fc2.n1100 fc2.n1099 0.032
R14628 fc2.n1211 fc2.n1071 0.032
R14629 fc2.n1289 fc2.n1259 0.032
R14630 fc2.n1367 fc2.n1337 0.032
R14631 fc2.n1045 fc2.n1044 0.032
R14632 fc2.n1233 fc2.n1232 0.032
R14633 fc2.n1311 fc2.n1310 0.032
R14634 fc2.n1389 fc2.n1388 0.032
R14635 fc2.n262 fc2.n261 0.031
R14636 fc2.n375 fc2.n374 0.031
R14637 fc2.n2179 fc2.n2178 0.031
R14638 fc2.n1779 fc2.n1777 0.031
R14639 fc2.n955 fc2.n952 0.031
R14640 fc2.n726 fc2.n723 0.031
R14641 fc2.n2338 fc2.n2335 0.031
R14642 fc2.n2098 fc2.n2095 0.031
R14643 fc2.n451 fc2.n448 0.031
R14644 fc2.n198 fc2.n195 0.031
R14645 fc2.n227 fc2.n226 0.031
R14646 fc2.n409 fc2.n408 0.031
R14647 fc2.n2131 fc2.n2130 0.031
R14648 fc2.n2382 fc2.n2381 0.031
R14649 fc2.n756 fc2.n755 0.031
R14650 fc2.n2527 fc2.n2526 0.031
R14651 fc2.n2601 fc2.n2600 0.031
R14652 fc2.n1935 fc2.n1934 0.031
R14653 fc2.n1154 fc2.n1153 0.031
R14654 fc2.n913 fc2.n912 0.031
R14655 fc2.n1728 fc2.n1727 0.031
R14656 fc2.n1581 fc2.n1580 0.031
R14657 fc2.n1208 fc2.n1207 0.031
R14658 fc2.n2299 fc2.n2298 0.031
R14659 fc2.n671 fc2.n670 0.031
R14660 fc2.n601 fc2.n600 0.031
R14661 fc2.n1620 fc2.n1619 0.031
R14662 fc2.n1657 fc2.n1656 0.031
R14663 fc2.n1286 fc2.n1285 0.031
R14664 fc2.n494 fc2.n493 0.031
R14665 fc2.n2043 fc2.n2042 0.031
R14666 fc2.n2226 fc2.n2225 0.031
R14667 fc2.n806 fc2.n805 0.031
R14668 fc2.n844 fc2.n843 0.031
R14669 fc2.n1829 fc2.n1828 0.031
R14670 fc2.n1867 fc2.n1866 0.031
R14671 fc2.n1364 fc2.n1363 0.031
R14672 fc2.t62 fc2.n340 0.031
R14673 fc2.t4 fc2.n2657 0.031
R14674 fc2.t10 fc2.n1110 0.031
R14675 fc2.t12 fc2.n1703 0.031
R14676 fc2.t52 fc2.n646 0.031
R14677 fc2.t98 fc2.n2019 0.031
R14678 fc2.t66 fc2.n149 0.031
R14679 fc2.n298 fc2.n294 0.031
R14680 fc2.n2613 fc2.n2587 0.031
R14681 fc2.n3307 fc2.n3306 0.031
R14682 fc2.n2672 fc2.n2671 0.031
R14683 fc2.n294 fc2.n293 0.031
R14684 fc2.n2587 fc2.n2586 0.031
R14685 fc2.n1050 fc2.n1049 0.03
R14686 fc2.n1238 fc2.n1237 0.03
R14687 fc2.n1316 fc2.n1315 0.03
R14688 fc2.n1394 fc2.n1393 0.03
R14689 fc2.t56 fc2.n3380 0.03
R14690 fc2.t56 fc2.n3365 0.03
R14691 fc2.n1985 fc2.n1979 0.03
R14692 fc2.n3755 fc2.n3747 0.03
R14693 fc2.n3755 fc2.n3752 0.03
R14694 fc2.n1092 fc2.n1083 0.029
R14695 fc2.n1690 fc2.n1681 0.029
R14696 fc2.n633 fc2.n624 0.029
R14697 fc2.n2006 fc2.n1997 0.029
R14698 fc2.n136 fc2.n127 0.029
R14699 fc2.n2651 fc2.n2650 0.029
R14700 fc2.n2571 fc2.n2570 0.028
R14701 fc2.n2707 fc2.n2706 0.028
R14702 fc2.n2504 fc2.n2500 0.028
R14703 fc2.n2686 fc2.n2685 0.028
R14704 fc2.n2629 fc2.n2628 0.028
R14705 fc2.n2799 fc2.n2798 0.028
R14706 fc2.n552 fc2.n551 0.028
R14707 fc2.n2437 fc2.n2436 0.028
R14708 fc2.n1010 fc2.n1009 0.028
R14709 fc2.n1539 fc2.n1538 0.028
R14710 fc2.n1521 fc2.n1520 0.028
R14711 fc2.n109 fc2.n2 0.028
R14712 fc2.n1082 fc2.n1081 0.028
R14713 fc2.n1482 fc2.n1481 0.028
R14714 fc2.n1029 fc2.n1026 0.028
R14715 fc2.n1680 fc2.n1679 0.028
R14716 fc2.n623 fc2.n622 0.028
R14717 fc2.n1996 fc2.n1995 0.028
R14718 fc2.n126 fc2.n125 0.028
R14719 fc2.n2649 fc2.n2648 0.028
R14720 fc2.n2767 fc2.n2766 0.027
R14721 fc2.t14 fc2.n25 0.027
R14722 fc2.n2740 fc2.n2732 0.027
R14723 fc2.n2718 fc2.n2710 0.027
R14724 fc2.n2575 fc2.n2555 0.027
R14725 fc2.n2507 fc2.n2488 0.027
R14726 fc2.n2766 fc2.n2761 0.027
R14727 fc2.n2540 fc2.n2531 0.027
R14728 fc2.n2608 fc2.n2605 0.027
R14729 fc2.n314 fc2.n311 0.027
R14730 fc2.n1938 fc2.n1914 0.027
R14731 fc2.n1251 fc2.n1222 0.027
R14732 fc2.n1584 fc2.n1558 0.027
R14733 fc2.n1731 fc2.n1709 0.027
R14734 fc2.n916 fc2.n891 0.027
R14735 fc2.n1329 fc2.n1300 0.027
R14736 fc2.n1660 fc2.n1634 0.027
R14737 fc2.n1623 fc2.n1595 0.027
R14738 fc2.n604 fc2.n578 0.027
R14739 fc2.n674 fc2.n652 0.027
R14740 fc2.n2302 fc2.n2273 0.027
R14741 fc2.n3581 fc2.n3454 0.027
R14742 fc2.n3982 fc2.n3969 0.027
R14743 fc2.n3681 fc2.n3594 0.027
R14744 fc2.n3859 fc2.n3846 0.027
R14745 fc2.n3777 fc2.n3765 0.027
R14746 fc2.n3741 fc2.n3730 0.027
R14747 fc2.n3777 fc2.n3775 0.027
R14748 fc2.n2472 fc2.n2458 0.027
R14749 fc2.n2472 fc2.n2466 0.027
R14750 fc2.t14 fc2.n22 0.027
R14751 fc2.t14 fc2.n43 0.026
R14752 fc2.t14 fc2.n36 0.026
R14753 fc2.n1963 fc2.n1960 0.026
R14754 fc2.n1511 fc2.n1510 0.025
R14755 fc2.n1105 fc2.n1104 0.025
R14756 fc2.n1063 fc2.n1023 0.025
R14757 fc2.n1698 fc2.n1697 0.025
R14758 fc2.n641 fc2.n640 0.025
R14759 fc2.n2014 fc2.n2013 0.025
R14760 fc2.n144 fc2.n143 0.025
R14761 fc2.n1529 fc2.n1511 0.025
R14762 fc2.n3349 fc2.n3348 0.025
R14763 fc2.n3438 fc2.n3433 0.025
R14764 fc2.n1966 fc2.n1965 0.025
R14765 fc2.n527 fc2.n524 0.025
R14766 fc2.n16 fc2.n15 0.024
R14767 fc2.n2647 fc2.n2646 0.024
R14768 fc2.n2564 fc2.n2563 0.024
R14769 fc2.n2568 fc2.n2567 0.024
R14770 fc2.n259 fc2.n258 0.024
R14771 fc2.n370 fc2.n369 0.024
R14772 fc2.n373 fc2.n372 0.024
R14773 fc2.n2703 fc2.n2702 0.024
R14774 fc2.n2559 fc2.n2558 0.024
R14775 fc2.n1776 fc2.n1775 0.024
R14776 fc2.n954 fc2.n953 0.024
R14777 fc2.n951 fc2.n950 0.024
R14778 fc2.n725 fc2.n724 0.024
R14779 fc2.n2337 fc2.n2336 0.024
R14780 fc2.n2334 fc2.n2333 0.024
R14781 fc2.n2097 fc2.n2096 0.024
R14782 fc2.n450 fc2.n449 0.024
R14783 fc2.n447 fc2.n446 0.024
R14784 fc2.n197 fc2.n196 0.024
R14785 fc2.n2502 fc2.n2501 0.024
R14786 fc2.n2498 fc2.n2497 0.024
R14787 fc2.n2669 fc2.n2668 0.024
R14788 fc2.n2492 fc2.n2491 0.024
R14789 fc2.n224 fc2.n223 0.024
R14790 fc2.n404 fc2.n403 0.024
R14791 fc2.n407 fc2.n406 0.024
R14792 fc2.n2128 fc2.n2127 0.024
R14793 fc2.n2377 fc2.n2376 0.024
R14794 fc2.n2380 fc2.n2379 0.024
R14795 fc2.n2681 fc2.n2680 0.024
R14796 fc2.n2515 fc2.n2514 0.024
R14797 fc2.n2522 fc2.n2521 0.024
R14798 fc2.n2525 fc2.n2524 0.024
R14799 fc2.n2624 fc2.n2623 0.024
R14800 fc2.n2589 fc2.n2588 0.024
R14801 fc2.n2596 fc2.n2595 0.024
R14802 fc2.n2599 fc2.n2598 0.024
R14803 fc2.n1456 fc2.n1455 0.024
R14804 fc2.n1094 fc2.n1093 0.024
R14805 fc2.n1097 fc2.n1096 0.024
R14806 fc2.n1078 fc2.n1077 0.024
R14807 fc2.n1081 fc2.n1080 0.024
R14808 fc2.n1476 fc2.n1475 0.024
R14809 fc2.n1481 fc2.n1480 0.024
R14810 fc2.n1031 fc2.n1030 0.024
R14811 fc2.n1026 fc2.n1025 0.024
R14812 fc2.n1692 fc2.n1691 0.024
R14813 fc2.n1909 fc2.n1908 0.024
R14814 fc2.n1676 fc2.n1675 0.024
R14815 fc2.n1679 fc2.n1678 0.024
R14816 fc2.n1930 fc2.n1929 0.024
R14817 fc2.n1933 fc2.n1932 0.024
R14818 fc2.n1150 fc2.n1149 0.024
R14819 fc2.n1152 fc2.n1151 0.024
R14820 fc2.n635 fc2.n634 0.024
R14821 fc2.n886 fc2.n885 0.024
R14822 fc2.n620 fc2.n619 0.024
R14823 fc2.n622 fc2.n621 0.024
R14824 fc2.n908 fc2.n907 0.024
R14825 fc2.n911 fc2.n910 0.024
R14826 fc2.n1725 fc2.n1724 0.024
R14827 fc2.n1576 fc2.n1575 0.024
R14828 fc2.n1579 fc2.n1578 0.024
R14829 fc2.n1204 fc2.n1203 0.024
R14830 fc2.n1206 fc2.n1205 0.024
R14831 fc2.n2008 fc2.n2007 0.024
R14832 fc2.n2268 fc2.n2267 0.024
R14833 fc2.n1994 fc2.n1993 0.024
R14834 fc2.n2294 fc2.n2293 0.024
R14835 fc2.n2297 fc2.n2296 0.024
R14836 fc2.n668 fc2.n667 0.024
R14837 fc2.n596 fc2.n595 0.024
R14838 fc2.n599 fc2.n598 0.024
R14839 fc2.n1617 fc2.n1616 0.024
R14840 fc2.n1652 fc2.n1651 0.024
R14841 fc2.n1655 fc2.n1654 0.024
R14842 fc2.n1282 fc2.n1281 0.024
R14843 fc2.n1284 fc2.n1283 0.024
R14844 fc2.n138 fc2.n137 0.024
R14845 fc2.n463 fc2.n462 0.024
R14846 fc2.n124 fc2.n123 0.024
R14847 fc2.n489 fc2.n488 0.024
R14848 fc2.n492 fc2.n491 0.024
R14849 fc2.n2040 fc2.n2039 0.024
R14850 fc2.n2221 fc2.n2220 0.024
R14851 fc2.n2224 fc2.n2223 0.024
R14852 fc2.n803 fc2.n802 0.024
R14853 fc2.n839 fc2.n838 0.024
R14854 fc2.n842 fc2.n841 0.024
R14855 fc2.n1826 fc2.n1825 0.024
R14856 fc2.n1862 fc2.n1861 0.024
R14857 fc2.n1865 fc2.n1864 0.024
R14858 fc2.n1360 fc2.n1359 0.024
R14859 fc2.n1362 fc2.n1361 0.024
R14860 fc2.n75 fc2.n74 0.024
R14861 fc2.n105 fc2.n104 0.024
R14862 fc2.n104 fc2.n103 0.024
R14863 fc2.n2452 fc2.n2451 0.023
R14864 fc2.n2190 fc2.n2189 0.023
R14865 fc2.n1963 fc2.n1959 0.023
R14866 fc2.n566 fc2.n565 0.023
R14867 fc2.n119 fc2.n118 0.023
R14868 fc2.n1487 fc2.n1484 0.023
R14869 fc2.n1695 fc2.n1694 0.023
R14870 fc2.n1034 fc2.n1033 0.023
R14871 fc2.n638 fc2.n637 0.023
R14872 fc2.n1219 fc2.n1218 0.023
R14873 fc2.n2011 fc2.n2010 0.023
R14874 fc2.n1297 fc2.n1296 0.023
R14875 fc2.n141 fc2.n140 0.023
R14876 fc2.n1375 fc2.n1374 0.023
R14877 fc2.n3576 fc2.n3575 0.023
R14878 fc2.n3578 fc2.n3577 0.023
R14879 fc2.n3452 fc2.n3451 0.023
R14880 fc2.n3450 fc2.n3449 0.023
R14881 fc2.n3977 fc2.n3974 0.023
R14882 fc2.n3979 fc2.n3978 0.023
R14883 fc2.n3967 fc2.n3966 0.023
R14884 fc2.n3965 fc2.n3962 0.023
R14885 fc2.n3676 fc2.n3675 0.023
R14886 fc2.n3678 fc2.n3677 0.023
R14887 fc2.n3592 fc2.n3591 0.023
R14888 fc2.n3590 fc2.n3589 0.023
R14889 fc2.n3854 fc2.n3851 0.023
R14890 fc2.n3856 fc2.n3855 0.023
R14891 fc2.n3844 fc2.n3843 0.023
R14892 fc2.n3842 fc2.n3839 0.023
R14893 fc2.n3726 fc2.n3725 0.023
R14894 fc2.n3728 fc2.n3727 0.023
R14895 fc2.n3736 fc2.n3735 0.023
R14896 fc2.n3738 fc2.n3737 0.023
R14897 fc2.n526 fc2.n525 0.023
R14898 fc2.n2555 fc2.n2554 0.023
R14899 fc2.n2488 fc2.n2487 0.023
R14900 fc2.n2531 fc2.n2530 0.023
R14901 fc2.n2605 fc2.n2604 0.023
R14902 fc2.n311 fc2.n310 0.023
R14903 fc2.n1914 fc2.n1913 0.023
R14904 fc2.n891 fc2.n890 0.023
R14905 fc2.n2273 fc2.n2272 0.023
R14906 fc2.n1048 fc2.n1047 0.023
R14907 fc2.n1236 fc2.n1235 0.023
R14908 fc2.n1314 fc2.n1313 0.023
R14909 fc2.n1392 fc2.n1391 0.023
R14910 fc2.n2736 fc2.n2735 0.022
R14911 fc2.n3404 fc2.n3403 0.022
R14912 fc2.n111 fc2.n110 0.022
R14913 fc2.n524 fc2.n523 0.022
R14914 fc2.n2572 fc2.n2571 0.021
R14915 fc2.n2708 fc2.n2707 0.021
R14916 fc2.n2505 fc2.n2504 0.021
R14917 fc2.n3402 fc2.n3401 0.021
R14918 fc2.n3759 fc2.n3757 0.021
R14919 fc2.n345 fc2.n344 0.021
R14920 fc2.n241 fc2.n240 0.021
R14921 fc2.n177 fc2.n176 0.021
R14922 fc2.n422 fc2.n421 0.021
R14923 fc2.n2078 fc2.n2077 0.021
R14924 fc2.n2309 fc2.n2308 0.021
R14925 fc2.n706 fc2.n705 0.021
R14926 fc2.n926 fc2.n925 0.021
R14927 fc2.n2765 fc2.n2764 0.021
R14928 fc2.n1165 fc2.n1164 0.021
R14929 fc2.n1800 fc2.n1799 0.021
R14930 fc2.n987 fc2.n986 0.021
R14931 fc2.n777 fc2.n776 0.021
R14932 fc2.n2414 fc2.n2413 0.021
R14933 fc2.n2150 fc2.n2149 0.021
R14934 fc2.n2352 fc2.n2351 0.021
R14935 fc2.n2111 fc2.n2110 0.021
R14936 fc2.n1215 fc2.n1214 0.021
R14937 fc2.n1552 fc2.n1551 0.021
R14938 fc2.n1707 fc2.n1706 0.021
R14939 fc2.n1293 fc2.n1292 0.021
R14940 fc2.n1628 fc2.n1627 0.021
R14941 fc2.n1593 fc2.n1592 0.021
R14942 fc2.n572 fc2.n571 0.021
R14943 fc2.n650 fc2.n649 0.021
R14944 fc2.n1371 fc2.n1370 0.021
R14945 fc2.n1837 fc2.n1836 0.021
R14946 fc2.n1669 fc2.n1668 0.021
R14947 fc2.n814 fc2.n813 0.021
R14948 fc2.n613 fc2.n612 0.021
R14949 fc2.n2196 fc2.n2195 0.021
R14950 fc2.n2023 fc2.n2022 0.021
R14951 fc2.n1418 fc2.n1417 0.021
R14952 fc2.n1113 fc2.n1112 0.021
R14953 fc2.n1881 fc2.n1880 0.021
R14954 fc2.n1740 fc2.n1739 0.021
R14955 fc2.n858 fc2.n857 0.021
R14956 fc2.n683 fc2.n682 0.021
R14957 fc2.n2243 fc2.n2242 0.021
R14958 fc2.n2055 fc2.n2054 0.021
R14959 fc2.n509 fc2.n508 0.021
R14960 fc2.n153 fc2.n152 0.021
R14961 fc2.n2471 fc2.n2470 0.021
R14962 fc2.n165 fc2.n164 0.021
R14963 fc2.n532 fc2.n531 0.021
R14964 fc2.n2066 fc2.n2065 0.021
R14965 fc2.n2260 fc2.n2259 0.021
R14966 fc2.n694 fc2.n693 0.021
R14967 fc2.n875 fc2.n874 0.021
R14968 fc2.n1751 fc2.n1750 0.021
R14969 fc2.n1898 fc2.n1897 0.021
R14970 fc2.n1124 fc2.n1123 0.021
R14971 fc2.n1437 fc2.n1436 0.021
R14972 fc2.n321 fc2.n317 0.021
R14973 fc2.n2396 fc2.n2392 0.021
R14974 fc2.n969 fc2.n965 0.021
R14975 fc2.n1950 fc2.n1946 0.021
R14976 fc2.n3339 fc2.n3338 0.021
R14977 fc2.n3339 fc2.n3315 0.021
R14978 fc2.n177 fc2.n174 0.021
R14979 fc2.n2078 fc2.n2075 0.021
R14980 fc2.n706 fc2.n703 0.021
R14981 fc2.n165 fc2.n162 0.021
R14982 fc2.n2066 fc2.n2064 0.021
R14983 fc2.n2260 fc2.n2258 0.021
R14984 fc2.n694 fc2.n692 0.021
R14985 fc2.n875 fc2.n873 0.021
R14986 fc2.n1751 fc2.n1749 0.021
R14987 fc2.n1898 fc2.n1896 0.021
R14988 fc2.n1124 fc2.n1122 0.021
R14989 fc2.n1437 fc2.n1433 0.021
R14990 fc2.n1912 fc2.n1911 0.021
R14991 fc2.n889 fc2.n888 0.021
R14992 fc2.n2271 fc2.n2270 0.021
R14993 fc2.n2457 fc2.n2456 0.021
R14994 fc2.n241 fc2.n239 0.021
R14995 fc2.n1800 fc2.n1798 0.021
R14996 fc2.n777 fc2.n775 0.021
R14997 fc2.n2111 fc2.n2109 0.021
R14998 fc2.n1669 fc2.n1667 0.021
R14999 fc2.n613 fc2.n611 0.021
R15000 fc2.n2023 fc2.n2021 0.021
R15001 fc2.n1113 fc2.n1111 0.021
R15002 fc2.n1740 fc2.n1738 0.021
R15003 fc2.n683 fc2.n681 0.021
R15004 fc2.n2055 fc2.n2053 0.021
R15005 fc2.n153 fc2.n151 0.021
R15006 fc2.n1462 fc2.n1461 0.019
R15007 fc2.n109 fc2.n54 0.019
R15008 fc2.n349 fc2.n348 0.019
R15009 fc2.n425 fc2.n423 0.019
R15010 fc2.n2312 fc2.n2310 0.019
R15011 fc2.n929 fc2.n927 0.019
R15012 fc2.n980 fc2.n979 0.019
R15013 fc2.n2407 fc2.n2406 0.019
R15014 fc2.n2356 fc2.n2355 0.019
R15015 fc2.n1053 fc2.n1052 0.019
R15016 fc2.n1555 fc2.n1554 0.019
R15017 fc2.n1241 fc2.n1240 0.019
R15018 fc2.n1631 fc2.n1630 0.019
R15019 fc2.n575 fc2.n574 0.019
R15020 fc2.n1319 fc2.n1318 0.019
R15021 fc2.n3346 fc2.n3345 0.019
R15022 fc2.n1841 fc2.n1840 0.019
R15023 fc2.n818 fc2.n817 0.019
R15024 fc2.n2200 fc2.n2199 0.019
R15025 fc2.n1397 fc2.n1396 0.019
R15026 fc2.n1422 fc2.n1421 0.019
R15027 fc2.n1885 fc2.n1884 0.019
R15028 fc2.n862 fc2.n861 0.019
R15029 fc2.n2247 fc2.n2246 0.019
R15030 fc2.n513 fc2.n512 0.019
R15031 fc2.n1102 fc2.n1101 0.019
R15032 fc2.n1105 fc2.n1102 0.019
R15033 fc2.n1063 fc2.n1034 0.019
R15034 fc2.n1698 fc2.n1695 0.019
R15035 fc2.n641 fc2.n638 0.019
R15036 fc2.n2014 fc2.n2011 0.019
R15037 fc2.n144 fc2.n141 0.019
R15038 fc2.n3435 fc2.n3434 0.019
R15039 fc2.n1222 fc2.n1221 0.019
R15040 fc2.n1300 fc2.n1299 0.019
R15041 fc2.n1459 fc2.n1458 0.019
R15042 fc2.n252 fc2.n251 0.019
R15043 fc2.n362 fc2.n361 0.019
R15044 fc2.n2170 fc2.n2169 0.019
R15045 fc2.n1770 fc2.n1769 0.019
R15046 fc2.n942 fc2.n941 0.019
R15047 fc2.n717 fc2.n716 0.019
R15048 fc2.n2325 fc2.n2324 0.019
R15049 fc2.n2089 fc2.n2088 0.019
R15050 fc2.n438 fc2.n437 0.019
R15051 fc2.n188 fc2.n187 0.019
R15052 fc2.n396 fc2.n395 0.019
R15053 fc2.n2122 fc2.n2121 0.019
R15054 fc2.n2369 fc2.n2368 0.019
R15055 fc2.n747 fc2.n746 0.019
R15056 fc2.n218 fc2.n217 0.019
R15057 fc2.n1924 fc2.n1923 0.019
R15058 fc2.n1144 fc2.n1143 0.019
R15059 fc2.n1057 fc2.n1043 0.019
R15060 fc2.n901 fc2.n900 0.019
R15061 fc2.n1719 fc2.n1718 0.019
R15062 fc2.n1568 fc2.n1567 0.019
R15063 fc2.n1198 fc2.n1197 0.019
R15064 fc2.n1245 fc2.n1231 0.019
R15065 fc2.n2286 fc2.n2285 0.019
R15066 fc2.n662 fc2.n661 0.019
R15067 fc2.n588 fc2.n587 0.019
R15068 fc2.n1611 fc2.n1610 0.019
R15069 fc2.n1644 fc2.n1643 0.019
R15070 fc2.n1276 fc2.n1275 0.019
R15071 fc2.n1323 fc2.n1309 0.019
R15072 fc2.n471 fc2.n470 0.019
R15073 fc2.n481 fc2.n480 0.019
R15074 fc2.n2034 fc2.n2033 0.019
R15075 fc2.n2213 fc2.n2212 0.019
R15076 fc2.n797 fc2.n796 0.019
R15077 fc2.n831 fc2.n830 0.019
R15078 fc2.n1820 fc2.n1819 0.019
R15079 fc2.n1854 fc2.n1853 0.019
R15080 fc2.n1354 fc2.n1353 0.019
R15081 fc2.n1401 fc2.n1387 0.019
R15082 fc2.n1217 fc2.n1216 0.018
R15083 fc2.n1295 fc2.n1294 0.018
R15084 fc2.n1373 fc2.n1372 0.018
R15085 fc2.n2806 fc2.n2805 0.018
R15086 fc2.n2444 fc2.n2443 0.018
R15087 fc2.n1017 fc2.n1016 0.018
R15088 fc2.n1367 fc2.n1338 0.018
R15089 fc2.n2806 fc2.n2453 0.018
R15090 fc2.n2444 fc2.n2191 0.018
R15091 fc2.n1017 fc2.n567 0.018
R15092 fc2.n559 fc2.n120 0.018
R15093 fc2.n348 fc2.n347 0.018
R15094 fc2.n979 fc2.n978 0.018
R15095 fc2.n2406 fc2.n2405 0.018
R15096 fc2.n2355 fc2.n2354 0.018
R15097 fc2.n3345 fc2.n3344 0.018
R15098 fc2.n1840 fc2.n1839 0.018
R15099 fc2.n817 fc2.n816 0.018
R15100 fc2.n2199 fc2.n2198 0.018
R15101 fc2.n1421 fc2.n1420 0.018
R15102 fc2.n1884 fc2.n1883 0.018
R15103 fc2.n861 fc2.n860 0.018
R15104 fc2.n2246 fc2.n2245 0.018
R15105 fc2.n512 fc2.n511 0.018
R15106 fc2.t56 fc2.n3349 0.017
R15107 fc2.t56 fc2.n3438 0.017
R15108 fc2.n1378 fc2.n1377 0.017
R15109 fc2.n1782 fc2.n1760 0.017
R15110 fc2.n1986 fc2.n1545 0.017
R15111 fc2.n467 fc2.n466 0.017
R15112 fc2.n1071 fc2.n1070 0.017
R15113 fc2.n1259 fc2.n1258 0.017
R15114 fc2.n1337 fc2.n1336 0.017
R15115 fc2.n1467 fc2.n1466 0.017
R15116 fc2.n1478 fc2.n1477 0.017
R15117 fc2.n1028 fc2.n1027 0.017
R15118 fc2.n1101 fc2.n1100 0.017
R15119 fc2.n1530 fc2.n1018 0.017
R15120 fc2.n559 fc2.n558 0.017
R15121 fc2.n1484 fc2.n1483 0.017
R15122 fc2.n1054 fc2.n1053 0.016
R15123 fc2.n1242 fc2.n1241 0.016
R15124 fc2.n1320 fc2.n1319 0.016
R15125 fc2.n1398 fc2.n1397 0.016
R15126 fc2.n3209 fc2.n3208 0.016
R15127 fc2.n3219 fc2.n3218 0.016
R15128 fc2.n3229 fc2.n3228 0.016
R15129 fc2.n3239 fc2.n3238 0.016
R15130 fc2.n3249 fc2.n3248 0.016
R15131 fc2.n3259 fc2.n3258 0.016
R15132 fc2.n3269 fc2.n3268 0.016
R15133 fc2.n3279 fc2.n3278 0.016
R15134 fc2.n3289 fc2.n3288 0.016
R15135 fc2.n3299 fc2.n3298 0.016
R15136 fc2.n3069 fc2.n3064 0.016
R15137 fc2.n2998 fc2.n2993 0.016
R15138 fc2.n2967 fc2.n2966 0.016
R15139 fc2.n2955 fc2.n2951 0.016
R15140 fc2.n2904 fc2.n2899 0.016
R15141 fc2.n2813 fc2.n2808 0.016
R15142 fc2.n1033 fc2.n1032 0.016
R15143 fc2.n1694 fc2.n1693 0.016
R15144 fc2.n637 fc2.n636 0.016
R15145 fc2.n2010 fc2.n2009 0.016
R15146 fc2.n140 fc2.n139 0.016
R15147 fc2.n2739 fc2.n2738 0.016
R15148 fc2.n2573 fc2.n2572 0.016
R15149 fc2.n350 fc2.n349 0.016
R15150 fc2.n2709 fc2.n2708 0.016
R15151 fc2.n426 fc2.n425 0.016
R15152 fc2.n2313 fc2.n2312 0.016
R15153 fc2.n930 fc2.n929 0.016
R15154 fc2.n2506 fc2.n2505 0.016
R15155 fc2.n2759 fc2.n2758 0.016
R15156 fc2.n981 fc2.n980 0.016
R15157 fc2.n2408 fc2.n2407 0.016
R15158 fc2.n2357 fc2.n2356 0.016
R15159 fc2.n2529 fc2.n2528 0.016
R15160 fc2.n309 fc2.n308 0.016
R15161 fc2.n2603 fc2.n2602 0.016
R15162 fc2.n1215 fc2.n1213 0.016
R15163 fc2.n1556 fc2.n1555 0.016
R15164 fc2.n1293 fc2.n1291 0.016
R15165 fc2.n1632 fc2.n1631 0.016
R15166 fc2.n576 fc2.n575 0.016
R15167 fc2.n3347 fc2.n3342 0.016
R15168 fc2.n1842 fc2.n1841 0.016
R15169 fc2.n819 fc2.n818 0.016
R15170 fc2.n2201 fc2.n2200 0.016
R15171 fc2.n3756 fc2.n3755 0.016
R15172 fc2.n3755 fc2.n3754 0.016
R15173 fc2.n1423 fc2.n1422 0.016
R15174 fc2.n1886 fc2.n1885 0.016
R15175 fc2.n863 fc2.n862 0.016
R15176 fc2.n2248 fc2.n2247 0.016
R15177 fc2.n514 fc2.n513 0.016
R15178 fc2.n3432 fc2.n3429 0.016
R15179 fc2.n1964 fc2.n1963 0.016
R15180 fc2.n3169 fc2.n3168 0.016
R15181 fc2.n3149 fc2.n3148 0.016
R15182 fc2.n3129 fc2.n3128 0.016
R15183 fc2.n3109 fc2.n3108 0.016
R15184 fc2.n3058 fc2.n3057 0.016
R15185 fc2.n3038 fc2.n3037 0.016
R15186 fc2.n2944 fc2.n2943 0.016
R15187 fc2.n2893 fc2.n2892 0.016
R15188 fc2.n2873 fc2.n2872 0.016
R15189 fc2.n2853 fc2.n2852 0.016
R15190 fc2.n3172 fc2.n3070 0.016
R15191 fc2.n3159 fc2.n3152 0.016
R15192 fc2.n3139 fc2.n3132 0.016
R15193 fc2.n3119 fc2.n3112 0.016
R15194 fc2.n3061 fc2.n2999 0.016
R15195 fc2.n3048 fc2.n3041 0.016
R15196 fc2.n2947 fc2.n2905 0.016
R15197 fc2.n2896 fc2.n2814 0.016
R15198 fc2.n2883 fc2.n2876 0.016
R15199 fc2.n2863 fc2.n2856 0.016
R15200 fc2.n3568 fc2.n3567 0.016
R15201 fc2.n3557 fc2.n3556 0.016
R15202 fc2.n3547 fc2.n3546 0.016
R15203 fc2.n3537 fc2.n3536 0.016
R15204 fc2.n3527 fc2.n3526 0.016
R15205 fc2.n3517 fc2.n3516 0.016
R15206 fc2.n3507 fc2.n3506 0.016
R15207 fc2.n3497 fc2.n3496 0.016
R15208 fc2.n3487 fc2.n3486 0.016
R15209 fc2.n3958 fc2.n3957 0.016
R15210 fc2.n3948 fc2.n3947 0.016
R15211 fc2.n3938 fc2.n3937 0.016
R15212 fc2.n3928 fc2.n3927 0.016
R15213 fc2.n3918 fc2.n3917 0.016
R15214 fc2.n3908 fc2.n3907 0.016
R15215 fc2.n3898 fc2.n3897 0.016
R15216 fc2.n3668 fc2.n3667 0.016
R15217 fc2.n3657 fc2.n3656 0.016
R15218 fc2.n3647 fc2.n3646 0.016
R15219 fc2.n3637 fc2.n3636 0.016
R15220 fc2.n3627 fc2.n3626 0.016
R15221 fc2.n3835 fc2.n3834 0.016
R15222 fc2.n3825 fc2.n3824 0.016
R15223 fc2.n3815 fc2.n3814 0.016
R15224 fc2.n3696 fc2.n3687 0.016
R15225 fc2.n3317 fc2.n3316 0.015
R15226 fc2.n1558 fc2.n1557 0.015
R15227 fc2.n1634 fc2.n1633 0.015
R15228 fc2.n578 fc2.n577 0.015
R15229 fc2.n3358 fc2.n3357 0.015
R15230 fc2.n3456 fc2.n3455 0.015
R15231 fc2.n3466 fc2.n3465 0.015
R15232 fc2.n3885 fc2.n3884 0.015
R15233 fc2.n3875 fc2.n3874 0.015
R15234 fc2.n3596 fc2.n3595 0.015
R15235 fc2.n3606 fc2.n3605 0.015
R15236 fc2.n3802 fc2.n3801 0.015
R15237 fc2.n3792 fc2.n3791 0.015
R15238 fc2.n3718 fc2.n3717 0.015
R15239 fc2.n3698 fc2.n3697 0.015
R15240 fc2.n3301 fc2.n3178 0.015
R15241 fc2.n3303 fc2.n3302 0.015
R15242 fc2.n529 fc2.n528 0.015
R15243 fc2.n2694 fc2.n2686 0.014
R15244 fc2.t4 fc2.n2629 0.014
R15245 fc2.t14 fc2.n44 0.014
R15246 fc2.t14 fc2.n39 0.014
R15247 fc2.n2761 fc2.n2760 0.014
R15248 fc2.n2452 fc2.n2447 0.014
R15249 fc2.n2450 fc2.n2449 0.014
R15250 fc2.n2190 fc2.n2186 0.014
R15251 fc2.n264 fc2.n263 0.014
R15252 fc2.n377 fc2.n376 0.014
R15253 fc2.n2181 fc2.n2180 0.014
R15254 fc2.n2188 fc2.n2187 0.014
R15255 fc2.n1781 fc2.n1780 0.014
R15256 fc2.n957 fc2.n956 0.014
R15257 fc2.n728 fc2.n727 0.014
R15258 fc2.n2340 fc2.n2339 0.014
R15259 fc2.n2100 fc2.n2099 0.014
R15260 fc2.n453 fc2.n452 0.014
R15261 fc2.n200 fc2.n199 0.014
R15262 fc2.n566 fc2.n562 0.014
R15263 fc2.n229 fc2.n228 0.014
R15264 fc2.n411 fc2.n410 0.014
R15265 fc2.n2133 fc2.n2132 0.014
R15266 fc2.n2384 fc2.n2383 0.014
R15267 fc2.n758 fc2.n757 0.014
R15268 fc2.n564 fc2.n563 0.014
R15269 fc2.n119 fc2.n114 0.014
R15270 fc2.n117 fc2.n116 0.014
R15271 fc2.n3445 fc2.n2807 0.014
R15272 fc2.n3445 fc2.n3308 0.014
R15273 fc2.n1455 fc2.n1454 0.014
R15274 fc2.n1937 fc2.n1936 0.014
R15275 fc2.n1156 fc2.n1155 0.014
R15276 fc2.n915 fc2.n914 0.014
R15277 fc2.n1730 fc2.n1729 0.014
R15278 fc2.n1583 fc2.n1582 0.014
R15279 fc2.n1210 fc2.n1209 0.014
R15280 fc2.n2301 fc2.n2300 0.014
R15281 fc2.n673 fc2.n672 0.014
R15282 fc2.n603 fc2.n602 0.014
R15283 fc2.n1622 fc2.n1621 0.014
R15284 fc2.n1659 fc2.n1658 0.014
R15285 fc2.n1288 fc2.n1287 0.014
R15286 fc2.n496 fc2.n495 0.014
R15287 fc2.n2045 fc2.n2044 0.014
R15288 fc2.n2228 fc2.n2227 0.014
R15289 fc2.n808 fc2.n807 0.014
R15290 fc2.n846 fc2.n845 0.014
R15291 fc2.n1831 fc2.n1830 0.014
R15292 fc2.n1869 fc2.n1868 0.014
R15293 fc2.n1366 fc2.n1365 0.014
R15294 fc2.n3584 fc2.n3446 0.014
R15295 fc2.n3684 fc2.n3586 0.014
R15296 fc2.n3744 fc2.n3686 0.014
R15297 fc2.n352 fc2.n351 0.014
R15298 fc2.n428 fc2.n427 0.014
R15299 fc2.n2315 fc2.n2314 0.014
R15300 fc2.n932 fc2.n931 0.014
R15301 fc2.n983 fc2.n982 0.014
R15302 fc2.n2410 fc2.n2409 0.014
R15303 fc2.n2359 fc2.n2358 0.014
R15304 fc2.n1844 fc2.n1843 0.014
R15305 fc2.n821 fc2.n820 0.014
R15306 fc2.n2203 fc2.n2202 0.014
R15307 fc2.n1425 fc2.n1424 0.014
R15308 fc2.n1888 fc2.n1887 0.014
R15309 fc2.n865 fc2.n864 0.014
R15310 fc2.n2250 fc2.n2249 0.014
R15311 fc2.n516 fc2.n515 0.014
R15312 fc2.n3337 fc2.n3321 0.014
R15313 fc2.n3337 fc2.n3328 0.014
R15314 fc2.n1211 fc2.n1072 0.014
R15315 fc2.n1289 fc2.n1260 0.014
R15316 fc2.n1062 fc2.n1061 0.014
R15317 fc2.n1250 fc2.n1249 0.014
R15318 fc2.n1328 fc2.n1327 0.014
R15319 fc2.n1406 fc2.n1405 0.014
R15320 fc2.n314 fc2.n121 0.013
R15321 fc2.n3415 fc2.n3414 0.013
R15322 fc2.n1494 fc2.n1488 0.013
R15323 fc2.n3415 fc2.n3412 0.013
R15324 fc2.n3404 fc2.n3399 0.013
R15325 fc2.n3387 fc2.n3385 0.013
R15326 fc2.n3375 fc2.n3372 0.013
R15327 fc2.n3347 fc2.n3346 0.013
R15328 fc2.n1371 fc2.n1369 0.013
R15329 fc2.n3360 fc2.n3356 0.013
R15330 fc2.t56 fc2.n3427 0.013
R15331 fc2.n532 fc2.n530 0.013
R15332 fc2.n3432 fc2.n3431 0.013
R15333 fc2.n73 fc2.n72 0.013
R15334 fc2.n102 fc2.n101 0.013
R15335 fc2.n1464 fc2.n1450 0.012
R15336 fc2.n1173 fc2.n1172 0.012
R15337 fc2.n1050 fc2.n1048 0.012
R15338 fc2.n1238 fc2.n1236 0.012
R15339 fc2.n1316 fc2.n1314 0.012
R15340 fc2.n1394 fc2.n1392 0.012
R15341 fc2.n2738 fc2.n2737 0.012
R15342 fc2.n263 fc2.n262 0.012
R15343 fc2.n376 fc2.n375 0.012
R15344 fc2.n2180 fc2.n2179 0.012
R15345 fc2.n1780 fc2.n1779 0.012
R15346 fc2.n956 fc2.n955 0.012
R15347 fc2.n727 fc2.n726 0.012
R15348 fc2.n2339 fc2.n2338 0.012
R15349 fc2.n2099 fc2.n2098 0.012
R15350 fc2.n452 fc2.n451 0.012
R15351 fc2.n199 fc2.n198 0.012
R15352 fc2.n228 fc2.n227 0.012
R15353 fc2.n410 fc2.n409 0.012
R15354 fc2.n2132 fc2.n2131 0.012
R15355 fc2.n2383 fc2.n2382 0.012
R15356 fc2.n757 fc2.n756 0.012
R15357 fc2.n2528 fc2.n2527 0.012
R15358 fc2.n308 fc2.n307 0.012
R15359 fc2.n2602 fc2.n2601 0.012
R15360 fc2.n1936 fc2.n1935 0.012
R15361 fc2.n1155 fc2.n1154 0.012
R15362 fc2.n914 fc2.n913 0.012
R15363 fc2.n1729 fc2.n1728 0.012
R15364 fc2.n1582 fc2.n1581 0.012
R15365 fc2.n1209 fc2.n1208 0.012
R15366 fc2.n2300 fc2.n2299 0.012
R15367 fc2.n672 fc2.n671 0.012
R15368 fc2.n602 fc2.n601 0.012
R15369 fc2.n1621 fc2.n1620 0.012
R15370 fc2.n1658 fc2.n1657 0.012
R15371 fc2.n1287 fc2.n1286 0.012
R15372 fc2.n495 fc2.n494 0.012
R15373 fc2.n2044 fc2.n2043 0.012
R15374 fc2.n2227 fc2.n2226 0.012
R15375 fc2.n807 fc2.n806 0.012
R15376 fc2.n845 fc2.n844 0.012
R15377 fc2.n1830 fc2.n1829 0.012
R15378 fc2.n1868 fc2.n1867 0.012
R15379 fc2.n1365 fc2.n1364 0.012
R15380 fc2.n265 fc2.n264 0.012
R15381 fc2.n378 fc2.n377 0.012
R15382 fc2.n2182 fc2.n2181 0.012
R15383 fc2.n378 fc2.n345 0.012
R15384 fc2.n265 fc2.n241 0.012
R15385 fc2.n1981 fc2.n1980 0.012
R15386 fc2.n201 fc2.n177 0.012
R15387 fc2.n454 fc2.n422 0.012
R15388 fc2.n2101 fc2.n2078 0.012
R15389 fc2.n2341 fc2.n2309 0.012
R15390 fc2.n729 fc2.n706 0.012
R15391 fc2.n958 fc2.n926 0.012
R15392 fc2.n1782 fc2.n1781 0.012
R15393 fc2.n958 fc2.n957 0.012
R15394 fc2.n729 fc2.n728 0.012
R15395 fc2.n2341 fc2.n2340 0.012
R15396 fc2.n2101 fc2.n2100 0.012
R15397 fc2.n454 fc2.n453 0.012
R15398 fc2.n201 fc2.n200 0.012
R15399 fc2.n281 fc2.n273 0.012
R15400 fc2.n335 fc2.n321 0.012
R15401 fc2.n2151 fc2.n2142 0.012
R15402 fc2.n2415 fc2.n2396 0.012
R15403 fc2.n778 fc2.n767 0.012
R15404 fc2.n988 fc2.n969 0.012
R15405 fc2.n1801 fc2.n1790 0.012
R15406 fc2.n1966 fc2.n1950 0.012
R15407 fc2.n1179 fc2.n1165 0.012
R15408 fc2.n1801 fc2.n1800 0.012
R15409 fc2.n988 fc2.n987 0.012
R15410 fc2.n778 fc2.n777 0.012
R15411 fc2.n2415 fc2.n2414 0.012
R15412 fc2.n2151 fc2.n2150 0.012
R15413 fc2.n412 fc2.n411 0.012
R15414 fc2.n2134 fc2.n2133 0.012
R15415 fc2.n2385 fc2.n2384 0.012
R15416 fc2.n759 fc2.n758 0.012
R15417 fc2.n2385 fc2.n2352 0.012
R15418 fc2.n2134 fc2.n2111 0.012
R15419 fc2.n231 fc2.n229 0.012
R15420 fc2.n1449 fc2.n1447 0.012
R15421 fc2.n1490 fc2.n1489 0.012
R15422 fc2.n1488 fc2.n1487 0.012
R15423 fc2.n1938 fc2.n1937 0.012
R15424 fc2.n1157 fc2.n1156 0.012
R15425 fc2.n916 fc2.n915 0.012
R15426 fc2.n1731 fc2.n1730 0.012
R15427 fc2.n1584 fc2.n1583 0.012
R15428 fc2.n1211 fc2.n1210 0.012
R15429 fc2.n2302 fc2.n2301 0.012
R15430 fc2.n674 fc2.n673 0.012
R15431 fc2.n604 fc2.n603 0.012
R15432 fc2.n1623 fc2.n1622 0.012
R15433 fc2.n1660 fc2.n1659 0.012
R15434 fc2.n1289 fc2.n1288 0.012
R15435 fc2.n1407 fc2.n1371 0.012
R15436 fc2.n1870 fc2.n1837 0.012
R15437 fc2.n1832 fc2.n1669 0.012
R15438 fc2.n847 fc2.n814 0.012
R15439 fc2.n809 fc2.n613 0.012
R15440 fc2.n2229 fc2.n2196 0.012
R15441 fc2.n2046 fc2.n2023 0.012
R15442 fc2.n497 fc2.n467 0.012
R15443 fc2.n497 fc2.n496 0.012
R15444 fc2.n2046 fc2.n2045 0.012
R15445 fc2.n2229 fc2.n2228 0.012
R15446 fc2.n809 fc2.n808 0.012
R15447 fc2.n847 fc2.n846 0.012
R15448 fc2.n1832 fc2.n1831 0.012
R15449 fc2.n1870 fc2.n1869 0.012
R15450 fc2.n1367 fc2.n1366 0.012
R15451 fc2.n3454 fc2.n3453 0.012
R15452 fc2.n3969 fc2.n3968 0.012
R15453 fc2.n3594 fc2.n3593 0.012
R15454 fc2.n3846 fc2.n3845 0.012
R15455 fc2.n3730 fc2.n3729 0.012
R15456 fc2.n1438 fc2.n1418 0.012
R15457 fc2.n1125 fc2.n1113 0.012
R15458 fc2.n1899 fc2.n1881 0.012
R15459 fc2.n1752 fc2.n1740 0.012
R15460 fc2.n876 fc2.n858 0.012
R15461 fc2.n695 fc2.n683 0.012
R15462 fc2.n2261 fc2.n2243 0.012
R15463 fc2.n2067 fc2.n2055 0.012
R15464 fc2.n533 fc2.n509 0.012
R15465 fc2.n166 fc2.n153 0.012
R15466 fc2.n166 fc2.n165 0.012
R15467 fc2.n533 fc2.n532 0.012
R15468 fc2.n2067 fc2.n2066 0.012
R15469 fc2.n2261 fc2.n2260 0.012
R15470 fc2.n695 fc2.n694 0.012
R15471 fc2.n876 fc2.n875 0.012
R15472 fc2.n1752 fc2.n1751 0.012
R15473 fc2.n1899 fc2.n1898 0.012
R15474 fc2.n1125 fc2.n1124 0.012
R15475 fc2.n1438 fc2.n1437 0.012
R15476 fc2.n1464 fc2.n1463 0.012
R15477 fc2.n3326 fc2.n3325 0.012
R15478 fc2.n3324 fc2.n3323 0.012
R15479 fc2.n3319 fc2.n3318 0.012
R15480 fc2.n1984 fc2.n1982 0.012
R15481 fc2.n1220 fc2.n1219 0.012
R15482 fc2.n1298 fc2.n1297 0.012
R15483 fc2.n1376 fc2.n1375 0.012
R15484 fc2.n71 fc2.n70 0.012
R15485 fc2.n69 fc2.n68 0.012
R15486 fc2.n67 fc2.n66 0.012
R15487 fc2.n100 fc2.n99 0.012
R15488 fc2.n98 fc2.n97 0.012
R15489 fc2.n96 fc2.n95 0.012
R15490 fc2.n94 fc2.n93 0.012
R15491 fc2.n1529 fc2.n1528 0.011
R15492 fc2.n3189 fc2.n3188 0.011
R15493 fc2.n3172 fc2.n3171 0.011
R15494 fc2.n3160 fc2.n3159 0.011
R15495 fc2.n3140 fc2.n3139 0.011
R15496 fc2.n3120 fc2.n3119 0.011
R15497 fc2.n3100 fc2.n3099 0.011
R15498 fc2.n3090 fc2.n3089 0.011
R15499 fc2.n3061 fc2.n3060 0.011
R15500 fc2.n3049 fc2.n3048 0.011
R15501 fc2.n3029 fc2.n3028 0.011
R15502 fc2.n3019 fc2.n3018 0.011
R15503 fc2.n2976 fc2.n2975 0.011
R15504 fc2.n2985 fc2.n2984 0.011
R15505 fc2.n2947 fc2.n2946 0.011
R15506 fc2.n2935 fc2.n2934 0.011
R15507 fc2.n2925 fc2.n2924 0.011
R15508 fc2.n2896 fc2.n2895 0.011
R15509 fc2.n2884 fc2.n2883 0.011
R15510 fc2.n2864 fc2.n2863 0.011
R15511 fc2.n2844 fc2.n2843 0.011
R15512 fc2.n2834 fc2.n2833 0.011
R15513 fc2.n3487 fc2.n3479 0.011
R15514 fc2.n3497 fc2.n3489 0.011
R15515 fc2.n3507 fc2.n3499 0.011
R15516 fc2.n3517 fc2.n3509 0.011
R15517 fc2.n3527 fc2.n3519 0.011
R15518 fc2.n3537 fc2.n3529 0.011
R15519 fc2.n3547 fc2.n3539 0.011
R15520 fc2.n3557 fc2.n3549 0.011
R15521 fc2.n3568 fc2.n3560 0.011
R15522 fc2.n3899 fc2.n3898 0.011
R15523 fc2.n3909 fc2.n3908 0.011
R15524 fc2.n3919 fc2.n3918 0.011
R15525 fc2.n3929 fc2.n3928 0.011
R15526 fc2.n3939 fc2.n3938 0.011
R15527 fc2.n3949 fc2.n3948 0.011
R15528 fc2.n3959 fc2.n3958 0.011
R15529 fc2.n3627 fc2.n3619 0.011
R15530 fc2.n3637 fc2.n3629 0.011
R15531 fc2.n3647 fc2.n3639 0.011
R15532 fc2.n3657 fc2.n3649 0.011
R15533 fc2.n3668 fc2.n3660 0.011
R15534 fc2.n3816 fc2.n3815 0.011
R15535 fc2.n3826 fc2.n3825 0.011
R15536 fc2.n3836 fc2.n3835 0.011
R15537 fc2.n3696 fc2.n3695 0.011
R15538 fc2.n3200 fc2.n3199 0.011
R15539 fc2.n3210 fc2.n3209 0.011
R15540 fc2.n3220 fc2.n3219 0.011
R15541 fc2.n3230 fc2.n3229 0.011
R15542 fc2.n3240 fc2.n3239 0.011
R15543 fc2.n3250 fc2.n3249 0.011
R15544 fc2.n3260 fc2.n3259 0.011
R15545 fc2.n3270 fc2.n3269 0.011
R15546 fc2.n3280 fc2.n3279 0.011
R15547 fc2.n3290 fc2.n3289 0.011
R15548 fc2.n3300 fc2.n3299 0.011
R15549 fc2.n3411 fc2.n3410 0.011
R15550 fc2.n1962 fc2.n1961 0.011
R15551 fc2.t56 fc2.n3392 0.011
R15552 fc2.n65 fc2.n64 0.011
R15553 fc2.n527 fc2.n526 0.011
R15554 fc2.n1461 fc2.n1457 0.011
R15555 fc2.n2652 fc2.n2645 0.011
R15556 fc2.n3170 fc2.n3169 0.01
R15557 fc2.n3150 fc2.n3149 0.01
R15558 fc2.n3130 fc2.n3129 0.01
R15559 fc2.n3110 fc2.n3109 0.01
R15560 fc2.n3059 fc2.n3058 0.01
R15561 fc2.n3039 fc2.n3038 0.01
R15562 fc2.n2945 fc2.n2944 0.01
R15563 fc2.n2894 fc2.n2893 0.01
R15564 fc2.n2874 fc2.n2873 0.01
R15565 fc2.n2854 fc2.n2853 0.01
R15566 fc2.n1221 fc2.n1220 0.01
R15567 fc2.n1299 fc2.n1298 0.01
R15568 fc2.n1105 fc2.n1092 0.01
R15569 fc2.n1698 fc2.n1690 0.01
R15570 fc2.n641 fc2.n633 0.01
R15571 fc2.n2014 fc2.n2006 0.01
R15572 fc2.n144 fc2.n136 0.01
R15573 fc2.n2652 fc2.n2651 0.01
R15574 fc2.n1494 fc2.n1467 0.01
R15575 fc2.n3311 fc2.n3310 0.01
R15576 fc2.n3312 fc2.n3311 0.01
R15577 fc2.n3313 fc2.n3312 0.01
R15578 fc2.n3444 fc2.n3313 0.01
R15579 fc2.n3310 fc2.n3309 0.01
R15580 fc2.n3069 fc2.n3068 0.01
R15581 fc2.n2998 fc2.n2997 0.01
R15582 fc2.n2967 fc2.n2962 0.01
R15583 fc2.n2904 fc2.n2903 0.01
R15584 fc2.n2813 fc2.n2812 0.01
R15585 fc2.n1436 fc2.n1435 0.01
R15586 fc2.n705 fc2.n704 0.01
R15587 fc2.n2077 fc2.n2076 0.01
R15588 fc2.n176 fc2.n175 0.01
R15589 fc2.n1706 fc2.n1705 0.01
R15590 fc2.n1592 fc2.n1591 0.01
R15591 fc2.n649 fc2.n648 0.01
R15592 fc2.n1463 fc2.n1462 0.01
R15593 fc2.n3708 fc2.n3707 0.009
R15594 fc2.n1377 fc2.n1376 0.009
R15595 fc2.n2740 fc2.n2739 0.009
R15596 fc2.n2718 fc2.n2709 0.009
R15597 fc2.n2575 fc2.n2573 0.009
R15598 fc2.n2507 fc2.n2506 0.009
R15599 fc2.n2765 fc2.n2763 0.009
R15600 fc2.n2766 fc2.n2765 0.009
R15601 fc2.n2540 fc2.n2529 0.009
R15602 fc2.n2608 fc2.n2603 0.009
R15603 fc2.n314 fc2.n309 0.009
R15604 fc2.n1938 fc2.n1912 0.009
R15605 fc2.n1055 fc2.n1050 0.009
R15606 fc2.n1046 fc2.n1045 0.009
R15607 fc2.n1251 fc2.n1215 0.009
R15608 fc2.n1584 fc2.n1552 0.009
R15609 fc2.n1552 fc2.n1550 0.009
R15610 fc2.n1731 fc2.n1707 0.009
R15611 fc2.n916 fc2.n889 0.009
R15612 fc2.n1243 fc2.n1238 0.009
R15613 fc2.n1234 fc2.n1233 0.009
R15614 fc2.n1329 fc2.n1293 0.009
R15615 fc2.n1660 fc2.n1628 0.009
R15616 fc2.n1628 fc2.n1626 0.009
R15617 fc2.n1623 fc2.n1593 0.009
R15618 fc2.n604 fc2.n572 0.009
R15619 fc2.n572 fc2.n570 0.009
R15620 fc2.n674 fc2.n650 0.009
R15621 fc2.n2302 fc2.n2271 0.009
R15622 fc2.n1321 fc2.n1316 0.009
R15623 fc2.n1312 fc2.n1311 0.009
R15624 fc2.n3346 fc2.n3343 0.009
R15625 fc2.n3348 fc2.n3347 0.009
R15626 fc2.n1399 fc2.n1394 0.009
R15627 fc2.n1390 fc2.n1389 0.009
R15628 fc2.n2472 fc2.n2457 0.009
R15629 fc2.n2472 fc2.n2471 0.009
R15630 fc2.n3431 fc2.n3430 0.009
R15631 fc2.n3433 fc2.n3432 0.009
R15632 fc2.n1063 fc2.n1062 0.009
R15633 fc2.n1251 fc2.n1250 0.009
R15634 fc2.n1329 fc2.n1328 0.009
R15635 fc2.n1407 fc2.n1406 0.009
R15636 fc2.n2575 fc2.n2547 0.009
R15637 fc2.n2507 fc2.n2480 0.009
R15638 fc2.n412 fc2.n386 0.009
R15639 fc2.n2540 fc2.n2539 0.009
R15640 fc2.n2608 fc2.n2607 0.009
R15641 fc2.n3477 fc2.n3476 0.009
R15642 fc2.n3888 fc2.n3887 0.009
R15643 fc2.n3617 fc2.n3616 0.009
R15644 fc2.n3805 fc2.n3804 0.009
R15645 fc2.n3985 fc2.n3984 0.009
R15646 fc2.n3862 fc2.n3861 0.009
R15647 fc2.n3984 fc2.n3864 0.009
R15648 fc2.n3861 fc2.n3781 0.009
R15649 fc2.n759 fc2.n737 0.008
R15650 fc2.n1178 fc2.n1177 0.008
R15651 fc2.n1493 fc2.n1492 0.008
R15652 fc2.n345 fc2.n343 0.008
R15653 fc2.n422 fc2.n420 0.008
R15654 fc2.n2309 fc2.n2307 0.008
R15655 fc2.n926 fc2.n924 0.008
R15656 fc2.n273 fc2.n272 0.008
R15657 fc2.n321 fc2.n320 0.008
R15658 fc2.n2142 fc2.n2141 0.008
R15659 fc2.n2396 fc2.n2395 0.008
R15660 fc2.n767 fc2.n766 0.008
R15661 fc2.n969 fc2.n968 0.008
R15662 fc2.n1790 fc2.n1789 0.008
R15663 fc2.n1950 fc2.n1949 0.008
R15664 fc2.n987 fc2.n985 0.008
R15665 fc2.n2414 fc2.n2412 0.008
R15666 fc2.n2352 fc2.n2350 0.008
R15667 fc2.n1060 fc2.n1059 0.008
R15668 fc2.n1248 fc2.n1247 0.008
R15669 fc2.n1326 fc2.n1325 0.008
R15670 fc2.n1837 fc2.n1835 0.008
R15671 fc2.n814 fc2.n812 0.008
R15672 fc2.n2196 fc2.n2194 0.008
R15673 fc2.n1404 fc2.n1403 0.008
R15674 fc2.n1418 fc2.n1416 0.008
R15675 fc2.n1881 fc2.n1879 0.008
R15676 fc2.n858 fc2.n856 0.008
R15677 fc2.n2243 fc2.n2241 0.008
R15678 fc2.n509 fc2.n507 0.008
R15679 fc2.n3387 fc2.n3386 0.008
R15680 fc2.n3375 fc2.n3374 0.008
R15681 fc2.n1219 fc2.n1217 0.008
R15682 fc2.n1297 fc2.n1295 0.008
R15683 fc2.n1375 fc2.n1373 0.008
R15684 fc2.n3477 fc2.n3468 0.008
R15685 fc2.n3889 fc2.n3888 0.008
R15686 fc2.n3617 fc2.n3608 0.008
R15687 fc2.n3806 fc2.n3805 0.008
R15688 fc2.n3708 fc2.n3700 0.008
R15689 fc2.n3988 fc2.n3987 0.008
R15690 fc2.n1985 fc2.n1984 0.007
R15691 fc2.n3464 fc2.n3458 0.007
R15692 fc2.n3464 fc2.n3463 0.007
R15693 fc2.n3873 fc2.n3868 0.007
R15694 fc2.n3873 fc2.n3872 0.007
R15695 fc2.n3604 fc2.n3598 0.007
R15696 fc2.n3604 fc2.n3603 0.007
R15697 fc2.n3790 fc2.n3785 0.007
R15698 fc2.n3790 fc2.n3789 0.007
R15699 fc2.n3719 fc2.n3715 0.007
R15700 fc2.n3719 fc2.n3710 0.007
R15701 fc2.n1057 fc2.n1056 0.007
R15702 fc2.n1245 fc2.n1244 0.007
R15703 fc2.n1323 fc2.n1322 0.007
R15704 fc2.n1401 fc2.n1400 0.007
R15705 fc2.n1511 fc2.n1507 0.007
R15706 fc2.n2777 fc2.n2776 0.007
R15707 fc2.n2182 fc2.n1988 0.007
R15708 fc2.n281 fc2.n280 0.007
R15709 fc2.n231 fc2.n208 0.007
R15710 fc2.n2185 fc2.n2184 0.006
R15711 fc2.n2573 fc2.n2562 0.006
R15712 fc2.n264 fc2.n257 0.006
R15713 fc2.n377 fc2.n368 0.006
R15714 fc2.n2181 fc2.n2174 0.006
R15715 fc2.n1781 fc2.n1774 0.006
R15716 fc2.n957 fc2.n948 0.006
R15717 fc2.n728 fc2.n721 0.006
R15718 fc2.n2340 fc2.n2331 0.006
R15719 fc2.n2100 fc2.n2093 0.006
R15720 fc2.n453 fc2.n444 0.006
R15721 fc2.n200 fc2.n193 0.006
R15722 fc2.n2506 fc2.n2495 0.006
R15723 fc2.n561 fc2.n560 0.006
R15724 fc2.n229 fc2.n222 0.006
R15725 fc2.n411 fc2.n402 0.006
R15726 fc2.n2133 fc2.n2126 0.006
R15727 fc2.n2384 fc2.n2375 0.006
R15728 fc2.n758 fc2.n751 0.006
R15729 fc2.n2529 fc2.n2520 0.006
R15730 fc2.n309 fc2.n305 0.006
R15731 fc2.n2603 fc2.n2594 0.006
R15732 fc2.n1937 fc2.n1928 0.006
R15733 fc2.n1156 fc2.n1148 0.006
R15734 fc2.n915 fc2.n906 0.006
R15735 fc2.n1730 fc2.n1723 0.006
R15736 fc2.n1583 fc2.n1574 0.006
R15737 fc2.n1210 fc2.n1202 0.006
R15738 fc2.n2301 fc2.n2292 0.006
R15739 fc2.n673 fc2.n666 0.006
R15740 fc2.n603 fc2.n594 0.006
R15741 fc2.n1622 fc2.n1615 0.006
R15742 fc2.n1659 fc2.n1650 0.006
R15743 fc2.n1288 fc2.n1280 0.006
R15744 fc2.n496 fc2.n487 0.006
R15745 fc2.n2045 fc2.n2038 0.006
R15746 fc2.n2228 fc2.n2219 0.006
R15747 fc2.n808 fc2.n801 0.006
R15748 fc2.n846 fc2.n837 0.006
R15749 fc2.n1831 fc2.n1824 0.006
R15750 fc2.n1869 fc2.n1860 0.006
R15751 fc2.n1366 fc2.n1358 0.006
R15752 fc2.n3427 fc2.n3426 0.006
R15753 fc2.n2570 fc2.n2569 0.006
R15754 fc2.n2706 fc2.n2705 0.006
R15755 fc2.n2500 fc2.n2499 0.006
R15756 fc2.n2667 fc2.n2666 0.006
R15757 fc2.n2684 fc2.n2683 0.006
R15758 fc2.n2627 fc2.n2626 0.006
R15759 fc2.n1099 fc2.n1098 0.006
R15760 fc2.n3176 fc2.n3175 0.006
R15761 fc2.n2760 fc2.n2759 0.006
R15762 fc2.n3099 fc2.n3092 0.006
R15763 fc2.n3028 fc2.n3021 0.006
R15764 fc2.n2976 fc2.n2968 0.006
R15765 fc2.n2934 fc2.n2927 0.006
R15766 fc2.n2843 fc2.n2836 0.006
R15767 fc2.n1062 fc2.n1057 0.006
R15768 fc2.n1250 fc2.n1245 0.006
R15769 fc2.n1328 fc2.n1323 0.006
R15770 fc2.n1406 fc2.n1401 0.006
R15771 fc2.n3089 fc2.n3082 0.005
R15772 fc2.n3018 fc2.n3011 0.005
R15773 fc2.n2985 fc2.n2977 0.005
R15774 fc2.n2924 fc2.n2917 0.005
R15775 fc2.n2833 fc2.n2826 0.005
R15776 fc2.n335 fc2.n334 0.005
R15777 fc2.n1557 fc2.n1556 0.005
R15778 fc2.n1633 fc2.n1632 0.005
R15779 fc2.n577 fc2.n576 0.005
R15780 fc2.n2447 fc2.n2446 0.005
R15781 fc2.n2186 fc2.n2185 0.005
R15782 fc2.n2561 fc2.n2557 0.005
R15783 fc2.n255 fc2.n254 0.005
R15784 fc2.n366 fc2.n365 0.005
R15785 fc2.n2172 fc2.n2171 0.005
R15786 fc2.n1772 fc2.n1771 0.005
R15787 fc2.n946 fc2.n943 0.005
R15788 fc2.n719 fc2.n718 0.005
R15789 fc2.n2329 fc2.n2326 0.005
R15790 fc2.n2091 fc2.n2090 0.005
R15791 fc2.n442 fc2.n439 0.005
R15792 fc2.n191 fc2.n190 0.005
R15793 fc2.n2494 fc2.n2490 0.005
R15794 fc2.n562 fc2.n561 0.005
R15795 fc2.n220 fc2.n219 0.005
R15796 fc2.n400 fc2.n399 0.005
R15797 fc2.n2124 fc2.n2123 0.005
R15798 fc2.n2373 fc2.n2372 0.005
R15799 fc2.n749 fc2.n748 0.005
R15800 fc2.n2519 fc2.n2518 0.005
R15801 fc2.n114 fc2.n113 0.005
R15802 fc2.n304 fc2.n303 0.005
R15803 fc2.n2593 fc2.n2592 0.005
R15804 fc2.n1926 fc2.n1925 0.005
R15805 fc2.n1146 fc2.n1145 0.005
R15806 fc2.n904 fc2.n903 0.005
R15807 fc2.n1721 fc2.n1720 0.005
R15808 fc2.n1572 fc2.n1571 0.005
R15809 fc2.n1200 fc2.n1199 0.005
R15810 fc2.n2290 fc2.n2289 0.005
R15811 fc2.n664 fc2.n663 0.005
R15812 fc2.n592 fc2.n591 0.005
R15813 fc2.n1613 fc2.n1612 0.005
R15814 fc2.n1648 fc2.n1647 0.005
R15815 fc2.n1278 fc2.n1277 0.005
R15816 fc2.n485 fc2.n484 0.005
R15817 fc2.n2036 fc2.n2035 0.005
R15818 fc2.n2217 fc2.n2216 0.005
R15819 fc2.n799 fc2.n798 0.005
R15820 fc2.n835 fc2.n834 0.005
R15821 fc2.n1822 fc2.n1821 0.005
R15822 fc2.n1858 fc2.n1857 0.005
R15823 fc2.n1356 fc2.n1355 0.005
R15824 fc2.n3584 fc2.n3583 0.005
R15825 fc2.n3684 fc2.n3683 0.005
R15826 fc2.n3744 fc2.n3743 0.005
R15827 fc2.n109 fc2.n108 0.005
R15828 fc2.n2777 fc2.n2767 0.005
R15829 fc2.n3199 fc2.n3198 0.005
R15830 fc2.n3360 fc2.n3359 0.005
R15831 fc2.n3437 fc2.n3435 0.005
R15832 fc2.n1177 fc2.n1175 0.005
R15833 fc2.n1709 fc2.n1708 0.005
R15834 fc2.n1595 fc2.n1594 0.005
R15835 fc2.n652 fc2.n651 0.005
R15836 fc2.n1056 fc2.n1055 0.005
R15837 fc2.n1244 fc2.n1243 0.005
R15838 fc2.n1322 fc2.n1321 0.005
R15839 fc2.n1400 fc2.n1399 0.005
R15840 fc2.n58 fc2.n57 0.004
R15841 fc2.n87 fc2.n86 0.004
R15842 fc2.n3964 fc2.n3963 0.004
R15843 fc2.n3976 fc2.n3975 0.004
R15844 fc2.n60 fc2.n59 0.004
R15845 fc2.n89 fc2.n88 0.004
R15846 fc2.n3841 fc2.n3840 0.004
R15847 fc2.n3853 fc2.n3852 0.004
R15848 fc2.n62 fc2.n61 0.004
R15849 fc2.n91 fc2.n90 0.004
R15850 fc2.n301 fc2.n300 0.004
R15851 fc2.n2611 fc2.n2610 0.004
R15852 fc2.n2461 fc2.n2460 0.004
R15853 fc2.n157 fc2.n156 0.004
R15854 fc2.n519 fc2.n518 0.004
R15855 fc2.n2059 fc2.n2058 0.004
R15856 fc2.n2253 fc2.n2252 0.004
R15857 fc2.n687 fc2.n686 0.004
R15858 fc2.n868 fc2.n867 0.004
R15859 fc2.n1744 fc2.n1743 0.004
R15860 fc2.n1891 fc2.n1890 0.004
R15861 fc2.n1117 fc2.n1116 0.004
R15862 fc2.n1428 fc2.n1427 0.004
R15863 fc2.n2728 fc2.n2727 0.004
R15864 fc2.n2790 fc2.n2789 0.004
R15865 fc2.n2717 fc2.n2716 0.004
R15866 fc2.n2550 fc2.n2549 0.004
R15867 fc2.n245 fc2.n244 0.004
R15868 fc2.n355 fc2.n354 0.004
R15869 fc2.n1991 fc2.n1990 0.004
R15870 fc2.n2428 fc2.n2427 0.004
R15871 fc2.n1547 fc2.n1546 0.004
R15872 fc2.n1763 fc2.n1762 0.004
R15873 fc2.n935 fc2.n934 0.004
R15874 fc2.n710 fc2.n709 0.004
R15875 fc2.n2318 fc2.n2317 0.004
R15876 fc2.n2082 fc2.n2081 0.004
R15877 fc2.n431 fc2.n430 0.004
R15878 fc2.n181 fc2.n180 0.004
R15879 fc2.n2483 fc2.n2482 0.004
R15880 fc2.n2662 fc2.n2661 0.004
R15881 fc2.n2620 fc2.n2619 0.004
R15882 fc2.n2770 fc2.n2769 0.004
R15883 fc2.n279 fc2.n278 0.004
R15884 fc2.n331 fc2.n330 0.004
R15885 fc2.n2148 fc2.n2147 0.004
R15886 fc2.n2403 fc2.n2402 0.004
R15887 fc2.n773 fc2.n772 0.004
R15888 fc2.n976 fc2.n975 0.004
R15889 fc2.n1796 fc2.n1795 0.004
R15890 fc2.n1956 fc2.n1955 0.004
R15891 fc2.n1171 fc2.n1170 0.004
R15892 fc2.n1020 fc2.n1019 0.004
R15893 fc2.n2693 fc2.n2692 0.004
R15894 fc2.n2538 fc2.n2537 0.004
R15895 fc2.n211 fc2.n210 0.004
R15896 fc2.n389 fc2.n388 0.004
R15897 fc2.n2115 fc2.n2114 0.004
R15898 fc2.n2362 fc2.n2361 0.004
R15899 fc2.n740 fc2.n739 0.004
R15900 fc2.n1001 fc2.n1000 0.004
R15901 fc2.n1470 fc2.n1469 0.004
R15902 fc2.n1917 fc2.n1916 0.004
R15903 fc2.n1137 fc2.n1136 0.004
R15904 fc2.n1037 fc2.n1036 0.004
R15905 fc2.n894 fc2.n893 0.004
R15906 fc2.n1712 fc2.n1711 0.004
R15907 fc2.n1561 fc2.n1560 0.004
R15908 fc2.n1075 fc2.n1074 0.004
R15909 fc2.n1225 fc2.n1224 0.004
R15910 fc2.n2276 fc2.n2275 0.004
R15911 fc2.n655 fc2.n654 0.004
R15912 fc2.n581 fc2.n580 0.004
R15913 fc2.n1598 fc2.n1597 0.004
R15914 fc2.n1637 fc2.n1636 0.004
R15915 fc2.n1263 fc2.n1262 0.004
R15916 fc2.n1303 fc2.n1302 0.004
R15917 fc2.n474 fc2.n473 0.004
R15918 fc2.n2027 fc2.n2026 0.004
R15919 fc2.n2206 fc2.n2205 0.004
R15920 fc2.n617 fc2.n616 0.004
R15921 fc2.n824 fc2.n823 0.004
R15922 fc2.n1673 fc2.n1672 0.004
R15923 fc2.n1847 fc2.n1846 0.004
R15924 fc2.n1341 fc2.n1340 0.004
R15925 fc2.n1381 fc2.n1380 0.004
R15926 fc2.n293 fc2.n292 0.004
R15927 fc2.n2586 fc2.n2585 0.004
R15928 fc2.n164 fc2.n163 0.004
R15929 fc2.n2673 fc2.n2672 0.004
R15930 fc2.n3404 fc2.n3402 0.004
R15931 fc2.n1061 fc2.n1060 0.004
R15932 fc2.n1249 fc2.n1248 0.004
R15933 fc2.n1327 fc2.n1326 0.004
R15934 fc2.n1405 fc2.n1404 0.004
R15935 fc2.n3582 fc2.n3581 0.004
R15936 fc2.n3682 fc2.n3681 0.004
R15937 fc2.n3742 fc2.n3741 0.004
R15938 fc2.n351 fc2.n350 0.004
R15939 fc2.n427 fc2.n426 0.004
R15940 fc2.n2314 fc2.n2313 0.004
R15941 fc2.n931 fc2.n930 0.004
R15942 fc2.n982 fc2.n981 0.004
R15943 fc2.n2409 fc2.n2408 0.004
R15944 fc2.n2358 fc2.n2357 0.004
R15945 fc2.n1843 fc2.n1842 0.004
R15946 fc2.n820 fc2.n819 0.004
R15947 fc2.n2202 fc2.n2201 0.004
R15948 fc2.n1424 fc2.n1423 0.004
R15949 fc2.n1887 fc2.n1886 0.004
R15950 fc2.n864 fc2.n863 0.004
R15951 fc2.n2249 fc2.n2248 0.004
R15952 fc2.n515 fc2.n514 0.004
R15953 fc2.n2614 fc2.n2583 0.004
R15954 fc2.n297 fc2.n296 0.004
R15955 fc2.n2261 fc2.n2239 0.004
R15956 fc2.n876 fc2.n854 0.004
R15957 fc2.n1899 fc2.n1877 0.004
R15958 fc2.n1438 fc2.n1414 0.004
R15959 fc2.t4 fc2.n2655 0.004
R15960 fc2.t14 fc2.n47 0.004
R15961 fc2.t14 fc2.n41 0.004
R15962 fc2.t14 fc2.n27 0.004
R15963 fc2.t14 fc2.n20 0.004
R15964 fc2.t14 fc2.n34 0.004
R15965 fc2.t56 fc2.n3341 0.004
R15966 fc2.t10 fc2.n1108 0.004
R15967 fc2.t12 fc2.n1701 0.004
R15968 fc2.t52 fc2.n644 0.004
R15969 fc2.t98 fc2.n2017 0.004
R15970 fc2.t66 fc2.n147 0.004
R15971 fc2.n533 fc2.n505 0.004
R15972 fc2.t56 fc2.n3425 0.004
R15973 fc2.t56 fc2.n3408 0.004
R15974 fc2.t56 fc2.n3391 0.004
R15975 fc2.t56 fc2.n3379 0.004
R15976 fc2.t56 fc2.n3364 0.004
R15977 fc2.n2955 fc2.n2950 0.004
R15978 fc2.n1958 fc2.n1957 0.004
R15979 fc2.n1749 fc2.n1748 0.004
R15980 fc2.n1896 fc2.n1895 0.004
R15981 fc2.n1433 fc2.n1432 0.004
R15982 fc2.t14 fc2.n7 0.004
R15983 fc2.t62 fc2.n541 0.004
R15984 fc2.n1986 fc2.n1985 0.004
R15985 fc2.n2775 fc2.n2774 0.004
R15986 fc2.n319 fc2.n318 0.004
R15987 fc2.n2394 fc2.n2393 0.004
R15988 fc2.n967 fc2.n966 0.004
R15989 fc2.n1946 fc2.n1945 0.004
R15990 fc2.n1948 fc2.n1947 0.004
R15991 fc2.n2987 fc2.n2986 0.003
R15992 fc2.n3079 fc2.n3078 0.003
R15993 fc2.n3008 fc2.n3007 0.003
R15994 fc2.n2957 fc2.n2956 0.003
R15995 fc2.n2914 fc2.n2913 0.003
R15996 fc2.n2823 fc2.n2822 0.003
R15997 fc2.n3767 fc2.n3766 0.003
R15998 fc2.n3572 fc2.n3571 0.003
R15999 fc2.n3971 fc2.n3970 0.003
R16000 fc2.n3672 fc2.n3671 0.003
R16001 fc2.n3848 fc2.n3847 0.003
R16002 fc2.n3732 fc2.n3731 0.003
R16003 fc2.n3294 fc2.n3292 0.003
R16004 fc2.n3284 fc2.n3282 0.003
R16005 fc2.n3274 fc2.n3272 0.003
R16006 fc2.n3264 fc2.n3262 0.003
R16007 fc2.n3254 fc2.n3252 0.003
R16008 fc2.n3244 fc2.n3242 0.003
R16009 fc2.n3234 fc2.n3232 0.003
R16010 fc2.n3224 fc2.n3222 0.003
R16011 fc2.n3214 fc2.n3212 0.003
R16012 fc2.n3204 fc2.n3202 0.003
R16013 fc2.n3193 fc2.n3191 0.003
R16014 fc2.n3184 fc2.n3182 0.003
R16015 fc2.n3085 fc2.n3084 0.003
R16016 fc2.n3095 fc2.n3094 0.003
R16017 fc2.n3115 fc2.n3114 0.003
R16018 fc2.n3135 fc2.n3134 0.003
R16019 fc2.n3155 fc2.n3154 0.003
R16020 fc2.n3073 fc2.n3072 0.003
R16021 fc2.n3164 fc2.n3162 0.003
R16022 fc2.n3144 fc2.n3142 0.003
R16023 fc2.n3124 fc2.n3122 0.003
R16024 fc2.n3104 fc2.n3102 0.003
R16025 fc2.n3014 fc2.n3013 0.003
R16026 fc2.n3024 fc2.n3023 0.003
R16027 fc2.n3044 fc2.n3043 0.003
R16028 fc2.n3002 fc2.n3001 0.003
R16029 fc2.n3053 fc2.n3051 0.003
R16030 fc2.n3033 fc2.n3031 0.003
R16031 fc2.n2980 fc2.n2979 0.003
R16032 fc2.n2971 fc2.n2970 0.003
R16033 fc2.n2920 fc2.n2919 0.003
R16034 fc2.n2930 fc2.n2929 0.003
R16035 fc2.n2908 fc2.n2907 0.003
R16036 fc2.n2939 fc2.n2937 0.003
R16037 fc2.n2829 fc2.n2828 0.003
R16038 fc2.n2839 fc2.n2838 0.003
R16039 fc2.n2859 fc2.n2858 0.003
R16040 fc2.n2879 fc2.n2878 0.003
R16041 fc2.n2817 fc2.n2816 0.003
R16042 fc2.n2888 fc2.n2886 0.003
R16043 fc2.n2868 fc2.n2866 0.003
R16044 fc2.n2848 fc2.n2846 0.003
R16045 fc2.n3690 fc2.n3689 0.003
R16046 fc2.n3563 fc2.n3561 0.003
R16047 fc2.n3552 fc2.n3550 0.003
R16048 fc2.n3542 fc2.n3540 0.003
R16049 fc2.n3532 fc2.n3530 0.003
R16050 fc2.n3522 fc2.n3520 0.003
R16051 fc2.n3512 fc2.n3510 0.003
R16052 fc2.n3502 fc2.n3500 0.003
R16053 fc2.n3492 fc2.n3490 0.003
R16054 fc2.n3482 fc2.n3480 0.003
R16055 fc2.n3471 fc2.n3469 0.003
R16056 fc2.n3953 fc2.n3951 0.003
R16057 fc2.n3943 fc2.n3941 0.003
R16058 fc2.n3933 fc2.n3931 0.003
R16059 fc2.n3923 fc2.n3921 0.003
R16060 fc2.n3913 fc2.n3911 0.003
R16061 fc2.n3903 fc2.n3901 0.003
R16062 fc2.n3893 fc2.n3891 0.003
R16063 fc2.n3880 fc2.n3878 0.003
R16064 fc2.n3663 fc2.n3661 0.003
R16065 fc2.n3652 fc2.n3650 0.003
R16066 fc2.n3642 fc2.n3640 0.003
R16067 fc2.n3632 fc2.n3630 0.003
R16068 fc2.n3622 fc2.n3620 0.003
R16069 fc2.n3611 fc2.n3609 0.003
R16070 fc2.n3830 fc2.n3828 0.003
R16071 fc2.n3820 fc2.n3818 0.003
R16072 fc2.n3810 fc2.n3808 0.003
R16073 fc2.n3797 fc2.n3795 0.003
R16074 fc2.n3703 fc2.n3701 0.003
R16075 fc2.n3297 fc2.n3295 0.003
R16076 fc2.n3287 fc2.n3285 0.003
R16077 fc2.n3277 fc2.n3275 0.003
R16078 fc2.n3267 fc2.n3265 0.003
R16079 fc2.n3257 fc2.n3255 0.003
R16080 fc2.n3247 fc2.n3245 0.003
R16081 fc2.n3237 fc2.n3235 0.003
R16082 fc2.n3227 fc2.n3225 0.003
R16083 fc2.n3217 fc2.n3215 0.003
R16084 fc2.n3207 fc2.n3205 0.003
R16085 fc2.n3196 fc2.n3194 0.003
R16086 fc2.n3187 fc2.n3185 0.003
R16087 fc2.n3088 fc2.n3086 0.003
R16088 fc2.n3098 fc2.n3096 0.003
R16089 fc2.n3118 fc2.n3116 0.003
R16090 fc2.n3138 fc2.n3136 0.003
R16091 fc2.n3158 fc2.n3156 0.003
R16092 fc2.n3076 fc2.n3074 0.003
R16093 fc2.n3067 fc2.n3066 0.003
R16094 fc2.n3167 fc2.n3165 0.003
R16095 fc2.n3147 fc2.n3145 0.003
R16096 fc2.n3127 fc2.n3125 0.003
R16097 fc2.n3107 fc2.n3105 0.003
R16098 fc2.n3017 fc2.n3015 0.003
R16099 fc2.n3027 fc2.n3025 0.003
R16100 fc2.n3047 fc2.n3045 0.003
R16101 fc2.n3005 fc2.n3003 0.003
R16102 fc2.n2996 fc2.n2995 0.003
R16103 fc2.n3056 fc2.n3054 0.003
R16104 fc2.n3036 fc2.n3034 0.003
R16105 fc2.n2983 fc2.n2981 0.003
R16106 fc2.n2974 fc2.n2972 0.003
R16107 fc2.n2964 fc2.n2963 0.003
R16108 fc2.n2954 fc2.n2953 0.003
R16109 fc2.n2923 fc2.n2921 0.003
R16110 fc2.n2933 fc2.n2931 0.003
R16111 fc2.n2911 fc2.n2909 0.003
R16112 fc2.n2902 fc2.n2901 0.003
R16113 fc2.n2942 fc2.n2940 0.003
R16114 fc2.n2832 fc2.n2830 0.003
R16115 fc2.n2842 fc2.n2840 0.003
R16116 fc2.n2862 fc2.n2860 0.003
R16117 fc2.n2882 fc2.n2880 0.003
R16118 fc2.n2820 fc2.n2818 0.003
R16119 fc2.n2811 fc2.n2810 0.003
R16120 fc2.n2891 fc2.n2889 0.003
R16121 fc2.n2871 fc2.n2869 0.003
R16122 fc2.n2851 fc2.n2849 0.003
R16123 fc2.n3693 fc2.n3691 0.003
R16124 fc2.n3461 fc2.n3460 0.003
R16125 fc2.n3566 fc2.n3564 0.003
R16126 fc2.n3555 fc2.n3553 0.003
R16127 fc2.n3545 fc2.n3543 0.003
R16128 fc2.n3535 fc2.n3533 0.003
R16129 fc2.n3525 fc2.n3523 0.003
R16130 fc2.n3515 fc2.n3513 0.003
R16131 fc2.n3505 fc2.n3503 0.003
R16132 fc2.n3495 fc2.n3493 0.003
R16133 fc2.n3485 fc2.n3483 0.003
R16134 fc2.n3474 fc2.n3472 0.003
R16135 fc2.n3871 fc2.n3870 0.003
R16136 fc2.n3956 fc2.n3954 0.003
R16137 fc2.n3946 fc2.n3944 0.003
R16138 fc2.n3936 fc2.n3934 0.003
R16139 fc2.n3926 fc2.n3924 0.003
R16140 fc2.n3916 fc2.n3914 0.003
R16141 fc2.n3906 fc2.n3904 0.003
R16142 fc2.n3896 fc2.n3894 0.003
R16143 fc2.n3883 fc2.n3881 0.003
R16144 fc2.n3601 fc2.n3600 0.003
R16145 fc2.n3666 fc2.n3664 0.003
R16146 fc2.n3655 fc2.n3653 0.003
R16147 fc2.n3645 fc2.n3643 0.003
R16148 fc2.n3635 fc2.n3633 0.003
R16149 fc2.n3625 fc2.n3623 0.003
R16150 fc2.n3614 fc2.n3612 0.003
R16151 fc2.n3788 fc2.n3787 0.003
R16152 fc2.n3833 fc2.n3831 0.003
R16153 fc2.n3823 fc2.n3821 0.003
R16154 fc2.n3813 fc2.n3811 0.003
R16155 fc2.n3800 fc2.n3798 0.003
R16156 fc2.n3706 fc2.n3704 0.003
R16157 fc2.n3712 fc2.n3711 0.003
R16158 fc2.n3749 fc2.n3748 0.003
R16159 fc2.n290 fc2.n289 0.003
R16160 fc2.n2617 fc2.n2616 0.003
R16161 fc2.n333 fc2.n332 0.003
R16162 fc2.n1530 fc2.n1529 0.003
R16163 fc2.n2475 fc2.n2474 0.003
R16164 fc2.n172 fc2.n171 0.003
R16165 fc2.n536 fc2.n535 0.003
R16166 fc2.n2073 fc2.n2072 0.003
R16167 fc2.n2264 fc2.n2263 0.003
R16168 fc2.n701 fc2.n700 0.003
R16169 fc2.n882 fc2.n881 0.003
R16170 fc2.n1758 fc2.n1757 0.003
R16171 fc2.n1905 fc2.n1904 0.003
R16172 fc2.n1131 fc2.n1130 0.003
R16173 fc2.n1444 fc2.n1443 0.003
R16174 fc2.n2743 fc2.n2742 0.003
R16175 fc2.n2786 fc2.n2785 0.003
R16176 fc2.n2721 fc2.n2720 0.003
R16177 fc2.n2578 fc2.n2577 0.003
R16178 fc2.n268 fc2.n267 0.003
R16179 fc2.n384 fc2.n383 0.003
R16180 fc2.n2163 fc2.n2162 0.003
R16181 fc2.n2424 fc2.n2423 0.003
R16182 fc2.n1977 fc2.n1976 0.003
R16183 fc2.n1785 fc2.n1784 0.003
R16184 fc2.n961 fc2.n960 0.003
R16185 fc2.n732 fc2.n731 0.003
R16186 fc2.n2344 fc2.n2343 0.003
R16187 fc2.n2104 fc2.n2103 0.003
R16188 fc2.n460 fc2.n459 0.003
R16189 fc2.n204 fc2.n203 0.003
R16190 fc2.n2510 fc2.n2509 0.003
R16191 fc2.n2676 fc2.n2675 0.003
R16192 fc2.n2754 fc2.n2753 0.003
R16193 fc2.n2780 fc2.n2779 0.003
R16194 fc2.n284 fc2.n283 0.003
R16195 fc2.n338 fc2.n337 0.003
R16196 fc2.n2154 fc2.n2153 0.003
R16197 fc2.n2418 fc2.n2417 0.003
R16198 fc2.n781 fc2.n780 0.003
R16199 fc2.n991 fc2.n990 0.003
R16200 fc2.n1804 fc2.n1803 0.003
R16201 fc2.n1969 fc2.n1968 0.003
R16202 fc2.n1182 fc2.n1181 0.003
R16203 fc2.n1505 fc2.n1504 0.003
R16204 fc2.n2697 fc2.n2696 0.003
R16205 fc2.n2543 fc2.n2542 0.003
R16206 fc2.n234 fc2.n233 0.003
R16207 fc2.n418 fc2.n417 0.003
R16208 fc2.n2137 fc2.n2136 0.003
R16209 fc2.n2388 fc2.n2387 0.003
R16210 fc2.n762 fc2.n761 0.003
R16211 fc2.n997 fc2.n996 0.003
R16212 fc2.n1497 fc2.n1496 0.003
R16213 fc2.n1941 fc2.n1940 0.003
R16214 fc2.n1160 fc2.n1159 0.003
R16215 fc2.n1069 fc2.n1068 0.003
R16216 fc2.n919 fc2.n918 0.003
R16217 fc2.n1737 fc2.n1736 0.003
R16218 fc2.n1590 fc2.n1589 0.003
R16219 fc2.n1191 fc2.n1190 0.003
R16220 fc2.n1257 fc2.n1256 0.003
R16221 fc2.n2305 fc2.n2304 0.003
R16222 fc2.n680 fc2.n679 0.003
R16223 fc2.n610 fc2.n609 0.003
R16224 fc2.n1604 fc2.n1603 0.003
R16225 fc2.n1666 fc2.n1665 0.003
R16226 fc2.n1269 fc2.n1268 0.003
R16227 fc2.n1335 fc2.n1334 0.003
R16228 fc2.n503 fc2.n502 0.003
R16229 fc2.n2052 fc2.n2051 0.003
R16230 fc2.n2235 fc2.n2234 0.003
R16231 fc2.n790 fc2.n789 0.003
R16232 fc2.n853 fc2.n852 0.003
R16233 fc2.n1813 fc2.n1812 0.003
R16234 fc2.n1876 fc2.n1875 0.003
R16235 fc2.n1347 fc2.n1346 0.003
R16236 fc2.n1413 fc2.n1412 0.003
R16237 fc2.n2472 fc2.n2464 0.003
R16238 fc2.n166 fc2.n160 0.003
R16239 fc2.n533 fc2.n522 0.003
R16240 fc2.n2067 fc2.n2062 0.003
R16241 fc2.n2261 fc2.n2256 0.003
R16242 fc2.n695 fc2.n690 0.003
R16243 fc2.n876 fc2.n871 0.003
R16244 fc2.n1752 fc2.n1747 0.003
R16245 fc2.n1899 fc2.n1894 0.003
R16246 fc2.n1125 fc2.n1120 0.003
R16247 fc2.n1438 fc2.n1431 0.003
R16248 fc2.n2740 fc2.n2731 0.003
R16249 fc2.n2718 fc2.n2714 0.003
R16250 fc2.n2575 fc2.n2553 0.003
R16251 fc2.n265 fc2.n248 0.003
R16252 fc2.n378 fc2.n358 0.003
R16253 fc2.n2182 fc2.n2166 0.003
R16254 fc2.n1782 fc2.n1766 0.003
R16255 fc2.n958 fc2.n938 0.003
R16256 fc2.n729 fc2.n713 0.003
R16257 fc2.n2341 fc2.n2321 0.003
R16258 fc2.n2101 fc2.n2085 0.003
R16259 fc2.n454 fc2.n434 0.003
R16260 fc2.n201 fc2.n184 0.003
R16261 fc2.n2507 fc2.n2486 0.003
R16262 fc2.n2673 fc2.n2665 0.003
R16263 fc2.n2766 fc2.n2757 0.003
R16264 fc2.n2777 fc2.n2773 0.003
R16265 fc2.n281 fc2.n276 0.003
R16266 fc2.n335 fc2.n325 0.003
R16267 fc2.n2151 fc2.n2145 0.003
R16268 fc2.n2415 fc2.n2400 0.003
R16269 fc2.n778 fc2.n770 0.003
R16270 fc2.n988 fc2.n973 0.003
R16271 fc2.n1801 fc2.n1793 0.003
R16272 fc2.n1966 fc2.n1953 0.003
R16273 fc2.n1179 fc2.n1168 0.003
R16274 fc2.n2694 fc2.n2690 0.003
R16275 fc2.n2540 fc2.n2535 0.003
R16276 fc2.n231 fc2.n214 0.003
R16277 fc2.n412 fc2.n392 0.003
R16278 fc2.n2134 fc2.n2118 0.003
R16279 fc2.n2385 fc2.n2365 0.003
R16280 fc2.n759 fc2.n743 0.003
R16281 fc2.n1494 fc2.n1473 0.003
R16282 fc2.n1938 fc2.n1920 0.003
R16283 fc2.n1157 fc2.n1140 0.003
R16284 fc2.n1063 fc2.n1040 0.003
R16285 fc2.n916 fc2.n897 0.003
R16286 fc2.n1731 fc2.n1715 0.003
R16287 fc2.n1584 fc2.n1564 0.003
R16288 fc2.n1211 fc2.n1194 0.003
R16289 fc2.n1251 fc2.n1228 0.003
R16290 fc2.n2302 fc2.n2282 0.003
R16291 fc2.n674 fc2.n658 0.003
R16292 fc2.n604 fc2.n584 0.003
R16293 fc2.n1623 fc2.n1607 0.003
R16294 fc2.n1660 fc2.n1640 0.003
R16295 fc2.n1289 fc2.n1272 0.003
R16296 fc2.n1329 fc2.n1306 0.003
R16297 fc2.n497 fc2.n477 0.003
R16298 fc2.n2046 fc2.n2030 0.003
R16299 fc2.n2229 fc2.n2209 0.003
R16300 fc2.n809 fc2.n793 0.003
R16301 fc2.n847 fc2.n827 0.003
R16302 fc2.n1832 fc2.n1816 0.003
R16303 fc2.n1870 fc2.n1850 0.003
R16304 fc2.n1367 fc2.n1350 0.003
R16305 fc2.n1407 fc2.n1384 0.003
R16306 fc2.n1179 fc2.n1178 0.003
R16307 fc2.n166 fc2.n150 0.003
R16308 fc2.n2446 fc2.n2445 0.003
R16309 fc2.n113 fc2.n112 0.003
R16310 fc2.t4 fc2.n2634 0.003
R16311 fc2.t4 fc2.n2632 0.003
R16312 fc2.t14 fc2.n9 0.003
R16313 fc2.t56 fc2.n3442 0.003
R16314 fc2.n528 fc2.n527 0.003
R16315 fc2.n3958 fc2.n3950 0.003
R16316 fc2.n3948 fc2.n3940 0.003
R16317 fc2.n3938 fc2.n3930 0.003
R16318 fc2.n3928 fc2.n3920 0.003
R16319 fc2.n3918 fc2.n3910 0.003
R16320 fc2.n3908 fc2.n3900 0.003
R16321 fc2.n3898 fc2.n3890 0.003
R16322 fc2.n3835 fc2.n3827 0.003
R16323 fc2.n3825 fc2.n3817 0.003
R16324 fc2.n3815 fc2.n3807 0.003
R16325 fc2.n3299 fc2.n3291 0.003
R16326 fc2.n3289 fc2.n3281 0.003
R16327 fc2.n3279 fc2.n3271 0.003
R16328 fc2.n3269 fc2.n3261 0.003
R16329 fc2.n3259 fc2.n3251 0.003
R16330 fc2.n3249 fc2.n3241 0.003
R16331 fc2.n3239 fc2.n3231 0.003
R16332 fc2.n3229 fc2.n3221 0.003
R16333 fc2.n3219 fc2.n3211 0.003
R16334 fc2.n3209 fc2.n3201 0.003
R16335 fc2.n3199 fc2.n3190 0.003
R16336 fc2.n3888 fc2.n3877 0.003
R16337 fc2.n3805 fc2.n3794 0.003
R16338 fc2.n3188 fc2.n3181 0.003
R16339 fc2.n3318 fc2.n3317 0.003
R16340 fc2.n3089 fc2.n3077 0.003
R16341 fc2.n3099 fc2.n3091 0.003
R16342 fc2.n3109 fc2.n3101 0.003
R16343 fc2.n3119 fc2.n3111 0.003
R16344 fc2.n3129 fc2.n3121 0.003
R16345 fc2.n3139 fc2.n3131 0.003
R16346 fc2.n3149 fc2.n3141 0.003
R16347 fc2.n3159 fc2.n3151 0.003
R16348 fc2.n3169 fc2.n3161 0.003
R16349 fc2.n3018 fc2.n3006 0.003
R16350 fc2.n3028 fc2.n3020 0.003
R16351 fc2.n3038 fc2.n3030 0.003
R16352 fc2.n3048 fc2.n3040 0.003
R16353 fc2.n3058 fc2.n3050 0.003
R16354 fc2.n2924 fc2.n2912 0.003
R16355 fc2.n2934 fc2.n2926 0.003
R16356 fc2.n2944 fc2.n2936 0.003
R16357 fc2.n2833 fc2.n2821 0.003
R16358 fc2.n2843 fc2.n2835 0.003
R16359 fc2.n2853 fc2.n2845 0.003
R16360 fc2.n2863 fc2.n2855 0.003
R16361 fc2.n2873 fc2.n2865 0.003
R16362 fc2.n2883 fc2.n2875 0.003
R16363 fc2.n2893 fc2.n2885 0.003
R16364 fc2.n72 fc2.n71 0.003
R16365 fc2.n101 fc2.n100 0.003
R16366 fc2.n70 fc2.n69 0.003
R16367 fc2.n99 fc2.n98 0.003
R16368 fc2.n68 fc2.n67 0.003
R16369 fc2.n97 fc2.n96 0.003
R16370 fc2.n66 fc2.n65 0.003
R16371 fc2.n95 fc2.n94 0.003
R16372 fc2.n93 fc2.n92 0.003
R16373 fc2.n3174 fc2.n3069 0.002
R16374 fc2.n3063 fc2.n2998 0.002
R16375 fc2.n2949 fc2.n2904 0.002
R16376 fc2.n2898 fc2.n2813 0.002
R16377 fc2.n3320 fc2.n3319 0.002
R16378 fc2.n3327 fc2.n3326 0.002
R16379 fc2.n3325 fc2.n3324 0.002
R16380 fc2.n3323 fc2.n3322 0.002
R16381 fc2.n3371 fc2.n3370 0.002
R16382 fc2.n3355 fc2.n3354 0.002
R16383 fc2.n2608 fc2.n2606 0.002
R16384 fc2.n2540 fc2.n2532 0.002
R16385 fc2.n231 fc2.n230 0.002
R16386 fc2.n315 fc2.n314 0.002
R16387 fc2.n2575 fc2.n2574 0.002
R16388 fc2.n2562 fc2.n2561 0.002
R16389 fc2.n256 fc2.n255 0.002
R16390 fc2.n367 fc2.n366 0.002
R16391 fc2.n2173 fc2.n2172 0.002
R16392 fc2.n1773 fc2.n1772 0.002
R16393 fc2.n947 fc2.n946 0.002
R16394 fc2.n720 fc2.n719 0.002
R16395 fc2.n2330 fc2.n2329 0.002
R16396 fc2.n2092 fc2.n2091 0.002
R16397 fc2.n443 fc2.n442 0.002
R16398 fc2.n192 fc2.n191 0.002
R16399 fc2.n2495 fc2.n2494 0.002
R16400 fc2.n1509 fc2.n1508 0.002
R16401 fc2.n1510 fc2.n1509 0.002
R16402 fc2.n221 fc2.n220 0.002
R16403 fc2.n401 fc2.n400 0.002
R16404 fc2.n2125 fc2.n2124 0.002
R16405 fc2.n2374 fc2.n2373 0.002
R16406 fc2.n750 fc2.n749 0.002
R16407 fc2.n2520 fc2.n2519 0.002
R16408 fc2.n305 fc2.n304 0.002
R16409 fc2.n2594 fc2.n2593 0.002
R16410 fc2.n1927 fc2.n1926 0.002
R16411 fc2.n1147 fc2.n1146 0.002
R16412 fc2.n905 fc2.n904 0.002
R16413 fc2.n1722 fc2.n1721 0.002
R16414 fc2.n1573 fc2.n1572 0.002
R16415 fc2.n1201 fc2.n1200 0.002
R16416 fc2.n2291 fc2.n2290 0.002
R16417 fc2.n665 fc2.n664 0.002
R16418 fc2.n593 fc2.n592 0.002
R16419 fc2.n1614 fc2.n1613 0.002
R16420 fc2.n1649 fc2.n1648 0.002
R16421 fc2.n1279 fc2.n1278 0.002
R16422 fc2.n486 fc2.n485 0.002
R16423 fc2.n2037 fc2.n2036 0.002
R16424 fc2.n2218 fc2.n2217 0.002
R16425 fc2.n800 fc2.n799 0.002
R16426 fc2.n836 fc2.n835 0.002
R16427 fc2.n1823 fc2.n1822 0.002
R16428 fc2.n1859 fc2.n1858 0.002
R16429 fc2.n1357 fc2.n1356 0.002
R16430 fc2.n3581 fc2.n3570 0.002
R16431 fc2.n3681 fc2.n3670 0.002
R16432 fc2.n64 fc2.n63 0.002
R16433 fc2.n3741 fc2.n3722 0.002
R16434 fc2 fc2.n3445 0.002
R16435 fc2.n2 fc2.n0 0.002
R16436 fc2.n2694 fc2.n2687 0.002
R16437 fc2.t4 fc2.n2630 0.002
R16438 fc2.n80 fc2.n79 0.002
R16439 fc2.n1531 fc2.n1530 0.002
R16440 fc2.n3173 fc2.n3172 0.002
R16441 fc2.n3062 fc2.n3061 0.002
R16442 fc2.n2948 fc2.n2947 0.002
R16443 fc2.n2897 fc2.n2896 0.002
R16444 fc2.n3983 fc2.n3982 0.002
R16445 fc2.n3860 fc2.n3859 0.002
R16446 fc2.n3778 fc2.n3777 0.002
R16447 fc2.n1987 fc2.n1986 0.002
R16448 fc2.n3304 fc2.n3176 0.002
R16449 fc2.n109 fc2.n53 0.002
R16450 fc2.n3781 fc2.n3779 0.002
R16451 fc2.n3987 fc2.n3985 0.002
R16452 fc2.n3864 fc2.n3862 0.002
R16453 fc2.n53 fc2.t14 0.001
R16454 fc2.n2801 fc2.n2800 0.001
R16455 fc2.n554 fc2.n553 0.001
R16456 fc2.n2439 fc2.n2438 0.001
R16457 fc2.n1012 fc2.n1011 0.001
R16458 fc2.n1541 fc2.n1540 0.001
R16459 fc2.n1523 fc2.n1522 0.001
R16460 fc2.n3304 fc2.n3301 0.001
R16461 fc2.n3304 fc2.n3303 0.001
R16462 fc2.n3991 fc2.n3988 0.001
R16463 fc2.n3443 fc2.t56 0.001
R16464 fc2.t14 fc2.n16 0.001
R16465 fc2.t14 fc2.n29 0.001
R16466 fc2.t14 fc2.n52 0.001
R16467 fc2.t56 fc2.n3420 0.001
R16468 fc2.n314 fc2.n313 0.001
R16469 fc2.n2642 fc2.n2641 0.001
R16470 fc2.n133 fc2.n132 0.001
R16471 fc2.n2003 fc2.n2002 0.001
R16472 fc2.n630 fc2.n629 0.001
R16473 fc2.n1687 fc2.n1686 0.001
R16474 fc2.n1089 fc2.n1088 0.001
R16475 fc2.n1910 fc2.n1909 0.001
R16476 fc2.n887 fc2.n886 0.001
R16477 fc2.n2269 fc2.n2268 0.001
R16478 fc2.n465 fc2.n463 0.001
R16479 fc2.n3340 fc2.n3339 0.001
R16480 fc2.n1106 fc2.n1105 0.001
R16481 fc2.n1699 fc2.n1698 0.001
R16482 fc2.n642 fc2.n641 0.001
R16483 fc2.n2015 fc2.n2014 0.001
R16484 fc2.n145 fc2.n144 0.001
R16485 fc2.n2653 fc2.n2652 0.001
R16486 fc2.n559 fc2.n542 0.001
R16487 fc2.n2567 fc2.n2566 0.001
R16488 fc2.n257 fc2.n256 0.001
R16489 fc2.n364 fc2.n363 0.001
R16490 fc2.n368 fc2.n367 0.001
R16491 fc2.n372 fc2.n371 0.001
R16492 fc2.n2174 fc2.n2173 0.001
R16493 fc2.n2560 fc2.n2559 0.001
R16494 fc2.n1774 fc2.n1773 0.001
R16495 fc2.n950 fc2.n949 0.001
R16496 fc2.n948 fc2.n947 0.001
R16497 fc2.n945 fc2.n944 0.001
R16498 fc2.n721 fc2.n720 0.001
R16499 fc2.n2333 fc2.n2332 0.001
R16500 fc2.n2331 fc2.n2330 0.001
R16501 fc2.n2328 fc2.n2327 0.001
R16502 fc2.n2093 fc2.n2092 0.001
R16503 fc2.n446 fc2.n445 0.001
R16504 fc2.n444 fc2.n443 0.001
R16505 fc2.n441 fc2.n440 0.001
R16506 fc2.n193 fc2.n192 0.001
R16507 fc2.n2497 fc2.n2496 0.001
R16508 fc2.n2493 fc2.n2492 0.001
R16509 fc2.n222 fc2.n221 0.001
R16510 fc2.n398 fc2.n397 0.001
R16511 fc2.n402 fc2.n401 0.001
R16512 fc2.n406 fc2.n405 0.001
R16513 fc2.n2126 fc2.n2125 0.001
R16514 fc2.n2371 fc2.n2370 0.001
R16515 fc2.n2375 fc2.n2374 0.001
R16516 fc2.n2379 fc2.n2378 0.001
R16517 fc2.n751 fc2.n750 0.001
R16518 fc2.n2516 fc2.n2515 0.001
R16519 fc2.n2524 fc2.n2523 0.001
R16520 fc2.n2590 fc2.n2589 0.001
R16521 fc2.n2598 fc2.n2597 0.001
R16522 fc2.t56 fc2.n3417 0.001
R16523 fc2.n1492 fc2.n1491 0.001
R16524 fc2.n1480 fc2.n1479 0.001
R16525 fc2.t56 fc2.n3423 0.001
R16526 fc2.n1025 fc2.n1024 0.001
R16527 fc2.n1678 fc2.n1677 0.001
R16528 fc2.n1928 fc2.n1927 0.001
R16529 fc2.n1932 fc2.n1931 0.001
R16530 fc2.n1148 fc2.n1147 0.001
R16531 fc2.t56 fc2.n3406 0.001
R16532 fc2.n906 fc2.n905 0.001
R16533 fc2.n910 fc2.n909 0.001
R16534 fc2.n1723 fc2.n1722 0.001
R16535 fc2.n1570 fc2.n1569 0.001
R16536 fc2.n1574 fc2.n1573 0.001
R16537 fc2.n1578 fc2.n1577 0.001
R16538 fc2.n1202 fc2.n1201 0.001
R16539 fc2.t56 fc2.n3389 0.001
R16540 fc2.n2288 fc2.n2287 0.001
R16541 fc2.n2292 fc2.n2291 0.001
R16542 fc2.n2296 fc2.n2295 0.001
R16543 fc2.n666 fc2.n665 0.001
R16544 fc2.n590 fc2.n589 0.001
R16545 fc2.n594 fc2.n593 0.001
R16546 fc2.n598 fc2.n597 0.001
R16547 fc2.n1615 fc2.n1614 0.001
R16548 fc2.n1646 fc2.n1645 0.001
R16549 fc2.n1650 fc2.n1649 0.001
R16550 fc2.n1654 fc2.n1653 0.001
R16551 fc2.n1280 fc2.n1279 0.001
R16552 fc2.t56 fc2.n3377 0.001
R16553 fc2.n483 fc2.n482 0.001
R16554 fc2.n487 fc2.n486 0.001
R16555 fc2.n491 fc2.n490 0.001
R16556 fc2.n2038 fc2.n2037 0.001
R16557 fc2.n2215 fc2.n2214 0.001
R16558 fc2.n2219 fc2.n2218 0.001
R16559 fc2.n2223 fc2.n2222 0.001
R16560 fc2.n801 fc2.n800 0.001
R16561 fc2.n833 fc2.n832 0.001
R16562 fc2.n837 fc2.n836 0.001
R16563 fc2.n841 fc2.n840 0.001
R16564 fc2.n1824 fc2.n1823 0.001
R16565 fc2.n1856 fc2.n1855 0.001
R16566 fc2.n1860 fc2.n1859 0.001
R16567 fc2.n1864 fc2.n1863 0.001
R16568 fc2.n1358 fc2.n1357 0.001
R16569 fc2.t56 fc2.n3362 0.001
R16570 fc2.n3577 fc2.n3576 0.001
R16571 fc2.n3451 fc2.n3450 0.001
R16572 fc2.n3978 fc2.n3977 0.001
R16573 fc2.n3966 fc2.n3965 0.001
R16574 fc2.n3677 fc2.n3676 0.001
R16575 fc2.n3591 fc2.n3590 0.001
R16576 fc2.n3855 fc2.n3854 0.001
R16577 fc2.n3843 fc2.n3842 0.001
R16578 fc2.n3727 fc2.n3726 0.001
R16579 fc2.n3737 fc2.n3736 0.001
R16580 fc2.n2468 fc2.n2467 0.001
R16581 fc2.n81 fc2.n80 0.001
R16582 fc2.n108 fc2.n107 0.001
R16583 fc2.n298 fc2.n297 0.001
R16584 fc2.t38 fc2.n2614 0.001
R16585 fc2.n2614 fc2.n2613 0.001
R16586 fc2.t56 fc2.n3397 0.001
R16587 fc2.t56 fc2.n3383 0.001
R16588 fc2.t56 fc2.n3368 0.001
R16589 fc2.t56 fc2.n3352 0.001
R16590 fc2.n542 fc2.t62 0.001
R16591 fc2.t4 fc2.n2653 0.001
R16592 fc2.t10 fc2.n1106 0.001
R16593 fc2.t12 fc2.n1699 0.001
R16594 fc2.t52 fc2.n642 0.001
R16595 fc2.t98 fc2.n2015 0.001
R16596 fc2.t66 fc2.n145 0.001
R16597 fc2.t56 fc2.n3340 0.001
R16598 fc2.n465 fc2.n464 0.001
R16599 fc2.t14 fc2.n32 0.001
R16600 fc2.t14 fc2.n5 0.001
R16601 fc2.n2641 fc2.n2640 0.001
R16602 fc2.n132 fc2.n131 0.001
R16603 fc2.n2002 fc2.n2001 0.001
R16604 fc2.n629 fc2.n628 0.001
R16605 fc2.n1686 fc2.n1685 0.001
R16606 fc2.n1088 fc2.n1087 0.001
R16607 fc2.t14 fc2.n12 0.001
R16608 fc2.n1157 fc2.n1133 0.001
R16609 fc2.n1731 fc2.n1704 0.001
R16610 fc2.n674 fc2.n647 0.001
R16611 fc2.n2046 fc2.n2020 0.001
R16612 fc2.n2740 fc2.n2725 0.001
R16613 fc2.n2718 fc2.n2711 0.001
R16614 fc2.n2673 fc2.n2659 0.001
R16615 fc2.n1584 fc2.n1548 0.001
R16616 fc2.n604 fc2.n568 0.001
R16617 fc2.n2229 fc2.n2192 0.001
R16618 fc2.n3336 fc2.n3335 0.001
R16619 fc2.n1063 fc2.n1021 0.001
R16620 fc2.n1251 fc2.n1212 0.001
R16621 fc2.n1329 fc2.n1290 0.001
R16622 fc2.n1660 fc2.n1624 0.001
R16623 fc2.n1407 fc2.n1368 0.001
R16624 fc2.n1870 fc2.n1833 0.001
R16625 fc2.n847 fc2.n810 0.001
R16626 fc2.n265 fc2.n238 0.001
R16627 fc2.n378 fc2.n341 0.001
R16628 fc2.n2183 fc2.n2182 0.001
R16629 fc2.n412 fc2.n385 0.001
R16630 fc2.n2134 fc2.n2108 0.001
R16631 fc2.n2385 fc2.n2348 0.001
R16632 fc2.n759 fc2.n736 0.001
R16633 fc2.n2464 fc2.n2463 0.001
R16634 fc2.n160 fc2.n159 0.001
R16635 fc2.n522 fc2.n521 0.001
R16636 fc2.n2062 fc2.n2061 0.001
R16637 fc2.n2256 fc2.n2255 0.001
R16638 fc2.n690 fc2.n689 0.001
R16639 fc2.n871 fc2.n870 0.001
R16640 fc2.n1747 fc2.n1746 0.001
R16641 fc2.n1894 fc2.n1893 0.001
R16642 fc2.n1120 fc2.n1119 0.001
R16643 fc2.n1431 fc2.n1430 0.001
R16644 fc2.n2731 fc2.n2730 0.001
R16645 fc2.n2714 fc2.n2713 0.001
R16646 fc2.n2553 fc2.n2552 0.001
R16647 fc2.n248 fc2.n247 0.001
R16648 fc2.n358 fc2.n357 0.001
R16649 fc2.n2166 fc2.n2165 0.001
R16650 fc2.n1766 fc2.n1765 0.001
R16651 fc2.n938 fc2.n937 0.001
R16652 fc2.n713 fc2.n712 0.001
R16653 fc2.n2321 fc2.n2320 0.001
R16654 fc2.n2085 fc2.n2084 0.001
R16655 fc2.n434 fc2.n433 0.001
R16656 fc2.n184 fc2.n183 0.001
R16657 fc2.n2486 fc2.n2485 0.001
R16658 fc2.n2665 fc2.n2664 0.001
R16659 fc2.n2757 fc2.n2756 0.001
R16660 fc2.n2773 fc2.n2772 0.001
R16661 fc2.n276 fc2.n275 0.001
R16662 fc2.n325 fc2.n324 0.001
R16663 fc2.n2145 fc2.n2144 0.001
R16664 fc2.n2400 fc2.n2399 0.001
R16665 fc2.n770 fc2.n769 0.001
R16666 fc2.n973 fc2.n972 0.001
R16667 fc2.n1793 fc2.n1792 0.001
R16668 fc2.n1953 fc2.n1952 0.001
R16669 fc2.n1168 fc2.n1167 0.001
R16670 fc2.n2690 fc2.n2689 0.001
R16671 fc2.n2535 fc2.n2534 0.001
R16672 fc2.n214 fc2.n213 0.001
R16673 fc2.n392 fc2.n391 0.001
R16674 fc2.n2118 fc2.n2117 0.001
R16675 fc2.n2365 fc2.n2364 0.001
R16676 fc2.n743 fc2.n742 0.001
R16677 fc2.n1473 fc2.n1472 0.001
R16678 fc2.n1920 fc2.n1919 0.001
R16679 fc2.n1140 fc2.n1139 0.001
R16680 fc2.n1040 fc2.n1039 0.001
R16681 fc2.n897 fc2.n896 0.001
R16682 fc2.n1715 fc2.n1714 0.001
R16683 fc2.n1564 fc2.n1563 0.001
R16684 fc2.n1194 fc2.n1193 0.001
R16685 fc2.n1228 fc2.n1227 0.001
R16686 fc2.n2282 fc2.n2281 0.001
R16687 fc2.n658 fc2.n657 0.001
R16688 fc2.n584 fc2.n583 0.001
R16689 fc2.n1607 fc2.n1606 0.001
R16690 fc2.n1640 fc2.n1639 0.001
R16691 fc2.n1272 fc2.n1271 0.001
R16692 fc2.n1306 fc2.n1305 0.001
R16693 fc2.n477 fc2.n476 0.001
R16694 fc2.n2030 fc2.n2029 0.001
R16695 fc2.n2209 fc2.n2208 0.001
R16696 fc2.n793 fc2.n792 0.001
R16697 fc2.n827 fc2.n826 0.001
R16698 fc2.n1816 fc2.n1815 0.001
R16699 fc2.n1850 fc2.n1849 0.001
R16700 fc2.n1350 fc2.n1349 0.001
R16701 fc2.n1384 fc2.n1383 0.001
R16702 fc2.n79 fc2.n78 0.001
R16703 fc2.n2800 fc2.n2799 0.001
R16704 fc2.n553 fc2.n552 0.001
R16705 fc2.n2438 fc2.n2437 0.001
R16706 fc2.n1011 fc2.n1010 0.001
R16707 fc2.n1540 fc2.n1539 0.001
R16708 fc2.n1522 fc2.n1521 0.001
R16709 fc2.n2990 fc2.n2985 0.001
R16710 fc2.n2991 fc2.n2976 0.001
R16711 fc2.n3569 fc2.n3568 0.001
R16712 fc2.n3558 fc2.n3557 0.001
R16713 fc2.n3548 fc2.n3547 0.001
R16714 fc2.n3538 fc2.n3537 0.001
R16715 fc2.n3528 fc2.n3527 0.001
R16716 fc2.n3518 fc2.n3517 0.001
R16717 fc2.n3508 fc2.n3507 0.001
R16718 fc2.n3498 fc2.n3497 0.001
R16719 fc2.n3488 fc2.n3487 0.001
R16720 fc2.n3478 fc2.n3477 0.001
R16721 fc2.n3669 fc2.n3668 0.001
R16722 fc2.n3658 fc2.n3657 0.001
R16723 fc2.n3648 fc2.n3647 0.001
R16724 fc2.n3638 fc2.n3637 0.001
R16725 fc2.n3628 fc2.n3627 0.001
R16726 fc2.n3618 fc2.n3617 0.001
R16727 fc2.n3720 fc2.n3708 0.001
R16728 fc2.n3721 fc2.n3696 0.001
R16729 fc2.n3335 fc2.n3332 0.001
R16730 fc2.n3335 fc2.n3334 0.001
R16731 fc2.n3335 fc2.n3331 0.001
R16732 fc2.n3335 fc2.n3333 0.001
R16733 fc2.n3335 fc2.n3330 0.001
R16734 fc2.n1517 fc2.n1516 0.001
R16735 fc2.n1091 fc2.n1090 0.001
R16736 fc2.n1689 fc2.n1688 0.001
R16737 fc2.n632 fc2.n631 0.001
R16738 fc2.n2005 fc2.n2004 0.001
R16739 fc2.n135 fc2.n134 0.001
R16740 fc2.n2644 fc2.n2643 0.001
R16741 fc2.n3304 fc2.n3177 0.001
R16742 fc2.n3299 fc2.n3297 0.001
R16743 fc2.n3289 fc2.n3287 0.001
R16744 fc2.n3279 fc2.n3277 0.001
R16745 fc2.n3269 fc2.n3267 0.001
R16746 fc2.n3259 fc2.n3257 0.001
R16747 fc2.n3249 fc2.n3247 0.001
R16748 fc2.n3239 fc2.n3237 0.001
R16749 fc2.n3229 fc2.n3227 0.001
R16750 fc2.n3219 fc2.n3217 0.001
R16751 fc2.n3209 fc2.n3207 0.001
R16752 fc2.n3199 fc2.n3196 0.001
R16753 fc2.n3188 fc2.n3187 0.001
R16754 fc2.n3089 fc2.n3088 0.001
R16755 fc2.n3099 fc2.n3098 0.001
R16756 fc2.n3119 fc2.n3118 0.001
R16757 fc2.n3139 fc2.n3138 0.001
R16758 fc2.n3159 fc2.n3158 0.001
R16759 fc2.n3172 fc2.n3076 0.001
R16760 fc2.n3069 fc2.n3067 0.001
R16761 fc2.n3169 fc2.n3167 0.001
R16762 fc2.n3149 fc2.n3147 0.001
R16763 fc2.n3129 fc2.n3127 0.001
R16764 fc2.n3109 fc2.n3107 0.001
R16765 fc2.n3018 fc2.n3017 0.001
R16766 fc2.n3028 fc2.n3027 0.001
R16767 fc2.n3048 fc2.n3047 0.001
R16768 fc2.n3061 fc2.n3005 0.001
R16769 fc2.n2998 fc2.n2996 0.001
R16770 fc2.n3058 fc2.n3056 0.001
R16771 fc2.n3038 fc2.n3036 0.001
R16772 fc2.n2985 fc2.n2983 0.001
R16773 fc2.n2976 fc2.n2974 0.001
R16774 fc2.n2967 fc2.n2964 0.001
R16775 fc2.n2955 fc2.n2954 0.001
R16776 fc2.n2924 fc2.n2923 0.001
R16777 fc2.n2934 fc2.n2933 0.001
R16778 fc2.n2947 fc2.n2911 0.001
R16779 fc2.n2904 fc2.n2902 0.001
R16780 fc2.n2944 fc2.n2942 0.001
R16781 fc2.n2833 fc2.n2832 0.001
R16782 fc2.n2843 fc2.n2842 0.001
R16783 fc2.n2863 fc2.n2862 0.001
R16784 fc2.n2883 fc2.n2882 0.001
R16785 fc2.n2896 fc2.n2820 0.001
R16786 fc2.n2813 fc2.n2811 0.001
R16787 fc2.n2893 fc2.n2891 0.001
R16788 fc2.n2873 fc2.n2871 0.001
R16789 fc2.n2853 fc2.n2851 0.001
R16790 fc2.n3696 fc2.n3693 0.001
R16791 fc2.n3464 fc2.n3461 0.001
R16792 fc2.n3568 fc2.n3566 0.001
R16793 fc2.n3557 fc2.n3555 0.001
R16794 fc2.n3547 fc2.n3545 0.001
R16795 fc2.n3537 fc2.n3535 0.001
R16796 fc2.n3527 fc2.n3525 0.001
R16797 fc2.n3517 fc2.n3515 0.001
R16798 fc2.n3507 fc2.n3505 0.001
R16799 fc2.n3497 fc2.n3495 0.001
R16800 fc2.n3487 fc2.n3485 0.001
R16801 fc2.n3477 fc2.n3474 0.001
R16802 fc2.n3873 fc2.n3871 0.001
R16803 fc2.n3958 fc2.n3956 0.001
R16804 fc2.n3948 fc2.n3946 0.001
R16805 fc2.n3938 fc2.n3936 0.001
R16806 fc2.n3928 fc2.n3926 0.001
R16807 fc2.n3918 fc2.n3916 0.001
R16808 fc2.n3908 fc2.n3906 0.001
R16809 fc2.n3898 fc2.n3896 0.001
R16810 fc2.n3888 fc2.n3883 0.001
R16811 fc2.n3604 fc2.n3601 0.001
R16812 fc2.n3668 fc2.n3666 0.001
R16813 fc2.n3657 fc2.n3655 0.001
R16814 fc2.n3647 fc2.n3645 0.001
R16815 fc2.n3637 fc2.n3635 0.001
R16816 fc2.n3627 fc2.n3625 0.001
R16817 fc2.n3617 fc2.n3614 0.001
R16818 fc2.n3790 fc2.n3788 0.001
R16819 fc2.n3835 fc2.n3833 0.001
R16820 fc2.n3825 fc2.n3823 0.001
R16821 fc2.n3815 fc2.n3813 0.001
R16822 fc2.n3805 fc2.n3800 0.001
R16823 fc2.n3708 fc2.n3706 0.001
R16824 fc2.n3719 fc2.n3712 0.001
R16825 fc2.n3755 fc2.n3749 0.001
R16826 fc2.n3299 fc2.n3294 0.001
R16827 fc2.n3289 fc2.n3284 0.001
R16828 fc2.n3279 fc2.n3274 0.001
R16829 fc2.n3269 fc2.n3264 0.001
R16830 fc2.n3259 fc2.n3254 0.001
R16831 fc2.n3249 fc2.n3244 0.001
R16832 fc2.n3239 fc2.n3234 0.001
R16833 fc2.n3229 fc2.n3224 0.001
R16834 fc2.n3219 fc2.n3214 0.001
R16835 fc2.n3209 fc2.n3204 0.001
R16836 fc2.n3199 fc2.n3193 0.001
R16837 fc2.n3188 fc2.n3184 0.001
R16838 fc2.n3089 fc2.n3085 0.001
R16839 fc2.n3099 fc2.n3095 0.001
R16840 fc2.n3119 fc2.n3115 0.001
R16841 fc2.n3139 fc2.n3135 0.001
R16842 fc2.n3159 fc2.n3155 0.001
R16843 fc2.n3172 fc2.n3073 0.001
R16844 fc2.n3169 fc2.n3164 0.001
R16845 fc2.n3149 fc2.n3144 0.001
R16846 fc2.n3129 fc2.n3124 0.001
R16847 fc2.n3109 fc2.n3104 0.001
R16848 fc2.n3018 fc2.n3014 0.001
R16849 fc2.n3028 fc2.n3024 0.001
R16850 fc2.n3048 fc2.n3044 0.001
R16851 fc2.n3061 fc2.n3002 0.001
R16852 fc2.n3058 fc2.n3053 0.001
R16853 fc2.n3038 fc2.n3033 0.001
R16854 fc2.n2985 fc2.n2980 0.001
R16855 fc2.n2976 fc2.n2971 0.001
R16856 fc2.n2924 fc2.n2920 0.001
R16857 fc2.n2934 fc2.n2930 0.001
R16858 fc2.n2947 fc2.n2908 0.001
R16859 fc2.n2944 fc2.n2939 0.001
R16860 fc2.n2833 fc2.n2829 0.001
R16861 fc2.n2843 fc2.n2839 0.001
R16862 fc2.n2863 fc2.n2859 0.001
R16863 fc2.n2883 fc2.n2879 0.001
R16864 fc2.n2896 fc2.n2817 0.001
R16865 fc2.n2893 fc2.n2888 0.001
R16866 fc2.n2873 fc2.n2868 0.001
R16867 fc2.n2853 fc2.n2848 0.001
R16868 fc2.n3696 fc2.n3690 0.001
R16869 fc2.n3568 fc2.n3563 0.001
R16870 fc2.n3557 fc2.n3552 0.001
R16871 fc2.n3547 fc2.n3542 0.001
R16872 fc2.n3537 fc2.n3532 0.001
R16873 fc2.n3527 fc2.n3522 0.001
R16874 fc2.n3517 fc2.n3512 0.001
R16875 fc2.n3507 fc2.n3502 0.001
R16876 fc2.n3497 fc2.n3492 0.001
R16877 fc2.n3487 fc2.n3482 0.001
R16878 fc2.n3477 fc2.n3471 0.001
R16879 fc2.n3958 fc2.n3953 0.001
R16880 fc2.n3948 fc2.n3943 0.001
R16881 fc2.n3938 fc2.n3933 0.001
R16882 fc2.n3928 fc2.n3923 0.001
R16883 fc2.n3918 fc2.n3913 0.001
R16884 fc2.n3908 fc2.n3903 0.001
R16885 fc2.n3898 fc2.n3893 0.001
R16886 fc2.n3888 fc2.n3880 0.001
R16887 fc2.n3668 fc2.n3663 0.001
R16888 fc2.n3657 fc2.n3652 0.001
R16889 fc2.n3647 fc2.n3642 0.001
R16890 fc2.n3637 fc2.n3632 0.001
R16891 fc2.n3627 fc2.n3622 0.001
R16892 fc2.n3617 fc2.n3611 0.001
R16893 fc2.n3835 fc2.n3830 0.001
R16894 fc2.n3825 fc2.n3820 0.001
R16895 fc2.n3815 fc2.n3810 0.001
R16896 fc2.n3805 fc2.n3797 0.001
R16897 fc2.n3708 fc2.n3703 0.001
R16898 fc2.n3777 fc2.n3767 0.001
R16899 fc2.n3581 fc2.n3572 0.001
R16900 fc2.n3982 fc2.n3971 0.001
R16901 fc2.n3681 fc2.n3672 0.001
R16902 fc2.n3859 fc2.n3848 0.001
R16903 fc2.n3741 fc2.n3732 0.001
R16904 fc2.n3081 fc2.n3079 0.001
R16905 fc2.n3010 fc2.n3008 0.001
R16906 fc2.n2959 fc2.n2957 0.001
R16907 fc2.n2916 fc2.n2914 0.001
R16908 fc2.n2825 fc2.n2823 0.001
R16909 fc2.n3180 fc2.n3179 0.001
R16910 fc2.n2989 fc2.n2987 0.001
R16911 fc2.n298 fc2.n290 0.001
R16912 fc2.n302 fc2.n298 0.001
R16913 fc2.n290 fc2.t66 0.001
R16914 fc2.n2613 fc2.n2612 0.001
R16915 fc2.t38 fc2.n2617 0.001
R16916 fc2.t38 fc2.n2475 0.001
R16917 fc2.t38 fc2.n2478 0.001
R16918 fc2.t66 fc2.n172 0.001
R16919 fc2.t66 fc2.n169 0.001
R16920 fc2.n169 fc2.n166 0.001
R16921 fc2.t62 fc2.n536 0.001
R16922 fc2.t62 fc2.n539 0.001
R16923 fc2.t98 fc2.n2073 0.001
R16924 fc2.t98 fc2.n2070 0.001
R16925 fc2.n2070 fc2.n2067 0.001
R16926 fc2.t23 fc2.n2264 0.001
R16927 fc2.t23 fc2.n2238 0.001
R16928 fc2.t52 fc2.n701 0.001
R16929 fc2.t52 fc2.n698 0.001
R16930 fc2.n698 fc2.n695 0.001
R16931 fc2.t47 fc2.n882 0.001
R16932 fc2.t47 fc2.n879 0.001
R16933 fc2.n879 fc2.n876 0.001
R16934 fc2.t12 fc2.n1758 0.001
R16935 fc2.t12 fc2.n1755 0.001
R16936 fc2.n1755 fc2.n1752 0.001
R16937 fc2.t28 fc2.n1905 0.001
R16938 fc2.t28 fc2.n1902 0.001
R16939 fc2.n1902 fc2.n1899 0.001
R16940 fc2.t10 fc2.n1131 0.001
R16941 fc2.t10 fc2.n1128 0.001
R16942 fc2.n1128 fc2.n1125 0.001
R16943 fc2.t94 fc2.n1444 0.001
R16944 fc2.t94 fc2.n1441 0.001
R16945 fc2.n1441 fc2.n1438 0.001
R16946 fc2.n2992 fc2.n2967 0.001
R16947 fc2.n2960 fc2.n2955 0.001
R16948 fc2.t4 fc2.n2743 0.001
R16949 fc2.t4 fc2.n2746 0.001
R16950 fc2.n2786 fc2.t38 0.001
R16951 fc2.n2806 fc2.n2788 0.001
R16952 fc2.t4 fc2.n2721 0.001
R16953 fc2.t4 fc2.n2724 0.001
R16954 fc2.t38 fc2.n2578 0.001
R16955 fc2.t38 fc2.n2581 0.001
R16956 fc2.t66 fc2.n268 0.001
R16957 fc2.t66 fc2.n271 0.001
R16958 fc2.t62 fc2.n384 0.001
R16959 fc2.t62 fc2.n381 0.001
R16960 fc2.n381 fc2.n378 0.001
R16961 fc2.n2160 fc2.t98 0.001
R16962 fc2.n2182 fc2.n2160 0.001
R16963 fc2.n2424 fc2.t23 0.001
R16964 fc2.n2444 fc2.n2426 0.001
R16965 fc2.n1974 fc2.t28 0.001
R16966 fc2.n1986 fc2.n1974 0.001
R16967 fc2.t12 fc2.n1785 0.001
R16968 fc2.t12 fc2.n1788 0.001
R16969 fc2.t47 fc2.n961 0.001
R16970 fc2.t47 fc2.n964 0.001
R16971 fc2.t52 fc2.n732 0.001
R16972 fc2.t52 fc2.n735 0.001
R16973 fc2.t23 fc2.n2344 0.001
R16974 fc2.t23 fc2.n2347 0.001
R16975 fc2.t98 fc2.n2104 0.001
R16976 fc2.t98 fc2.n2107 0.001
R16977 fc2.t62 fc2.n460 0.001
R16978 fc2.t62 fc2.n457 0.001
R16979 fc2.n457 fc2.n454 0.001
R16980 fc2.t66 fc2.n204 0.001
R16981 fc2.t66 fc2.n207 0.001
R16982 fc2.t38 fc2.n2510 0.001
R16983 fc2.t38 fc2.n2513 0.001
R16984 fc2.t4 fc2.n2676 0.001
R16985 fc2.t4 fc2.n2679 0.001
R16986 fc2.n2751 fc2.t4 0.001
R16987 fc2.n2766 fc2.n2751 0.001
R16988 fc2.t38 fc2.n2780 0.001
R16989 fc2.t38 fc2.n2783 0.001
R16990 fc2.t66 fc2.n284 0.001
R16991 fc2.t66 fc2.n287 0.001
R16992 fc2.t62 fc2.n338 0.001
R16993 fc2.n335 fc2.n328 0.001
R16994 fc2.t98 fc2.n2154 0.001
R16995 fc2.t98 fc2.n2157 0.001
R16996 fc2.t23 fc2.n2418 0.001
R16997 fc2.t23 fc2.n2421 0.001
R16998 fc2.t52 fc2.n781 0.001
R16999 fc2.t52 fc2.n784 0.001
R17000 fc2.t47 fc2.n991 0.001
R17001 fc2.t47 fc2.n994 0.001
R17002 fc2.t12 fc2.n1804 0.001
R17003 fc2.t12 fc2.n1807 0.001
R17004 fc2.t28 fc2.n1969 0.001
R17005 fc2.t28 fc2.n1972 0.001
R17006 fc2.t10 fc2.n1182 0.001
R17007 fc2.t10 fc2.n1185 0.001
R17008 fc2.n1502 fc2.t94 0.001
R17009 fc2.n1530 fc2.n1502 0.001
R17010 fc2.t4 fc2.n2697 0.001
R17011 fc2.t4 fc2.n2700 0.001
R17012 fc2.t38 fc2.n2543 0.001
R17013 fc2.t38 fc2.n2546 0.001
R17014 fc2.t66 fc2.n234 0.001
R17015 fc2.t66 fc2.n237 0.001
R17016 fc2.t62 fc2.n418 0.001
R17017 fc2.t62 fc2.n415 0.001
R17018 fc2.n415 fc2.n412 0.001
R17019 fc2.t98 fc2.n2137 0.001
R17020 fc2.t98 fc2.n2140 0.001
R17021 fc2.t23 fc2.n2388 0.001
R17022 fc2.t23 fc2.n2391 0.001
R17023 fc2.t52 fc2.n762 0.001
R17024 fc2.t52 fc2.n765 0.001
R17025 fc2.n997 fc2.t47 0.001
R17026 fc2.n1017 fc2.n999 0.001
R17027 fc2.t94 fc2.n1497 0.001
R17028 fc2.t94 fc2.n1500 0.001
R17029 fc2.t28 fc2.n1941 0.001
R17030 fc2.t28 fc2.n1944 0.001
R17031 fc2.t10 fc2.n1160 0.001
R17032 fc2.t10 fc2.n1163 0.001
R17033 fc2.t94 fc2.n1069 0.001
R17034 fc2.t94 fc2.n1066 0.001
R17035 fc2.n1066 fc2.n1063 0.001
R17036 fc2.t47 fc2.n919 0.001
R17037 fc2.t47 fc2.n922 0.001
R17038 fc2.t12 fc2.n1737 0.001
R17039 fc2.t12 fc2.n1734 0.001
R17040 fc2.n1734 fc2.n1731 0.001
R17041 fc2.t28 fc2.n1590 0.001
R17042 fc2.t28 fc2.n1587 0.001
R17043 fc2.n1587 fc2.n1584 0.001
R17044 fc2.n1188 fc2.t10 0.001
R17045 fc2.n1211 fc2.n1188 0.001
R17046 fc2.t94 fc2.n1257 0.001
R17047 fc2.t94 fc2.n1254 0.001
R17048 fc2.n1254 fc2.n1251 0.001
R17049 fc2.t23 fc2.n2305 0.001
R17050 fc2.n2302 fc2.n2279 0.001
R17051 fc2.t52 fc2.n680 0.001
R17052 fc2.t52 fc2.n677 0.001
R17053 fc2.n677 fc2.n674 0.001
R17054 fc2.t47 fc2.n610 0.001
R17055 fc2.t47 fc2.n607 0.001
R17056 fc2.n607 fc2.n604 0.001
R17057 fc2.n1623 fc2.n1601 0.001
R17058 fc2.t28 fc2.n1666 0.001
R17059 fc2.t28 fc2.n1663 0.001
R17060 fc2.n1663 fc2.n1660 0.001
R17061 fc2.n1289 fc2.n1266 0.001
R17062 fc2.t94 fc2.n1335 0.001
R17063 fc2.t94 fc2.n1332 0.001
R17064 fc2.n1332 fc2.n1329 0.001
R17065 fc2.t62 fc2.n503 0.001
R17066 fc2.t62 fc2.n500 0.001
R17067 fc2.n500 fc2.n497 0.001
R17068 fc2.t98 fc2.n2052 0.001
R17069 fc2.t98 fc2.n2049 0.001
R17070 fc2.n2049 fc2.n2046 0.001
R17071 fc2.t23 fc2.n2235 0.001
R17072 fc2.t23 fc2.n2232 0.001
R17073 fc2.n2232 fc2.n2229 0.001
R17074 fc2.n787 fc2.t52 0.001
R17075 fc2.n809 fc2.n787 0.001
R17076 fc2.t47 fc2.n853 0.001
R17077 fc2.t47 fc2.n850 0.001
R17078 fc2.n850 fc2.n847 0.001
R17079 fc2.n1810 fc2.t12 0.001
R17080 fc2.n1832 fc2.n1810 0.001
R17081 fc2.t28 fc2.n1876 0.001
R17082 fc2.t28 fc2.n1873 0.001
R17083 fc2.n1873 fc2.n1870 0.001
R17084 fc2.n1367 fc2.n1344 0.001
R17085 fc2.t94 fc2.n1413 0.001
R17086 fc2.t94 fc2.n1410 0.001
R17087 fc2.n1410 fc2.n1407 0.001
R17088 fc2.n2264 fc2.n2261 0.001
R17089 fc2.n536 fc2.n533 0.001
R17090 fc2.n2475 fc2.n2472 0.001
R17091 fc2.n809 fc2.n790 0.001
R17092 fc2.n1832 fc2.n1813 0.001
R17093 fc2.n1367 fc2.n1347 0.001
R17094 fc2.n2305 fc2.n2302 0.001
R17095 fc2.n1623 fc2.n1604 0.001
R17096 fc2.n1289 fc2.n1269 0.001
R17097 fc2.n919 fc2.n916 0.001
R17098 fc2.n1211 fc2.n1191 0.001
R17099 fc2.n1941 fc2.n1938 0.001
R17100 fc2.n1160 fc2.n1157 0.001
R17101 fc2.n1497 fc2.n1494 0.001
R17102 fc2.n1182 fc2.n1179 0.001
R17103 fc2.n2766 fc2.n2754 0.001
R17104 fc2.n961 fc2.n958 0.001
R17105 fc2.n732 fc2.n729 0.001
R17106 fc2.n2344 fc2.n2341 0.001
R17107 fc2.n2104 fc2.n2101 0.001
R17108 fc2.n204 fc2.n201 0.001
R17109 fc2.n2510 fc2.n2507 0.001
R17110 fc2.n2676 fc2.n2673 0.001
R17111 fc2.n1785 fc2.n1782 0.001
R17112 fc2.n1986 fc2.n1977 0.001
R17113 fc2.n1017 fc2.n997 0.001
R17114 fc2.n2388 fc2.n2385 0.001
R17115 fc2.n2137 fc2.n2134 0.001
R17116 fc2.n234 fc2.n231 0.001
R17117 fc2.n2543 fc2.n2540 0.001
R17118 fc2.n2697 fc2.n2694 0.001
R17119 fc2.n762 fc2.n759 0.001
R17120 fc2.n2444 fc2.n2424 0.001
R17121 fc2.n268 fc2.n265 0.001
R17122 fc2.n2578 fc2.n2575 0.001
R17123 fc2.n2721 fc2.n2718 0.001
R17124 fc2.n2182 fc2.n2163 0.001
R17125 fc2.n2806 fc2.n2786 0.001
R17126 fc2.n2743 fc2.n2740 0.001
R17127 fc2.n284 fc2.n281 0.001
R17128 fc2.n338 fc2.n335 0.001
R17129 fc2.n2154 fc2.n2151 0.001
R17130 fc2.n2418 fc2.n2415 0.001
R17131 fc2.n781 fc2.n778 0.001
R17132 fc2.n991 fc2.n988 0.001
R17133 fc2.n1804 fc2.n1801 0.001
R17134 fc2.n1969 fc2.n1966 0.001
R17135 fc2.n2780 fc2.n2777 0.001
R17136 fc2.n1530 fc2.n1505 0.001
R17137 fc2.n2802 fc2.n2801 0.001
R17138 fc2.n555 fc2.n554 0.001
R17139 fc2.n2440 fc2.n2439 0.001
R17140 fc2.n1013 fc2.n1012 0.001
R17141 fc2.n1542 fc2.n1541 0.001
R17142 fc2.n1524 fc2.n1523 0.001
R17143 fc2.n82 fc2.n81 0.001
R17144 fc2.n2803 fc2.n2802 0.001
R17145 fc2.n556 fc2.n555 0.001
R17146 fc2.n2441 fc2.n2440 0.001
R17147 fc2.n1014 fc2.n1013 0.001
R17148 fc2.n1543 fc2.n1542 0.001
R17149 fc2.n1015 fc2.n1004 0.001
R17150 fc2.n2442 fc2.n2431 0.001
R17151 fc2.n557 fc2.n546 0.001
R17152 fc2.n2804 fc2.n2793 0.001
R17153 fc2.n1525 fc2.n1524 0.001
R17154 fc2.n106 fc2.n85 0.001
R17155 fc2.n314 fc2.n302 0.001
R17156 fc2.n2612 fc2.n2608 0.001
R17157 VN.n1714 VN.n1712 169.353
R17158 VN.n1137 VN.n1136 169.353
R17159 VN.n833 VN.n832 169.353
R17160 VN.n523 VN.n522 169.353
R17161 VN.n1735 VN.n1734 169.353
R17162 VN.n499 VN.n498 169.353
R17163 VN.n1714 VN.n1713 169.353
R17164 VN.n497 VN.n496 137.98
R17165 VN.n1733 VN.n1732 137.98
R17166 VN.n521 VN.n520 137.98
R17167 VN.n831 VN.n830 137.98
R17168 VN.n1135 VN.n1134 137.98
R17169 VN.n1711 VN.n1710 137.98
R17170 VN.n1203 VN.n1202 135.611
R17171 VN.n977 VN.n976 135.611
R17172 VN.n654 VN.n653 135.611
R17173 VN.n1862 VN.n1861 135.611
R17174 VN.n153 VN.n152 135.611
R17175 VN.n307 VN.n306 135.611
R17176 VN.n1716 VN.t24 118.651
R17177 VN.n1205 VN.t15 118.651
R17178 VN.n1139 VN.t30 118.651
R17179 VN.n979 VN.t47 118.651
R17180 VN.n835 VN.t91 118.651
R17181 VN.n656 VN.t74 118.651
R17182 VN.n525 VN.t33 118.651
R17183 VN.n1864 VN.t45 118.651
R17184 VN.n1737 VN.t9 118.651
R17185 VN.n155 VN.t81 118.651
R17186 VN.n501 VN.t93 118.651
R17187 VN.n309 VN.t26 118.651
R17188 VN.t5 VN.n1669 114.696
R17189 VN.t50 VN.n1293 114.696
R17190 VN.t11 VN.n1389 114.696
R17191 VN.t22 VN.n1069 114.696
R17192 VN.t37 VN.n930 114.696
R17193 VN.t13 VN.n727 114.696
R17194 VN.t17 VN.n587 114.696
R17195 VN.t2 VN.n1912 114.696
R17196 VN.t39 VN.n1776 114.696
R17197 VN.t20 VN.n209 114.696
R17198 VN.t42 VN.n469 114.696
R17199 VN.t7 VN.n274 114.696
R17200 VN.t52 VN.n11 114.696
R17201 VN.n1214 VN.n1213 91.65
R17202 VN.n298 VN.n297 91.65
R17203 VN.n666 VN.n665 91.65
R17204 VN.n1873 VN.n1872 91.65
R17205 VN.n165 VN.n164 91.65
R17206 VN.n989 VN.n988 91.65
R17207 VN.n491 VN.n490 91.389
R17208 VN.n2007 VN.n2006 91.389
R17209 VN.n1701 VN.n1700 91.389
R17210 VN.n1431 VN.n1430 91.389
R17211 VN.n1126 VN.n1125 91.389
R17212 VN.n802 VN.n801 91.389
R17213 VN.n1556 VN.n1555 87.222
R17214 VN.n1600 VN.n1599 87.222
R17215 VN.n1568 VN.n1567 87.222
R17216 VN.n1581 VN.n1580 87.222
R17217 VN.n1590 VN.n1589 87.222
R17218 VN.n1603 VN.n1602 87.222
R17219 VN.n101 VN.n100 86.961
R17220 VN.n56 VN.n55 86.961
R17221 VN.n66 VN.n65 86.961
R17222 VN.n74 VN.n73 86.961
R17223 VN.n82 VN.n81 86.961
R17224 VN.n44 VN.n43 86.961
R17225 VN.n1669 VN.t0 21.258
R17226 VN.n967 VN.t259 3.904
R17227 VN.n969 VN.n968 3.904
R17228 VN.n10 VN.t62 3.904
R17229 VN.n9 VN.t106 3.904
R17230 VN.n491 VN.t188 3.904
R17231 VN.n439 VN.t102 3.904
R17232 VN.n101 VN.t354 3.904
R17233 VN.n99 VN.t297 3.904
R17234 VN.n282 VN.n281 3.904
R17235 VN.n290 VN.t58 3.904
R17236 VN.n293 VN.t97 3.904
R17237 VN.n285 VN.n284 3.904
R17238 VN.n477 VN.n476 3.904
R17239 VN.n485 VN.t290 3.904
R17240 VN.n488 VN.t228 3.904
R17241 VN.n480 VN.n479 3.904
R17242 VN.n189 VN.n188 3.904
R17243 VN.n207 VN.t54 3.904
R17244 VN.n204 VN.t95 3.904
R17245 VN.n192 VN.n191 3.904
R17246 VN.n2007 VN.t310 3.904
R17247 VN.n2009 VN.t224 3.904
R17248 VN.n1215 VN.t353 3.904
R17249 VN.n1680 VN.n1679 3.904
R17250 VN.n1695 VN.t233 3.904
R17251 VN.n1698 VN.t4 3.904
R17252 VN.n1683 VN.n1682 3.904
R17253 VN.n1554 VN.t256 3.904
R17254 VN.n1596 VN.t373 3.904
R17255 VN.n1656 VN.n1655 3.904
R17256 VN.n1667 VN.t121 3.904
R17257 VN.n1664 VN.t171 3.904
R17258 VN.n1659 VN.n1658 3.904
R17259 VN.n1371 VN.n1370 3.904
R17260 VN.n1387 VN.t249 3.904
R17261 VN.n1384 VN.t175 3.904
R17262 VN.n1368 VN.n1367 3.904
R17263 VN.n295 VN.t220 3.904
R17264 VN.n447 VN.n446 3.904
R17265 VN.n467 VN.t43 3.904
R17266 VN.n464 VN.t266 3.904
R17267 VN.n444 VN.n443 3.904
R17268 VN.n174 VN.n173 3.904
R17269 VN.n183 VN.t119 3.904
R17270 VN.n180 VN.t136 3.904
R17271 VN.n171 VN.n170 3.904
R17272 VN.n1757 VN.n1756 3.904
R17273 VN.n1774 VN.t335 3.904
R17274 VN.n1771 VN.t197 3.904
R17275 VN.n1754 VN.n1753 3.904
R17276 VN.n1901 VN.n1900 3.904
R17277 VN.n1910 VN.t3 3.904
R17278 VN.n1907 VN.t34 3.904
R17279 VN.n1898 VN.n1897 3.904
R17280 VN.n568 VN.n567 3.904
R17281 VN.n585 VN.t250 3.904
R17282 VN.n582 VN.t117 3.904
R17283 VN.n565 VN.n564 3.904
R17284 VN.n716 VN.n715 3.904
R17285 VN.n725 VN.t316 3.904
R17286 VN.n722 VN.t348 3.904
R17287 VN.n713 VN.n712 3.904
R17288 VN.n911 VN.n910 3.904
R17289 VN.n928 VN.t181 3.904
R17290 VN.n925 VN.t180 3.904
R17291 VN.n908 VN.n907 3.904
R17292 VN.n1057 VN.n1056 3.904
R17293 VN.n1067 VN.t382 3.904
R17294 VN.n1064 VN.t31 3.904
R17295 VN.n1054 VN.n1053 3.904
R17296 VN.n1280 VN.n1279 3.904
R17297 VN.n1291 VN.t378 3.904
R17298 VN.n1288 VN.t25 3.904
R17299 VN.n1283 VN.n1282 3.904
R17300 VN.n1562 VN.t384 3.904
R17301 VN.n1479 VN.n1478 3.904
R17302 VN.n1504 VN.t341 3.904
R17303 VN.n1501 VN.t186 3.904
R17304 VN.n1482 VN.n1481 3.904
R17305 VN.n1161 VN.n1160 3.904
R17306 VN.n1173 VN.t385 3.904
R17307 VN.n1170 VN.t252 3.904
R17308 VN.n1158 VN.n1157 3.904
R17309 VN.n940 VN.n939 3.904
R17310 VN.n956 VN.t173 3.904
R17311 VN.n959 VN.t318 3.904
R17312 VN.n937 VN.n936 3.904
R17313 VN.n667 VN.t340 3.904
R17314 VN.n998 VN.n997 3.904
R17315 VN.n1008 VN.t161 3.904
R17316 VN.n1005 VN.t185 3.904
R17317 VN.n995 VN.n994 3.904
R17318 VN.n1237 VN.n1236 3.904
R17319 VN.n1255 VN.t84 3.904
R17320 VN.n1252 VN.t104 3.904
R17321 VN.n1240 VN.n1239 3.904
R17322 VN.n1192 VN.n1191 3.904
R17323 VN.n1311 VN.t264 3.904
R17324 VN.n1314 VN.t294 3.904
R17325 VN.n1317 VN.n1316 3.904
R17326 VN.n1608 VN.n1607 3.904
R17327 VN.n1624 VN.t368 3.904
R17328 VN.n1621 VN.t57 3.904
R17329 VN.n1611 VN.n1610 3.904
R17330 VN.n1572 VN.t262 3.904
R17331 VN.n1874 VN.t300 3.904
R17332 VN.n601 VN.n600 3.904
R17333 VN.n609 VN.t138 3.904
R17334 VN.n612 VN.t344 3.904
R17335 VN.n598 VN.n597 3.904
R17336 VN.n681 VN.n680 3.904
R17337 VN.n689 VN.t202 3.904
R17338 VN.n686 VN.t219 3.904
R17339 VN.n678 VN.n677 3.904
R17340 VN.n855 VN.n854 3.904
R17341 VN.n873 VN.t38 3.904
R17342 VN.n870 VN.t210 3.904
R17343 VN.n852 VN.n851 3.904
R17344 VN.n1022 VN.n1021 3.904
R17345 VN.n1030 VN.t23 3.904
R17346 VN.n1027 VN.t56 3.904
R17347 VN.n1019 VN.n1018 3.904
R17348 VN.n1188 VN.n1187 3.904
R17349 VN.n1342 VN.t263 3.904
R17350 VN.n1339 VN.t60 3.904
R17351 VN.n1185 VN.n1184 3.904
R17352 VN.n1587 VN.t137 3.904
R17353 VN.n1262 VN.n1261 3.904
R17354 VN.n1274 VN.t139 3.904
R17355 VN.n1271 VN.t163 3.904
R17356 VN.n1265 VN.n1264 3.904
R17357 VN.n1351 VN.n1350 3.904
R17358 VN.n1363 VN.t372 3.904
R17359 VN.n1360 VN.t304 3.904
R17360 VN.n1354 VN.n1353 3.904
R17361 VN.n1036 VN.n1035 3.904
R17362 VN.n1049 VN.t140 3.904
R17363 VN.n1046 VN.t170 3.904
R17364 VN.n1039 VN.n1038 3.904
R17365 VN.n882 VN.n881 3.904
R17366 VN.n894 VN.t284 3.904
R17367 VN.n891 VN.t308 3.904
R17368 VN.n885 VN.n884 3.904
R17369 VN.n695 VN.n694 3.904
R17370 VN.n708 VN.t69 3.904
R17371 VN.n705 VN.t92 3.904
R17372 VN.n698 VN.n697 3.904
R17373 VN.n539 VN.n538 3.904
R17374 VN.n551 VN.t374 3.904
R17375 VN.n548 VN.t243 3.904
R17376 VN.n542 VN.n541 3.904
R17377 VN.n1880 VN.n1879 3.904
R17378 VN.n1893 VN.t154 3.904
R17379 VN.n1890 VN.t172 3.904
R17380 VN.n1883 VN.n1882 3.904
R17381 VN.n1788 VN.n1787 3.904
R17382 VN.n1797 VN.t96 3.904
R17383 VN.n1800 VN.t305 3.904
R17384 VN.n1791 VN.n1790 3.904
R17385 VN.n166 VN.t261 3.904
R17386 VN.n1634 VN.n1633 3.904
R17387 VN.n1646 VN.t247 3.904
R17388 VN.n1643 VN.t299 3.904
R17389 VN.n1637 VN.n1636 3.904
R17390 VN.n1601 VN.t128 3.904
R17391 VN.n1457 VN.n1456 3.904
R17392 VN.n1468 VN.t107 3.904
R17393 VN.n1465 VN.t285 3.904
R17394 VN.n1460 VN.n1459 3.904
R17395 VN.n1396 VN.n1395 3.904
R17396 VN.n1408 VN.t144 3.904
R17397 VN.n1411 VN.t358 3.904
R17398 VN.n1393 VN.n1392 3.904
R17399 VN.n990 VN.t312 3.904
R17400 VN.n1221 VN.n1220 3.904
R17401 VN.n1232 VN.t215 3.904
R17402 VN.n1229 VN.t231 3.904
R17403 VN.n1224 VN.n1223 3.904
R17404 VN.n1701 VN.t379 3.904
R17405 VN.n1703 VN.t32 3.904
R17406 VN.n1296 VN.n1295 3.904
R17407 VN.n1305 VN.t255 3.904
R17408 VN.n1308 VN.t278 3.904
R17409 VN.n1299 VN.n1298 3.904
R17410 VN.n1416 VN.n1415 3.904
R17411 VN.n1425 VN.t124 3.904
R17412 VN.n1428 VN.t41 3.904
R17413 VN.n1419 VN.n1418 3.904
R17414 VN.n1090 VN.n1089 3.904
R17415 VN.n1103 VN.t49 3.904
R17416 VN.n1106 VN.t48 3.904
R17417 VN.n1093 VN.n1092 3.904
R17418 VN.n731 VN.n730 3.904
R17419 VN.n740 VN.t191 3.904
R17420 VN.n743 VN.t225 3.904
R17421 VN.n734 VN.n733 3.904
R17422 VN.n616 VN.n615 3.904
R17423 VN.n629 VN.t55 3.904
R17424 VN.n632 VN.t355 3.904
R17425 VN.n619 VN.n618 3.904
R17426 VN.n1916 VN.n1915 3.904
R17427 VN.n1925 VN.t193 3.904
R17428 VN.n1928 VN.t229 3.904
R17429 VN.n1919 VN.n1918 3.904
R17430 VN.n1804 VN.n1803 3.904
R17431 VN.n1817 VN.t209 3.904
R17432 VN.n1820 VN.t360 3.904
R17433 VN.n1807 VN.n1806 3.904
R17434 VN.n407 VN.n406 3.904
R17435 VN.n410 VN.t356 3.904
R17436 VN.n413 VN.t371 3.904
R17437 VN.n416 VN.n415 3.904
R17438 VN.n424 VN.n423 3.904
R17439 VN.n437 VN.t287 3.904
R17440 VN.n385 VN.t151 3.904
R17441 VN.n427 VN.n426 3.904
R17442 VN.n389 VN.n388 3.904
R17443 VN.n392 VN.t71 3.904
R17444 VN.n395 VN.t94 3.904
R17445 VN.n398 VN.n397 3.904
R17446 VN.n56 VN.t177 3.904
R17447 VN.n50 VN.t377 3.904
R17448 VN.n1431 VN.t380 3.904
R17449 VN.n1433 VN.t286 3.904
R17450 VN.n1073 VN.n1072 3.904
R17451 VN.n1081 VN.t131 3.904
R17452 VN.n1084 VN.t157 3.904
R17453 VN.n1076 VN.n1075 3.904
R17454 VN.n1114 VN.n1113 3.904
R17455 VN.n1118 VN.t293 3.904
R17456 VN.n1121 VN.t292 3.904
R17457 VN.n1111 VN.n1110 3.904
R17458 VN.n66 VN.t68 3.904
R17459 VN.n61 VN.t254 3.904
R17460 VN.n376 VN.n375 3.904
R17461 VN.n373 VN.t315 3.904
R17462 VN.n370 VN.t332 3.904
R17463 VN.n272 VN.n271 3.904
R17464 VN.n251 VN.n250 3.904
R17465 VN.n248 VN.t159 3.904
R17466 VN.n382 VN.t241 3.904
R17467 VN.n245 VN.n244 3.904
R17468 VN.n265 VN.n264 3.904
R17469 VN.n262 VN.t66 3.904
R17470 VN.n259 VN.t108 3.904
R17471 VN.n256 VN.n255 3.904
R17472 VN.n1828 VN.n1827 3.904
R17473 VN.n1832 VN.t302 3.904
R17474 VN.n1835 VN.t236 3.904
R17475 VN.n1825 VN.n1824 3.904
R17476 VN.n1936 VN.n1935 3.904
R17477 VN.n1941 VN.t65 3.904
R17478 VN.n1944 VN.t103 3.904
R17479 VN.n1933 VN.n1932 3.904
R17480 VN.n640 VN.n639 3.904
R17481 VN.n779 VN.t298 3.904
R17482 VN.n782 VN.t234 3.904
R17483 VN.n637 VN.n636 3.904
R17484 VN.n774 VN.n773 3.904
R17485 VN.n771 VN.t59 3.904
R17486 VN.n768 VN.t98 3.904
R17487 VN.n645 VN.n644 3.904
R17488 VN.n1126 VN.t189 3.904
R17489 VN.n1123 VN.t162 3.904
R17490 VN.n748 VN.n747 3.904
R17491 VN.n762 VN.t303 3.904
R17492 VN.n765 VN.t337 3.904
R17493 VN.n751 VN.n750 3.904
R17494 VN.n790 VN.n789 3.904
R17495 VN.n794 VN.t169 3.904
R17496 VN.n797 VN.t109 3.904
R17497 VN.n787 VN.n786 3.904
R17498 VN.n74 VN.t244 3.904
R17499 VN.n68 VN.t127 3.904
R17500 VN.n323 VN.n322 3.904
R17501 VN.n328 VN.t314 3.904
R17502 VN.n331 VN.t345 3.904
R17503 VN.n320 VN.n319 3.904
R17504 VN.n137 VN.n136 3.904
R17505 VN.n240 VN.t178 3.904
R17506 VN.n129 VN.t114 3.904
R17507 VN.n134 VN.n133 3.904
R17508 VN.n234 VN.n233 3.904
R17509 VN.n231 VN.t311 3.904
R17510 VN.n228 VN.t342 3.904
R17511 VN.n142 VN.n141 3.904
R17512 VN.n1843 VN.n1842 3.904
R17513 VN.n1979 VN.t174 3.904
R17514 VN.n1982 VN.t112 3.904
R17515 VN.n1840 VN.n1839 3.904
R17516 VN.n1974 VN.n1973 3.904
R17517 VN.n1971 VN.t307 3.904
R17518 VN.n1968 VN.t339 3.904
R17519 VN.n1848 VN.n1847 3.904
R17520 VN.n802 VN.t63 3.904
R17521 VN.n799 VN.t343 3.904
R17522 VN.n1947 VN.n1946 3.904
R17523 VN.n1962 VN.t179 3.904
R17524 VN.n1965 VN.t217 3.904
R17525 VN.n1950 VN.n1949 3.904
R17526 VN.n1992 VN.n1991 3.904
R17527 VN.n2001 VN.t40 3.904
R17528 VN.n2004 VN.t347 3.904
R17529 VN.n1995 VN.n1994 3.904
R17530 VN.n82 VN.t116 3.904
R17531 VN.n79 VN.t53 3.904
R17532 VN.n336 VN.n335 3.904
R17533 VN.n344 VN.t190 3.904
R17534 VN.n347 VN.t222 3.904
R17535 VN.n339 VN.n338 3.904
R17536 VN.n115 VN.n114 3.904
R17537 VN.n126 VN.t44 3.904
R17538 VN.n123 VN.t351 3.904
R17539 VN.n118 VN.n117 3.904
R17540 VN.n214 VN.n213 3.904
R17541 VN.n222 VN.t184 3.904
R17542 VN.n225 VN.t221 3.904
R17543 VN.n217 VN.n216 3.904
R17544 VN.n44 VN.t232 3.904
R17545 VN.n42 VN.t167 3.904
R17546 VN.n356 VN.n355 3.904
R17547 VN.n364 VN.t301 3.904
R17548 VN.n367 VN.t336 3.904
R17549 VN.n359 VN.n358 3.904
R17550 VN.n962 VN.t282 3.904
R17551 VN.n1087 VN.n1086 3.904
R17552 VN.n967 VN.n966 3.643
R17553 VN.n969 VN.t230 3.643
R17554 VN.n106 VN.t240 3.643
R17555 VN.n98 VN.t203 3.643
R17556 VN.n282 VN.t8 3.643
R17557 VN.n290 VN.n289 3.643
R17558 VN.n293 VN.n292 3.643
R17559 VN.n285 VN.t327 3.643
R17560 VN.n477 VN.t196 3.643
R17561 VN.n485 VN.n484 3.643
R17562 VN.n488 VN.n487 3.643
R17563 VN.n480 VN.t363 3.643
R17564 VN.n189 VN.t36 3.643
R17565 VN.n207 VN.n206 3.643
R17566 VN.n204 VN.n203 3.643
R17567 VN.n192 VN.t198 3.643
R17568 VN.n2011 VN.t361 3.643
R17569 VN.n1214 VN.t309 3.643
R17570 VN.n1194 VN.t111 3.643
R17571 VN.n1680 VN.t134 3.643
R17572 VN.n1695 VN.n1694 3.643
R17573 VN.n1698 VN.n1697 3.643
R17574 VN.n1683 VN.t239 3.643
R17575 VN.n1556 VN.t388 3.643
R17576 VN.n1553 VN.t226 3.643
R17577 VN.n1600 VN.t143 3.643
R17578 VN.n1595 VN.t364 3.643
R17579 VN.n1656 VN.t386 3.643
R17580 VN.n1667 VN.n1666 3.643
R17581 VN.n1664 VN.n1663 3.643
R17582 VN.n1659 VN.t313 3.643
R17583 VN.n1371 VN.t146 3.643
R17584 VN.n1387 VN.n1386 3.643
R17585 VN.n1384 VN.n1383 3.643
R17586 VN.n1368 VN.t317 3.643
R17587 VN.n298 VN.t168 3.643
R17588 VN.n299 VN.t295 3.643
R17589 VN.n447 VN.t322 3.643
R17590 VN.n467 VN.n466 3.643
R17591 VN.n464 VN.n463 3.643
R17592 VN.n444 VN.t105 3.643
R17593 VN.n174 VN.t90 3.643
R17594 VN.n183 VN.n182 3.643
R17595 VN.n180 VN.n179 3.643
R17596 VN.n171 VN.t257 3.643
R17597 VN.n1757 VN.t238 3.643
R17598 VN.n1774 VN.n1773 3.643
R17599 VN.n1771 VN.n1770 3.643
R17600 VN.n1754 VN.t10 3.643
R17601 VN.n1901 VN.t367 3.643
R17602 VN.n1910 VN.n1909 3.643
R17603 VN.n1907 VN.n1906 3.643
R17604 VN.n1898 VN.t160 3.643
R17605 VN.n568 VN.t87 3.643
R17606 VN.n585 VN.n584 3.643
R17607 VN.n582 VN.n581 3.643
R17608 VN.n565 VN.t258 3.643
R17609 VN.n716 VN.t281 3.643
R17610 VN.n725 VN.n724 3.643
R17611 VN.n722 VN.n721 3.643
R17612 VN.n713 VN.t89 3.643
R17613 VN.n911 VN.t83 3.643
R17614 VN.n928 VN.n927 3.643
R17615 VN.n925 VN.n924 3.643
R17616 VN.n908 VN.t253 3.643
R17617 VN.n1057 VN.t352 3.643
R17618 VN.n1067 VN.n1066 3.643
R17619 VN.n1064 VN.n1063 3.643
R17620 VN.n1054 VN.t150 3.643
R17621 VN.n1280 VN.t349 3.643
R17622 VN.n1291 VN.n1290 3.643
R17623 VN.n1288 VN.n1287 3.643
R17624 VN.n1283 VN.t148 3.643
R17625 VN.n1568 VN.t153 3.643
R17626 VN.n1561 VN.t357 3.643
R17627 VN.n1479 VN.t6 3.643
R17628 VN.n1504 VN.n1503 3.643
R17629 VN.n1501 VN.n1500 3.643
R17630 VN.n1482 VN.t326 3.643
R17631 VN.n1161 VN.t283 3.643
R17632 VN.n1173 VN.n1172 3.643
R17633 VN.n1170 VN.n1169 3.643
R17634 VN.n1158 VN.t88 3.643
R17635 VN.n940 VN.t77 3.643
R17636 VN.n956 VN.n955 3.643
R17637 VN.n959 VN.n958 3.643
R17638 VN.n937 VN.t227 3.643
R17639 VN.n666 VN.t296 3.643
R17640 VN.n647 VN.t99 3.643
R17641 VN.n998 VN.t141 3.643
R17642 VN.n1008 VN.n1007 3.643
R17643 VN.n1005 VN.n1004 3.643
R17644 VN.n995 VN.t306 3.643
R17645 VN.n1237 VN.t51 3.643
R17646 VN.n1255 VN.n1254 3.643
R17647 VN.n1252 VN.n1251 3.643
R17648 VN.n1240 VN.t223 3.643
R17649 VN.n1192 VN.t237 3.643
R17650 VN.n1311 VN.n1310 3.643
R17651 VN.n1314 VN.n1313 3.643
R17652 VN.n1317 VN.t16 3.643
R17653 VN.n1608 VN.t270 3.643
R17654 VN.n1624 VN.n1623 3.643
R17655 VN.n1621 VN.n1620 3.643
R17656 VN.n1611 VN.t200 3.643
R17657 VN.n1581 VN.t1 3.643
R17658 VN.n1571 VN.t235 3.643
R17659 VN.n1873 VN.t260 3.643
R17660 VN.n1850 VN.t46 3.643
R17661 VN.n601 VN.t18 3.643
R17662 VN.n609 VN.n608 3.643
R17663 VN.n612 VN.n611 3.643
R17664 VN.n598 VN.t183 3.643
R17665 VN.n681 VN.t165 3.643
R17666 VN.n689 VN.n688 3.643
R17667 VN.n686 VN.n685 3.643
R17668 VN.n678 VN.t338 3.643
R17669 VN.n855 VN.t319 3.643
R17670 VN.n873 VN.n872 3.643
R17671 VN.n870 VN.n869 3.643
R17672 VN.n852 VN.t120 3.643
R17673 VN.n1022 VN.t383 3.643
R17674 VN.n1030 VN.n1029 3.643
R17675 VN.n1027 VN.n1026 3.643
R17676 VN.n1019 VN.t176 3.643
R17677 VN.n1188 VN.t12 3.643
R17678 VN.n1342 VN.n1341 3.643
R17679 VN.n1339 VN.n1338 3.643
R17680 VN.n1185 VN.t205 3.643
R17681 VN.n1590 VN.t269 3.643
R17682 VN.n1586 VN.t110 3.643
R17683 VN.n1262 VN.t113 3.643
R17684 VN.n1274 VN.n1273 3.643
R17685 VN.n1271 VN.n1270 3.643
R17686 VN.n1265 VN.t272 3.643
R17687 VN.n1351 VN.t271 3.643
R17688 VN.n1363 VN.n1362 3.643
R17689 VN.n1360 VN.n1359 3.643
R17690 VN.n1354 VN.t73 3.643
R17691 VN.n1036 VN.t115 3.643
R17692 VN.n1049 VN.n1048 3.643
R17693 VN.n1046 VN.n1045 3.643
R17694 VN.n1039 VN.t276 3.643
R17695 VN.n882 VN.t213 3.643
R17696 VN.n894 VN.n893 3.643
R17697 VN.n891 VN.n890 3.643
R17698 VN.n885 VN.t376 3.643
R17699 VN.n695 VN.t28 3.643
R17700 VN.n708 VN.n707 3.643
R17701 VN.n705 VN.n704 3.643
R17702 VN.n698 VN.t214 3.643
R17703 VN.n539 VN.t273 3.643
R17704 VN.n551 VN.n550 3.643
R17705 VN.n548 VN.n547 3.643
R17706 VN.n542 VN.t76 3.643
R17707 VN.n1880 VN.t133 3.643
R17708 VN.n1893 VN.n1892 3.643
R17709 VN.n1890 VN.n1889 3.643
R17710 VN.n1883 VN.t291 3.643
R17711 VN.n1788 VN.t362 3.643
R17712 VN.n1797 VN.n1796 3.643
R17713 VN.n1800 VN.n1799 3.643
R17714 VN.n1791 VN.t142 3.643
R17715 VN.n165 VN.t218 3.643
R17716 VN.n144 VN.t381 3.643
R17717 VN.n1634 VN.t145 3.643
R17718 VN.n1646 VN.n1645 3.643
R17719 VN.n1643 VN.n1642 3.643
R17720 VN.n1637 VN.t67 3.643
R17721 VN.n1603 VN.t265 3.643
R17722 VN.n1604 VN.t101 3.643
R17723 VN.n1457 VN.t369 3.643
R17724 VN.n1468 VN.n1467 3.643
R17725 VN.n1465 VN.n1464 3.643
R17726 VN.n1460 VN.t132 3.643
R17727 VN.n1396 VN.t35 3.643
R17728 VN.n1408 VN.n1407 3.643
R17729 VN.n1411 VN.n1410 3.643
R17730 VN.n1393 VN.t195 3.643
R17731 VN.n989 VN.t267 3.643
R17732 VN.n970 VN.t64 3.643
R17733 VN.n1221 VN.t182 3.643
R17734 VN.n1232 VN.n1231 3.643
R17735 VN.n1229 VN.n1228 3.643
R17736 VN.n1224 VN.t346 3.643
R17737 VN.n1547 VN.t350 3.643
R17738 VN.n1525 VN.t147 3.643
R17739 VN.n1705 VN.t187 3.643
R17740 VN.n1296 VN.t245 3.643
R17741 VN.n1305 VN.n1304 3.643
R17742 VN.n1308 VN.n1307 3.643
R17743 VN.n1299 VN.t389 3.643
R17744 VN.n1416 VN.t387 3.643
R17745 VN.n1425 VN.n1424 3.643
R17746 VN.n1428 VN.n1427 3.643
R17747 VN.n1419 VN.t192 3.643
R17748 VN.n1090 VN.t325 3.643
R17749 VN.n1103 VN.n1102 3.643
R17750 VN.n1106 VN.n1105 3.643
R17751 VN.n1093 VN.t126 3.643
R17752 VN.n731 VN.t156 3.643
R17753 VN.n740 VN.n739 3.643
R17754 VN.n743 VN.n742 3.643
R17755 VN.n734 VN.t330 3.643
R17756 VN.n616 VN.t329 3.643
R17757 VN.n629 VN.n628 3.643
R17758 VN.n632 VN.n631 3.643
R17759 VN.n619 VN.t130 3.643
R17760 VN.n1916 VN.t158 3.643
R17761 VN.n1925 VN.n1924 3.643
R17762 VN.n1928 VN.n1927 3.643
R17763 VN.n1919 VN.t334 3.643
R17764 VN.n1804 VN.t333 3.643
R17765 VN.n1817 VN.n1816 3.643
R17766 VN.n1820 VN.n1819 3.643
R17767 VN.n1807 VN.t135 3.643
R17768 VN.n407 VN.t331 3.643
R17769 VN.n410 VN.n409 3.643
R17770 VN.n413 VN.n412 3.643
R17771 VN.n416 VN.t129 3.643
R17772 VN.n424 VN.t194 3.643
R17773 VN.n437 VN.n436 3.643
R17774 VN.n385 VN.n384 3.643
R17775 VN.n427 VN.t359 3.643
R17776 VN.n389 VN.t29 3.643
R17777 VN.n392 VN.n391 3.643
R17778 VN.n395 VN.n394 3.643
R17779 VN.n398 VN.t164 3.643
R17780 VN.n49 VN.t274 3.643
R17781 VN.n1435 VN.t61 3.643
R17782 VN.n1073 VN.t122 3.643
R17783 VN.n1081 VN.n1080 3.643
R17784 VN.n1084 VN.n1083 3.643
R17785 VN.n1076 VN.t268 3.643
R17786 VN.n1114 VN.t199 3.643
R17787 VN.n1118 VN.n1117 3.643
R17788 VN.n1121 VN.n1120 3.643
R17789 VN.n1111 VN.t365 3.643
R17790 VN.n62 VN.t149 3.643
R17791 VN.n376 VN.t280 3.643
R17792 VN.n373 VN.n372 3.643
R17793 VN.n370 VN.n369 3.643
R17794 VN.n272 VN.t27 3.643
R17795 VN.n251 VN.t211 3.643
R17796 VN.n248 VN.n247 3.643
R17797 VN.n382 VN.n381 3.643
R17798 VN.n245 VN.t375 3.643
R17799 VN.n265 VN.t21 3.643
R17800 VN.n262 VN.n261 3.643
R17801 VN.n259 VN.n258 3.643
R17802 VN.n256 VN.t212 3.643
R17803 VN.n1828 VN.t207 3.643
R17804 VN.n1832 VN.n1831 3.643
R17805 VN.n1835 VN.n1834 3.643
R17806 VN.n1825 VN.t370 3.643
R17807 VN.n1936 VN.t19 3.643
R17808 VN.n1941 VN.n1940 3.643
R17809 VN.n1944 VN.n1943 3.643
R17810 VN.n1933 VN.t208 3.643
R17811 VN.n640 VN.t204 3.643
R17812 VN.n779 VN.n778 3.643
R17813 VN.n782 VN.n781 3.643
R17814 VN.n637 VN.t366 3.643
R17815 VN.n774 VN.t14 3.643
R17816 VN.n771 VN.n770 3.643
R17817 VN.n768 VN.n767 3.643
R17818 VN.n645 VN.t206 3.643
R17819 VN.n840 VN.t242 3.643
R17820 VN.n748 VN.t289 3.643
R17821 VN.n762 VN.n761 3.643
R17822 VN.n765 VN.n764 3.643
R17823 VN.n751 VN.t75 3.643
R17824 VN.n790 VN.t72 3.643
R17825 VN.n794 VN.n793 3.643
R17826 VN.n797 VN.n796 3.643
R17827 VN.n787 VN.t246 3.643
R17828 VN.n69 VN.t86 3.643
R17829 VN.n323 VN.t279 3.643
R17830 VN.n328 VN.n327 3.643
R17831 VN.n331 VN.n330 3.643
R17832 VN.n320 VN.t216 3.643
R17833 VN.n137 VN.t80 3.643
R17834 VN.n240 VN.n239 3.643
R17835 VN.n129 VN.n128 3.643
R17836 VN.n134 VN.t251 3.643
R17837 VN.n234 VN.t277 3.643
R17838 VN.n231 VN.n230 3.643
R17839 VN.n228 VN.n227 3.643
R17840 VN.n142 VN.t82 3.643
R17841 VN.n1843 VN.t78 3.643
R17842 VN.n1979 VN.n1978 3.643
R17843 VN.n1982 VN.n1981 3.643
R17844 VN.n1840 VN.t248 3.643
R17845 VN.n1974 VN.t275 3.643
R17846 VN.n1971 VN.n1970 3.643
R17847 VN.n1968 VN.n1967 3.643
R17848 VN.n1848 VN.t79 3.643
R17849 VN.n530 VN.t118 3.643
R17850 VN.n1947 VN.t166 3.643
R17851 VN.n1962 VN.n1961 3.643
R17852 VN.n1965 VN.n1964 3.643
R17853 VN.n1950 VN.t321 3.643
R17854 VN.n1992 VN.t320 3.643
R17855 VN.n2001 VN.n2000 3.643
R17856 VN.n2004 VN.n2003 3.643
R17857 VN.n1995 VN.t123 3.643
R17858 VN.n78 VN.t328 3.643
R17859 VN.n336 VN.t155 3.643
R17860 VN.n344 VN.n343 3.643
R17861 VN.n347 VN.n346 3.643
R17862 VN.n339 VN.t85 3.643
R17863 VN.n115 VN.t323 3.643
R17864 VN.n126 VN.n125 3.643
R17865 VN.n123 VN.n122 3.643
R17866 VN.n118 VN.t125 3.643
R17867 VN.n214 VN.t152 3.643
R17868 VN.n222 VN.n221 3.643
R17869 VN.n225 VN.n224 3.643
R17870 VN.n217 VN.t324 3.643
R17871 VN.n45 VN.t70 3.643
R17872 VN.n356 VN.t288 3.643
R17873 VN.n364 VN.n363 3.643
R17874 VN.n367 VN.n366 3.643
R17875 VN.n359 VN.t201 3.643
R17876 VN.n962 VN.n961 3.643
R17877 VN.n1087 VN.t390 3.643
R17878 VN.n1205 VN.n1203 2.799
R17879 VN.n979 VN.n977 2.799
R17880 VN.n656 VN.n654 2.799
R17881 VN.n1864 VN.n1862 2.799
R17882 VN.n155 VN.n153 2.799
R17883 VN.n309 VN.n307 2.799
R17884 VN.n1529 VN.n1528 2.645
R17885 VN.n1199 VN.n1198 2.645
R17886 VN.n973 VN.n972 2.645
R17887 VN.n650 VN.n649 2.645
R17888 VN.n1858 VN.n1857 2.645
R17889 VN.n149 VN.n148 2.645
R17890 VN.n511 VN.n510 0.21
R17891 VN.n7 VN.n4 0.178
R17892 VN.n1709 VN.n1708 0.172
R17893 VN.n1531 VN.n1527 0.164
R17894 VN VN.n105 0.138
R17895 VN.n1794 VN.n1793 0.133
R17896 VN.n545 VN.n544 0.133
R17897 VN.n888 VN.n887 0.133
R17898 VN.n1357 VN.n1356 0.133
R17899 VN.n1422 VN.n1421 0.133
R17900 VN.n1729 VN.n1442 0.114
R17901 VN.n1728 VN.n1721 0.111
R17902 VN.n1730 VN.n1132 0.111
R17903 VN.n1731 VN.n808 0.111
R17904 VN.n48 VN.n47 0.11
R17905 VN.n2029 VN.n2028 0.11
R17906 VN.n2030 VN.n508 0.11
R17907 VN.n758 VN.n753 0.106
R17908 VN.n200 VN.n195 0.106
R17909 VN.n1495 VN.n1490 0.104
R17910 VN.n1182 VN.n1181 0.097
R17911 VN.n849 VN.n848 0.097
R17912 VN.n595 VN.n594 0.097
R17913 VN.n1494 VN.n1491 0.097
R17914 VN.n2021 VN.n2020 0.095
R17915 VN.n60 VN.n59 0.093
R17916 VN.n303 VN.n302 0.093
R17917 VN.n147 VN.n146 0.093
R17918 VN.n16 VN.n15 0.092
R17919 VN.n92 VN.n91 0.092
R17920 VN.n41 VN.n40 0.087
R17921 VN.n58 VN.n57 0.085
R17922 VN.n1718 VN.n1716 0.082
R17923 VN.n1142 VN.n1139 0.082
R17924 VN.n838 VN.n835 0.082
R17925 VN.n528 VN.n525 0.082
R17926 VN.n1740 VN.n1737 0.082
R17927 VN.n506 VN.n501 0.082
R17928 VN.n590 VN.n589 0.08
R17929 VN.n844 VN.n843 0.08
R17930 VN.n1177 VN.n1176 0.08
R17931 VN.n1543 VN.n1535 0.08
R17932 VN.n1543 VN.n1533 0.08
R17933 VN.n104 VN.n103 0.079
R17934 VN.n1323 VN.n1322 0.077
R17935 VN.n1014 VN.n1013 0.077
R17936 VN.n673 VN.n672 0.077
R17937 VN.n1869 VN.n1868 0.076
R17938 VN.n822 VN.n821 0.075
R17939 VN.n314 VN.n313 0.074
R17940 VN.n661 VN.n660 0.074
R17941 VN.n160 VN.n159 0.074
R17942 VN.n984 VN.n983 0.074
R17943 VN.n1210 VN.n1209 0.074
R17944 VN.n64 VN.n63 0.073
R17945 VN.n72 VN.n71 0.073
R17946 VN.n77 VN.n76 0.073
R17947 VN.n756 VN.n755 0.07
R17948 VN.n198 VN.n197 0.07
R17949 VN.t52 VN.n54 0.068
R17950 VN.n1543 VN.n1542 0.067
R17951 VN.n1593 VN.n1591 0.067
R17952 VN.n1593 VN.n1592 0.067
R17953 VN.n1559 VN.n1557 0.067
R17954 VN.n1584 VN.n1582 0.067
R17955 VN.n1584 VN.n1583 0.067
R17956 VN.n1575 VN.n1573 0.067
R17957 VN.n1575 VN.n1574 0.067
R17958 VN.n1559 VN.n1558 0.067
R17959 VN.n1718 VN.n1717 0.067
R17960 VN.n838 VN.n829 0.067
R17961 VN.n838 VN.n827 0.067
R17962 VN.n528 VN.n519 0.067
R17963 VN.n528 VN.n518 0.067
R17964 VN.n506 VN.n495 0.067
R17965 VN.n506 VN.n505 0.067
R17966 VN.n1718 VN.n1707 0.067
R17967 VN.n1619 VN.n1618 0.066
R17968 VN.n1720 VN.n1719 0.065
R17969 VN.n1741 VN.n1740 0.063
R17970 VN.n1382 VN.n1381 0.063
R17971 VN.n923 VN.n922 0.063
R17972 VN.n580 VN.n579 0.063
R17973 VN.n1769 VN.n1768 0.063
R17974 VN.n1662 VN.n1649 0.063
R17975 VN.n1168 VN.n1167 0.063
R17976 VN.n1358 VN.n1345 0.063
R17977 VN.n889 VN.n876 0.063
R17978 VN.n546 VN.n533 0.063
R17979 VN.n1641 VN.n1627 0.063
R17980 VN.n1463 VN.n1448 0.063
R17981 VN.n1693 VN.n1692 0.063
R17982 VN.n1243 VN.n1242 0.062
R17983 VN.n1594 VN.n1593 0.062
R17984 VN.n1560 VN.n1559 0.062
R17985 VN.n1549 VN.n1548 0.062
R17986 VN.n1585 VN.n1584 0.062
R17987 VN.n1576 VN.n1575 0.061
R17988 VN.n8 VN.n7 0.061
R17989 VN.n1524 VN.n1523 0.06
R17990 VN.n1640 VN.n1639 0.059
R17991 VN.n458 VN.n457 0.059
R17992 VN.n1778 VN.n1777 0.059
R17993 VN.n507 VN.n506 0.058
R17994 VN.n810 VN.n809 0.058
R17995 VN.n1720 VN.n1718 0.058
R17996 VN.n1546 VN.n1525 0.055
R17997 VN.n2010 VN.n2009 0.055
R17998 VN.n1704 VN.n1703 0.055
R17999 VN.n1434 VN.n1433 0.055
R18000 VN.n1124 VN.n1123 0.055
R18001 VN.n800 VN.n799 0.055
R18002 VN.n492 VN.n106 0.054
R18003 VN.n1212 VN.n1194 0.054
R18004 VN.n316 VN.n299 0.054
R18005 VN.n664 VN.n647 0.054
R18006 VN.n1871 VN.n1850 0.054
R18007 VN.n163 VN.n144 0.054
R18008 VN.n987 VN.n970 0.054
R18009 VN.n294 VN.n293 0.054
R18010 VN.n489 VN.n488 0.054
R18011 VN.n205 VN.n204 0.054
R18012 VN.n1699 VN.n1698 0.054
R18013 VN.n1665 VN.n1664 0.054
R18014 VN.n1385 VN.n1384 0.054
R18015 VN.n465 VN.n464 0.054
R18016 VN.n181 VN.n180 0.054
R18017 VN.n1772 VN.n1771 0.054
R18018 VN.n1908 VN.n1907 0.054
R18019 VN.n583 VN.n582 0.054
R18020 VN.n723 VN.n722 0.054
R18021 VN.n926 VN.n925 0.054
R18022 VN.n1065 VN.n1064 0.054
R18023 VN.n1289 VN.n1288 0.054
R18024 VN.n1502 VN.n1501 0.054
R18025 VN.n1171 VN.n1170 0.054
R18026 VN.n960 VN.n959 0.054
R18027 VN.n1006 VN.n1005 0.054
R18028 VN.n1253 VN.n1252 0.054
R18029 VN.n1315 VN.n1314 0.054
R18030 VN.n1622 VN.n1621 0.054
R18031 VN.n613 VN.n612 0.054
R18032 VN.n687 VN.n686 0.054
R18033 VN.n871 VN.n870 0.054
R18034 VN.n1028 VN.n1027 0.054
R18035 VN.n1340 VN.n1339 0.054
R18036 VN.n1272 VN.n1271 0.054
R18037 VN.n1361 VN.n1360 0.054
R18038 VN.n1047 VN.n1046 0.054
R18039 VN.n892 VN.n891 0.054
R18040 VN.n706 VN.n705 0.054
R18041 VN.n549 VN.n548 0.054
R18042 VN.n1891 VN.n1890 0.054
R18043 VN.n1801 VN.n1800 0.054
R18044 VN.n1644 VN.n1643 0.054
R18045 VN.n1466 VN.n1465 0.054
R18046 VN.n1412 VN.n1411 0.054
R18047 VN.n1230 VN.n1229 0.054
R18048 VN.n1309 VN.n1308 0.054
R18049 VN.n1429 VN.n1428 0.054
R18050 VN.n1107 VN.n1106 0.054
R18051 VN.n744 VN.n743 0.054
R18052 VN.n633 VN.n632 0.054
R18053 VN.n1929 VN.n1928 0.054
R18054 VN.n1821 VN.n1820 0.054
R18055 VN.n414 VN.n413 0.054
R18056 VN.n386 VN.n385 0.054
R18057 VN.n396 VN.n395 0.054
R18058 VN.n1085 VN.n1084 0.054
R18059 VN.n1122 VN.n1121 0.054
R18060 VN.n371 VN.n370 0.054
R18061 VN.n383 VN.n382 0.054
R18062 VN.n260 VN.n259 0.054
R18063 VN.n1836 VN.n1835 0.054
R18064 VN.n1945 VN.n1944 0.054
R18065 VN.n783 VN.n782 0.054
R18066 VN.n769 VN.n768 0.054
R18067 VN.n766 VN.n765 0.054
R18068 VN.n798 VN.n797 0.054
R18069 VN.n332 VN.n331 0.054
R18070 VN.n130 VN.n129 0.054
R18071 VN.n229 VN.n228 0.054
R18072 VN.n1983 VN.n1982 0.054
R18073 VN.n1969 VN.n1968 0.054
R18074 VN.n1966 VN.n1965 0.054
R18075 VN.n2005 VN.n2004 0.054
R18076 VN.n348 VN.n347 0.054
R18077 VN.n124 VN.n123 0.054
R18078 VN.n226 VN.n225 0.054
R18079 VN.n368 VN.n367 0.054
R18080 VN.n102 VN.n9 0.053
R18081 VN.t22 VN.n962 0.052
R18082 VN.n1208 VN.n1207 0.052
R18083 VN.n982 VN.n981 0.052
R18084 VN.n659 VN.n658 0.052
R18085 VN.n1867 VN.n1866 0.052
R18086 VN.n158 VN.n157 0.052
R18087 VN.n312 VN.n311 0.052
R18088 VN.n1145 VN.n1144 0.052
R18089 VN.n755 VN.n754 0.052
R18090 VN.n1130 VN.n1129 0.052
R18091 VN.n806 VN.n805 0.052
R18092 VN.n2026 VN.n2025 0.052
R18093 VN.n197 VN.n196 0.052
R18094 VN.t22 VN.n1087 0.051
R18095 VN.n952 VN.n950 0.051
R18096 VN.n1404 VN.n1402 0.051
R18097 VN.n1672 VN.n1671 0.051
R18098 VN.n20 VN.n19 0.051
R18099 VN.n22 VN.n21 0.051
R18100 VN.n88 VN.n87 0.051
R18101 VN.n435 VN.n421 0.051
R18102 VN.n380 VN.n268 0.051
R18103 VN.n1423 VN.n1413 0.051
R18104 VN.n238 VN.n237 0.051
R18105 VN.n462 VN.n461 0.05
R18106 VN.n954 VN.n953 0.05
R18107 VN.n1795 VN.n1781 0.05
R18108 VN.n1406 VN.n1405 0.05
R18109 VN.n1693 VN.n1674 0.05
R18110 VN.n1337 VN.n1325 0.05
R18111 VN.n1652 VN.n1651 0.05
R18112 VN.n1017 VN.n1016 0.049
R18113 VN.n676 VN.n675 0.049
R18114 VN.n1321 VN.n1320 0.049
R18115 VN.n511 VN.n509 0.049
R18116 VN.n1959 VN.n1958 0.048
R18117 VN.n1143 VN.n1142 0.048
R18118 VN.n839 VN.n838 0.048
R18119 VN.n529 VN.n528 0.048
R18120 VN.n288 VN.n286 0.047
R18121 VN.n483 VN.n481 0.047
R18122 VN.n202 VN.n193 0.047
R18123 VN.n2028 VN.n2012 0.047
R18124 VN.n1693 VN.n1684 0.047
R18125 VN.n1662 VN.n1660 0.047
R18126 VN.n1382 VN.n1369 0.047
R18127 VN.n462 VN.n445 0.047
R18128 VN.n178 VN.n172 0.047
R18129 VN.n1769 VN.n1755 0.047
R18130 VN.n1905 VN.n1899 0.047
R18131 VN.n580 VN.n566 0.047
R18132 VN.n720 VN.n714 0.047
R18133 VN.n923 VN.n909 0.047
R18134 VN.n1062 VN.n1055 0.047
R18135 VN.n1286 VN.n1284 0.047
R18136 VN.n1499 VN.n1483 0.047
R18137 VN.n1168 VN.n1159 0.047
R18138 VN.n954 VN.n938 0.047
R18139 VN.n1003 VN.n996 0.047
R18140 VN.n1250 VN.n1241 0.047
R18141 VN.n1324 VN.n1318 0.047
R18142 VN.n1619 VN.n1612 0.047
R18143 VN.n607 VN.n599 0.047
R18144 VN.n684 VN.n679 0.047
R18145 VN.n868 VN.n853 0.047
R18146 VN.n1025 VN.n1020 0.047
R18147 VN.n1337 VN.n1186 0.047
R18148 VN.n1269 VN.n1266 0.047
R18149 VN.n1358 VN.n1355 0.047
R18150 VN.n1044 VN.n1040 0.047
R18151 VN.n889 VN.n886 0.047
R18152 VN.n703 VN.n699 0.047
R18153 VN.n546 VN.n543 0.047
R18154 VN.n1888 VN.n1884 0.047
R18155 VN.n1795 VN.n1792 0.047
R18156 VN.n1641 VN.n1638 0.047
R18157 VN.n1463 VN.n1461 0.047
R18158 VN.n1406 VN.n1394 0.047
R18159 VN.n1227 VN.n1225 0.047
R18160 VN.n1721 VN.n1706 0.047
R18161 VN.n1303 VN.n1300 0.047
R18162 VN.n1423 VN.n1420 0.047
R18163 VN.n1101 VN.n1094 0.047
R18164 VN.n738 VN.n735 0.047
R18165 VN.n627 VN.n620 0.047
R18166 VN.n1923 VN.n1920 0.047
R18167 VN.n1815 VN.n1808 0.047
R18168 VN.n420 VN.n417 0.047
R18169 VN.n435 VN.n428 0.047
R18170 VN.n403 VN.n399 0.047
R18171 VN.n1441 VN.n1436 0.047
R18172 VN.n1079 VN.n1077 0.047
R18173 VN.n1116 VN.n1112 0.047
R18174 VN.n378 VN.n273 0.047
R18175 VN.n380 VN.n246 0.047
R18176 VN.n267 VN.n257 0.047
R18177 VN.n1830 VN.n1826 0.047
R18178 VN.n1939 VN.n1934 0.047
R18179 VN.n777 VN.n638 0.047
R18180 VN.n776 VN.n646 0.047
R18181 VN.n1132 VN.n841 0.047
R18182 VN.n760 VN.n752 0.047
R18183 VN.n792 VN.n788 0.047
R18184 VN.n326 VN.n321 0.047
R18185 VN.n238 VN.n135 0.047
R18186 VN.n236 VN.n143 0.047
R18187 VN.n1977 VN.n1841 0.047
R18188 VN.n1976 VN.n1849 0.047
R18189 VN.n808 VN.n531 0.047
R18190 VN.n1960 VN.n1951 0.047
R18191 VN.n1999 VN.n1996 0.047
R18192 VN.n342 VN.n340 0.047
R18193 VN.n121 VN.n119 0.047
R18194 VN.n220 VN.n218 0.047
R18195 VN.n362 VN.n360 0.047
R18196 VN.n1155 VN.n1154 0.047
R18197 VN.n1101 VN.t22 0.046
R18198 VN.n777 VN.n776 0.046
R18199 VN.n1977 VN.n1976 0.045
R18200 VN.n1998 VN.n1997 0.045
R18201 VN.n84 VN.n83 0.045
R18202 VN.n86 VN.n85 0.045
R18203 VN.n1244 VN.n1243 0.045
R18204 VN.n1518 VN.n1517 0.045
R18205 VN.n1334 VN.n1326 0.045
R18206 VN.n865 VN.n857 0.045
R18207 VN.n812 VN.n811 0.045
R18208 VN.n13 VN.n12 0.045
R18209 VN.n435 VN.n404 0.044
R18210 VN.n380 VN.n379 0.044
R18211 VN.n48 VN.n46 0.044
R18212 VN.n1566 VN.n1565 0.044
R18213 VN.n1452 VN.n1451 0.044
R18214 VN.n1473 VN.n1472 0.044
R18215 VN.n461 VN.n460 0.043
R18216 VN.n1781 VN.n1780 0.043
R18217 VN.n1164 VN.n1163 0.043
R18218 VN.n1455 VN.n1454 0.043
R18219 VN.n1347 VN.n1346 0.042
R18220 VN.n1765 VN.n1760 0.042
R18221 VN.n576 VN.n571 0.042
R18222 VN.n919 VN.n914 0.042
R18223 VN.n1378 VN.n1373 0.042
R18224 VN.n1606 VN.n1605 0.042
R18225 VN.n1632 VN.n1631 0.042
R18226 VN.n535 VN.n534 0.042
R18227 VN.n878 VN.n877 0.042
R18228 VN.n305 VN.n304 0.042
R18229 VN.n1629 VN.n1628 0.041
R18230 VN.n935 VN.n934 0.041
R18231 VN.n1446 VN.n1445 0.041
R18232 VN.n1544 VN.n1531 0.04
R18233 VN.n1208 VN.n1199 0.04
R18234 VN.n982 VN.n973 0.04
R18235 VN.n659 VN.n650 0.04
R18236 VN.n1867 VN.n1858 0.04
R18237 VN.n158 VN.n149 0.04
R18238 VN.n30 VN.n29 0.04
R18239 VN.n28 VN.n27 0.04
R18240 VN.n26 VN.n25 0.04
R18241 VN.n71 VN.n70 0.039
R18242 VN.n76 VN.n75 0.039
R18243 VN.n1530 VN.n1529 0.039
R18244 VN.n2017 VN.n2016 0.039
R18245 VN.n813 VN.n812 0.039
R18246 VN.n818 VN.n817 0.039
R18247 VN.n90 VN.n89 0.039
R18248 VN.n1207 VN.n1200 0.039
R18249 VN.n981 VN.n974 0.039
R18250 VN.n658 VN.n651 0.039
R18251 VN.n1866 VN.n1859 0.039
R18252 VN.n157 VN.n150 0.039
R18253 VN.n303 VN.n301 0.038
R18254 VN.n147 VN.n145 0.038
R18255 VN.n1751 VN.n1750 0.038
R18256 VN.n562 VN.n561 0.038
R18257 VN.n905 VN.n904 0.038
R18258 VN.n1688 VN.n1687 0.038
R18259 VN.n1728 VN.n1727 0.038
R18260 VN.n1686 VN.n1685 0.038
R18261 VN.n1206 VN.n1201 0.037
R18262 VN.n980 VN.n975 0.037
R18263 VN.n657 VN.n652 0.037
R18264 VN.n1865 VN.n1860 0.037
R18265 VN.n156 VN.n151 0.037
R18266 VN.n3 VN.n0 0.037
R18267 VN.n606 VN.n604 0.037
R18268 VN.n2017 VN.n2014 0.037
R18269 VN.n2016 VN.n2015 0.037
R18270 VN.n1337 VN.n1183 0.037
R18271 VN.n868 VN.n850 0.037
R18272 VN.n607 VN.n596 0.037
R18273 VN.n818 VN.n815 0.037
R18274 VN.n817 VN.n816 0.037
R18275 VN.n112 VN.n111 0.037
R18276 VN.n1989 VN.n1988 0.037
R18277 VN.n1196 VN.n1195 0.036
R18278 VN.n1721 VN.n1446 0.036
R18279 VN.n1033 VN.n1032 0.036
R18280 VN.n692 VN.n691 0.036
R18281 VN.n1877 VN.n1876 0.036
R18282 VN.n1259 VN.n1257 0.036
R18283 VN.n1219 VN.n1218 0.036
R18284 VN.n474 VN.n473 0.035
R18285 VN.n440 VN.n439 0.035
R18286 VN.n1216 VN.n1215 0.035
R18287 VN.n296 VN.n295 0.035
R18288 VN.n668 VN.n667 0.035
R18289 VN.n1875 VN.n1874 0.035
R18290 VN.n167 VN.n166 0.035
R18291 VN.n991 VN.n990 0.035
R18292 VN.n2018 VN.n2017 0.035
R18293 VN.n1751 VN.n1746 0.035
R18294 VN.n562 VN.n557 0.035
R18295 VN.n905 VN.n900 0.035
R18296 VN.n954 VN.n935 0.035
R18297 VN.n1493 VN.n1492 0.035
R18298 VN.n811 VN.n810 0.035
R18299 VN.n819 VN.n818 0.035
R18300 VN.t52 VN.n99 0.035
R18301 VN.t100 VN.n1554 0.035
R18302 VN.t100 VN.n1596 0.035
R18303 VN.t100 VN.n1562 0.035
R18304 VN.t100 VN.n1572 0.035
R18305 VN.t100 VN.n1587 0.035
R18306 VN.t100 VN.n1601 0.035
R18307 VN.t52 VN.n50 0.035
R18308 VN.t52 VN.n61 0.035
R18309 VN.t52 VN.n68 0.035
R18310 VN.t52 VN.n79 0.035
R18311 VN.t52 VN.n42 0.035
R18312 VN.n53 VN.n52 0.035
R18313 VN.n516 VN.n515 0.034
R18314 VN.n1552 VN.n1551 0.034
R18315 VN.n403 VN.n400 0.034
R18316 VN.n435 VN.n430 0.034
R18317 VN.n1815 VN.n1810 0.034
R18318 VN.n627 VN.n622 0.034
R18319 VN.n1101 VN.n1096 0.034
R18320 VN.n1441 VN.n1133 0.034
R18321 VN.n1132 VN.n1131 0.034
R18322 VN.n808 VN.n807 0.034
R18323 VN.n2028 VN.n2027 0.034
R18324 VN.n661 VN.n648 0.034
R18325 VN.n984 VN.n971 0.034
R18326 VN.n1210 VN.n1197 0.034
R18327 VN.n18 VN.n17 0.034
R18328 VN.n94 VN.n93 0.034
R18329 VN.t52 VN.n98 0.034
R18330 VN.t100 VN.n1553 0.034
R18331 VN.t100 VN.n1595 0.034
R18332 VN.t100 VN.n1561 0.034
R18333 VN.t100 VN.n1571 0.034
R18334 VN.t100 VN.n1586 0.034
R18335 VN.t100 VN.n1604 0.034
R18336 VN.t52 VN.n49 0.034
R18337 VN.t52 VN.n62 0.034
R18338 VN.t52 VN.n69 0.034
R18339 VN.t52 VN.n78 0.034
R18340 VN.t52 VN.n45 0.034
R18341 VN.n1544 VN.n1543 0.033
R18342 VN.n314 VN.n303 0.032
R18343 VN.n160 VN.n147 0.032
R18344 VN.n1012 VN.n1011 0.032
R18345 VN.n671 VN.n670 0.032
R18346 VN.n1852 VN.n1851 0.032
R18347 VN.t42 VN.n440 0.031
R18348 VN.t50 VN.n1216 0.031
R18349 VN.t7 VN.n296 0.031
R18350 VN.t13 VN.n668 0.031
R18351 VN.t2 VN.n1875 0.031
R18352 VN.t20 VN.n167 0.031
R18353 VN.t22 VN.n991 0.031
R18354 VN.n1746 VN.n1745 0.031
R18355 VN.n557 VN.n556 0.031
R18356 VN.n900 VN.n899 0.031
R18357 VN.n1444 VN.n1443 0.031
R18358 VN.n433 VN.n432 0.031
R18359 VN.n1813 VN.n1812 0.031
R18360 VN.n625 VN.n624 0.031
R18361 VN.n1099 VN.n1098 0.031
R18362 VN.n1399 VN.n1398 0.03
R18363 VN.n862 VN.n861 0.03
R18364 VN.n1331 VN.n1330 0.03
R18365 VN.n1676 VN.n1675 0.03
R18366 VN.n947 VN.n942 0.029
R18367 VN.n1378 VN.n1377 0.029
R18368 VN.n1060 VN.n1059 0.029
R18369 VN.n919 VN.n918 0.029
R18370 VN.n576 VN.n575 0.029
R18371 VN.n1765 VN.n1764 0.029
R18372 VN.n1001 VN.n1000 0.029
R18373 VN.n861 VN.n860 0.029
R18374 VN.n1330 VN.n1329 0.029
R18375 VN.n1509 VN.n1508 0.029
R18376 VN.n1746 VN.n1743 0.028
R18377 VN.n557 VN.n554 0.028
R18378 VN.n900 VN.n897 0.028
R18379 VN.n1180 VN.n1179 0.028
R18380 VN.n1182 VN.n1180 0.028
R18381 VN.n847 VN.n846 0.028
R18382 VN.n849 VN.n847 0.028
R18383 VN.n593 VN.n592 0.028
R18384 VN.n595 VN.n593 0.028
R18385 VN.n455 VN.n454 0.028
R18386 VN.n947 VN.n946 0.028
R18387 VN.n1156 VN.n1155 0.028
R18388 VN.n1716 VN.n1711 0.028
R18389 VN.n1139 VN.n1135 0.028
R18390 VN.n835 VN.n831 0.028
R18391 VN.n525 VN.n521 0.028
R18392 VN.n1737 VN.n1733 0.028
R18393 VN.n501 VN.n497 0.028
R18394 VN.n112 VN.n110 0.027
R18395 VN.n1989 VN.n1987 0.027
R18396 VN.n1619 VN.n1614 0.027
R18397 VN.n1441 VN.n1440 0.027
R18398 VN.n1098 VN.n1097 0.027
R18399 VN.n1096 VN.n1095 0.027
R18400 VN.n624 VN.n623 0.027
R18401 VN.n622 VN.n621 0.027
R18402 VN.n1812 VN.n1811 0.027
R18403 VN.n1810 VN.n1809 0.027
R18404 VN.n432 VN.n431 0.027
R18405 VN.n430 VN.n429 0.027
R18406 VN.n1382 VN.n1379 0.026
R18407 VN.n1062 VN.n1061 0.026
R18408 VN.n923 VN.n920 0.026
R18409 VN.n720 VN.n719 0.026
R18410 VN.n580 VN.n577 0.026
R18411 VN.n1905 VN.n1904 0.026
R18412 VN.n1769 VN.n1766 0.026
R18413 VN.n178 VN.n177 0.026
R18414 VN.n462 VN.n456 0.026
R18415 VN.n1286 VN.n1278 0.026
R18416 VN.n1168 VN.n1165 0.026
R18417 VN.n1003 VN.n1002 0.026
R18418 VN.n954 VN.n948 0.026
R18419 VN.n1014 VN.n1012 0.026
R18420 VN.n673 VN.n671 0.026
R18421 VN.n1358 VN.n1348 0.026
R18422 VN.n889 VN.n879 0.026
R18423 VN.n546 VN.n536 0.026
R18424 VN.n1795 VN.n1785 0.026
R18425 VN.n1887 VN.n1886 0.026
R18426 VN.n702 VN.n701 0.026
R18427 VN.n1043 VN.n1042 0.026
R18428 VN.n1641 VN.n1630 0.026
R18429 VN.n1406 VN.n1400 0.026
R18430 VN.n1693 VN.n1689 0.026
R18431 VN.n1693 VN.n1677 0.026
R18432 VN.n202 VN.n186 0.026
R18433 VN.n353 VN.n352 0.026
R18434 VN.n279 VN.n278 0.026
R18435 VN.n1486 VN.n1485 0.026
R18436 VN.t100 VN.n1522 0.025
R18437 VN.n1475 VN.n1474 0.025
R18438 VN.n1579 VN.n1578 0.024
R18439 VN.n1141 VN.n1140 0.024
R18440 VN.n837 VN.n836 0.024
R18441 VN.n527 VN.n526 0.024
R18442 VN.n1739 VN.n1738 0.024
R18443 VN.n503 VN.n502 0.024
R18444 VN.n6 VN.n5 0.024
R18445 VN.n1155 VN.n1150 0.024
R18446 VN.n1337 VN.n1178 0.024
R18447 VN.n868 VN.n845 0.024
R18448 VN.n607 VN.n591 0.024
R18449 VN.n1440 VN.n1439 0.024
R18450 VN.n1578 VN.n1577 0.024
R18451 VN.n195 VN.n194 0.023
R18452 VN.n2026 VN.n2013 0.023
R18453 VN.n97 VN.n86 0.023
R18454 VN.n1689 VN.n1686 0.023
R18455 VN.n1248 VN.n1244 0.023
R18456 VN.n1476 VN.n1473 0.023
R18457 VN.t100 VN.n1579 0.023
R18458 VN.n1853 VN.n1852 0.023
R18459 VN.n591 VN.n590 0.023
R18460 VN.n845 VN.n844 0.023
R18461 VN.n1178 VN.n1177 0.023
R18462 VN.n1337 VN.n1182 0.023
R18463 VN.n868 VN.n849 0.023
R18464 VN.n607 VN.n595 0.023
R18465 VN.n1321 VN.n1319 0.023
R18466 VN.n1453 VN.n1450 0.023
R18467 VN.n53 VN.n51 0.023
R18468 VN.n1145 VN.n1143 0.023
R18469 VN.n1438 VN.n1437 0.023
R18470 VN.n1130 VN.n1128 0.023
R18471 VN.n815 VN.n814 0.023
R18472 VN.n806 VN.n804 0.023
R18473 VN.n24 VN.n13 0.023
R18474 VN.n1150 VN.n1148 0.023
R18475 VN.n1472 VN.n1471 0.023
R18476 VN.n460 VN.n459 0.022
R18477 VN.n863 VN.n859 0.022
R18478 VN.n1332 VN.n1328 0.022
R18479 VN.n1780 VN.n1779 0.022
R18480 VN.n1512 VN.n1507 0.022
R18481 VN.n1495 VN.n1494 0.022
R18482 VN.n822 VN.n820 0.022
R18483 VN.n952 VN.n951 0.022
R18484 VN.n1404 VN.n1403 0.022
R18485 VN.n1672 VN.n1670 0.022
R18486 VN.n1784 VN.n1783 0.022
R18487 VN.n455 VN.n450 0.021
R18488 VN.n1377 VN.n1376 0.021
R18489 VN.n918 VN.n917 0.021
R18490 VN.n914 VN.n913 0.021
R18491 VN.n575 VN.n574 0.021
R18492 VN.n571 VN.n570 0.021
R18493 VN.n1764 VN.n1763 0.021
R18494 VN.n1760 VN.n1759 0.021
R18495 VN.n454 VN.n453 0.021
R18496 VN.n1651 VN.n1650 0.021
R18497 VN.n946 VN.n945 0.021
R18498 VN.n1856 VN.n1855 0.021
R18499 VN.n1745 VN.n1744 0.021
R18500 VN.n556 VN.n555 0.021
R18501 VN.n899 VN.n898 0.021
R18502 VN.n1649 VN.n1648 0.021
R18503 VN.n953 VN.n952 0.021
R18504 VN.n606 VN.n605 0.021
R18505 VN.n1405 VN.n1404 0.021
R18506 VN.n1448 VN.n1447 0.021
R18507 VN.n1674 VN.n1672 0.021
R18508 VN.n60 VN.n58 0.021
R18509 VN.n1496 VN.n1489 0.021
R18510 VN.n512 VN.n511 0.021
R18511 VN.n1247 VN.n1245 0.02
R18512 VN.n23 VN.n14 0.02
R18513 VN.n96 VN.n90 0.02
R18514 VN.n473 VN.n472 0.02
R18515 VN.n461 VN.n458 0.02
R18516 VN.n1150 VN.n1149 0.02
R18517 VN.n953 VN.n949 0.02
R18518 VN.n1781 VN.n1778 0.02
R18519 VN.n1510 VN.n1509 0.02
R18520 VN.n1405 VN.n1401 0.02
R18521 VN.n1674 VN.n1673 0.02
R18522 VN.n1716 VN.n1715 0.019
R18523 VN.n1139 VN.n1138 0.019
R18524 VN.n835 VN.n834 0.019
R18525 VN.n525 VN.n524 0.019
R18526 VN.n1737 VN.n1736 0.019
R18527 VN.n501 VN.n500 0.019
R18528 VN.t100 VN.n1566 0.019
R18529 VN.n1017 VN.n1015 0.019
R18530 VN.n676 VN.n674 0.019
R18531 VN.n1519 VN.n1518 0.019
R18532 VN.n867 VN.n866 0.019
R18533 VN.n1336 VN.n1335 0.019
R18534 VN.n1616 VN.n1615 0.018
R18535 VN.n1473 VN.n1470 0.018
R18536 VN.n1450 VN.n1449 0.018
R18537 VN.n1956 VN.n1955 0.018
R18538 VN.n1570 VN.n1569 0.018
R18539 VN.n1954 VN.n1953 0.017
R18540 VN.n1498 VN.n1497 0.017
R18541 VN.n350 VN.n349 0.017
R18542 VN.n276 VN.n275 0.017
R18543 VN.n1960 VN.n1957 0.017
R18544 VN.n2023 VN.n2022 0.017
R18545 VN.n2022 VN.n2021 0.017
R18546 VN.n825 VN.n824 0.017
R18547 VN.n823 VN.n822 0.016
R18548 VN.n1148 VN.n1147 0.015
R18549 VN.n110 VN.n109 0.015
R18550 VN.n1987 VN.n1986 0.015
R18551 VN.n450 VN.n449 0.015
R18552 VN.n865 VN.n864 0.015
R18553 VN.n864 VN.n863 0.015
R18554 VN.n863 VN.n862 0.015
R18555 VN.n1334 VN.n1333 0.015
R18556 VN.n1333 VN.n1332 0.015
R18557 VN.n1332 VN.n1331 0.015
R18558 VN.n1783 VN.n1782 0.015
R18559 VN.n1513 VN.n1512 0.015
R18560 VN.n1512 VN.n1511 0.015
R18561 VN.t52 VN.n53 0.015
R18562 VN.n1132 VN.n839 0.015
R18563 VN.n109 VN.n108 0.015
R18564 VN.n1986 VN.n1985 0.015
R18565 VN.n808 VN.n529 0.015
R18566 VN.n829 VN.n828 0.015
R18567 VN.n505 VN.n504 0.015
R18568 VN.n827 VN.n826 0.015
R18569 VN.n495 VN.n494 0.015
R18570 VN.n1748 VN.n1747 0.015
R18571 VN.n559 VN.n558 0.015
R18572 VN.n902 VN.n901 0.015
R18573 VN.n1516 VN.n1515 0.014
R18574 VN.n515 VN.n513 0.014
R18575 VN.n121 VN.n112 0.014
R18576 VN.n1999 VN.n1989 0.014
R18577 VN.n759 VN.n758 0.014
R18578 VN.n201 VN.n200 0.014
R18579 VN.n1752 VN.n1751 0.013
R18580 VN.n563 VN.n562 0.013
R18581 VN.n906 VN.n905 0.013
R18582 VN.n604 VN.n603 0.013
R18583 VN.n1489 VN.n1488 0.013
R18584 VN.n1535 VN.n1534 0.013
R18585 VN.n1533 VN.n1532 0.013
R18586 VN.n758 VN.n757 0.013
R18587 VN.n200 VN.n199 0.013
R18588 VN.t100 VN.n1520 0.012
R18589 VN.n529 VN.n517 0.012
R18590 VN.n2019 VN.n2018 0.012
R18591 VN.n1749 VN.n1748 0.012
R18592 VN.n560 VN.n559 0.012
R18593 VN.n903 VN.n902 0.012
R18594 VN.n1662 VN.n1653 0.012
R18595 VN.n1153 VN.n1152 0.012
R18596 VN.n1494 VN.n1493 0.012
R18597 VN.n1463 VN.n1453 0.012
R18598 VN.n757 VN.n756 0.012
R18599 VN.n820 VN.n819 0.012
R18600 VN.n21 VN.n20 0.012
R18601 VN.n89 VN.n88 0.012
R18602 VN.n199 VN.n198 0.012
R18603 VN.n1499 VN.n1486 0.011
R18604 VN.n288 VN.n279 0.011
R18605 VN.n362 VN.n353 0.011
R18606 VN.n1960 VN.n1954 0.01
R18607 VN.n1259 VN.n1258 0.01
R18608 VN.n933 VN.n932 0.01
R18609 VN.n1476 VN.n1475 0.01
R18610 VN.n1025 VN.n1017 0.01
R18611 VN.n684 VN.n676 0.01
R18612 VN.n1888 VN.n1885 0.01
R18613 VN.n703 VN.n700 0.01
R18614 VN.n1044 VN.n1041 0.01
R18615 VN.n1269 VN.n1267 0.01
R18616 VN.n1511 VN.n1510 0.01
R18617 VN.n1324 VN.n1321 0.01
R18618 VN.n1499 VN.n1498 0.01
R18619 VN.n1303 VN.n1301 0.01
R18620 VN.n1441 VN.n1438 0.01
R18621 VN.n1441 VN.n1145 0.01
R18622 VN.n1132 VN.n1130 0.01
R18623 VN.n808 VN.n806 0.01
R18624 VN.n362 VN.n350 0.01
R18625 VN.n288 VN.n276 0.01
R18626 VN.n2028 VN.n2026 0.01
R18627 VN.n1619 VN.n1516 0.01
R18628 VN.n1453 VN.n1452 0.01
R18629 VN.n2021 VN.n2019 0.01
R18630 VN.n1870 VN.n1856 0.01
R18631 VN.n508 VN.n493 0.009
R18632 VN.n2024 VN.n2023 0.009
R18633 VN.n607 VN.n606 0.009
R18634 VN.t52 VN.n60 0.009
R18635 VN.n1729 VN.n1728 0.009
R18636 VN.n1730 VN.n1729 0.009
R18637 VN.n1731 VN.n1730 0.009
R18638 VN.n2029 VN.n1731 0.009
R18639 VN.n2030 VN.n2029 0.009
R18640 VN.n2028 VN.n1741 0.009
R18641 VN.n1497 VN.n1496 0.008
R18642 VN.n23 VN.n22 0.008
R18643 VN.n96 VN.n95 0.008
R18644 VN.n1750 VN.n1749 0.008
R18645 VN.n561 VN.n560 0.008
R18646 VN.n904 VN.n903 0.008
R18647 VN.n1381 VN.n1380 0.008
R18648 VN.n916 VN.n915 0.008
R18649 VN.n922 VN.n921 0.008
R18650 VN.n573 VN.n572 0.008
R18651 VN.n579 VN.n578 0.008
R18652 VN.n1762 VN.n1761 0.008
R18653 VN.n1768 VN.n1767 0.008
R18654 VN.n452 VN.n451 0.008
R18655 VN.n1375 VN.n1374 0.008
R18656 VN.n1167 VN.n1166 0.008
R18657 VN.n944 VN.n943 0.008
R18658 VN.n1025 VN.n1014 0.008
R18659 VN.n684 VN.n673 0.008
R18660 VN.n1345 VN.n1344 0.008
R18661 VN.n876 VN.n875 0.008
R18662 VN.n533 VN.n532 0.008
R18663 VN.n1888 VN.n1887 0.008
R18664 VN.n703 VN.n702 0.008
R18665 VN.n1044 VN.n1043 0.008
R18666 VN.n1269 VN.n1268 0.008
R18667 VN.n1627 VN.n1626 0.008
R18668 VN.n1324 VN.n1323 0.008
R18669 VN.n1692 VN.n1690 0.008
R18670 VN.n1723 VN.n1722 0.008
R18671 VN.n1724 VN.n1723 0.008
R18672 VN.n1725 VN.n1724 0.008
R18673 VN.n1726 VN.n1725 0.008
R18674 VN.n1727 VN.n1726 0.008
R18675 VN.n1303 VN.n1302 0.008
R18676 VN.n1721 VN.n1444 0.008
R18677 VN.n1960 VN.n1959 0.008
R18678 VN VN.n2030 0.008
R18679 VN.n471 VN.n470 0.008
R18680 VN.n1618 VN.n1617 0.008
R18681 VN.n1618 VN.n1616 0.007
R18682 VN.n1249 VN.n1248 0.007
R18683 VN.t100 VN.n1552 0.007
R18684 VN.n1515 VN.n1514 0.007
R18685 VN.t52 VN.n67 0.006
R18686 VN.t52 VN.n80 0.006
R18687 VN.n1376 VN.n1375 0.006
R18688 VN.n917 VN.n916 0.006
R18689 VN.n574 VN.n573 0.006
R18690 VN.n1763 VN.n1762 0.006
R18691 VN.n453 VN.n452 0.006
R18692 VN.n945 VN.n944 0.006
R18693 VN.n1692 VN.n1691 0.006
R18694 VN.n472 VN.n471 0.006
R18695 VN.n1250 VN.n1249 0.006
R18696 VN.n1248 VN.n1247 0.006
R18697 VN.n24 VN.n23 0.006
R18698 VN.n97 VN.n96 0.006
R18699 VN.n1247 VN.n1246 0.006
R18700 VN.n1499 VN.n1476 0.006
R18701 VN.n1154 VN.n1153 0.005
R18702 VN.t100 VN.n1564 0.005
R18703 VN.n22 VN.n18 0.005
R18704 VN.n95 VN.n94 0.005
R18705 VN.t100 VN.n1576 0.005
R18706 VN.n286 VN.n285 0.004
R18707 VN.n481 VN.n480 0.004
R18708 VN.n193 VN.n192 0.004
R18709 VN.n2012 VN.n2011 0.004
R18710 VN.n1684 VN.n1683 0.004
R18711 VN.n1660 VN.n1659 0.004
R18712 VN.n1369 VN.n1368 0.004
R18713 VN.n445 VN.n444 0.004
R18714 VN.n172 VN.n171 0.004
R18715 VN.n1755 VN.n1754 0.004
R18716 VN.n1899 VN.n1898 0.004
R18717 VN.n566 VN.n565 0.004
R18718 VN.n714 VN.n713 0.004
R18719 VN.n909 VN.n908 0.004
R18720 VN.n1055 VN.n1054 0.004
R18721 VN.n1284 VN.n1283 0.004
R18722 VN.n1483 VN.n1482 0.004
R18723 VN.n1159 VN.n1158 0.004
R18724 VN.n938 VN.n937 0.004
R18725 VN.n996 VN.n995 0.004
R18726 VN.n1241 VN.n1240 0.004
R18727 VN.n1318 VN.n1317 0.004
R18728 VN.n1612 VN.n1611 0.004
R18729 VN.n599 VN.n598 0.004
R18730 VN.n679 VN.n678 0.004
R18731 VN.n853 VN.n852 0.004
R18732 VN.n1020 VN.n1019 0.004
R18733 VN.n1186 VN.n1185 0.004
R18734 VN.n1266 VN.n1265 0.004
R18735 VN.n1355 VN.n1354 0.004
R18736 VN.n1040 VN.n1039 0.004
R18737 VN.n886 VN.n885 0.004
R18738 VN.n699 VN.n698 0.004
R18739 VN.n543 VN.n542 0.004
R18740 VN.n1884 VN.n1883 0.004
R18741 VN.n1792 VN.n1791 0.004
R18742 VN.n1638 VN.n1637 0.004
R18743 VN.n1461 VN.n1460 0.004
R18744 VN.n1394 VN.n1393 0.004
R18745 VN.n1225 VN.n1224 0.004
R18746 VN.n1706 VN.n1705 0.004
R18747 VN.n1300 VN.n1299 0.004
R18748 VN.n1420 VN.n1419 0.004
R18749 VN.n1094 VN.n1093 0.004
R18750 VN.n735 VN.n734 0.004
R18751 VN.n620 VN.n619 0.004
R18752 VN.n1920 VN.n1919 0.004
R18753 VN.n1808 VN.n1807 0.004
R18754 VN.n417 VN.n416 0.004
R18755 VN.n428 VN.n427 0.004
R18756 VN.n399 VN.n398 0.004
R18757 VN.n1436 VN.n1435 0.004
R18758 VN.n1077 VN.n1076 0.004
R18759 VN.n1112 VN.n1111 0.004
R18760 VN.n273 VN.n272 0.004
R18761 VN.n246 VN.n245 0.004
R18762 VN.n257 VN.n256 0.004
R18763 VN.n1826 VN.n1825 0.004
R18764 VN.n1934 VN.n1933 0.004
R18765 VN.n638 VN.n637 0.004
R18766 VN.n646 VN.n645 0.004
R18767 VN.n841 VN.n840 0.004
R18768 VN.n752 VN.n751 0.004
R18769 VN.n788 VN.n787 0.004
R18770 VN.n321 VN.n320 0.004
R18771 VN.n135 VN.n134 0.004
R18772 VN.n143 VN.n142 0.004
R18773 VN.n1841 VN.n1840 0.004
R18774 VN.n1849 VN.n1848 0.004
R18775 VN.n531 VN.n530 0.004
R18776 VN.n1951 VN.n1950 0.004
R18777 VN.n1996 VN.n1995 0.004
R18778 VN.n340 VN.n339 0.004
R18779 VN.n119 VN.n118 0.004
R18780 VN.n218 VN.n217 0.004
R18781 VN.n360 VN.n359 0.004
R18782 VN.n1641 VN.n1640 0.004
R18783 VN.t100 VN.n1570 0.004
R18784 VN.n1662 VN.n1661 0.004
R18785 VN.n1463 VN.n1462 0.004
R18786 VN.t100 VN.n1585 0.004
R18787 VN.n1211 VN.n1196 0.004
R18788 VN.n663 VN.n662 0.004
R18789 VN.n859 VN.n858 0.004
R18790 VN.n1328 VN.n1327 0.004
R18791 VN.n1507 VN.n1506 0.004
R18792 VN.n315 VN.n314 0.004
R18793 VN.n663 VN.n661 0.004
R18794 VN.n1044 VN.n1033 0.004
R18795 VN.n703 VN.n692 0.004
R18796 VN.n1888 VN.n1877 0.004
R18797 VN.n162 VN.n160 0.004
R18798 VN.n1269 VN.n1259 0.004
R18799 VN.n986 VN.n984 0.004
R18800 VN.n1211 VN.n1210 0.004
R18801 VN.n1152 VN.n1151 0.004
R18802 VN.n1870 VN.n1853 0.004
R18803 VN.n867 VN.n865 0.004
R18804 VN.n1336 VN.n1334 0.004
R18805 VN.n1488 VN.n1487 0.004
R18806 VN.n825 VN.n813 0.004
R18807 VN.n1132 VN.n825 0.004
R18808 VN.n211 VN.n210 0.004
R18809 VN.n517 VN.n516 0.004
R18810 VN.n808 VN.n512 0.004
R18811 VN.t52 VN.n64 0.004
R18812 VN.t52 VN.n72 0.004
R18813 VN.t52 VN.n77 0.004
R18814 VN.t50 VN.n1214 0.004
R18815 VN.t100 VN.n1556 0.004
R18816 VN.t100 VN.n1600 0.004
R18817 VN.t7 VN.n298 0.004
R18818 VN.t100 VN.n1568 0.004
R18819 VN.t13 VN.n666 0.004
R18820 VN.t100 VN.n1581 0.004
R18821 VN.t2 VN.n1873 0.004
R18822 VN.t100 VN.n1590 0.004
R18823 VN.t20 VN.n165 0.004
R18824 VN.t100 VN.n1603 0.004
R18825 VN.t22 VN.n989 0.004
R18826 VN.t100 VN.n1547 0.004
R18827 VN.t52 VN.n101 0.004
R18828 VN.t52 VN.n56 0.004
R18829 VN.t52 VN.n66 0.004
R18830 VN.t52 VN.n74 0.004
R18831 VN.t52 VN.n82 0.004
R18832 VN.t52 VN.n44 0.004
R18833 VN.t100 VN.n1598 0.004
R18834 VN.t52 VN.n48 0.004
R18835 VN.t42 VN.n491 0.004
R18836 VN.t100 VN.n1524 0.004
R18837 VN.t100 VN.n1594 0.004
R18838 VN.t100 VN.n1560 0.004
R18839 VN.t100 VN.n1549 0.004
R18840 VN.n162 VN.n161 0.004
R18841 VN.n1003 VN.n993 0.004
R18842 VN.n291 VN.n290 0.003
R18843 VN.n486 VN.n485 0.003
R18844 VN.n208 VN.n207 0.003
R18845 VN.n2008 VN.n2007 0.003
R18846 VN.n1696 VN.n1695 0.003
R18847 VN.n1668 VN.n1667 0.003
R18848 VN.n1388 VN.n1387 0.003
R18849 VN.n468 VN.n467 0.003
R18850 VN.n184 VN.n183 0.003
R18851 VN.n1775 VN.n1774 0.003
R18852 VN.n1911 VN.n1910 0.003
R18853 VN.n586 VN.n585 0.003
R18854 VN.n726 VN.n725 0.003
R18855 VN.n929 VN.n928 0.003
R18856 VN.n1068 VN.n1067 0.003
R18857 VN.n1292 VN.n1291 0.003
R18858 VN.n1505 VN.n1504 0.003
R18859 VN.n1174 VN.n1173 0.003
R18860 VN.n957 VN.n956 0.003
R18861 VN.n1009 VN.n1008 0.003
R18862 VN.n1256 VN.n1255 0.003
R18863 VN.n1312 VN.n1311 0.003
R18864 VN.n1625 VN.n1624 0.003
R18865 VN.n610 VN.n609 0.003
R18866 VN.n690 VN.n689 0.003
R18867 VN.n874 VN.n873 0.003
R18868 VN.n1031 VN.n1030 0.003
R18869 VN.n1343 VN.n1342 0.003
R18870 VN.n1275 VN.n1274 0.003
R18871 VN.n1364 VN.n1363 0.003
R18872 VN.n1050 VN.n1049 0.003
R18873 VN.n895 VN.n894 0.003
R18874 VN.n709 VN.n708 0.003
R18875 VN.n552 VN.n551 0.003
R18876 VN.n1894 VN.n1893 0.003
R18877 VN.n1798 VN.n1797 0.003
R18878 VN.n1647 VN.n1646 0.003
R18879 VN.n1469 VN.n1468 0.003
R18880 VN.n1409 VN.n1408 0.003
R18881 VN.n1233 VN.n1232 0.003
R18882 VN.n1702 VN.n1701 0.003
R18883 VN.n1306 VN.n1305 0.003
R18884 VN.n1426 VN.n1425 0.003
R18885 VN.n1104 VN.n1103 0.003
R18886 VN.n741 VN.n740 0.003
R18887 VN.n630 VN.n629 0.003
R18888 VN.n1926 VN.n1925 0.003
R18889 VN.n1818 VN.n1817 0.003
R18890 VN.n411 VN.n410 0.003
R18891 VN.n438 VN.n437 0.003
R18892 VN.n393 VN.n392 0.003
R18893 VN.n1432 VN.n1431 0.003
R18894 VN.n1082 VN.n1081 0.003
R18895 VN.n1119 VN.n1118 0.003
R18896 VN.n374 VN.n373 0.003
R18897 VN.n249 VN.n248 0.003
R18898 VN.n263 VN.n262 0.003
R18899 VN.n1833 VN.n1832 0.003
R18900 VN.n1942 VN.n1941 0.003
R18901 VN.n780 VN.n779 0.003
R18902 VN.n772 VN.n771 0.003
R18903 VN.n1127 VN.n1126 0.003
R18904 VN.n763 VN.n762 0.003
R18905 VN.n795 VN.n794 0.003
R18906 VN.n329 VN.n328 0.003
R18907 VN.n241 VN.n240 0.003
R18908 VN.n232 VN.n231 0.003
R18909 VN.n1980 VN.n1979 0.003
R18910 VN.n1972 VN.n1971 0.003
R18911 VN.n803 VN.n802 0.003
R18912 VN.n1963 VN.n1962 0.003
R18913 VN.n2002 VN.n2001 0.003
R18914 VN.n345 VN.n344 0.003
R18915 VN.n127 VN.n126 0.003
R18916 VN.n223 VN.n222 0.003
R18917 VN.n365 VN.n364 0.003
R18918 VN.n288 VN.n283 0.003
R18919 VN.n483 VN.n478 0.003
R18920 VN.n202 VN.n190 0.003
R18921 VN.n1693 VN.n1681 0.003
R18922 VN.n1662 VN.n1657 0.003
R18923 VN.n1382 VN.n1372 0.003
R18924 VN.n462 VN.n448 0.003
R18925 VN.n178 VN.n175 0.003
R18926 VN.n1769 VN.n1758 0.003
R18927 VN.n1905 VN.n1902 0.003
R18928 VN.n580 VN.n569 0.003
R18929 VN.n720 VN.n717 0.003
R18930 VN.n923 VN.n912 0.003
R18931 VN.n1062 VN.n1058 0.003
R18932 VN.n1286 VN.n1281 0.003
R18933 VN.n1499 VN.n1480 0.003
R18934 VN.n1168 VN.n1162 0.003
R18935 VN.n954 VN.n941 0.003
R18936 VN.n1003 VN.n999 0.003
R18937 VN.n1250 VN.n1238 0.003
R18938 VN.n1324 VN.n1193 0.003
R18939 VN.n1619 VN.n1609 0.003
R18940 VN.n607 VN.n602 0.003
R18941 VN.n684 VN.n682 0.003
R18942 VN.n868 VN.n856 0.003
R18943 VN.n1025 VN.n1023 0.003
R18944 VN.n1337 VN.n1189 0.003
R18945 VN.n1269 VN.n1263 0.003
R18946 VN.n1358 VN.n1352 0.003
R18947 VN.n1044 VN.n1037 0.003
R18948 VN.n889 VN.n883 0.003
R18949 VN.n703 VN.n696 0.003
R18950 VN.n546 VN.n540 0.003
R18951 VN.n1888 VN.n1881 0.003
R18952 VN.n1795 VN.n1789 0.003
R18953 VN.n1641 VN.n1635 0.003
R18954 VN.n1463 VN.n1458 0.003
R18955 VN.n1406 VN.n1397 0.003
R18956 VN.n1227 VN.n1222 0.003
R18957 VN.n1303 VN.n1297 0.003
R18958 VN.n1423 VN.n1417 0.003
R18959 VN.n1101 VN.n1091 0.003
R18960 VN.n738 VN.n732 0.003
R18961 VN.n627 VN.n617 0.003
R18962 VN.n1923 VN.n1917 0.003
R18963 VN.n1815 VN.n1805 0.003
R18964 VN.n420 VN.n408 0.003
R18965 VN.n435 VN.n425 0.003
R18966 VN.n403 VN.n390 0.003
R18967 VN.n1079 VN.n1074 0.003
R18968 VN.n1116 VN.n1115 0.003
R18969 VN.n378 VN.n377 0.003
R18970 VN.n380 VN.n252 0.003
R18971 VN.n267 VN.n266 0.003
R18972 VN.n1830 VN.n1829 0.003
R18973 VN.n1939 VN.n1937 0.003
R18974 VN.n777 VN.n641 0.003
R18975 VN.n776 VN.n775 0.003
R18976 VN.n760 VN.n749 0.003
R18977 VN.n792 VN.n791 0.003
R18978 VN.n326 VN.n324 0.003
R18979 VN.n238 VN.n138 0.003
R18980 VN.n236 VN.n235 0.003
R18981 VN.n1977 VN.n1844 0.003
R18982 VN.n1976 VN.n1975 0.003
R18983 VN.n1960 VN.n1948 0.003
R18984 VN.n1999 VN.n1993 0.003
R18985 VN.n342 VN.n337 0.003
R18986 VN.n121 VN.n116 0.003
R18987 VN.n220 VN.n215 0.003
R18988 VN.n362 VN.n357 0.003
R18989 VN.n1721 VN.n1720 0.003
R18990 VN.n1522 VN.n1521 0.003
R18991 VN.n105 VN.n8 0.003
R18992 VN.n105 VN.n104 0.003
R18993 VN.n1870 VN.n1869 0.003
R18994 VN.n1689 VN.n1688 0.003
R18995 VN.n1855 VN.n1854 0.003
R18996 VN.n868 VN.n867 0.003
R18997 VN.n1337 VN.n1336 0.003
R18998 VN.n220 VN.n211 0.003
R18999 VN.n508 VN.n507 0.003
R19000 VN.n1227 VN.n1219 0.003
R19001 VN.t22 VN.n969 0.003
R19002 VN.t22 VN.n967 0.003
R19003 VN.t52 VN.n10 0.003
R19004 VN.n315 VN.n300 0.003
R19005 VN.n986 VN.n985 0.003
R19006 VN.n1785 VN.n1784 0.003
R19007 VN.n483 VN.n474 0.003
R19008 VN.t52 VN.n41 0.003
R19009 VN.t52 VN.n84 0.003
R19010 VN.n1653 VN.n1652 0.003
R19011 VN.n1514 VN.n1513 0.003
R19012 VN.n108 VN.n107 0.003
R19013 VN.n1985 VN.n1984 0.003
R19014 VN.n1619 VN.n1606 0.002
R19015 VN.n1324 VN.n1190 0.002
R19016 VN.n1337 VN.n1175 0.002
R19017 VN.n1025 VN.n1010 0.002
R19018 VN.n868 VN.n842 0.002
R19019 VN.n684 VN.n669 0.002
R19020 VN.n1888 VN.n1878 0.002
R19021 VN.n546 VN.n537 0.002
R19022 VN.n703 VN.n693 0.002
R19023 VN.n889 VN.n880 0.002
R19024 VN.n1044 VN.n1034 0.002
R19025 VN.n1641 VN.n1632 0.002
R19026 VN.n1269 VN.n1260 0.002
R19027 VN.n1358 VN.n1349 0.002
R19028 VN.n1227 VN.n1217 0.002
R19029 VN.n1463 VN.n1455 0.002
R19030 VN.n403 VN.n387 0.002
R19031 VN.n435 VN.n422 0.002
R19032 VN.n420 VN.n405 0.002
R19033 VN.n1815 VN.n1802 0.002
R19034 VN.n1923 VN.n1914 0.002
R19035 VN.n627 VN.n614 0.002
R19036 VN.n738 VN.n729 0.002
R19037 VN.n1423 VN.n1414 0.002
R19038 VN.t22 VN.n963 0.002
R19039 VN.n1101 VN.n1088 0.002
R19040 VN.n378 VN.n269 0.002
R19041 VN.n380 VN.n242 0.002
R19042 VN.n267 VN.n253 0.002
R19043 VN.n1830 VN.n1822 0.002
R19044 VN.n1939 VN.n1930 0.002
R19045 VN.n777 VN.n634 0.002
R19046 VN.n776 VN.n642 0.002
R19047 VN.n1116 VN.n1108 0.002
R19048 VN.n1079 VN.n1071 0.002
R19049 VN.n326 VN.n317 0.002
R19050 VN.n238 VN.n131 0.002
R19051 VN.n236 VN.n139 0.002
R19052 VN.n1977 VN.n1837 0.002
R19053 VN.n1976 VN.n1845 0.002
R19054 VN.n792 VN.n784 0.002
R19055 VN.n760 VN.n746 0.002
R19056 VN.n220 VN.n212 0.002
R19057 VN.n121 VN.n113 0.002
R19058 VN.n342 VN.n334 0.002
R19059 VN.n1960 VN.n1952 0.002
R19060 VN.n1999 VN.n1990 0.002
R19061 VN.n202 VN.n187 0.002
R19062 VN.n483 VN.n475 0.002
R19063 VN.n288 VN.n280 0.002
R19064 VN.n607 VN.n588 0.002
R19065 VN.n1795 VN.n1786 0.002
R19066 VN.n1406 VN.n1390 0.002
R19067 VN.n824 VN.n823 0.002
R19068 VN.n1496 VN.n1495 0.002
R19069 VN.n17 VN.n16 0.002
R19070 VN.n93 VN.n92 0.002
R19071 VN.n32 VN.n31 0.002
R19072 VN.n35 VN.n34 0.002
R19073 VN.n38 VN.n37 0.002
R19074 VN.t100 VN.n1588 0.002
R19075 VN.n1423 VN.n1422 0.002
R19076 VN.n1677 VN.n1676 0.002
R19077 VN.n456 VN.n455 0.002
R19078 VN.n948 VN.n947 0.002
R19079 VN.n1382 VN.n1366 0.002
R19080 VN.n1116 VN.n1109 0.002
R19081 VN.n792 VN.n785 0.002
R19082 VN.n220 VN.n219 0.002
R19083 VN.n121 VN.n120 0.002
R19084 VN.n342 VN.n341 0.002
R19085 VN.n202 VN.n201 0.002
R19086 VN.n483 VN.n482 0.002
R19087 VN.n288 VN.n287 0.002
R19088 VN.n1400 VN.n1399 0.002
R19089 VN.n178 VN.n169 0.002
R19090 VN.n1769 VN.n1752 0.002
R19091 VN.n1905 VN.n1896 0.002
R19092 VN.n580 VN.n563 0.002
R19093 VN.n720 VN.n711 0.002
R19094 VN.n923 VN.n906 0.002
R19095 VN.n1062 VN.n1052 0.002
R19096 VN.n1286 VN.n1285 0.002
R19097 VN.n1227 VN.n1226 0.002
R19098 VN.n378 VN.n270 0.002
R19099 VN.n380 VN.n243 0.002
R19100 VN.n267 VN.n254 0.002
R19101 VN.n1830 VN.n1823 0.002
R19102 VN.n1939 VN.n1931 0.002
R19103 VN.n777 VN.n635 0.002
R19104 VN.n776 VN.n643 0.002
R19105 VN.n1079 VN.n1078 0.002
R19106 VN.n326 VN.n318 0.002
R19107 VN.n238 VN.n132 0.002
R19108 VN.n236 VN.n140 0.002
R19109 VN.n1977 VN.n1838 0.002
R19110 VN.n1976 VN.n1846 0.002
R19111 VN.n760 VN.n759 0.002
R19112 VN.n1999 VN.n1998 0.002
R19113 VN.n362 VN.n361 0.002
R19114 VN.n1619 VN.n1519 0.002
R19115 VN.n1960 VN.n1956 0.002
R19116 VN.n1541 VN.n1540 0.002
R19117 VN.t52 VN.n24 0.002
R19118 VN.t52 VN.n97 0.002
R19119 VN.n462 VN.n442 0.002
R19120 VN.n1406 VN.n1391 0.002
R19121 VN.n1545 VN.n1544 0.002
R19122 VN.n1795 VN.n1794 0.002
R19123 VN.n546 VN.n545 0.002
R19124 VN.n889 VN.n888 0.002
R19125 VN.n1358 VN.n1357 0.002
R19126 VN.n760 VN.n745 0.002
R19127 VN.n237 VN.n236 0.002
R19128 VN.n326 VN.n325 0.002
R19129 VN.n342 VN.n333 0.002
R19130 VN.n684 VN.n683 0.002
R19131 VN.n1025 VN.n1024 0.002
R19132 VN.n1325 VN.n1324 0.002
R19133 VN.n738 VN.n728 0.002
R19134 VN.n1923 VN.n1913 0.002
R19135 VN.n421 VN.n420 0.002
R19136 VN.n404 VN.n403 0.002
R19137 VN.n1079 VN.n1070 0.002
R19138 VN.n1939 VN.n1938 0.002
R19139 VN.n268 VN.n267 0.002
R19140 VN.n379 VN.n378 0.002
R19141 VN.n1693 VN.n1678 0.002
R19142 VN.n462 VN.n441 0.002
R19143 VN.n178 VN.n168 0.002
R19144 VN.n1769 VN.n1742 0.002
R19145 VN.n1905 VN.n1895 0.002
R19146 VN.n580 VN.n553 0.002
R19147 VN.n720 VN.n710 0.002
R19148 VN.n923 VN.n896 0.002
R19149 VN.n1062 VN.n1051 0.002
R19150 VN.n1382 VN.n1365 0.002
R19151 VN.n1286 VN.n1276 0.002
R19152 VN.n1662 VN.n1654 0.002
R19153 VN.n954 VN.n931 0.002
R19154 VN.n1003 VN.n992 0.002
R19155 VN.n1168 VN.n1146 0.002
R19156 VN.n1250 VN.n1234 0.002
R19157 VN.n1499 VN.n1477 0.002
R19158 VN.n362 VN.n354 0.002
R19159 VN.n105 VN.n102 0.002
R19160 VN.n1630 VN.n1629 0.002
R19161 VN.n40 VN.n33 0.001
R19162 VN.n40 VN.n36 0.001
R19163 VN.n40 VN.n39 0.001
R19164 VN.n2 VN.n1 0.001
R19165 VN.n1165 VN.n1164 0.001
R19166 VN.n1546 VN.n1545 0.001
R19167 VN.t100 VN.n1546 0.001
R19168 VN.n536 VN.n535 0.001
R19169 VN.n879 VN.n878 0.001
R19170 VN.n102 VN.t52 0.001
R19171 VN.n515 VN.n514 0.001
R19172 VN.n1168 VN.n1156 0.001
R19173 VN.n2025 VN.n2024 0.001
R19174 VN.n1379 VN.n1378 0.001
R19175 VN.n1061 VN.n1060 0.001
R19176 VN.n920 VN.n919 0.001
R19177 VN.n719 VN.n718 0.001
R19178 VN.n577 VN.n576 0.001
R19179 VN.n1904 VN.n1903 0.001
R19180 VN.n1766 VN.n1765 0.001
R19181 VN.n177 VN.n176 0.001
R19182 VN.n1278 VN.n1277 0.001
R19183 VN.n1002 VN.n1001 0.001
R19184 VN.n1348 VN.n1347 0.001
R19185 VN.n1303 VN.n1294 0.001
R19186 VN.t100 VN.n1550 0.001
R19187 VN.n1605 VN.t100 0.001
R19188 VN.t100 VN.n1597 0.001
R19189 VN.t100 VN.n1563 0.001
R19190 VN.n1207 VN.n1206 0.001
R19191 VN.n981 VN.n980 0.001
R19192 VN.n658 VN.n657 0.001
R19193 VN.n1866 VN.n1865 0.001
R19194 VN.n157 VN.n156 0.001
R19195 VN.n4 VN.n3 0.001
R19196 VN.n316 VN.n315 0.001
R19197 VN.n664 VN.n663 0.001
R19198 VN.n1871 VN.n1870 0.001
R19199 VN.n163 VN.n162 0.001
R19200 VN.n987 VN.n986 0.001
R19201 VN.n1212 VN.n1211 0.001
R19202 VN.n508 VN.n492 0.001
R19203 VN.n1541 VN.n1539 0.001
R19204 VN.n954 VN.n933 0.001
R19205 VN.n1485 VN.n1484 0.001
R19206 VN.n403 VN.n402 0.001
R19207 VN.n435 VN.n434 0.001
R19208 VN.n420 VN.n419 0.001
R19209 VN.n1815 VN.n1814 0.001
R19210 VN.n1923 VN.n1922 0.001
R19211 VN.n627 VN.n626 0.001
R19212 VN.n738 VN.n737 0.001
R19213 VN.n1101 VN.n1100 0.001
R19214 VN.t22 VN.n965 0.001
R19215 VN.n352 VN.n351 0.001
R19216 VN.n278 VN.n277 0.001
R19217 VN.n1205 VN.n1204 0.001
R19218 VN.n979 VN.n978 0.001
R19219 VN.n656 VN.n655 0.001
R19220 VN.n1864 VN.n1863 0.001
R19221 VN.n155 VN.n154 0.001
R19222 VN.n309 VN.n308 0.001
R19223 VN.n492 VN.t42 0.001
R19224 VN.t50 VN.n1212 0.001
R19225 VN.t7 VN.n316 0.001
R19226 VN.t13 VN.n664 0.001
R19227 VN.t2 VN.n1871 0.001
R19228 VN.t20 VN.n163 0.001
R19229 VN.t22 VN.n987 0.001
R19230 VN.n1442 VN.n1441 0.001
R19231 VN.n3 VN.n2 0.001
R19232 VN.n1206 VN.n1205 0.001
R19233 VN.n980 VN.n979 0.001
R19234 VN.n657 VN.n656 0.001
R19235 VN.n1865 VN.n1864 0.001
R19236 VN.n156 VN.n155 0.001
R19237 VN.n311 VN.n305 0.001
R19238 VN.n40 VN.n30 0.001
R19239 VN.n186 VN.n185 0.001
R19240 VN.n1250 VN.n1235 0.001
R19241 VN.n1542 VN.n1541 0.001
R19242 VN.n1715 VN.n1714 0.001
R19243 VN.n1138 VN.n1137 0.001
R19244 VN.n834 VN.n833 0.001
R19245 VN.n524 VN.n523 0.001
R19246 VN.n1736 VN.n1735 0.001
R19247 VN.n500 VN.n499 0.001
R19248 VN.n1614 VN.n1613 0.001
R19249 VN.n1541 VN.n1536 0.001
R19250 VN.n1541 VN.n1537 0.001
R19251 VN.n283 VN.n282 0.001
R19252 VN.n478 VN.n477 0.001
R19253 VN.n190 VN.n189 0.001
R19254 VN.n1681 VN.n1680 0.001
R19255 VN.n1657 VN.n1656 0.001
R19256 VN.n1372 VN.n1371 0.001
R19257 VN.n448 VN.n447 0.001
R19258 VN.n175 VN.n174 0.001
R19259 VN.n1758 VN.n1757 0.001
R19260 VN.n1902 VN.n1901 0.001
R19261 VN.n569 VN.n568 0.001
R19262 VN.n717 VN.n716 0.001
R19263 VN.n912 VN.n911 0.001
R19264 VN.n1058 VN.n1057 0.001
R19265 VN.n1281 VN.n1280 0.001
R19266 VN.n1480 VN.n1479 0.001
R19267 VN.n1162 VN.n1161 0.001
R19268 VN.n941 VN.n940 0.001
R19269 VN.n999 VN.n998 0.001
R19270 VN.n1238 VN.n1237 0.001
R19271 VN.n1193 VN.n1192 0.001
R19272 VN.n1609 VN.n1608 0.001
R19273 VN.n602 VN.n601 0.001
R19274 VN.n682 VN.n681 0.001
R19275 VN.n856 VN.n855 0.001
R19276 VN.n1023 VN.n1022 0.001
R19277 VN.n1189 VN.n1188 0.001
R19278 VN.n1263 VN.n1262 0.001
R19279 VN.n1352 VN.n1351 0.001
R19280 VN.n1037 VN.n1036 0.001
R19281 VN.n883 VN.n882 0.001
R19282 VN.n696 VN.n695 0.001
R19283 VN.n540 VN.n539 0.001
R19284 VN.n1881 VN.n1880 0.001
R19285 VN.n1789 VN.n1788 0.001
R19286 VN.n1635 VN.n1634 0.001
R19287 VN.n1458 VN.n1457 0.001
R19288 VN.n1397 VN.n1396 0.001
R19289 VN.n1222 VN.n1221 0.001
R19290 VN.n1297 VN.n1296 0.001
R19291 VN.n1417 VN.n1416 0.001
R19292 VN.n1091 VN.n1090 0.001
R19293 VN.n732 VN.n731 0.001
R19294 VN.n617 VN.n616 0.001
R19295 VN.n1917 VN.n1916 0.001
R19296 VN.n1805 VN.n1804 0.001
R19297 VN.n408 VN.n407 0.001
R19298 VN.n425 VN.n424 0.001
R19299 VN.n390 VN.n389 0.001
R19300 VN.n1074 VN.n1073 0.001
R19301 VN.n1115 VN.n1114 0.001
R19302 VN.n377 VN.n376 0.001
R19303 VN.n252 VN.n251 0.001
R19304 VN.n266 VN.n265 0.001
R19305 VN.n1829 VN.n1828 0.001
R19306 VN.n1937 VN.n1936 0.001
R19307 VN.n641 VN.n640 0.001
R19308 VN.n775 VN.n774 0.001
R19309 VN.n749 VN.n748 0.001
R19310 VN.n791 VN.n790 0.001
R19311 VN.n324 VN.n323 0.001
R19312 VN.n138 VN.n137 0.001
R19313 VN.n235 VN.n234 0.001
R19314 VN.n1844 VN.n1843 0.001
R19315 VN.n1975 VN.n1974 0.001
R19316 VN.n1948 VN.n1947 0.001
R19317 VN.n1993 VN.n1992 0.001
R19318 VN.n337 VN.n336 0.001
R19319 VN.n116 VN.n115 0.001
R19320 VN.n215 VN.n214 0.001
R19321 VN.n357 VN.n356 0.001
R19322 VN.n33 VN.n32 0.001
R19323 VN.n36 VN.n35 0.001
R19324 VN.n39 VN.n38 0.001
R19325 VN.n1541 VN.n1538 0.001
R19326 VN.n313 VN.n312 0.001
R19327 VN.n159 VN.n158 0.001
R19328 VN.n1868 VN.n1867 0.001
R19329 VN.n660 VN.n659 0.001
R19330 VN.n983 VN.n982 0.001
R19331 VN.n1209 VN.n1208 0.001
R19332 VN.t7 VN.n291 0.001
R19333 VN.t7 VN.n294 0.001
R19334 VN.t42 VN.n486 0.001
R19335 VN.t42 VN.n489 0.001
R19336 VN.t20 VN.n208 0.001
R19337 VN.t20 VN.n205 0.001
R19338 VN.n205 VN.n202 0.001
R19339 VN.n2008 VN.t39 0.001
R19340 VN.n2028 VN.n2010 0.001
R19341 VN.t5 VN.n1696 0.001
R19342 VN.t5 VN.n1699 0.001
R19343 VN.t5 VN.n1668 0.001
R19344 VN.t5 VN.n1665 0.001
R19345 VN.n1665 VN.n1662 0.001
R19346 VN.t11 VN.n1388 0.001
R19347 VN.t11 VN.n1385 0.001
R19348 VN.n1385 VN.n1382 0.001
R19349 VN.t42 VN.n468 0.001
R19350 VN.t42 VN.n465 0.001
R19351 VN.n465 VN.n462 0.001
R19352 VN.t20 VN.n184 0.001
R19353 VN.t20 VN.n181 0.001
R19354 VN.n181 VN.n178 0.001
R19355 VN.t39 VN.n1775 0.001
R19356 VN.t39 VN.n1772 0.001
R19357 VN.n1772 VN.n1769 0.001
R19358 VN.t2 VN.n1911 0.001
R19359 VN.t2 VN.n1908 0.001
R19360 VN.n1908 VN.n1905 0.001
R19361 VN.t17 VN.n586 0.001
R19362 VN.t17 VN.n583 0.001
R19363 VN.n583 VN.n580 0.001
R19364 VN.t13 VN.n726 0.001
R19365 VN.t13 VN.n723 0.001
R19366 VN.n723 VN.n720 0.001
R19367 VN.t37 VN.n929 0.001
R19368 VN.t37 VN.n926 0.001
R19369 VN.n926 VN.n923 0.001
R19370 VN.t22 VN.n1068 0.001
R19371 VN.t22 VN.n1065 0.001
R19372 VN.n1065 VN.n1062 0.001
R19373 VN.t50 VN.n1292 0.001
R19374 VN.t50 VN.n1289 0.001
R19375 VN.n1289 VN.n1286 0.001
R19376 VN.t5 VN.n1505 0.001
R19377 VN.t5 VN.n1502 0.001
R19378 VN.n1502 VN.n1499 0.001
R19379 VN.t11 VN.n1174 0.001
R19380 VN.t11 VN.n1171 0.001
R19381 VN.n1171 VN.n1168 0.001
R19382 VN.t37 VN.n957 0.001
R19383 VN.t37 VN.n960 0.001
R19384 VN.t22 VN.n1009 0.001
R19385 VN.t22 VN.n1006 0.001
R19386 VN.n1006 VN.n1003 0.001
R19387 VN.t50 VN.n1256 0.001
R19388 VN.t50 VN.n1253 0.001
R19389 VN.n1253 VN.n1250 0.001
R19390 VN.n1312 VN.t50 0.001
R19391 VN.n1324 VN.n1315 0.001
R19392 VN.t5 VN.n1625 0.001
R19393 VN.t5 VN.n1622 0.001
R19394 VN.n1622 VN.n1619 0.001
R19395 VN.t17 VN.n610 0.001
R19396 VN.t17 VN.n613 0.001
R19397 VN.t13 VN.n690 0.001
R19398 VN.t13 VN.n687 0.001
R19399 VN.n687 VN.n684 0.001
R19400 VN.t37 VN.n874 0.001
R19401 VN.t37 VN.n871 0.001
R19402 VN.n871 VN.n868 0.001
R19403 VN.t22 VN.n1031 0.001
R19404 VN.t22 VN.n1028 0.001
R19405 VN.n1028 VN.n1025 0.001
R19406 VN.t11 VN.n1343 0.001
R19407 VN.t11 VN.n1340 0.001
R19408 VN.n1340 VN.n1337 0.001
R19409 VN.t50 VN.n1275 0.001
R19410 VN.t50 VN.n1272 0.001
R19411 VN.n1272 VN.n1269 0.001
R19412 VN.t11 VN.n1364 0.001
R19413 VN.t11 VN.n1361 0.001
R19414 VN.n1361 VN.n1358 0.001
R19415 VN.t22 VN.n1050 0.001
R19416 VN.t22 VN.n1047 0.001
R19417 VN.n1047 VN.n1044 0.001
R19418 VN.t37 VN.n895 0.001
R19419 VN.t37 VN.n892 0.001
R19420 VN.n892 VN.n889 0.001
R19421 VN.t13 VN.n709 0.001
R19422 VN.t13 VN.n706 0.001
R19423 VN.n706 VN.n703 0.001
R19424 VN.t17 VN.n552 0.001
R19425 VN.t17 VN.n549 0.001
R19426 VN.n549 VN.n546 0.001
R19427 VN.t2 VN.n1894 0.001
R19428 VN.t2 VN.n1891 0.001
R19429 VN.n1891 VN.n1888 0.001
R19430 VN.t39 VN.n1798 0.001
R19431 VN.t39 VN.n1801 0.001
R19432 VN.t5 VN.n1647 0.001
R19433 VN.t5 VN.n1644 0.001
R19434 VN.n1644 VN.n1641 0.001
R19435 VN.t5 VN.n1469 0.001
R19436 VN.t5 VN.n1466 0.001
R19437 VN.n1466 VN.n1463 0.001
R19438 VN.t11 VN.n1409 0.001
R19439 VN.t11 VN.n1412 0.001
R19440 VN.t50 VN.n1233 0.001
R19441 VN.t50 VN.n1230 0.001
R19442 VN.n1230 VN.n1227 0.001
R19443 VN.n1702 VN.t5 0.001
R19444 VN.n1721 VN.n1704 0.001
R19445 VN.t50 VN.n1306 0.001
R19446 VN.t50 VN.n1309 0.001
R19447 VN.t11 VN.n1426 0.001
R19448 VN.t11 VN.n1429 0.001
R19449 VN.t37 VN.n1104 0.001
R19450 VN.t37 VN.n1107 0.001
R19451 VN.t13 VN.n741 0.001
R19452 VN.t13 VN.n744 0.001
R19453 VN.t17 VN.n630 0.001
R19454 VN.t17 VN.n633 0.001
R19455 VN.t2 VN.n1926 0.001
R19456 VN.t2 VN.n1929 0.001
R19457 VN.t39 VN.n1818 0.001
R19458 VN.t39 VN.n1821 0.001
R19459 VN.n420 VN.n414 0.001
R19460 VN.t42 VN.n438 0.001
R19461 VN.t42 VN.n386 0.001
R19462 VN.n403 VN.n396 0.001
R19463 VN.n402 VN.n401 0.001
R19464 VN.n434 VN.n433 0.001
R19465 VN.n419 VN.n418 0.001
R19466 VN.n1814 VN.n1813 0.001
R19467 VN.n1922 VN.n1921 0.001
R19468 VN.n626 VN.n625 0.001
R19469 VN.n737 VN.n736 0.001
R19470 VN.n1100 VN.n1099 0.001
R19471 VN.n965 VN.n964 0.001
R19472 VN.n1432 VN.t11 0.001
R19473 VN.n1441 VN.n1434 0.001
R19474 VN.t22 VN.n1082 0.001
R19475 VN.t22 VN.n1085 0.001
R19476 VN.t37 VN.n1119 0.001
R19477 VN.t37 VN.n1122 0.001
R19478 VN.n371 VN.t7 0.001
R19479 VN.n378 VN.n371 0.001
R19480 VN.t42 VN.n383 0.001
R19481 VN.n383 VN.n380 0.001
R19482 VN.n267 VN.n260 0.001
R19483 VN.t39 VN.n1833 0.001
R19484 VN.t39 VN.n1836 0.001
R19485 VN.t2 VN.n1942 0.001
R19486 VN.t2 VN.n1945 0.001
R19487 VN.t17 VN.n780 0.001
R19488 VN.t17 VN.n783 0.001
R19489 VN.n769 VN.t13 0.001
R19490 VN.n776 VN.n769 0.001
R19491 VN.n1124 VN.t37 0.001
R19492 VN.n1132 VN.n1124 0.001
R19493 VN.t13 VN.n763 0.001
R19494 VN.t13 VN.n766 0.001
R19495 VN.t17 VN.n795 0.001
R19496 VN.t17 VN.n798 0.001
R19497 VN.t7 VN.n329 0.001
R19498 VN.t7 VN.n332 0.001
R19499 VN.t42 VN.n241 0.001
R19500 VN.t42 VN.n130 0.001
R19501 VN.n229 VN.t20 0.001
R19502 VN.n236 VN.n229 0.001
R19503 VN.t39 VN.n1980 0.001
R19504 VN.t39 VN.n1983 0.001
R19505 VN.n1969 VN.t2 0.001
R19506 VN.n1976 VN.n1969 0.001
R19507 VN.n800 VN.t17 0.001
R19508 VN.n808 VN.n800 0.001
R19509 VN.t2 VN.n1963 0.001
R19510 VN.t2 VN.n1966 0.001
R19511 VN.t39 VN.n2002 0.001
R19512 VN.t39 VN.n2005 0.001
R19513 VN.t7 VN.n345 0.001
R19514 VN.t7 VN.n348 0.001
R19515 VN.t42 VN.n127 0.001
R19516 VN.t42 VN.n124 0.001
R19517 VN.n124 VN.n121 0.001
R19518 VN.t20 VN.n223 0.001
R19519 VN.t20 VN.n226 0.001
R19520 VN.n1527 VN.n1526 0.001
R19521 VN.n1531 VN.n1530 0.001
R19522 VN.n506 VN.n503 0.001
R19523 VN.n1740 VN.n1739 0.001
R19524 VN.n1718 VN.n1709 0.001
R19525 VN.n1142 VN.n1141 0.001
R19526 VN.n838 VN.n837 0.001
R19527 VN.n528 VN.n527 0.001
R19528 VN.n7 VN.n6 0.001
R19529 VN.n40 VN.n28 0.001
R19530 VN.n40 VN.n26 0.001
R19531 VN.n310 VN.n309 0.001
R19532 VN.n291 VN.n288 0.001
R19533 VN.n486 VN.n483 0.001
R19534 VN.n2028 VN.n2008 0.001
R19535 VN.n1798 VN.n1795 0.001
R19536 VN.n610 VN.n607 0.001
R19537 VN.n1324 VN.n1312 0.001
R19538 VN.n957 VN.n954 0.001
R19539 VN.n1409 VN.n1406 0.001
R19540 VN.n1696 VN.n1693 0.001
R19541 VN.n1721 VN.n1702 0.001
R19542 VN.n403 VN.n393 0.001
R19543 VN.n438 VN.n435 0.001
R19544 VN.n420 VN.n411 0.001
R19545 VN.n1818 VN.n1815 0.001
R19546 VN.n1926 VN.n1923 0.001
R19547 VN.n630 VN.n627 0.001
R19548 VN.n741 VN.n738 0.001
R19549 VN.n1104 VN.n1101 0.001
R19550 VN.n1426 VN.n1423 0.001
R19551 VN.n1306 VN.n1303 0.001
R19552 VN.n1441 VN.n1432 0.001
R19553 VN.n378 VN.n374 0.001
R19554 VN.n380 VN.n249 0.001
R19555 VN.n267 VN.n263 0.001
R19556 VN.n1833 VN.n1830 0.001
R19557 VN.n1942 VN.n1939 0.001
R19558 VN.n780 VN.n777 0.001
R19559 VN.n776 VN.n772 0.001
R19560 VN.n1119 VN.n1116 0.001
R19561 VN.n1082 VN.n1079 0.001
R19562 VN.n1132 VN.n1127 0.001
R19563 VN.n763 VN.n760 0.001
R19564 VN.n795 VN.n792 0.001
R19565 VN.n1976 VN.n1972 0.001
R19566 VN.n1980 VN.n1977 0.001
R19567 VN.n236 VN.n232 0.001
R19568 VN.n241 VN.n238 0.001
R19569 VN.n329 VN.n326 0.001
R19570 VN.n808 VN.n803 0.001
R19571 VN.n1963 VN.n1960 0.001
R19572 VN.n2002 VN.n1999 0.001
R19573 VN.n223 VN.n220 0.001
R19574 VN.n345 VN.n342 0.001
R19575 VN.n311 VN.n310 0.001
R19576 VN.t7 VN.n365 0.001
R19577 VN.t7 VN.n368 0.001
R19578 VN.n365 VN.n362 0.001
C0 fc2 out 529.67fF
C1 dw_2450_2450# VN 1715.16fF
C2 fc2 s3 2030.15fF
C3 fc2 s4 638.28fF
C4 s2 out 2148.21fF
C5 VN s4 2044.41fF
C6 VP fc1 1590.25fF
C7 dw_2450_21350# fc2 1760.90fF
C8 out s3 646.54fF
C9 dw_2450_2450# s4 43.87fF
C10 VP s1 6596.21fF
C11 fc2 VN 492.36fF
C12 fc1 s1 2132.03fF
C13 dw_2450_21350# out 734.48fF
C14 fc1 s2 6571.34fF
C15 dw_2450_21350# s3 78.08fF
C16 fc1 out 1693.92fF
C17 dw_2450_2450# fc2 723.90fF
C18 s4 a_400_38200# -247.75fF
C19 s3 a_400_38200# -237.90fF
C20 out a_400_38200# 1439.10fF
C21 s2 a_400_38200# -673.94fF
C22 s1 a_400_38200# -727.12fF
C23 VN a_400_38200# -812.84fF
C24 fc2 a_400_38200# -711.06fF
C25 fc1 a_400_38200# 2811.73fF
C26 VP a_400_38200# 1133.60fF
C27 dw_2450_2450# a_400_38200# 3796.15fF $ **FLOATING
C28 dw_2450_21350# a_400_38200# 3816.34fF $ **FLOATING
C29 VN.n0 a_400_38200# 10.39fF
C30 VN.n1 a_400_38200# 1.88fF
C31 VN.n2 a_400_38200# 17.23fF
C32 VN.n4 a_400_38200# 2.61fF
C33 VN.n5 a_400_38200# 0.84fF
C34 VN.n6 a_400_38200# 0.57fF
C35 VN.n7 a_400_38200# 10.72fF
C36 VN.n8 a_400_38200# 2.57fF
C37 VN.t106 a_400_38200# 0.03fF
C38 VN.n9 a_400_38200# 1.39fF
C39 VN.t62 a_400_38200# 0.03fF
C40 VN.n10 a_400_38200# 0.48fF
C41 VN.n11 a_400_38200# 9.61fF
C42 VN.n12 a_400_38200# 0.03fF
C43 VN.n13 a_400_38200# 0.03fF
C44 VN.n14 a_400_38200# 0.02fF
C45 VN.n15 a_400_38200# 0.05fF
C46 VN.n16 a_400_38200# 0.10fF
C47 VN.n17 a_400_38200# 0.32fF
C48 VN.n18 a_400_38200# 0.68fF
C49 VN.n19 a_400_38200# 0.03fF
C50 VN.n20 a_400_38200# 0.03fF
C51 VN.n21 a_400_38200# 0.03fF
C52 VN.n22 a_400_38200# 0.26fF
C53 VN.n23 a_400_38200# 0.16fF
C54 VN.n24 a_400_38200# 0.19fF
C55 VN.n25 a_400_38200# 1.34fF
C56 VN.n26 a_400_38200# 0.26fF
C57 VN.n27 a_400_38200# 1.34fF
C58 VN.n28 a_400_38200# 0.26fF
C59 VN.n29 a_400_38200# 1.35fF
C60 VN.n30 a_400_38200# 0.25fF
C61 VN.n32 a_400_38200# 1.60fF
C62 VN.n33 a_400_38200# 0.43fF
C63 VN.n35 a_400_38200# 1.60fF
C64 VN.n36 a_400_38200# 0.43fF
C65 VN.n38 a_400_38200# 1.83fF
C66 VN.n39 a_400_38200# 0.43fF
C67 VN.n40 a_400_38200# 68.86fF
C68 VN.n41 a_400_38200# 5.11fF
C69 VN.t167 a_400_38200# 0.03fF
C70 VN.n42 a_400_38200# 0.98fF
C71 VN.t232 a_400_38200# 0.03fF
C72 VN.n43 a_400_38200# 0.02fF
C73 VN.n44 a_400_38200# 0.40fF
C74 VN.t70 a_400_38200# 0.02fF
C75 VN.n45 a_400_38200# 0.97fF
C76 VN.n46 a_400_38200# 1.01fF
C77 VN.n47 a_400_38200# 4.45fF
C78 VN.n48 a_400_38200# 2.02fF
C79 VN.t274 a_400_38200# 0.02fF
C80 VN.n49 a_400_38200# 0.97fF
C81 VN.t377 a_400_38200# 0.03fF
C82 VN.n50 a_400_38200# 0.98fF
C83 VN.n51 a_400_38200# 2.32fF
C84 VN.n52 a_400_38200# 1.30fF
C85 VN.n53 a_400_38200# 0.36fF
C86 VN.n54 a_400_38200# 0.34fF
C87 VN.t177 a_400_38200# 0.03fF
C88 VN.n55 a_400_38200# 0.02fF
C89 VN.n56 a_400_38200# 0.40fF
C90 VN.n57 a_400_38200# 0.23fF
C91 VN.n58 a_400_38200# 2.39fF
C92 VN.n59 a_400_38200# 1.39fF
C93 VN.n60 a_400_38200# 0.34fF
C94 VN.t254 a_400_38200# 0.03fF
C95 VN.n61 a_400_38200# 0.98fF
C96 VN.t149 a_400_38200# 0.02fF
C97 VN.n62 a_400_38200# 0.97fF
C98 VN.n63 a_400_38200# 4.20fF
C99 VN.n64 a_400_38200# 3.05fF
C100 VN.t68 a_400_38200# 0.03fF
C101 VN.n65 a_400_38200# 0.02fF
C102 VN.n66 a_400_38200# 0.40fF
C103 VN.n67 a_400_38200# 2.65fF
C104 VN.t127 a_400_38200# 0.03fF
C105 VN.n68 a_400_38200# 0.98fF
C106 VN.t86 a_400_38200# 0.02fF
C107 VN.n69 a_400_38200# 0.97fF
C108 VN.n70 a_400_38200# 1.05fF
C109 VN.n71 a_400_38200# 3.93fF
C110 VN.n72 a_400_38200# 3.05fF
C111 VN.t244 a_400_38200# 0.03fF
C112 VN.n73 a_400_38200# 0.02fF
C113 VN.n74 a_400_38200# 0.40fF
C114 VN.n75 a_400_38200# 1.05fF
C115 VN.n76 a_400_38200# 3.93fF
C116 VN.n77 a_400_38200# 3.06fF
C117 VN.t328 a_400_38200# 0.02fF
C118 VN.n78 a_400_38200# 0.97fF
C119 VN.t53 a_400_38200# 0.03fF
C120 VN.n79 a_400_38200# 0.98fF
C121 VN.n80 a_400_38200# 2.65fF
C122 VN.t116 a_400_38200# 0.03fF
C123 VN.n81 a_400_38200# 0.02fF
C124 VN.n82 a_400_38200# 0.40fF
C125 VN.n83 a_400_38200# 4.31fF
C126 VN.n84 a_400_38200# 3.03fF
C127 VN.n85 a_400_38200# 0.03fF
C128 VN.n86 a_400_38200# 0.03fF
C129 VN.n87 a_400_38200# 0.03fF
C130 VN.n88 a_400_38200# 0.03fF
C131 VN.n89 a_400_38200# 0.03fF
C132 VN.n90 a_400_38200# 0.02fF
C133 VN.n91 a_400_38200# 0.05fF
C134 VN.n92 a_400_38200# 0.10fF
C135 VN.n93 a_400_38200# 0.32fF
C136 VN.n94 a_400_38200# 0.68fF
C137 VN.n95 a_400_38200# 0.26fF
C138 VN.n96 a_400_38200# 0.16fF
C139 VN.n97 a_400_38200# 0.19fF
C140 VN.t203 a_400_38200# 0.02fF
C141 VN.n98 a_400_38200# 0.97fF
C142 VN.t297 a_400_38200# 0.03fF
C143 VN.n99 a_400_38200# 0.98fF
C144 VN.t354 a_400_38200# 0.03fF
C145 VN.n100 a_400_38200# 0.02fF
C146 VN.n101 a_400_38200# 0.40fF
C147 VN.t52 a_400_38200# 70.80fF
C148 VN.n102 a_400_38200# 0.51fF
C149 VN.n103 a_400_38200# 4.84fF
C150 VN.n104 a_400_38200# 2.57fF
C151 VN.n105 a_400_38200# 5.82fF
C152 VN.t240 a_400_38200# 0.02fF
C153 VN.n106 a_400_38200# 1.33fF
C154 VN.n107 a_400_38200# 0.13fF
C155 VN.n108 a_400_38200# 0.13fF
C156 VN.n109 a_400_38200# 0.12fF
C157 VN.n110 a_400_38200# 0.39fF
C158 VN.n111 a_400_38200# 0.51fF
C159 VN.n112 a_400_38200# 1.24fF
C160 VN.n113 a_400_38200# 2.05fF
C161 VN.n114 a_400_38200# 0.13fF
C162 VN.t323 a_400_38200# 0.02fF
C163 VN.n115 a_400_38200# 0.15fF
C164 VN.t125 a_400_38200# 0.02fF
C165 VN.n117 a_400_38200# 0.26fF
C166 VN.n118 a_400_38200# 0.39fF
C167 VN.n119 a_400_38200# 0.66fF
C168 VN.n120 a_400_38200# 2.91fF
C169 VN.n121 a_400_38200# 4.29fF
C170 VN.t351 a_400_38200# 0.03fF
C171 VN.n122 a_400_38200# 0.26fF
C172 VN.n123 a_400_38200# 1.00fF
C173 VN.n124 a_400_38200# 0.05fF
C174 VN.t44 a_400_38200# 0.03fF
C175 VN.n125 a_400_38200# 0.13fF
C176 VN.n126 a_400_38200# 0.16fF
C177 VN.t114 a_400_38200# 0.03fF
C178 VN.n128 a_400_38200# 0.26fF
C179 VN.n129 a_400_38200# 1.00fF
C180 VN.n130 a_400_38200# 0.05fF
C181 VN.n131 a_400_38200# 2.05fF
C182 VN.n132 a_400_38200# 2.91fF
C183 VN.t251 a_400_38200# 0.02fF
C184 VN.n133 a_400_38200# 0.26fF
C185 VN.n134 a_400_38200# 0.39fF
C186 VN.n135 a_400_38200# 0.66fF
C187 VN.n136 a_400_38200# 0.13fF
C188 VN.t80 a_400_38200# 0.02fF
C189 VN.n137 a_400_38200# 0.15fF
C190 VN.n139 a_400_38200# 2.05fF
C191 VN.n140 a_400_38200# 2.91fF
C192 VN.t82 a_400_38200# 0.02fF
C193 VN.n141 a_400_38200# 0.26fF
C194 VN.n142 a_400_38200# 0.39fF
C195 VN.n143 a_400_38200# 0.66fF
C196 VN.t381 a_400_38200# 0.02fF
C197 VN.n144 a_400_38200# 1.33fF
C198 VN.n145 a_400_38200# 0.07fF
C199 VN.n146 a_400_38200# 0.11fF
C200 VN.n147 a_400_38200# 0.66fF
C201 VN.n148 a_400_38200# 0.39fF
C202 VN.n149 a_400_38200# 0.69fF
C203 VN.n150 a_400_38200# 1.26fF
C204 VN.n151 a_400_38200# 1.65fF
C205 VN.n152 a_400_38200# 0.65fF
C206 VN.n153 a_400_38200# 0.02fF
C207 VN.n154 a_400_38200# 1.06fF
C208 VN.t81 a_400_38200# 9.89fF
C209 VN.n155 a_400_38200# 10.65fF
C210 VN.n157 a_400_38200# 0.41fF
C211 VN.n158 a_400_38200# 0.25fF
C212 VN.n159 a_400_38200# 3.16fF
C213 VN.n160 a_400_38200# 2.64fF
C214 VN.n161 a_400_38200# 2.70fF
C215 VN.n162 a_400_38200# 4.68fF
C216 VN.n163 a_400_38200# 0.27fF
C217 VN.n164 a_400_38200# 0.01fF
C218 VN.t218 a_400_38200# 0.02fF
C219 VN.n165 a_400_38200# 0.28fF
C220 VN.t261 a_400_38200# 0.03fF
C221 VN.n166 a_400_38200# 1.04fF
C222 VN.n167 a_400_38200# 0.77fF
C223 VN.n168 a_400_38200# 2.06fF
C224 VN.n169 a_400_38200# 2.05fF
C225 VN.t257 a_400_38200# 0.02fF
C226 VN.n170 a_400_38200# 0.26fF
C227 VN.n171 a_400_38200# 0.39fF
C228 VN.n172 a_400_38200# 0.66fF
C229 VN.n173 a_400_38200# 0.13fF
C230 VN.t90 a_400_38200# 0.02fF
C231 VN.n174 a_400_38200# 0.15fF
C232 VN.n176 a_400_38200# 1.26fF
C233 VN.n177 a_400_38200# 0.24fF
C234 VN.n178 a_400_38200# 2.06fF
C235 VN.t136 a_400_38200# 0.03fF
C236 VN.n179 a_400_38200# 0.26fF
C237 VN.n180 a_400_38200# 1.00fF
C238 VN.n181 a_400_38200# 0.05fF
C239 VN.t119 a_400_38200# 0.03fF
C240 VN.n182 a_400_38200# 0.13fF
C241 VN.n183 a_400_38200# 0.16fF
C242 VN.n185 a_400_38200# 0.84fF
C243 VN.n186 a_400_38200# 0.48fF
C244 VN.n187 a_400_38200# 1.72fF
C245 VN.n188 a_400_38200# 0.13fF
C246 VN.t36 a_400_38200# 0.02fF
C247 VN.n189 a_400_38200# 0.15fF
C248 VN.t198 a_400_38200# 0.02fF
C249 VN.n191 a_400_38200# 0.26fF
C250 VN.n192 a_400_38200# 0.39fF
C251 VN.n193 a_400_38200# 0.66fF
C252 VN.n194 a_400_38200# 0.01fF
C253 VN.n195 a_400_38200# 0.07fF
C254 VN.n196 a_400_38200# 0.01fF
C255 VN.n197 a_400_38200# 0.02fF
C256 VN.n198 a_400_38200# 0.02fF
C257 VN.n199 a_400_38200# 0.26fF
C258 VN.n200 a_400_38200# 1.26fF
C259 VN.n201 a_400_38200# 1.46fF
C260 VN.n202 a_400_38200# 2.17fF
C261 VN.t95 a_400_38200# 0.03fF
C262 VN.n203 a_400_38200# 0.26fF
C263 VN.n204 a_400_38200# 1.00fF
C264 VN.n205 a_400_38200# 0.05fF
C265 VN.t54 a_400_38200# 0.03fF
C266 VN.n206 a_400_38200# 0.13fF
C267 VN.n207 a_400_38200# 0.16fF
C268 VN.n209 a_400_38200# 9.61fF
C269 VN.n210 a_400_38200# 0.10fF
C270 VN.n211 a_400_38200# 0.20fF
C271 VN.n212 a_400_38200# 2.05fF
C272 VN.n213 a_400_38200# 0.13fF
C273 VN.t152 a_400_38200# 0.02fF
C274 VN.n214 a_400_38200# 0.15fF
C275 VN.t324 a_400_38200# 0.02fF
C276 VN.n216 a_400_38200# 0.26fF
C277 VN.n217 a_400_38200# 0.39fF
C278 VN.n218 a_400_38200# 0.66fF
C279 VN.n219 a_400_38200# 2.90fF
C280 VN.n220 a_400_38200# 3.58fF
C281 VN.t184 a_400_38200# 0.03fF
C282 VN.n221 a_400_38200# 0.13fF
C283 VN.n222 a_400_38200# 0.16fF
C284 VN.t221 a_400_38200# 0.03fF
C285 VN.n224 a_400_38200# 0.26fF
C286 VN.n225 a_400_38200# 1.00fF
C287 VN.n226 a_400_38200# 0.05fF
C288 VN.t20 a_400_38200# 21.51fF
C289 VN.t342 a_400_38200# 0.03fF
C290 VN.n227 a_400_38200# 0.26fF
C291 VN.n228 a_400_38200# 1.00fF
C292 VN.n229 a_400_38200# 0.05fF
C293 VN.t311 a_400_38200# 0.03fF
C294 VN.n230 a_400_38200# 0.13fF
C295 VN.n231 a_400_38200# 0.16fF
C296 VN.n233 a_400_38200# 0.13fF
C297 VN.t277 a_400_38200# 0.02fF
C298 VN.n234 a_400_38200# 0.15fF
C299 VN.n236 a_400_38200# 2.51fF
C300 VN.n237 a_400_38200# 3.06fF
C301 VN.n238 a_400_38200# 5.64fF
C302 VN.t178 a_400_38200# 0.03fF
C303 VN.n239 a_400_38200# 0.13fF
C304 VN.n240 a_400_38200# 0.16fF
C305 VN.n242 a_400_38200# 2.05fF
C306 VN.n243 a_400_38200# 2.91fF
C307 VN.t375 a_400_38200# 0.02fF
C308 VN.n244 a_400_38200# 0.26fF
C309 VN.n245 a_400_38200# 0.39fF
C310 VN.n246 a_400_38200# 0.66fF
C311 VN.t159 a_400_38200# 0.03fF
C312 VN.n247 a_400_38200# 0.13fF
C313 VN.n248 a_400_38200# 0.16fF
C314 VN.n250 a_400_38200# 0.13fF
C315 VN.t211 a_400_38200# 0.02fF
C316 VN.n251 a_400_38200# 0.15fF
C317 VN.n253 a_400_38200# 2.05fF
C318 VN.n254 a_400_38200# 2.91fF
C319 VN.t212 a_400_38200# 0.02fF
C320 VN.n255 a_400_38200# 0.26fF
C321 VN.n256 a_400_38200# 0.39fF
C322 VN.n257 a_400_38200# 0.66fF
C323 VN.t108 a_400_38200# 0.03fF
C324 VN.n258 a_400_38200# 0.26fF
C325 VN.n259 a_400_38200# 1.00fF
C326 VN.n260 a_400_38200# 0.05fF
C327 VN.t66 a_400_38200# 0.03fF
C328 VN.n261 a_400_38200# 0.13fF
C329 VN.n262 a_400_38200# 0.16fF
C330 VN.n264 a_400_38200# 0.13fF
C331 VN.t21 a_400_38200# 0.02fF
C332 VN.n265 a_400_38200# 0.15fF
C333 VN.n267 a_400_38200# 2.51fF
C334 VN.n268 a_400_38200# 3.21fF
C335 VN.n269 a_400_38200# 2.12fF
C336 VN.n270 a_400_38200# 2.77fF
C337 VN.t27 a_400_38200# 0.02fF
C338 VN.n271 a_400_38200# 0.26fF
C339 VN.n272 a_400_38200# 0.39fF
C340 VN.n273 a_400_38200# 0.66fF
C341 VN.n274 a_400_38200# 9.61fF
C342 VN.n275 a_400_38200# 0.28fF
C343 VN.n276 a_400_38200# 0.13fF
C344 VN.n277 a_400_38200# 0.06fF
C345 VN.n278 a_400_38200# 0.19fF
C346 VN.n279 a_400_38200# 1.37fF
C347 VN.n280 a_400_38200# 3.02fF
C348 VN.n281 a_400_38200# 0.13fF
C349 VN.t8 a_400_38200# 0.02fF
C350 VN.n282 a_400_38200# 0.15fF
C351 VN.t327 a_400_38200# 0.02fF
C352 VN.n284 a_400_38200# 0.26fF
C353 VN.n285 a_400_38200# 0.39fF
C354 VN.n286 a_400_38200# 0.66fF
C355 VN.n287 a_400_38200# 2.85fF
C356 VN.n288 a_400_38200# 2.24fF
C357 VN.t58 a_400_38200# 0.03fF
C358 VN.n289 a_400_38200# 0.13fF
C359 VN.n290 a_400_38200# 0.16fF
C360 VN.t97 a_400_38200# 0.03fF
C361 VN.n292 a_400_38200# 0.26fF
C362 VN.n293 a_400_38200# 1.00fF
C363 VN.n294 a_400_38200# 0.05fF
C364 VN.t220 a_400_38200# 0.03fF
C365 VN.n295 a_400_38200# 1.04fF
C366 VN.n296 a_400_38200# 0.77fF
C367 VN.n297 a_400_38200# 0.01fF
C368 VN.t168 a_400_38200# 0.02fF
C369 VN.n298 a_400_38200# 0.28fF
C370 VN.t295 a_400_38200# 0.02fF
C371 VN.n299 a_400_38200# 1.33fF
C372 VN.n300 a_400_38200# 2.14fF
C373 VN.n301 a_400_38200# 0.07fF
C374 VN.n302 a_400_38200# 0.11fF
C375 VN.n303 a_400_38200# 0.66fF
C376 VN.n304 a_400_38200# 1.65fF
C377 VN.n305 a_400_38200# 1.01fF
C378 VN.n306 a_400_38200# 0.92fF
C379 VN.n307 a_400_38200# 0.02fF
C380 VN.n308 a_400_38200# 1.06fF
C381 VN.t26 a_400_38200# 9.89fF
C382 VN.n309 a_400_38200# 10.32fF
C383 VN.n311 a_400_38200# 1.33fF
C384 VN.n312 a_400_38200# 1.58fF
C385 VN.n313 a_400_38200# 3.16fF
C386 VN.n314 a_400_38200# 2.64fF
C387 VN.n315 a_400_38200# 4.20fF
C388 VN.n316 a_400_38200# 0.27fF
C389 VN.n317 a_400_38200# 2.12fF
C390 VN.n318 a_400_38200# 2.77fF
C391 VN.t216 a_400_38200# 0.02fF
C392 VN.n319 a_400_38200# 0.26fF
C393 VN.n320 a_400_38200# 0.39fF
C394 VN.n321 a_400_38200# 0.66fF
C395 VN.n322 a_400_38200# 0.13fF
C396 VN.t279 a_400_38200# 0.02fF
C397 VN.n323 a_400_38200# 0.15fF
C398 VN.n325 a_400_38200# 2.63fF
C399 VN.n326 a_400_38200# 2.51fF
C400 VN.t314 a_400_38200# 0.03fF
C401 VN.n327 a_400_38200# 0.13fF
C402 VN.n328 a_400_38200# 0.16fF
C403 VN.t345 a_400_38200# 0.03fF
C404 VN.n330 a_400_38200# 0.26fF
C405 VN.n331 a_400_38200# 1.00fF
C406 VN.n332 a_400_38200# 0.05fF
C407 VN.n333 a_400_38200# 2.63fF
C408 VN.n334 a_400_38200# 2.16fF
C409 VN.n335 a_400_38200# 0.13fF
C410 VN.t155 a_400_38200# 0.02fF
C411 VN.n336 a_400_38200# 0.15fF
C412 VN.t85 a_400_38200# 0.02fF
C413 VN.n338 a_400_38200# 0.26fF
C414 VN.n339 a_400_38200# 0.39fF
C415 VN.n340 a_400_38200# 0.66fF
C416 VN.n341 a_400_38200# 2.78fF
C417 VN.n342 a_400_38200# 2.52fF
C418 VN.t190 a_400_38200# 0.03fF
C419 VN.n343 a_400_38200# 0.13fF
C420 VN.n344 a_400_38200# 0.16fF
C421 VN.t222 a_400_38200# 0.03fF
C422 VN.n346 a_400_38200# 0.26fF
C423 VN.n347 a_400_38200# 1.00fF
C424 VN.n348 a_400_38200# 0.05fF
C425 VN.n349 a_400_38200# 0.28fF
C426 VN.n350 a_400_38200# 0.13fF
C427 VN.n351 a_400_38200# 0.06fF
C428 VN.n352 a_400_38200# 0.19fF
C429 VN.n353 a_400_38200# 1.25fF
C430 VN.n354 a_400_38200# 2.04fF
C431 VN.n355 a_400_38200# 0.13fF
C432 VN.t288 a_400_38200# 0.02fF
C433 VN.n356 a_400_38200# 0.15fF
C434 VN.t201 a_400_38200# 0.02fF
C435 VN.n358 a_400_38200# 0.26fF
C436 VN.n359 a_400_38200# 0.39fF
C437 VN.n360 a_400_38200# 0.66fF
C438 VN.n361 a_400_38200# 2.78fF
C439 VN.n362 a_400_38200# 2.12fF
C440 VN.t301 a_400_38200# 0.03fF
C441 VN.n363 a_400_38200# 0.13fF
C442 VN.n364 a_400_38200# 0.16fF
C443 VN.t336 a_400_38200# 0.03fF
C444 VN.n366 a_400_38200# 0.26fF
C445 VN.n367 a_400_38200# 1.00fF
C446 VN.n368 a_400_38200# 0.05fF
C447 VN.t7 a_400_38200# 21.51fF
C448 VN.t332 a_400_38200# 0.03fF
C449 VN.n369 a_400_38200# 0.26fF
C450 VN.n370 a_400_38200# 1.00fF
C451 VN.n371 a_400_38200# 0.05fF
C452 VN.t315 a_400_38200# 0.03fF
C453 VN.n372 a_400_38200# 0.13fF
C454 VN.n373 a_400_38200# 0.16fF
C455 VN.n375 a_400_38200# 0.13fF
C456 VN.t280 a_400_38200# 0.02fF
C457 VN.n376 a_400_38200# 0.15fF
C458 VN.n378 a_400_38200# 2.51fF
C459 VN.n379 a_400_38200# 1.93fF
C460 VN.n380 a_400_38200# 5.63fF
C461 VN.t241 a_400_38200# 0.03fF
C462 VN.n381 a_400_38200# 0.26fF
C463 VN.n382 a_400_38200# 1.00fF
C464 VN.n383 a_400_38200# 0.05fF
C465 VN.t151 a_400_38200# 0.03fF
C466 VN.n384 a_400_38200# 0.26fF
C467 VN.n385 a_400_38200# 1.00fF
C468 VN.n386 a_400_38200# 0.05fF
C469 VN.n387 a_400_38200# 2.12fF
C470 VN.n388 a_400_38200# 0.13fF
C471 VN.t29 a_400_38200# 0.02fF
C472 VN.n389 a_400_38200# 0.15fF
C473 VN.t71 a_400_38200# 0.03fF
C474 VN.n391 a_400_38200# 0.13fF
C475 VN.n392 a_400_38200# 0.16fF
C476 VN.t94 a_400_38200# 0.03fF
C477 VN.n394 a_400_38200# 0.26fF
C478 VN.n395 a_400_38200# 1.00fF
C479 VN.n396 a_400_38200# 0.05fF
C480 VN.t164 a_400_38200# 0.02fF
C481 VN.n397 a_400_38200# 0.26fF
C482 VN.n398 a_400_38200# 0.39fF
C483 VN.n399 a_400_38200# 0.66fF
C484 VN.n400 a_400_38200# 0.33fF
C485 VN.n401 a_400_38200# 1.19fF
C486 VN.n402 a_400_38200# 0.17fF
C487 VN.n403 a_400_38200# 2.29fF
C488 VN.n404 a_400_38200# 1.95fF
C489 VN.n405 a_400_38200# 2.05fF
C490 VN.n406 a_400_38200# 0.13fF
C491 VN.t331 a_400_38200# 0.02fF
C492 VN.n407 a_400_38200# 0.15fF
C493 VN.t356 a_400_38200# 0.03fF
C494 VN.n409 a_400_38200# 0.13fF
C495 VN.n410 a_400_38200# 0.16fF
C496 VN.t371 a_400_38200# 0.03fF
C497 VN.n412 a_400_38200# 0.26fF
C498 VN.n413 a_400_38200# 1.00fF
C499 VN.n414 a_400_38200# 0.05fF
C500 VN.t129 a_400_38200# 0.02fF
C501 VN.n415 a_400_38200# 0.26fF
C502 VN.n416 a_400_38200# 0.39fF
C503 VN.n417 a_400_38200# 0.66fF
C504 VN.n418 a_400_38200# 1.19fF
C505 VN.n419 a_400_38200# 0.17fF
C506 VN.n420 a_400_38200# 2.29fF
C507 VN.n421 a_400_38200# 3.21fF
C508 VN.n422 a_400_38200# 2.05fF
C509 VN.n423 a_400_38200# 0.13fF
C510 VN.t194 a_400_38200# 0.02fF
C511 VN.n424 a_400_38200# 0.15fF
C512 VN.t359 a_400_38200# 0.02fF
C513 VN.n426 a_400_38200# 0.26fF
C514 VN.n427 a_400_38200# 0.39fF
C515 VN.n428 a_400_38200# 0.66fF
C516 VN.n429 a_400_38200# 1.01fF
C517 VN.n430 a_400_38200# 0.35fF
C518 VN.n431 a_400_38200# 0.35fF
C519 VN.n432 a_400_38200# 1.01fF
C520 VN.n433 a_400_38200# 1.19fF
C521 VN.n434 a_400_38200# 0.17fF
C522 VN.n435 a_400_38200# 5.41fF
C523 VN.t287 a_400_38200# 0.03fF
C524 VN.n436 a_400_38200# 0.13fF
C525 VN.n437 a_400_38200# 0.16fF
C526 VN.t102 a_400_38200# 0.03fF
C527 VN.n439 a_400_38200# 1.04fF
C528 VN.n440 a_400_38200# 0.77fF
C529 VN.n441 a_400_38200# 1.92fF
C530 VN.n442 a_400_38200# 3.32fF
C531 VN.t105 a_400_38200# 0.02fF
C532 VN.n443 a_400_38200# 0.26fF
C533 VN.n444 a_400_38200# 0.39fF
C534 VN.n445 a_400_38200# 0.66fF
C535 VN.n446 a_400_38200# 0.13fF
C536 VN.t322 a_400_38200# 0.02fF
C537 VN.n447 a_400_38200# 0.15fF
C538 VN.n449 a_400_38200# 0.20fF
C539 VN.n450 a_400_38200# 0.22fF
C540 VN.n451 a_400_38200# 0.28fF
C541 VN.n452 a_400_38200# 0.10fF
C542 VN.n453 a_400_38200# 0.25fF
C543 VN.n454 a_400_38200# 0.72fF
C544 VN.n455 a_400_38200# 0.99fF
C545 VN.n456 a_400_38200# 0.25fF
C546 VN.n457 a_400_38200# 0.10fF
C547 VN.n458 a_400_38200# 0.23fF
C548 VN.n459 a_400_38200# 0.07fF
C549 VN.n460 a_400_38200# 0.06fF
C550 VN.n461 a_400_38200# 0.07fF
C551 VN.n462 a_400_38200# 2.17fF
C552 VN.t266 a_400_38200# 0.03fF
C553 VN.n463 a_400_38200# 0.26fF
C554 VN.n464 a_400_38200# 1.00fF
C555 VN.n465 a_400_38200# 0.05fF
C556 VN.t43 a_400_38200# 0.03fF
C557 VN.n466 a_400_38200# 0.13fF
C558 VN.n467 a_400_38200# 0.16fF
C559 VN.n469 a_400_38200# 9.61fF
C560 VN.n470 a_400_38200# 0.27fF
C561 VN.n471 a_400_38200# 0.10fF
C562 VN.n472 a_400_38200# 0.22fF
C563 VN.n473 a_400_38200# 0.85fF
C564 VN.n474 a_400_38200# 2.11fF
C565 VN.n475 a_400_38200# 2.05fF
C566 VN.n476 a_400_38200# 0.13fF
C567 VN.t196 a_400_38200# 0.02fF
C568 VN.n477 a_400_38200# 0.15fF
C569 VN.t363 a_400_38200# 0.02fF
C570 VN.n479 a_400_38200# 0.26fF
C571 VN.n480 a_400_38200# 0.39fF
C572 VN.n481 a_400_38200# 0.66fF
C573 VN.n482 a_400_38200# 2.91fF
C574 VN.n483 a_400_38200# 3.27fF
C575 VN.t290 a_400_38200# 0.03fF
C576 VN.n484 a_400_38200# 0.13fF
C577 VN.n485 a_400_38200# 0.16fF
C578 VN.t228 a_400_38200# 0.03fF
C579 VN.n487 a_400_38200# 0.26fF
C580 VN.n488 a_400_38200# 1.00fF
C581 VN.n489 a_400_38200# 0.05fF
C582 VN.t188 a_400_38200# 0.03fF
C583 VN.n490 a_400_38200# 0.01fF
C584 VN.n491 a_400_38200# 0.28fF
C585 VN.t42 a_400_38200# 21.51fF
C586 VN.n492 a_400_38200# 0.27fF
C587 VN.n493 a_400_38200# 3.18fF
C588 VN.n494 a_400_38200# 30.53fF
C589 VN.n495 a_400_38200# 44.05fF
C590 VN.n496 a_400_38200# 0.65fF
C591 VN.n497 a_400_38200# 0.48fF
C592 VN.n498 a_400_38200# 0.65fF
C593 VN.n499 a_400_38200# 2.08fF
C594 VN.n500 a_400_38200# 0.31fF
C595 VN.t93 a_400_38200# 9.89fF
C596 VN.n501 a_400_38200# 12.19fF
C597 VN.n502 a_400_38200# 0.84fF
C598 VN.n503 a_400_38200# 0.30fF
C599 VN.n504 a_400_38200# 30.53fF
C600 VN.n505 a_400_38200# 44.05fF
C601 VN.n506 a_400_38200# 4.91fF
C602 VN.n507 a_400_38200# 2.54fF
C603 VN.n508 a_400_38200# 4.99fF
C604 VN.n509 a_400_38200# 0.02fF
C605 VN.n510 a_400_38200# 0.03fF
C606 VN.n511 a_400_38200# 0.26fF
C607 VN.n512 a_400_38200# 0.14fF
C608 VN.n513 a_400_38200# 0.61fF
C609 VN.n514 a_400_38200# 0.03fF
C610 VN.n515 a_400_38200# 0.94fF
C611 VN.n516 a_400_38200# 0.24fF
C612 VN.n517 a_400_38200# 0.16fF
C613 VN.n518 a_400_38200# 30.53fF
C614 VN.n519 a_400_38200# 30.53fF
C615 VN.n520 a_400_38200# 0.65fF
C616 VN.n521 a_400_38200# 0.24fF
C617 VN.n522 a_400_38200# 0.65fF
C618 VN.n523 a_400_38200# 2.08fF
C619 VN.n524 a_400_38200# 0.31fF
C620 VN.t33 a_400_38200# 9.89fF
C621 VN.n525 a_400_38200# 12.19fF
C622 VN.n526 a_400_38200# 0.84fF
C623 VN.n527 a_400_38200# 0.30fF
C624 VN.n528 a_400_38200# 4.37fF
C625 VN.n529 a_400_38200# 1.24fF
C626 VN.t118 a_400_38200# 0.02fF
C627 VN.n530 a_400_38200# 0.70fF
C628 VN.n531 a_400_38200# 0.66fF
C629 VN.n532 a_400_38200# 0.27fF
C630 VN.n533 a_400_38200# 0.10fF
C631 VN.n534 a_400_38200# 0.23fF
C632 VN.n535 a_400_38200# 1.40fF
C633 VN.n536 a_400_38200# 0.58fF
C634 VN.n537 a_400_38200# 2.05fF
C635 VN.n538 a_400_38200# 0.13fF
C636 VN.t273 a_400_38200# 0.02fF
C637 VN.n539 a_400_38200# 0.15fF
C638 VN.t76 a_400_38200# 0.02fF
C639 VN.n541 a_400_38200# 0.26fF
C640 VN.n542 a_400_38200# 0.39fF
C641 VN.n543 a_400_38200# 0.66fF
C642 VN.n544 a_400_38200# 0.78fF
C643 VN.n545 a_400_38200# 1.72fF
C644 VN.n546 a_400_38200# 2.67fF
C645 VN.t243 a_400_38200# 0.03fF
C646 VN.n547 a_400_38200# 0.26fF
C647 VN.n548 a_400_38200# 1.00fF
C648 VN.n549 a_400_38200# 0.05fF
C649 VN.t374 a_400_38200# 0.03fF
C650 VN.n550 a_400_38200# 0.13fF
C651 VN.n551 a_400_38200# 0.16fF
C652 VN.n553 a_400_38200# 2.06fF
C653 VN.n554 a_400_38200# 0.06fF
C654 VN.n555 a_400_38200# 0.03fF
C655 VN.n556 a_400_38200# 0.04fF
C656 VN.n557 a_400_38200# 1.08fF
C657 VN.n558 a_400_38200# 0.02fF
C658 VN.n559 a_400_38200# 0.01fF
C659 VN.n560 a_400_38200# 0.02fF
C660 VN.n561 a_400_38200# 0.09fF
C661 VN.n562 a_400_38200# 0.39fF
C662 VN.n563 a_400_38200# 2.02fF
C663 VN.t258 a_400_38200# 0.02fF
C664 VN.n564 a_400_38200# 0.26fF
C665 VN.n565 a_400_38200# 0.39fF
C666 VN.n566 a_400_38200# 0.66fF
C667 VN.n567 a_400_38200# 0.13fF
C668 VN.t87 a_400_38200# 0.02fF
C669 VN.n568 a_400_38200# 0.15fF
C670 VN.n570 a_400_38200# 0.76fF
C671 VN.n571 a_400_38200# 0.25fF
C672 VN.n572 a_400_38200# 0.28fF
C673 VN.n573 a_400_38200# 0.10fF
C674 VN.n574 a_400_38200# 0.25fF
C675 VN.n575 a_400_38200# 0.76fF
C676 VN.n576 a_400_38200# 1.26fF
C677 VN.n577 a_400_38200# 0.24fF
C678 VN.n578 a_400_38200# 0.28fF
C679 VN.n579 a_400_38200# 0.10fF
C680 VN.n580 a_400_38200# 2.06fF
C681 VN.t117 a_400_38200# 0.03fF
C682 VN.n581 a_400_38200# 0.26fF
C683 VN.n582 a_400_38200# 1.00fF
C684 VN.n583 a_400_38200# 0.05fF
C685 VN.t250 a_400_38200# 0.03fF
C686 VN.n584 a_400_38200# 0.13fF
C687 VN.n585 a_400_38200# 0.16fF
C688 VN.n587 a_400_38200# 9.61fF
C689 VN.n588 a_400_38200# 2.60fF
C690 VN.n589 a_400_38200# 0.50fF
C691 VN.n590 a_400_38200# 0.24fF
C692 VN.n591 a_400_38200# 0.41fF
C693 VN.n592 a_400_38200# 0.17fF
C694 VN.n593 a_400_38200# 0.31fF
C695 VN.n594 a_400_38200# 0.23fF
C696 VN.n595 a_400_38200# 0.33fF
C697 VN.n596 a_400_38200# 0.22fF
C698 VN.t183 a_400_38200# 0.02fF
C699 VN.n597 a_400_38200# 0.26fF
C700 VN.n598 a_400_38200# 0.39fF
C701 VN.n599 a_400_38200# 0.66fF
C702 VN.n600 a_400_38200# 0.13fF
C703 VN.t18 a_400_38200# 0.02fF
C704 VN.n601 a_400_38200# 0.15fF
C705 VN.n603 a_400_38200# 0.21fF
C706 VN.n604 a_400_38200# 1.72fF
C707 VN.n605 a_400_38200# 2.41fF
C708 VN.n606 a_400_38200# 0.35fF
C709 VN.n607 a_400_38200# 2.61fF
C710 VN.t138 a_400_38200# 0.03fF
C711 VN.n608 a_400_38200# 0.13fF
C712 VN.n609 a_400_38200# 0.16fF
C713 VN.t344 a_400_38200# 0.03fF
C714 VN.n611 a_400_38200# 0.26fF
C715 VN.n612 a_400_38200# 1.00fF
C716 VN.n613 a_400_38200# 0.05fF
C717 VN.n614 a_400_38200# 2.05fF
C718 VN.n615 a_400_38200# 0.13fF
C719 VN.t329 a_400_38200# 0.02fF
C720 VN.n616 a_400_38200# 0.15fF
C721 VN.t130 a_400_38200# 0.02fF
C722 VN.n618 a_400_38200# 0.26fF
C723 VN.n619 a_400_38200# 0.39fF
C724 VN.n620 a_400_38200# 0.66fF
C725 VN.n621 a_400_38200# 1.01fF
C726 VN.n622 a_400_38200# 0.35fF
C727 VN.n623 a_400_38200# 0.35fF
C728 VN.n624 a_400_38200# 1.01fF
C729 VN.n625 a_400_38200# 1.19fF
C730 VN.n626 a_400_38200# 0.17fF
C731 VN.n627 a_400_38200# 5.41fF
C732 VN.t55 a_400_38200# 0.03fF
C733 VN.n628 a_400_38200# 0.13fF
C734 VN.n629 a_400_38200# 0.16fF
C735 VN.t355 a_400_38200# 0.03fF
C736 VN.n631 a_400_38200# 0.26fF
C737 VN.n632 a_400_38200# 1.00fF
C738 VN.n633 a_400_38200# 0.05fF
C739 VN.n634 a_400_38200# 2.05fF
C740 VN.n635 a_400_38200# 2.91fF
C741 VN.t366 a_400_38200# 0.02fF
C742 VN.n636 a_400_38200# 0.26fF
C743 VN.n637 a_400_38200# 0.39fF
C744 VN.n638 a_400_38200# 0.66fF
C745 VN.n639 a_400_38200# 0.13fF
C746 VN.t204 a_400_38200# 0.02fF
C747 VN.n640 a_400_38200# 0.15fF
C748 VN.n642 a_400_38200# 2.05fF
C749 VN.n643 a_400_38200# 2.92fF
C750 VN.t206 a_400_38200# 0.02fF
C751 VN.n644 a_400_38200# 0.26fF
C752 VN.n645 a_400_38200# 0.39fF
C753 VN.n646 a_400_38200# 0.66fF
C754 VN.t99 a_400_38200# 0.02fF
C755 VN.n647 a_400_38200# 1.33fF
C756 VN.n648 a_400_38200# 0.66fF
C757 VN.n649 a_400_38200# 0.39fF
C758 VN.n650 a_400_38200# 0.69fF
C759 VN.n651 a_400_38200# 1.26fF
C760 VN.n652 a_400_38200# 1.65fF
C761 VN.n653 a_400_38200# 0.65fF
C762 VN.n654 a_400_38200# 0.02fF
C763 VN.n655 a_400_38200# 1.06fF
C764 VN.t74 a_400_38200# 9.89fF
C765 VN.n656 a_400_38200# 10.65fF
C766 VN.n658 a_400_38200# 0.41fF
C767 VN.n659 a_400_38200# 0.25fF
C768 VN.n660 a_400_38200# 3.15fF
C769 VN.n661 a_400_38200# 2.68fF
C770 VN.n662 a_400_38200# 2.76fF
C771 VN.n663 a_400_38200# 4.30fF
C772 VN.n664 a_400_38200# 0.27fF
C773 VN.n665 a_400_38200# 0.01fF
C774 VN.t296 a_400_38200# 0.02fF
C775 VN.n666 a_400_38200# 0.28fF
C776 VN.t340 a_400_38200# 0.03fF
C777 VN.n667 a_400_38200# 1.04fF
C778 VN.n668 a_400_38200# 0.77fF
C779 VN.n669 a_400_38200# 2.05fF
C780 VN.n670 a_400_38200# 0.46fF
C781 VN.n671 a_400_38200# 0.52fF
C782 VN.n672 a_400_38200# 0.10fF
C783 VN.n673 a_400_38200# 0.36fF
C784 VN.n674 a_400_38200# 0.33fF
C785 VN.n675 a_400_38200# 0.84fF
C786 VN.n676 a_400_38200# 0.64fF
C787 VN.t338 a_400_38200# 0.02fF
C788 VN.n677 a_400_38200# 0.26fF
C789 VN.n678 a_400_38200# 0.39fF
C790 VN.n679 a_400_38200# 0.66fF
C791 VN.n680 a_400_38200# 0.13fF
C792 VN.t165 a_400_38200# 0.02fF
C793 VN.n681 a_400_38200# 0.15fF
C794 VN.n683 a_400_38200# 1.57fF
C795 VN.n684 a_400_38200# 2.35fF
C796 VN.t219 a_400_38200# 0.03fF
C797 VN.n685 a_400_38200# 0.26fF
C798 VN.n686 a_400_38200# 1.00fF
C799 VN.n687 a_400_38200# 0.05fF
C800 VN.t202 a_400_38200# 0.03fF
C801 VN.n688 a_400_38200# 0.13fF
C802 VN.n689 a_400_38200# 0.16fF
C803 VN.n691 a_400_38200# 0.85fF
C804 VN.n692 a_400_38200# 2.51fF
C805 VN.n693 a_400_38200# 2.05fF
C806 VN.n694 a_400_38200# 0.13fF
C807 VN.t28 a_400_38200# 0.02fF
C808 VN.n695 a_400_38200# 0.15fF
C809 VN.t214 a_400_38200# 0.02fF
C810 VN.n697 a_400_38200# 0.26fF
C811 VN.n698 a_400_38200# 0.39fF
C812 VN.n699 a_400_38200# 0.66fF
C813 VN.n700 a_400_38200# 1.51fF
C814 VN.n701 a_400_38200# 1.24fF
C815 VN.n702 a_400_38200# 0.38fF
C816 VN.n703 a_400_38200# 2.21fF
C817 VN.t92 a_400_38200# 0.03fF
C818 VN.n704 a_400_38200# 0.26fF
C819 VN.n705 a_400_38200# 1.00fF
C820 VN.n706 a_400_38200# 0.05fF
C821 VN.t69 a_400_38200# 0.03fF
C822 VN.n707 a_400_38200# 0.13fF
C823 VN.n708 a_400_38200# 0.16fF
C824 VN.n710 a_400_38200# 2.06fF
C825 VN.n711 a_400_38200# 2.05fF
C826 VN.t89 a_400_38200# 0.02fF
C827 VN.n712 a_400_38200# 0.26fF
C828 VN.n713 a_400_38200# 0.39fF
C829 VN.n714 a_400_38200# 0.66fF
C830 VN.n715 a_400_38200# 0.13fF
C831 VN.t281 a_400_38200# 0.02fF
C832 VN.n716 a_400_38200# 0.15fF
C833 VN.n718 a_400_38200# 1.26fF
C834 VN.n719 a_400_38200# 0.24fF
C835 VN.n720 a_400_38200# 2.06fF
C836 VN.t348 a_400_38200# 0.03fF
C837 VN.n721 a_400_38200# 0.26fF
C838 VN.n722 a_400_38200# 1.00fF
C839 VN.n723 a_400_38200# 0.05fF
C840 VN.t316 a_400_38200# 0.03fF
C841 VN.n724 a_400_38200# 0.13fF
C842 VN.n725 a_400_38200# 0.16fF
C843 VN.n727 a_400_38200# 9.61fF
C844 VN.n728 a_400_38200# 3.21fF
C845 VN.n729 a_400_38200# 2.05fF
C846 VN.n730 a_400_38200# 0.13fF
C847 VN.t156 a_400_38200# 0.02fF
C848 VN.n731 a_400_38200# 0.15fF
C849 VN.t330 a_400_38200# 0.02fF
C850 VN.n733 a_400_38200# 0.26fF
C851 VN.n734 a_400_38200# 0.39fF
C852 VN.n735 a_400_38200# 0.66fF
C853 VN.n736 a_400_38200# 1.19fF
C854 VN.n737 a_400_38200# 0.17fF
C855 VN.n738 a_400_38200# 2.29fF
C856 VN.t191 a_400_38200# 0.03fF
C857 VN.n739 a_400_38200# 0.13fF
C858 VN.n740 a_400_38200# 0.16fF
C859 VN.t225 a_400_38200# 0.03fF
C860 VN.n742 a_400_38200# 0.26fF
C861 VN.n743 a_400_38200# 1.00fF
C862 VN.n744 a_400_38200# 0.05fF
C863 VN.n745 a_400_38200# 2.97fF
C864 VN.n746 a_400_38200# 1.74fF
C865 VN.n747 a_400_38200# 0.13fF
C866 VN.t289 a_400_38200# 0.02fF
C867 VN.n748 a_400_38200# 0.15fF
C868 VN.t75 a_400_38200# 0.02fF
C869 VN.n750 a_400_38200# 0.26fF
C870 VN.n751 a_400_38200# 0.39fF
C871 VN.n752 a_400_38200# 0.66fF
C872 VN.n753 a_400_38200# 0.07fF
C873 VN.n754 a_400_38200# 0.01fF
C874 VN.n755 a_400_38200# 0.02fF
C875 VN.n756 a_400_38200# 0.02fF
C876 VN.n757 a_400_38200# 0.26fF
C877 VN.n758 a_400_38200# 1.27fF
C878 VN.n759 a_400_38200# 1.47fF
C879 VN.n760 a_400_38200# 2.51fF
C880 VN.t303 a_400_38200# 0.03fF
C881 VN.n761 a_400_38200# 0.13fF
C882 VN.n762 a_400_38200# 0.16fF
C883 VN.t337 a_400_38200# 0.03fF
C884 VN.n764 a_400_38200# 0.26fF
C885 VN.n765 a_400_38200# 1.00fF
C886 VN.n766 a_400_38200# 0.05fF
C887 VN.t13 a_400_38200# 21.51fF
C888 VN.t98 a_400_38200# 0.03fF
C889 VN.n767 a_400_38200# 0.26fF
C890 VN.n768 a_400_38200# 1.00fF
C891 VN.n769 a_400_38200# 0.05fF
C892 VN.t59 a_400_38200# 0.03fF
C893 VN.n770 a_400_38200# 0.13fF
C894 VN.n771 a_400_38200# 0.16fF
C895 VN.n773 a_400_38200# 0.13fF
C896 VN.t14 a_400_38200# 0.02fF
C897 VN.n774 a_400_38200# 0.15fF
C898 VN.n776 a_400_38200# 5.65fF
C899 VN.n777 a_400_38200# 5.33fF
C900 VN.t298 a_400_38200# 0.03fF
C901 VN.n778 a_400_38200# 0.13fF
C902 VN.n779 a_400_38200# 0.16fF
C903 VN.t234 a_400_38200# 0.03fF
C904 VN.n781 a_400_38200# 0.26fF
C905 VN.n782 a_400_38200# 1.00fF
C906 VN.n783 a_400_38200# 0.05fF
C907 VN.n784 a_400_38200# 2.05fF
C908 VN.n785 a_400_38200# 2.92fF
C909 VN.t246 a_400_38200# 0.02fF
C910 VN.n786 a_400_38200# 0.26fF
C911 VN.n787 a_400_38200# 0.39fF
C912 VN.n788 a_400_38200# 0.66fF
C913 VN.n789 a_400_38200# 0.13fF
C914 VN.t72 a_400_38200# 0.02fF
C915 VN.n790 a_400_38200# 0.15fF
C916 VN.n792 a_400_38200# 5.94fF
C917 VN.t169 a_400_38200# 0.03fF
C918 VN.n793 a_400_38200# 0.13fF
C919 VN.n794 a_400_38200# 0.16fF
C920 VN.t109 a_400_38200# 0.03fF
C921 VN.n796 a_400_38200# 0.26fF
C922 VN.n797 a_400_38200# 1.00fF
C923 VN.n798 a_400_38200# 0.05fF
C924 VN.t17 a_400_38200# 21.10fF
C925 VN.t343 a_400_38200# 0.03fF
C926 VN.n799 a_400_38200# 1.30fF
C927 VN.n800 a_400_38200# 0.05fF
C928 VN.t63 a_400_38200# 0.03fF
C929 VN.n801 a_400_38200# 0.01fF
C930 VN.n802 a_400_38200# 0.28fF
C931 VN.n804 a_400_38200# 1.64fF
C932 VN.n805 a_400_38200# 1.37fF
C933 VN.n806 a_400_38200# 0.30fF
C934 VN.n807 a_400_38200# 0.27fF
C935 VN.n808 a_400_38200# 4.79fF
C936 VN.n809 a_400_38200# 0.01fF
C937 VN.n810 a_400_38200# 0.02fF
C938 VN.n811 a_400_38200# 0.03fF
C939 VN.n812 a_400_38200# 0.04fF
C940 VN.n813 a_400_38200# 0.19fF
C941 VN.n814 a_400_38200# 0.01fF
C942 VN.n815 a_400_38200# 0.02fF
C943 VN.n816 a_400_38200# 0.01fF
C944 VN.n817 a_400_38200# 0.01fF
C945 VN.n818 a_400_38200# 0.01fF
C946 VN.n819 a_400_38200# 0.02fF
C947 VN.n820 a_400_38200# 0.03fF
C948 VN.n821 a_400_38200# 0.05fF
C949 VN.n822 a_400_38200# 0.04fF
C950 VN.n823 a_400_38200# 0.12fF
C951 VN.n824 a_400_38200# 0.41fF
C952 VN.n825 a_400_38200# 0.22fF
C953 VN.n826 a_400_38200# 30.53fF
C954 VN.n827 a_400_38200# 30.53fF
C955 VN.n828 a_400_38200# 30.53fF
C956 VN.n829 a_400_38200# 30.53fF
C957 VN.n830 a_400_38200# 0.65fF
C958 VN.n831 a_400_38200# 0.24fF
C959 VN.n832 a_400_38200# 0.65fF
C960 VN.n833 a_400_38200# 2.08fF
C961 VN.n834 a_400_38200# 0.31fF
C962 VN.t91 a_400_38200# 9.89fF
C963 VN.n835 a_400_38200# 12.19fF
C964 VN.n836 a_400_38200# 0.84fF
C965 VN.n837 a_400_38200# 0.30fF
C966 VN.n838 a_400_38200# 4.37fF
C967 VN.n839 a_400_38200# 1.47fF
C968 VN.t242 a_400_38200# 0.02fF
C969 VN.n840 a_400_38200# 0.70fF
C970 VN.n841 a_400_38200# 0.66fF
C971 VN.n842 a_400_38200# 2.05fF
C972 VN.n843 a_400_38200# 0.50fF
C973 VN.n844 a_400_38200# 0.24fF
C974 VN.n845 a_400_38200# 0.41fF
C975 VN.n846 a_400_38200# 0.17fF
C976 VN.n847 a_400_38200# 0.31fF
C977 VN.n848 a_400_38200# 0.23fF
C978 VN.n849 a_400_38200# 0.33fF
C979 VN.n850 a_400_38200# 0.22fF
C980 VN.t120 a_400_38200# 0.02fF
C981 VN.n851 a_400_38200# 0.26fF
C982 VN.n852 a_400_38200# 0.39fF
C983 VN.n853 a_400_38200# 0.66fF
C984 VN.n854 a_400_38200# 0.13fF
C985 VN.t319 a_400_38200# 0.02fF
C986 VN.n855 a_400_38200# 0.15fF
C987 VN.n857 a_400_38200# 0.05fF
C988 VN.n858 a_400_38200# 0.04fF
C989 VN.n859 a_400_38200# 0.03fF
C990 VN.n860 a_400_38200# 0.11fF
C991 VN.n861 a_400_38200# 0.40fF
C992 VN.n862 a_400_38200# 0.41fF
C993 VN.n863 a_400_38200# 0.12fF
C994 VN.n864 a_400_38200# 0.13fF
C995 VN.n865 a_400_38200# 0.08fF
C996 VN.n866 a_400_38200# 0.13fF
C997 VN.n867 a_400_38200# 0.20fF
C998 VN.n868 a_400_38200# 4.36fF
C999 VN.t210 a_400_38200# 0.03fF
C1000 VN.n869 a_400_38200# 0.26fF
C1001 VN.n870 a_400_38200# 1.00fF
C1002 VN.n871 a_400_38200# 0.05fF
C1003 VN.t38 a_400_38200# 0.03fF
C1004 VN.n872 a_400_38200# 0.13fF
C1005 VN.n873 a_400_38200# 0.16fF
C1006 VN.n875 a_400_38200# 0.27fF
C1007 VN.n876 a_400_38200# 0.10fF
C1008 VN.n877 a_400_38200# 0.23fF
C1009 VN.n878 a_400_38200# 1.40fF
C1010 VN.n879 a_400_38200# 0.58fF
C1011 VN.n880 a_400_38200# 2.05fF
C1012 VN.n881 a_400_38200# 0.13fF
C1013 VN.t213 a_400_38200# 0.02fF
C1014 VN.n882 a_400_38200# 0.15fF
C1015 VN.t376 a_400_38200# 0.02fF
C1016 VN.n884 a_400_38200# 0.26fF
C1017 VN.n885 a_400_38200# 0.39fF
C1018 VN.n886 a_400_38200# 0.66fF
C1019 VN.n887 a_400_38200# 0.78fF
C1020 VN.n888 a_400_38200# 1.72fF
C1021 VN.n889 a_400_38200# 2.67fF
C1022 VN.t308 a_400_38200# 0.03fF
C1023 VN.n890 a_400_38200# 0.26fF
C1024 VN.n891 a_400_38200# 1.00fF
C1025 VN.n892 a_400_38200# 0.05fF
C1026 VN.t284 a_400_38200# 0.03fF
C1027 VN.n893 a_400_38200# 0.13fF
C1028 VN.n894 a_400_38200# 0.16fF
C1029 VN.n896 a_400_38200# 2.06fF
C1030 VN.n897 a_400_38200# 0.06fF
C1031 VN.n898 a_400_38200# 0.03fF
C1032 VN.n899 a_400_38200# 0.04fF
C1033 VN.n900 a_400_38200# 1.08fF
C1034 VN.n901 a_400_38200# 0.02fF
C1035 VN.n902 a_400_38200# 0.01fF
C1036 VN.n903 a_400_38200# 0.02fF
C1037 VN.n904 a_400_38200# 0.09fF
C1038 VN.n905 a_400_38200# 0.39fF
C1039 VN.n906 a_400_38200# 2.02fF
C1040 VN.t253 a_400_38200# 0.02fF
C1041 VN.n907 a_400_38200# 0.26fF
C1042 VN.n908 a_400_38200# 0.39fF
C1043 VN.n909 a_400_38200# 0.66fF
C1044 VN.n910 a_400_38200# 0.13fF
C1045 VN.t83 a_400_38200# 0.02fF
C1046 VN.n911 a_400_38200# 0.15fF
C1047 VN.n913 a_400_38200# 0.76fF
C1048 VN.n914 a_400_38200# 0.25fF
C1049 VN.n915 a_400_38200# 0.28fF
C1050 VN.n916 a_400_38200# 0.10fF
C1051 VN.n917 a_400_38200# 0.25fF
C1052 VN.n918 a_400_38200# 0.76fF
C1053 VN.n919 a_400_38200# 1.26fF
C1054 VN.n920 a_400_38200# 0.24fF
C1055 VN.n921 a_400_38200# 0.28fF
C1056 VN.n922 a_400_38200# 0.10fF
C1057 VN.n923 a_400_38200# 2.06fF
C1058 VN.t180 a_400_38200# 0.03fF
C1059 VN.n924 a_400_38200# 0.26fF
C1060 VN.n925 a_400_38200# 1.00fF
C1061 VN.n926 a_400_38200# 0.05fF
C1062 VN.t181 a_400_38200# 0.03fF
C1063 VN.n927 a_400_38200# 0.13fF
C1064 VN.n928 a_400_38200# 0.16fF
C1065 VN.n930 a_400_38200# 9.61fF
C1066 VN.n931 a_400_38200# 1.87fF
C1067 VN.n932 a_400_38200# 0.72fF
C1068 VN.n933 a_400_38200# 0.76fF
C1069 VN.n934 a_400_38200# 0.79fF
C1070 VN.n935 a_400_38200# 0.40fF
C1071 VN.t227 a_400_38200# 0.02fF
C1072 VN.n936 a_400_38200# 0.26fF
C1073 VN.n937 a_400_38200# 0.39fF
C1074 VN.n938 a_400_38200# 0.66fF
C1075 VN.n939 a_400_38200# 0.13fF
C1076 VN.t77 a_400_38200# 0.02fF
C1077 VN.n940 a_400_38200# 0.15fF
C1078 VN.n942 a_400_38200# 0.34fF
C1079 VN.n943 a_400_38200# 0.28fF
C1080 VN.n944 a_400_38200# 0.10fF
C1081 VN.n945 a_400_38200# 0.25fF
C1082 VN.n946 a_400_38200# 0.72fF
C1083 VN.n947 a_400_38200# 1.04fF
C1084 VN.n948 a_400_38200# 0.25fF
C1085 VN.n949 a_400_38200# 0.23fF
C1086 VN.n950 a_400_38200# 0.22fF
C1087 VN.n951 a_400_38200# 0.07fF
C1088 VN.n952 a_400_38200# 0.10fF
C1089 VN.n953 a_400_38200# 0.10fF
C1090 VN.n954 a_400_38200# 1.83fF
C1091 VN.t173 a_400_38200# 0.03fF
C1092 VN.n955 a_400_38200# 0.13fF
C1093 VN.n956 a_400_38200# 0.16fF
C1094 VN.t318 a_400_38200# 0.03fF
C1095 VN.n958 a_400_38200# 0.26fF
C1096 VN.n959 a_400_38200# 1.00fF
C1097 VN.n960 a_400_38200# 0.05fF
C1098 VN.t282 a_400_38200# 0.03fF
C1099 VN.n961 a_400_38200# 0.26fF
C1100 VN.n962 a_400_38200# 1.01fF
C1101 VN.n963 a_400_38200# 2.05fF
C1102 VN.n964 a_400_38200# 1.69fF
C1103 VN.n965 a_400_38200# 0.17fF
C1104 VN.t259 a_400_38200# 0.03fF
C1105 VN.n966 a_400_38200# 0.13fF
C1106 VN.n967 a_400_38200# 0.16fF
C1107 VN.n968 a_400_38200# 0.13fF
C1108 VN.t230 a_400_38200# 0.02fF
C1109 VN.n969 a_400_38200# 0.15fF
C1110 VN.t64 a_400_38200# 0.02fF
C1111 VN.n970 a_400_38200# 1.33fF
C1112 VN.n971 a_400_38200# 0.66fF
C1113 VN.n972 a_400_38200# 0.39fF
C1114 VN.n973 a_400_38200# 0.69fF
C1115 VN.n974 a_400_38200# 1.26fF
C1116 VN.n975 a_400_38200# 1.65fF
C1117 VN.n976 a_400_38200# 0.65fF
C1118 VN.n977 a_400_38200# 0.02fF
C1119 VN.n978 a_400_38200# 1.06fF
C1120 VN.t47 a_400_38200# 9.89fF
C1121 VN.n979 a_400_38200# 10.65fF
C1122 VN.n981 a_400_38200# 0.41fF
C1123 VN.n982 a_400_38200# 0.25fF
C1124 VN.n983 a_400_38200# 3.16fF
C1125 VN.n984 a_400_38200# 2.68fF
C1126 VN.n985 a_400_38200# 2.14fF
C1127 VN.n986 a_400_38200# 4.67fF
C1128 VN.n987 a_400_38200# 0.27fF
C1129 VN.n988 a_400_38200# 0.01fF
C1130 VN.t267 a_400_38200# 0.02fF
C1131 VN.n989 a_400_38200# 0.28fF
C1132 VN.t312 a_400_38200# 0.03fF
C1133 VN.n990 a_400_38200# 1.04fF
C1134 VN.n991 a_400_38200# 0.77fF
C1135 VN.n992 a_400_38200# 2.06fF
C1136 VN.n993 a_400_38200# 1.89fF
C1137 VN.t306 a_400_38200# 0.02fF
C1138 VN.n994 a_400_38200# 0.26fF
C1139 VN.n995 a_400_38200# 0.39fF
C1140 VN.n996 a_400_38200# 0.66fF
C1141 VN.n997 a_400_38200# 0.13fF
C1142 VN.t141 a_400_38200# 0.02fF
C1143 VN.n998 a_400_38200# 0.15fF
C1144 VN.n1000 a_400_38200# 0.76fF
C1145 VN.n1001 a_400_38200# 1.26fF
C1146 VN.n1002 a_400_38200# 0.24fF
C1147 VN.n1003 a_400_38200# 2.66fF
C1148 VN.t185 a_400_38200# 0.03fF
C1149 VN.n1004 a_400_38200# 0.26fF
C1150 VN.n1005 a_400_38200# 1.00fF
C1151 VN.n1006 a_400_38200# 0.05fF
C1152 VN.t161 a_400_38200# 0.03fF
C1153 VN.n1007 a_400_38200# 0.13fF
C1154 VN.n1008 a_400_38200# 0.16fF
C1155 VN.n1010 a_400_38200# 2.05fF
C1156 VN.n1011 a_400_38200# 0.46fF
C1157 VN.n1012 a_400_38200# 0.52fF
C1158 VN.n1013 a_400_38200# 0.10fF
C1159 VN.n1014 a_400_38200# 0.36fF
C1160 VN.n1015 a_400_38200# 0.33fF
C1161 VN.n1016 a_400_38200# 0.84fF
C1162 VN.n1017 a_400_38200# 0.64fF
C1163 VN.t176 a_400_38200# 0.02fF
C1164 VN.n1018 a_400_38200# 0.26fF
C1165 VN.n1019 a_400_38200# 0.39fF
C1166 VN.n1020 a_400_38200# 0.66fF
C1167 VN.n1021 a_400_38200# 0.13fF
C1168 VN.t383 a_400_38200# 0.02fF
C1169 VN.n1022 a_400_38200# 0.15fF
C1170 VN.n1024 a_400_38200# 2.85fF
C1171 VN.n1025 a_400_38200# 2.35fF
C1172 VN.t56 a_400_38200# 0.03fF
C1173 VN.n1026 a_400_38200# 0.26fF
C1174 VN.n1027 a_400_38200# 1.00fF
C1175 VN.n1028 a_400_38200# 0.05fF
C1176 VN.t23 a_400_38200# 0.03fF
C1177 VN.n1029 a_400_38200# 0.13fF
C1178 VN.n1030 a_400_38200# 0.16fF
C1179 VN.n1032 a_400_38200# 0.85fF
C1180 VN.n1033 a_400_38200# 2.51fF
C1181 VN.n1034 a_400_38200# 2.05fF
C1182 VN.n1035 a_400_38200# 0.13fF
C1183 VN.t115 a_400_38200# 0.02fF
C1184 VN.n1036 a_400_38200# 0.15fF
C1185 VN.t276 a_400_38200# 0.02fF
C1186 VN.n1038 a_400_38200# 0.26fF
C1187 VN.n1039 a_400_38200# 0.39fF
C1188 VN.n1040 a_400_38200# 0.66fF
C1189 VN.n1041 a_400_38200# 1.51fF
C1190 VN.n1042 a_400_38200# 1.24fF
C1191 VN.n1043 a_400_38200# 0.38fF
C1192 VN.n1044 a_400_38200# 2.21fF
C1193 VN.t170 a_400_38200# 0.03fF
C1194 VN.n1045 a_400_38200# 0.26fF
C1195 VN.n1046 a_400_38200# 1.00fF
C1196 VN.n1047 a_400_38200# 0.05fF
C1197 VN.t140 a_400_38200# 0.03fF
C1198 VN.n1048 a_400_38200# 0.13fF
C1199 VN.n1049 a_400_38200# 0.16fF
C1200 VN.n1051 a_400_38200# 2.06fF
C1201 VN.n1052 a_400_38200# 2.92fF
C1202 VN.t150 a_400_38200# 0.02fF
C1203 VN.n1053 a_400_38200# 0.26fF
C1204 VN.n1054 a_400_38200# 0.39fF
C1205 VN.n1055 a_400_38200# 0.66fF
C1206 VN.n1056 a_400_38200# 0.13fF
C1207 VN.t352 a_400_38200# 0.02fF
C1208 VN.n1057 a_400_38200# 0.15fF
C1209 VN.n1059 a_400_38200# 0.76fF
C1210 VN.n1060 a_400_38200# 1.26fF
C1211 VN.n1061 a_400_38200# 0.24fF
C1212 VN.n1062 a_400_38200# 2.06fF
C1213 VN.t31 a_400_38200# 0.03fF
C1214 VN.n1063 a_400_38200# 0.26fF
C1215 VN.n1064 a_400_38200# 1.00fF
C1216 VN.n1065 a_400_38200# 0.05fF
C1217 VN.t382 a_400_38200# 0.03fF
C1218 VN.n1066 a_400_38200# 0.13fF
C1219 VN.n1067 a_400_38200# 0.16fF
C1220 VN.n1069 a_400_38200# 9.61fF
C1221 VN.n1070 a_400_38200# 2.97fF
C1222 VN.n1071 a_400_38200# 1.73fF
C1223 VN.n1072 a_400_38200# 0.13fF
C1224 VN.t122 a_400_38200# 0.02fF
C1225 VN.n1073 a_400_38200# 0.15fF
C1226 VN.t268 a_400_38200# 0.02fF
C1227 VN.n1075 a_400_38200# 0.26fF
C1228 VN.n1076 a_400_38200# 0.39fF
C1229 VN.n1077 a_400_38200# 0.66fF
C1230 VN.n1078 a_400_38200# 2.58fF
C1231 VN.n1079 a_400_38200# 2.51fF
C1232 VN.t131 a_400_38200# 0.03fF
C1233 VN.n1080 a_400_38200# 0.13fF
C1234 VN.n1081 a_400_38200# 0.16fF
C1235 VN.t157 a_400_38200# 0.03fF
C1236 VN.n1083 a_400_38200# 0.26fF
C1237 VN.n1084 a_400_38200# 1.00fF
C1238 VN.n1085 a_400_38200# 0.05fF
C1239 VN.n1086 a_400_38200# 0.26fF
C1240 VN.t390 a_400_38200# 0.02fF
C1241 VN.n1087 a_400_38200# 0.99fF
C1242 VN.t22 a_400_38200# 27.04fF
C1243 VN.n1088 a_400_38200# 2.05fF
C1244 VN.n1089 a_400_38200# 0.13fF
C1245 VN.t325 a_400_38200# 0.02fF
C1246 VN.n1090 a_400_38200# 0.15fF
C1247 VN.t126 a_400_38200# 0.02fF
C1248 VN.n1092 a_400_38200# 0.26fF
C1249 VN.n1093 a_400_38200# 0.39fF
C1250 VN.n1094 a_400_38200# 0.66fF
C1251 VN.n1095 a_400_38200# 1.01fF
C1252 VN.n1096 a_400_38200# 0.35fF
C1253 VN.n1097 a_400_38200# 0.35fF
C1254 VN.n1098 a_400_38200# 1.01fF
C1255 VN.n1099 a_400_38200# 1.19fF
C1256 VN.n1100 a_400_38200# 0.17fF
C1257 VN.n1101 a_400_38200# 5.11fF
C1258 VN.t49 a_400_38200# 0.03fF
C1259 VN.n1102 a_400_38200# 0.13fF
C1260 VN.n1103 a_400_38200# 0.16fF
C1261 VN.t48 a_400_38200# 0.03fF
C1262 VN.n1105 a_400_38200# 0.26fF
C1263 VN.n1106 a_400_38200# 1.00fF
C1264 VN.n1107 a_400_38200# 0.05fF
C1265 VN.n1108 a_400_38200# 2.05fF
C1266 VN.n1109 a_400_38200# 2.92fF
C1267 VN.t365 a_400_38200# 0.02fF
C1268 VN.n1110 a_400_38200# 0.26fF
C1269 VN.n1111 a_400_38200# 0.39fF
C1270 VN.n1112 a_400_38200# 0.66fF
C1271 VN.n1113 a_400_38200# 0.13fF
C1272 VN.t199 a_400_38200# 0.02fF
C1273 VN.n1114 a_400_38200# 0.15fF
C1274 VN.n1116 a_400_38200# 5.95fF
C1275 VN.t293 a_400_38200# 0.03fF
C1276 VN.n1117 a_400_38200# 0.13fF
C1277 VN.n1118 a_400_38200# 0.16fF
C1278 VN.t292 a_400_38200# 0.03fF
C1279 VN.n1120 a_400_38200# 0.26fF
C1280 VN.n1121 a_400_38200# 1.00fF
C1281 VN.n1122 a_400_38200# 0.05fF
C1282 VN.t37 a_400_38200# 21.10fF
C1283 VN.t162 a_400_38200# 0.03fF
C1284 VN.n1123 a_400_38200# 1.30fF
C1285 VN.n1124 a_400_38200# 0.05fF
C1286 VN.t189 a_400_38200# 0.03fF
C1287 VN.n1125 a_400_38200# 0.01fF
C1288 VN.n1126 a_400_38200# 0.28fF
C1289 VN.n1128 a_400_38200# 1.64fF
C1290 VN.n1129 a_400_38200# 1.42fF
C1291 VN.n1130 a_400_38200# 0.30fF
C1292 VN.n1131 a_400_38200# 0.27fF
C1293 VN.n1132 a_400_38200# 4.79fF
C1294 VN.n1133 a_400_38200# 0.27fF
C1295 VN.n1134 a_400_38200# 0.65fF
C1296 VN.n1135 a_400_38200# 0.24fF
C1297 VN.n1136 a_400_38200# 0.65fF
C1298 VN.n1137 a_400_38200# 2.08fF
C1299 VN.n1138 a_400_38200# 0.31fF
C1300 VN.t30 a_400_38200# 9.89fF
C1301 VN.n1139 a_400_38200# 12.19fF
C1302 VN.n1140 a_400_38200# 0.84fF
C1303 VN.n1141 a_400_38200# 0.30fF
C1304 VN.n1142 a_400_38200# 4.37fF
C1305 VN.n1143 a_400_38200# 1.64fF
C1306 VN.n1144 a_400_38200# 1.42fF
C1307 VN.n1145 a_400_38200# 0.30fF
C1308 VN.n1146 a_400_38200# 2.06fF
C1309 VN.n1147 a_400_38200# 0.04fF
C1310 VN.n1148 a_400_38200# 0.07fF
C1311 VN.n1149 a_400_38200# 0.06fF
C1312 VN.n1150 a_400_38200# 0.94fF
C1313 VN.n1151 a_400_38200# 0.01fF
C1314 VN.n1152 a_400_38200# 0.01fF
C1315 VN.n1153 a_400_38200# 0.01fF
C1316 VN.n1154 a_400_38200# 0.08fF
C1317 VN.n1155 a_400_38200# 0.75fF
C1318 VN.n1156 a_400_38200# 0.77fF
C1319 VN.t88 a_400_38200# 0.02fF
C1320 VN.n1157 a_400_38200# 0.26fF
C1321 VN.n1158 a_400_38200# 0.39fF
C1322 VN.n1159 a_400_38200# 0.66fF
C1323 VN.n1160 a_400_38200# 0.13fF
C1324 VN.t283 a_400_38200# 0.02fF
C1325 VN.n1161 a_400_38200# 0.15fF
C1326 VN.n1163 a_400_38200# 0.25fF
C1327 VN.n1164 a_400_38200# 1.04fF
C1328 VN.n1165 a_400_38200# 0.64fF
C1329 VN.n1166 a_400_38200# 0.28fF
C1330 VN.n1167 a_400_38200# 0.10fF
C1331 VN.n1168 a_400_38200# 2.52fF
C1332 VN.t252 a_400_38200# 0.03fF
C1333 VN.n1169 a_400_38200# 0.26fF
C1334 VN.n1170 a_400_38200# 1.00fF
C1335 VN.n1171 a_400_38200# 0.05fF
C1336 VN.t385 a_400_38200# 0.03fF
C1337 VN.n1172 a_400_38200# 0.13fF
C1338 VN.n1173 a_400_38200# 0.16fF
C1339 VN.n1175 a_400_38200# 2.05fF
C1340 VN.n1176 a_400_38200# 0.50fF
C1341 VN.n1177 a_400_38200# 0.24fF
C1342 VN.n1178 a_400_38200# 0.41fF
C1343 VN.n1179 a_400_38200# 0.17fF
C1344 VN.n1180 a_400_38200# 0.31fF
C1345 VN.n1181 a_400_38200# 0.23fF
C1346 VN.n1182 a_400_38200# 0.33fF
C1347 VN.n1183 a_400_38200# 0.22fF
C1348 VN.t205 a_400_38200# 0.02fF
C1349 VN.n1184 a_400_38200# 0.26fF
C1350 VN.n1185 a_400_38200# 0.39fF
C1351 VN.n1186 a_400_38200# 0.66fF
C1352 VN.n1187 a_400_38200# 0.13fF
C1353 VN.t12 a_400_38200# 0.02fF
C1354 VN.n1188 a_400_38200# 0.15fF
C1355 VN.n1190 a_400_38200# 2.05fF
C1356 VN.n1191 a_400_38200# 0.13fF
C1357 VN.t237 a_400_38200# 0.02fF
C1358 VN.n1192 a_400_38200# 0.15fF
C1359 VN.t111 a_400_38200# 0.02fF
C1360 VN.n1194 a_400_38200# 1.33fF
C1361 VN.n1195 a_400_38200# 0.86fF
C1362 VN.n1196 a_400_38200# 2.50fF
C1363 VN.n1197 a_400_38200# 0.66fF
C1364 VN.n1198 a_400_38200# 0.39fF
C1365 VN.n1199 a_400_38200# 0.69fF
C1366 VN.n1200 a_400_38200# 1.26fF
C1367 VN.n1201 a_400_38200# 1.65fF
C1368 VN.n1202 a_400_38200# 0.65fF
C1369 VN.n1203 a_400_38200# 0.02fF
C1370 VN.n1204 a_400_38200# 1.06fF
C1371 VN.t15 a_400_38200# 9.89fF
C1372 VN.n1205 a_400_38200# 10.65fF
C1373 VN.n1207 a_400_38200# 0.41fF
C1374 VN.n1208 a_400_38200# 0.25fF
C1375 VN.n1209 a_400_38200# 3.15fF
C1376 VN.n1210 a_400_38200# 2.68fF
C1377 VN.n1211 a_400_38200# 4.30fF
C1378 VN.n1212 a_400_38200# 0.27fF
C1379 VN.n1213 a_400_38200# 0.01fF
C1380 VN.t309 a_400_38200# 0.02fF
C1381 VN.n1214 a_400_38200# 0.28fF
C1382 VN.t353 a_400_38200# 0.03fF
C1383 VN.n1215 a_400_38200# 1.04fF
C1384 VN.n1216 a_400_38200# 0.77fF
C1385 VN.n1217 a_400_38200# 2.05fF
C1386 VN.n1218 a_400_38200# 0.85fF
C1387 VN.n1219 a_400_38200# 2.11fF
C1388 VN.n1220 a_400_38200# 0.13fF
C1389 VN.t182 a_400_38200# 0.02fF
C1390 VN.n1221 a_400_38200# 0.15fF
C1391 VN.t346 a_400_38200# 0.02fF
C1392 VN.n1223 a_400_38200# 0.26fF
C1393 VN.n1224 a_400_38200# 0.39fF
C1394 VN.n1225 a_400_38200# 0.66fF
C1395 VN.n1226 a_400_38200# 2.99fF
C1396 VN.n1227 a_400_38200# 3.24fF
C1397 VN.t231 a_400_38200# 0.03fF
C1398 VN.n1228 a_400_38200# 0.26fF
C1399 VN.n1229 a_400_38200# 1.00fF
C1400 VN.n1230 a_400_38200# 0.05fF
C1401 VN.t215 a_400_38200# 0.03fF
C1402 VN.n1231 a_400_38200# 0.13fF
C1403 VN.n1232 a_400_38200# 0.16fF
C1404 VN.n1234 a_400_38200# 2.06fF
C1405 VN.n1235 a_400_38200# 2.16fF
C1406 VN.n1236 a_400_38200# 0.13fF
C1407 VN.t51 a_400_38200# 0.02fF
C1408 VN.n1237 a_400_38200# 0.15fF
C1409 VN.t223 a_400_38200# 0.02fF
C1410 VN.n1239 a_400_38200# 0.26fF
C1411 VN.n1240 a_400_38200# 0.39fF
C1412 VN.n1241 a_400_38200# 0.66fF
C1413 VN.n1242 a_400_38200# 0.02fF
C1414 VN.n1243 a_400_38200# 0.03fF
C1415 VN.n1244 a_400_38200# 0.03fF
C1416 VN.n1245 a_400_38200# 0.02fF
C1417 VN.n1246 a_400_38200# 0.20fF
C1418 VN.n1247 a_400_38200# 0.12fF
C1419 VN.n1248 a_400_38200# 0.68fF
C1420 VN.n1249 a_400_38200# 0.95fF
C1421 VN.n1250 a_400_38200# 2.86fF
C1422 VN.t104 a_400_38200# 0.03fF
C1423 VN.n1251 a_400_38200# 0.26fF
C1424 VN.n1252 a_400_38200# 1.00fF
C1425 VN.n1253 a_400_38200# 0.05fF
C1426 VN.t84 a_400_38200# 0.03fF
C1427 VN.n1254 a_400_38200# 0.13fF
C1428 VN.n1255 a_400_38200# 0.16fF
C1429 VN.n1257 a_400_38200# 0.85fF
C1430 VN.n1258 a_400_38200# 1.31fF
C1431 VN.n1259 a_400_38200# 1.40fF
C1432 VN.n1260 a_400_38200# 2.05fF
C1433 VN.n1261 a_400_38200# 0.13fF
C1434 VN.t113 a_400_38200# 0.02fF
C1435 VN.n1262 a_400_38200# 0.15fF
C1436 VN.t272 a_400_38200# 0.02fF
C1437 VN.n1264 a_400_38200# 0.26fF
C1438 VN.n1265 a_400_38200# 0.39fF
C1439 VN.n1266 a_400_38200# 0.66fF
C1440 VN.n1267 a_400_38200# 1.36fF
C1441 VN.n1268 a_400_38200# 0.38fF
C1442 VN.n1269 a_400_38200# 2.21fF
C1443 VN.t163 a_400_38200# 0.03fF
C1444 VN.n1270 a_400_38200# 0.26fF
C1445 VN.n1271 a_400_38200# 1.00fF
C1446 VN.n1272 a_400_38200# 0.05fF
C1447 VN.t139 a_400_38200# 0.03fF
C1448 VN.n1273 a_400_38200# 0.13fF
C1449 VN.n1274 a_400_38200# 0.16fF
C1450 VN.n1276 a_400_38200# 2.06fF
C1451 VN.n1277 a_400_38200# 1.26fF
C1452 VN.n1278 a_400_38200# 0.24fF
C1453 VN.n1279 a_400_38200# 0.13fF
C1454 VN.t349 a_400_38200# 0.02fF
C1455 VN.n1280 a_400_38200# 0.15fF
C1456 VN.t148 a_400_38200# 0.02fF
C1457 VN.n1282 a_400_38200# 0.26fF
C1458 VN.n1283 a_400_38200# 0.39fF
C1459 VN.n1284 a_400_38200# 0.66fF
C1460 VN.n1285 a_400_38200# 2.98fF
C1461 VN.n1286 a_400_38200# 2.05fF
C1462 VN.t25 a_400_38200# 0.03fF
C1463 VN.n1287 a_400_38200# 0.26fF
C1464 VN.n1288 a_400_38200# 1.00fF
C1465 VN.n1289 a_400_38200# 0.05fF
C1466 VN.t378 a_400_38200# 0.03fF
C1467 VN.n1290 a_400_38200# 0.13fF
C1468 VN.n1291 a_400_38200# 0.16fF
C1469 VN.n1293 a_400_38200# 9.61fF
C1470 VN.n1294 a_400_38200# 2.11fF
C1471 VN.n1295 a_400_38200# 0.13fF
C1472 VN.t245 a_400_38200# 0.02fF
C1473 VN.n1296 a_400_38200# 0.15fF
C1474 VN.t389 a_400_38200# 0.02fF
C1475 VN.n1298 a_400_38200# 0.26fF
C1476 VN.n1299 a_400_38200# 0.39fF
C1477 VN.n1300 a_400_38200# 0.66fF
C1478 VN.n1301 a_400_38200# 1.71fF
C1479 VN.n1302 a_400_38200# 0.30fF
C1480 VN.n1303 a_400_38200# 2.29fF
C1481 VN.t255 a_400_38200# 0.03fF
C1482 VN.n1304 a_400_38200# 0.13fF
C1483 VN.n1305 a_400_38200# 0.16fF
C1484 VN.t278 a_400_38200# 0.03fF
C1485 VN.n1307 a_400_38200# 0.26fF
C1486 VN.n1308 a_400_38200# 1.00fF
C1487 VN.n1309 a_400_38200# 0.05fF
C1488 VN.t50 a_400_38200# 21.51fF
C1489 VN.t264 a_400_38200# 0.03fF
C1490 VN.n1310 a_400_38200# 0.13fF
C1491 VN.n1311 a_400_38200# 0.16fF
C1492 VN.t294 a_400_38200# 0.03fF
C1493 VN.n1313 a_400_38200# 0.26fF
C1494 VN.n1314 a_400_38200# 1.00fF
C1495 VN.n1315 a_400_38200# 0.05fF
C1496 VN.t16 a_400_38200# 0.02fF
C1497 VN.n1316 a_400_38200# 0.26fF
C1498 VN.n1317 a_400_38200# 0.39fF
C1499 VN.n1318 a_400_38200# 0.66fF
C1500 VN.n1319 a_400_38200# 0.99fF
C1501 VN.n1320 a_400_38200# 0.61fF
C1502 VN.n1321 a_400_38200# 1.06fF
C1503 VN.n1322 a_400_38200# 0.10fF
C1504 VN.n1323 a_400_38200# 0.36fF
C1505 VN.n1324 a_400_38200# 2.35fF
C1506 VN.n1325 a_400_38200# 2.85fF
C1507 VN.n1326 a_400_38200# 0.05fF
C1508 VN.n1327 a_400_38200# 0.04fF
C1509 VN.n1328 a_400_38200# 0.03fF
C1510 VN.n1329 a_400_38200# 0.11fF
C1511 VN.n1330 a_400_38200# 0.40fF
C1512 VN.n1331 a_400_38200# 0.41fF
C1513 VN.n1332 a_400_38200# 0.12fF
C1514 VN.n1333 a_400_38200# 0.13fF
C1515 VN.n1334 a_400_38200# 0.08fF
C1516 VN.n1335 a_400_38200# 0.13fF
C1517 VN.n1336 a_400_38200# 0.20fF
C1518 VN.n1337 a_400_38200# 4.36fF
C1519 VN.t60 a_400_38200# 0.03fF
C1520 VN.n1338 a_400_38200# 0.26fF
C1521 VN.n1339 a_400_38200# 1.00fF
C1522 VN.n1340 a_400_38200# 0.05fF
C1523 VN.t263 a_400_38200# 0.03fF
C1524 VN.n1341 a_400_38200# 0.13fF
C1525 VN.n1342 a_400_38200# 0.16fF
C1526 VN.n1344 a_400_38200# 0.27fF
C1527 VN.n1345 a_400_38200# 0.10fF
C1528 VN.n1346 a_400_38200# 0.23fF
C1529 VN.n1347 a_400_38200# 0.87fF
C1530 VN.n1348 a_400_38200# 0.48fF
C1531 VN.n1349 a_400_38200# 2.05fF
C1532 VN.n1350 a_400_38200# 0.13fF
C1533 VN.t271 a_400_38200# 0.02fF
C1534 VN.n1351 a_400_38200# 0.15fF
C1535 VN.t73 a_400_38200# 0.02fF
C1536 VN.n1353 a_400_38200# 0.26fF
C1537 VN.n1354 a_400_38200# 0.39fF
C1538 VN.n1355 a_400_38200# 0.66fF
C1539 VN.n1356 a_400_38200# 0.78fF
C1540 VN.n1357 a_400_38200# 1.72fF
C1541 VN.n1358 a_400_38200# 2.67fF
C1542 VN.t304 a_400_38200# 0.03fF
C1543 VN.n1359 a_400_38200# 0.26fF
C1544 VN.n1360 a_400_38200# 1.00fF
C1545 VN.n1361 a_400_38200# 0.05fF
C1546 VN.t372 a_400_38200# 0.03fF
C1547 VN.n1362 a_400_38200# 0.13fF
C1548 VN.n1363 a_400_38200# 0.16fF
C1549 VN.n1365 a_400_38200# 2.06fF
C1550 VN.n1366 a_400_38200# 2.91fF
C1551 VN.t317 a_400_38200# 0.02fF
C1552 VN.n1367 a_400_38200# 0.26fF
C1553 VN.n1368 a_400_38200# 0.39fF
C1554 VN.n1369 a_400_38200# 0.66fF
C1555 VN.n1370 a_400_38200# 0.13fF
C1556 VN.t146 a_400_38200# 0.02fF
C1557 VN.n1371 a_400_38200# 0.15fF
C1558 VN.n1373 a_400_38200# 0.25fF
C1559 VN.n1374 a_400_38200# 0.28fF
C1560 VN.n1375 a_400_38200# 0.10fF
C1561 VN.n1376 a_400_38200# 0.25fF
C1562 VN.n1377 a_400_38200# 0.76fF
C1563 VN.n1378 a_400_38200# 1.26fF
C1564 VN.n1379 a_400_38200# 0.24fF
C1565 VN.n1380 a_400_38200# 0.28fF
C1566 VN.n1381 a_400_38200# 0.10fF
C1567 VN.n1382 a_400_38200# 2.06fF
C1568 VN.t175 a_400_38200# 0.03fF
C1569 VN.n1383 a_400_38200# 0.26fF
C1570 VN.n1384 a_400_38200# 1.00fF
C1571 VN.n1385 a_400_38200# 0.05fF
C1572 VN.t249 a_400_38200# 0.03fF
C1573 VN.n1386 a_400_38200# 0.13fF
C1574 VN.n1387 a_400_38200# 0.16fF
C1575 VN.n1389 a_400_38200# 9.61fF
C1576 VN.n1390 a_400_38200# 2.55fF
C1577 VN.n1391 a_400_38200# 3.34fF
C1578 VN.t195 a_400_38200# 0.02fF
C1579 VN.n1392 a_400_38200# 0.26fF
C1580 VN.n1393 a_400_38200# 0.39fF
C1581 VN.n1394 a_400_38200# 0.66fF
C1582 VN.n1395 a_400_38200# 0.13fF
C1583 VN.t35 a_400_38200# 0.02fF
C1584 VN.n1396 a_400_38200# 0.15fF
C1585 VN.n1398 a_400_38200# 0.33fF
C1586 VN.n1399 a_400_38200# 0.76fF
C1587 VN.n1400 a_400_38200# 0.49fF
C1588 VN.n1401 a_400_38200# 0.23fF
C1589 VN.n1402 a_400_38200# 0.22fF
C1590 VN.n1403 a_400_38200# 0.07fF
C1591 VN.n1404 a_400_38200# 0.10fF
C1592 VN.n1405 a_400_38200# 0.10fF
C1593 VN.n1406 a_400_38200# 2.28fF
C1594 VN.t144 a_400_38200# 0.03fF
C1595 VN.n1407 a_400_38200# 0.13fF
C1596 VN.n1408 a_400_38200# 0.16fF
C1597 VN.t358 a_400_38200# 0.03fF
C1598 VN.n1410 a_400_38200# 0.26fF
C1599 VN.n1411 a_400_38200# 1.00fF
C1600 VN.n1412 a_400_38200# 0.05fF
C1601 VN.n1413 a_400_38200# 2.98fF
C1602 VN.n1414 a_400_38200# 2.05fF
C1603 VN.n1415 a_400_38200# 0.13fF
C1604 VN.t387 a_400_38200# 0.02fF
C1605 VN.n1416 a_400_38200# 0.15fF
C1606 VN.t192 a_400_38200# 0.02fF
C1607 VN.n1418 a_400_38200# 0.26fF
C1608 VN.n1419 a_400_38200# 0.39fF
C1609 VN.n1420 a_400_38200# 0.66fF
C1610 VN.n1421 a_400_38200# 0.77fF
C1611 VN.n1422 a_400_38200# 1.39fF
C1612 VN.n1423 a_400_38200# 6.51fF
C1613 VN.t124 a_400_38200# 0.03fF
C1614 VN.n1424 a_400_38200# 0.13fF
C1615 VN.n1425 a_400_38200# 0.16fF
C1616 VN.t41 a_400_38200# 0.03fF
C1617 VN.n1427 a_400_38200# 0.26fF
C1618 VN.n1428 a_400_38200# 1.00fF
C1619 VN.n1429 a_400_38200# 0.05fF
C1620 VN.t11 a_400_38200# 21.10fF
C1621 VN.t380 a_400_38200# 0.03fF
C1622 VN.n1430 a_400_38200# 0.01fF
C1623 VN.n1431 a_400_38200# 0.28fF
C1624 VN.t286 a_400_38200# 0.03fF
C1625 VN.n1433 a_400_38200# 1.30fF
C1626 VN.n1434 a_400_38200# 0.05fF
C1627 VN.t61 a_400_38200# 0.02fF
C1628 VN.n1435 a_400_38200# 0.70fF
C1629 VN.n1436 a_400_38200# 0.66fF
C1630 VN.n1437 a_400_38200# 1.64fF
C1631 VN.n1438 a_400_38200# 0.39fF
C1632 VN.n1439 a_400_38200# 1.42fF
C1633 VN.n1440 a_400_38200# 0.17fF
C1634 VN.n1441 a_400_38200# 1.81fF
C1635 VN.n1442 a_400_38200# 2.89fF
C1636 VN.n1443 a_400_38200# 1.28fF
C1637 VN.n1444 a_400_38200# 0.42fF
C1638 VN.n1445 a_400_38200# 1.32fF
C1639 VN.n1446 a_400_38200# 0.40fF
C1640 VN.n1447 a_400_38200# 0.20fF
C1641 VN.n1448 a_400_38200# 0.10fF
C1642 VN.n1449 a_400_38200# 1.03fF
C1643 VN.n1450 a_400_38200# 0.51fF
C1644 VN.n1451 a_400_38200# 0.23fF
C1645 VN.n1452 a_400_38200# 0.39fF
C1646 VN.n1453 a_400_38200# 0.58fF
C1647 VN.n1454 a_400_38200# 2.87fF
C1648 VN.n1455 a_400_38200# 1.64fF
C1649 VN.n1456 a_400_38200# 0.13fF
C1650 VN.t369 a_400_38200# 0.02fF
C1651 VN.n1457 a_400_38200# 0.15fF
C1652 VN.t132 a_400_38200# 0.02fF
C1653 VN.n1459 a_400_38200# 0.26fF
C1654 VN.n1460 a_400_38200# 0.39fF
C1655 VN.n1461 a_400_38200# 0.66fF
C1656 VN.n1462 a_400_38200# 2.70fF
C1657 VN.n1463 a_400_38200# 2.14fF
C1658 VN.t285 a_400_38200# 0.03fF
C1659 VN.n1464 a_400_38200# 0.26fF
C1660 VN.n1465 a_400_38200# 1.00fF
C1661 VN.n1466 a_400_38200# 0.05fF
C1662 VN.t107 a_400_38200# 0.03fF
C1663 VN.n1467 a_400_38200# 0.13fF
C1664 VN.n1468 a_400_38200# 0.16fF
C1665 VN.n1470 a_400_38200# 0.71fF
C1666 VN.n1471 a_400_38200# 0.27fF
C1667 VN.n1472 a_400_38200# 0.39fF
C1668 VN.n1473 a_400_38200# 0.48fF
C1669 VN.n1474 a_400_38200# 1.84fF
C1670 VN.n1475 a_400_38200# 0.52fF
C1671 VN.n1476 a_400_38200# 0.49fF
C1672 VN.n1477 a_400_38200# 2.01fF
C1673 VN.n1478 a_400_38200# 0.13fF
C1674 VN.t6 a_400_38200# 0.02fF
C1675 VN.n1479 a_400_38200# 0.15fF
C1676 VN.t326 a_400_38200# 0.02fF
C1677 VN.n1481 a_400_38200# 0.26fF
C1678 VN.n1482 a_400_38200# 0.39fF
C1679 VN.n1483 a_400_38200# 0.66fF
C1680 VN.n1484 a_400_38200# 0.05fF
C1681 VN.n1485 a_400_38200# 0.19fF
C1682 VN.n1486 a_400_38200# 1.72fF
C1683 VN.n1487 a_400_38200# 0.13fF
C1684 VN.n1488 a_400_38200# 0.28fF
C1685 VN.n1489 a_400_38200# 0.87fF
C1686 VN.n1490 a_400_38200# 0.03fF
C1687 VN.n1491 a_400_38200# 0.02fF
C1688 VN.n1492 a_400_38200# 0.01fF
C1689 VN.n1493 a_400_38200# 0.02fF
C1690 VN.n1494 a_400_38200# 0.03fF
C1691 VN.n1495 a_400_38200# 0.10fF
C1692 VN.n1496 a_400_38200# 0.07fF
C1693 VN.n1497 a_400_38200# 0.28fF
C1694 VN.n1498 a_400_38200# 0.13fF
C1695 VN.n1499 a_400_38200# 2.12fF
C1696 VN.t186 a_400_38200# 0.03fF
C1697 VN.n1500 a_400_38200# 0.26fF
C1698 VN.n1501 a_400_38200# 1.00fF
C1699 VN.n1502 a_400_38200# 0.05fF
C1700 VN.t341 a_400_38200# 0.03fF
C1701 VN.n1503 a_400_38200# 0.13fF
C1702 VN.n1504 a_400_38200# 0.16fF
C1703 VN.n1506 a_400_38200# 0.04fF
C1704 VN.n1507 a_400_38200# 0.03fF
C1705 VN.n1508 a_400_38200# 0.11fF
C1706 VN.n1509 a_400_38200# 0.27fF
C1707 VN.n1510 a_400_38200# 0.80fF
C1708 VN.n1511 a_400_38200# 0.16fF
C1709 VN.n1512 a_400_38200# 0.12fF
C1710 VN.n1513 a_400_38200# 0.13fF
C1711 VN.n1514 a_400_38200# 0.03fF
C1712 VN.n1515 a_400_38200# 0.08fF
C1713 VN.n1516 a_400_38200# 1.53fF
C1714 VN.n1517 a_400_38200# 0.05fF
C1715 VN.n1518 a_400_38200# 0.53fF
C1716 VN.n1519 a_400_38200# 0.41fF
C1717 VN.n1520 a_400_38200# 1.04fF
C1718 VN.n1521 a_400_38200# 0.37fF
C1719 VN.n1522 a_400_38200# 0.36fF
C1720 VN.n1523 a_400_38200# 5.87fF
C1721 VN.n1524 a_400_38200# 2.37fF
C1722 VN.t147 a_400_38200# 0.02fF
C1723 VN.n1525 a_400_38200# 1.42fF
C1724 VN.n1526 a_400_38200# 29.32fF
C1725 VN.n1527 a_400_38200# 2.42fF
C1726 VN.n1528 a_400_38200# 0.39fF
C1727 VN.n1529 a_400_38200# 0.68fF
C1728 VN.n1530 a_400_38200# 0.57fF
C1729 VN.n1531 a_400_38200# 4.00fF
C1730 VN.n1532 a_400_38200# 33.98fF
C1731 VN.n1533 a_400_38200# 53.30fF
C1732 VN.n1534 a_400_38200# 33.98fF
C1733 VN.n1535 a_400_38200# 53.30fF
C1734 VN.n1536 a_400_38200# 4.64fF
C1735 VN.n1537 a_400_38200# 4.61fF
C1736 VN.n1538 a_400_38200# 4.69fF
C1737 VN.n1539 a_400_38200# 4.67fF
C1738 VN.n1540 a_400_38200# 5.13fF
C1739 VN.n1541 a_400_38200# 53.06fF
C1740 VN.n1542 a_400_38200# 2.40fF
C1741 VN.n1543 a_400_38200# 13.88fF
C1742 VN.n1544 a_400_38200# 2.07fF
C1743 VN.n1545 a_400_38200# 9.82fF
C1744 VN.n1546 a_400_38200# 0.27fF
C1745 VN.t350 a_400_38200# 0.02fF
C1746 VN.n1547 a_400_38200# 0.48fF
C1747 VN.n1548 a_400_38200# 5.96fF
C1748 VN.n1549 a_400_38200# 2.00fF
C1749 VN.n1550 a_400_38200# 3.56fF
C1750 VN.n1551 a_400_38200# 0.34fF
C1751 VN.n1552 a_400_38200# 1.09fF
C1752 VN.t226 a_400_38200# 0.02fF
C1753 VN.n1553 a_400_38200# 0.97fF
C1754 VN.t256 a_400_38200# 0.03fF
C1755 VN.n1554 a_400_38200# 0.98fF
C1756 VN.n1555 a_400_38200# 0.02fF
C1757 VN.t388 a_400_38200# 0.02fF
C1758 VN.n1556 a_400_38200# 0.40fF
C1759 VN.n1557 a_400_38200# 33.98fF
C1760 VN.n1558 a_400_38200# 33.98fF
C1761 VN.n1559 a_400_38200# 5.75fF
C1762 VN.n1560 a_400_38200# 2.01fF
C1763 VN.t357 a_400_38200# 0.02fF
C1764 VN.n1561 a_400_38200# 0.97fF
C1765 VN.t384 a_400_38200# 0.03fF
C1766 VN.n1562 a_400_38200# 0.98fF
C1767 VN.n1563 a_400_38200# 3.57fF
C1768 VN.n1564 a_400_38200# 0.27fF
C1769 VN.n1565 a_400_38200# 1.15fF
C1770 VN.n1566 a_400_38200# 0.49fF
C1771 VN.n1567 a_400_38200# 0.02fF
C1772 VN.t153 a_400_38200# 0.02fF
C1773 VN.n1568 a_400_38200# 0.40fF
C1774 VN.n1569 a_400_38200# 0.40fF
C1775 VN.n1570 a_400_38200# 0.90fF
C1776 VN.t235 a_400_38200# 0.02fF
C1777 VN.n1571 a_400_38200# 0.97fF
C1778 VN.t262 a_400_38200# 0.03fF
C1779 VN.n1572 a_400_38200# 0.98fF
C1780 VN.n1573 a_400_38200# 33.98fF
C1781 VN.n1574 a_400_38200# 33.98fF
C1782 VN.n1575 a_400_38200# 6.27fF
C1783 VN.n1576 a_400_38200# 1.94fF
C1784 VN.n1577 a_400_38200# 1.24fF
C1785 VN.n1578 a_400_38200# 0.00fF
C1786 VN.n1579 a_400_38200# 0.43fF
C1787 VN.n1580 a_400_38200# 0.02fF
C1788 VN.t1 a_400_38200# 0.02fF
C1789 VN.n1581 a_400_38200# 0.40fF
C1790 VN.n1582 a_400_38200# 33.98fF
C1791 VN.n1583 a_400_38200# 33.98fF
C1792 VN.n1584 a_400_38200# 6.05fF
C1793 VN.n1585 a_400_38200# 1.96fF
C1794 VN.t110 a_400_38200# 0.02fF
C1795 VN.n1586 a_400_38200# 0.97fF
C1796 VN.t137 a_400_38200# 0.03fF
C1797 VN.n1587 a_400_38200# 0.98fF
C1798 VN.n1588 a_400_38200# 1.65fF
C1799 VN.n1589 a_400_38200# 0.02fF
C1800 VN.t269 a_400_38200# 0.02fF
C1801 VN.n1590 a_400_38200# 0.40fF
C1802 VN.n1591 a_400_38200# 110.74fF
C1803 VN.n1592 a_400_38200# 110.74fF
C1804 VN.n1593 a_400_38200# 6.31fF
C1805 VN.n1594 a_400_38200# 2.14fF
C1806 VN.t364 a_400_38200# 0.02fF
C1807 VN.n1595 a_400_38200# 0.97fF
C1808 VN.t373 a_400_38200# 0.03fF
C1809 VN.n1596 a_400_38200# 0.98fF
C1810 VN.n1597 a_400_38200# 3.57fF
C1811 VN.n1598 a_400_38200# 1.77fF
C1812 VN.n1599 a_400_38200# 0.02fF
C1813 VN.t143 a_400_38200# 0.02fF
C1814 VN.n1600 a_400_38200# 0.40fF
C1815 VN.t128 a_400_38200# 0.03fF
C1816 VN.n1601 a_400_38200# 0.98fF
C1817 VN.n1602 a_400_38200# 0.02fF
C1818 VN.t265 a_400_38200# 0.02fF
C1819 VN.n1603 a_400_38200# 0.40fF
C1820 VN.t101 a_400_38200# 0.02fF
C1821 VN.n1604 a_400_38200# 0.97fF
C1822 VN.t100 a_400_38200# 53.69fF
C1823 VN.n1605 a_400_38200# 2.87fF
C1824 VN.n1606 a_400_38200# 1.63fF
C1825 VN.n1607 a_400_38200# 0.13fF
C1826 VN.t270 a_400_38200# 0.02fF
C1827 VN.n1608 a_400_38200# 0.15fF
C1828 VN.t200 a_400_38200# 0.02fF
C1829 VN.n1610 a_400_38200# 0.26fF
C1830 VN.n1611 a_400_38200# 0.39fF
C1831 VN.n1612 a_400_38200# 0.66fF
C1832 VN.n1613 a_400_38200# 0.38fF
C1833 VN.n1614 a_400_38200# 0.59fF
C1834 VN.n1615 a_400_38200# 0.42fF
C1835 VN.n1616 a_400_38200# 0.19fF
C1836 VN.n1617 a_400_38200# 0.27fF
C1837 VN.n1618 a_400_38200# 0.10fF
C1838 VN.n1619 a_400_38200# 2.14fF
C1839 VN.t57 a_400_38200# 0.03fF
C1840 VN.n1620 a_400_38200# 0.26fF
C1841 VN.n1621 a_400_38200# 1.00fF
C1842 VN.n1622 a_400_38200# 0.05fF
C1843 VN.t368 a_400_38200# 0.03fF
C1844 VN.n1623 a_400_38200# 0.13fF
C1845 VN.n1624 a_400_38200# 0.16fF
C1846 VN.n1626 a_400_38200# 0.27fF
C1847 VN.n1627 a_400_38200# 0.10fF
C1848 VN.n1628 a_400_38200# 0.23fF
C1849 VN.n1629 a_400_38200# 1.89fF
C1850 VN.n1630 a_400_38200# 0.48fF
C1851 VN.n1631 a_400_38200# 2.87fF
C1852 VN.n1632 a_400_38200# 1.63fF
C1853 VN.n1633 a_400_38200# 0.13fF
C1854 VN.t145 a_400_38200# 0.02fF
C1855 VN.n1634 a_400_38200# 0.15fF
C1856 VN.t67 a_400_38200# 0.02fF
C1857 VN.n1636 a_400_38200# 0.26fF
C1858 VN.n1637 a_400_38200# 0.39fF
C1859 VN.n1638 a_400_38200# 0.66fF
C1860 VN.n1639 a_400_38200# 0.97fF
C1861 VN.n1640 a_400_38200# 3.34fF
C1862 VN.n1641 a_400_38200# 2.62fF
C1863 VN.t299 a_400_38200# 0.03fF
C1864 VN.n1642 a_400_38200# 0.26fF
C1865 VN.n1643 a_400_38200# 1.00fF
C1866 VN.n1644 a_400_38200# 0.05fF
C1867 VN.t247 a_400_38200# 0.03fF
C1868 VN.n1645 a_400_38200# 0.13fF
C1869 VN.n1646 a_400_38200# 0.16fF
C1870 VN.n1648 a_400_38200# 0.21fF
C1871 VN.n1649 a_400_38200# 0.10fF
C1872 VN.n1650 a_400_38200# 0.74fF
C1873 VN.n1651 a_400_38200# 0.30fF
C1874 VN.n1652 a_400_38200# 1.90fF
C1875 VN.n1653 a_400_38200# 0.23fF
C1876 VN.n1654 a_400_38200# 2.01fF
C1877 VN.n1655 a_400_38200# 0.13fF
C1878 VN.t386 a_400_38200# 0.02fF
C1879 VN.n1656 a_400_38200# 0.15fF
C1880 VN.t313 a_400_38200# 0.02fF
C1881 VN.n1658 a_400_38200# 0.26fF
C1882 VN.n1659 a_400_38200# 0.39fF
C1883 VN.n1660 a_400_38200# 0.66fF
C1884 VN.n1661 a_400_38200# 2.72fF
C1885 VN.n1662 a_400_38200# 2.03fF
C1886 VN.t171 a_400_38200# 0.03fF
C1887 VN.n1663 a_400_38200# 0.26fF
C1888 VN.n1664 a_400_38200# 1.00fF
C1889 VN.n1665 a_400_38200# 0.05fF
C1890 VN.t121 a_400_38200# 0.03fF
C1891 VN.n1666 a_400_38200# 0.13fF
C1892 VN.n1667 a_400_38200# 0.16fF
C1893 VN.t0 a_400_38200# 11.11fF
C1894 VN.n1669 a_400_38200# 9.61fF
C1895 VN.n1670 a_400_38200# 0.07fF
C1896 VN.n1671 a_400_38200# 0.22fF
C1897 VN.n1672 a_400_38200# 0.10fF
C1898 VN.n1673 a_400_38200# 0.23fF
C1899 VN.n1674 a_400_38200# 0.10fF
C1900 VN.n1675 a_400_38200# 0.33fF
C1901 VN.n1676 a_400_38200# 1.11fF
C1902 VN.n1677 a_400_38200# 0.49fF
C1903 VN.n1678 a_400_38200# 1.83fF
C1904 VN.n1679 a_400_38200# 0.13fF
C1905 VN.t134 a_400_38200# 0.02fF
C1906 VN.n1680 a_400_38200# 0.15fF
C1907 VN.t239 a_400_38200# 0.02fF
C1908 VN.n1682 a_400_38200# 0.26fF
C1909 VN.n1683 a_400_38200# 0.39fF
C1910 VN.n1684 a_400_38200# 0.66fF
C1911 VN.n1685 a_400_38200# 0.39fF
C1912 VN.n1686 a_400_38200# 0.44fF
C1913 VN.n1687 a_400_38200# 0.74fF
C1914 VN.n1688 a_400_38200# 0.43fF
C1915 VN.n1689 a_400_38200# 0.48fF
C1916 VN.n1690 a_400_38200# 0.27fF
C1917 VN.n1691 a_400_38200# 0.20fF
C1918 VN.n1692 a_400_38200# 0.10fF
C1919 VN.n1693 a_400_38200# 1.86fF
C1920 VN.t233 a_400_38200# 0.03fF
C1921 VN.n1694 a_400_38200# 0.13fF
C1922 VN.n1695 a_400_38200# 0.16fF
C1923 VN.t4 a_400_38200# 0.03fF
C1924 VN.n1697 a_400_38200# 0.26fF
C1925 VN.n1698 a_400_38200# 1.00fF
C1926 VN.n1699 a_400_38200# 0.05fF
C1927 VN.t5 a_400_38200# 21.10fF
C1928 VN.t379 a_400_38200# 0.03fF
C1929 VN.n1700 a_400_38200# 0.01fF
C1930 VN.n1701 a_400_38200# 0.28fF
C1931 VN.t32 a_400_38200# 0.03fF
C1932 VN.n1703 a_400_38200# 1.30fF
C1933 VN.n1704 a_400_38200# 0.05fF
C1934 VN.t187 a_400_38200# 0.02fF
C1935 VN.n1705 a_400_38200# 0.70fF
C1936 VN.n1706 a_400_38200# 0.66fF
C1937 VN.n1707 a_400_38200# 118.17fF
C1938 VN.n1708 a_400_38200# 0.23fF
C1939 VN.n1709 a_400_38200# 1.54fF
C1940 VN.n1710 a_400_38200# 0.65fF
C1941 VN.n1711 a_400_38200# 0.24fF
C1942 VN.n1712 a_400_38200# 0.96fF
C1943 VN.n1713 a_400_38200# 0.96fF
C1944 VN.n1714 a_400_38200# 2.08fF
C1945 VN.n1715 a_400_38200# 0.31fF
C1946 VN.t24 a_400_38200# 9.89fF
C1947 VN.n1716 a_400_38200# 12.19fF
C1948 VN.n1717 a_400_38200# 118.17fF
C1949 VN.n1718 a_400_38200# 4.63fF
C1950 VN.n1719 a_400_38200# 1.24fF
C1951 VN.n1720 a_400_38200# 1.96fF
C1952 VN.n1721 a_400_38200# 4.64fF
C1953 VN.n1722 a_400_38200# 57.57fF
C1954 VN.n1723 a_400_38200# 34.49fF
C1955 VN.n1724 a_400_38200# 34.49fF
C1956 VN.n1725 a_400_38200# 34.49fF
C1957 VN.n1726 a_400_38200# 34.49fF
C1958 VN.n1727 a_400_38200# 109.50fF
C1959 VN.n1728 a_400_38200# 118.26fF
C1960 VN.n1729 a_400_38200# 30.94fF
C1961 VN.n1730 a_400_38200# 30.87fF
C1962 VN.n1731 a_400_38200# 30.87fF
C1963 VN.n1732 a_400_38200# 0.65fF
C1964 VN.n1733 a_400_38200# 0.24fF
C1965 VN.n1734 a_400_38200# 0.65fF
C1966 VN.n1735 a_400_38200# 2.08fF
C1967 VN.n1736 a_400_38200# 0.31fF
C1968 VN.t9 a_400_38200# 9.89fF
C1969 VN.n1737 a_400_38200# 12.19fF
C1970 VN.n1738 a_400_38200# 0.84fF
C1971 VN.n1739 a_400_38200# 0.30fF
C1972 VN.n1740 a_400_38200# 4.65fF
C1973 VN.n1741 a_400_38200# 3.06fF
C1974 VN.n1742 a_400_38200# 2.06fF
C1975 VN.n1743 a_400_38200# 0.06fF
C1976 VN.n1744 a_400_38200# 0.03fF
C1977 VN.n1745 a_400_38200# 0.04fF
C1978 VN.n1746 a_400_38200# 1.08fF
C1979 VN.n1747 a_400_38200# 0.02fF
C1980 VN.n1748 a_400_38200# 0.01fF
C1981 VN.n1749 a_400_38200# 0.02fF
C1982 VN.n1750 a_400_38200# 0.09fF
C1983 VN.n1751 a_400_38200# 0.39fF
C1984 VN.n1752 a_400_38200# 2.02fF
C1985 VN.t10 a_400_38200# 0.02fF
C1986 VN.n1753 a_400_38200# 0.26fF
C1987 VN.n1754 a_400_38200# 0.39fF
C1988 VN.n1755 a_400_38200# 0.66fF
C1989 VN.n1756 a_400_38200# 0.13fF
C1990 VN.t238 a_400_38200# 0.02fF
C1991 VN.n1757 a_400_38200# 0.15fF
C1992 VN.n1759 a_400_38200# 0.76fF
C1993 VN.n1760 a_400_38200# 0.25fF
C1994 VN.n1761 a_400_38200# 0.28fF
C1995 VN.n1762 a_400_38200# 0.10fF
C1996 VN.n1763 a_400_38200# 0.25fF
C1997 VN.n1764 a_400_38200# 0.76fF
C1998 VN.n1765 a_400_38200# 1.26fF
C1999 VN.n1766 a_400_38200# 0.24fF
C2000 VN.n1767 a_400_38200# 0.28fF
C2001 VN.n1768 a_400_38200# 0.10fF
C2002 VN.n1769 a_400_38200# 2.06fF
C2003 VN.t197 a_400_38200# 0.03fF
C2004 VN.n1770 a_400_38200# 0.26fF
C2005 VN.n1771 a_400_38200# 1.00fF
C2006 VN.n1772 a_400_38200# 0.05fF
C2007 VN.t335 a_400_38200# 0.03fF
C2008 VN.n1773 a_400_38200# 0.13fF
C2009 VN.n1774 a_400_38200# 0.16fF
C2010 VN.n1776 a_400_38200# 9.61fF
C2011 VN.n1777 a_400_38200# 0.10fF
C2012 VN.n1778 a_400_38200# 0.23fF
C2013 VN.n1779 a_400_38200# 0.07fF
C2014 VN.n1780 a_400_38200# 0.06fF
C2015 VN.n1781 a_400_38200# 0.07fF
C2016 VN.n1782 a_400_38200# 0.20fF
C2017 VN.n1783 a_400_38200# 0.21fF
C2018 VN.n1784 a_400_38200# 1.13fF
C2019 VN.n1785 a_400_38200# 0.59fF
C2020 VN.n1786 a_400_38200# 2.55fF
C2021 VN.n1787 a_400_38200# 0.13fF
C2022 VN.t362 a_400_38200# 0.02fF
C2023 VN.n1788 a_400_38200# 0.15fF
C2024 VN.t142 a_400_38200# 0.02fF
C2025 VN.n1790 a_400_38200# 0.26fF
C2026 VN.n1791 a_400_38200# 0.39fF
C2027 VN.n1792 a_400_38200# 0.66fF
C2028 VN.n1793 a_400_38200# 0.78fF
C2029 VN.n1794 a_400_38200# 1.88fF
C2030 VN.n1795 a_400_38200# 2.66fF
C2031 VN.t96 a_400_38200# 0.03fF
C2032 VN.n1796 a_400_38200# 0.13fF
C2033 VN.n1797 a_400_38200# 0.16fF
C2034 VN.t305 a_400_38200# 0.03fF
C2035 VN.n1799 a_400_38200# 0.26fF
C2036 VN.n1800 a_400_38200# 1.00fF
C2037 VN.n1801 a_400_38200# 0.05fF
C2038 VN.n1802 a_400_38200# 2.05fF
C2039 VN.n1803 a_400_38200# 0.13fF
C2040 VN.t333 a_400_38200# 0.02fF
C2041 VN.n1804 a_400_38200# 0.15fF
C2042 VN.t135 a_400_38200# 0.02fF
C2043 VN.n1806 a_400_38200# 0.26fF
C2044 VN.n1807 a_400_38200# 0.39fF
C2045 VN.n1808 a_400_38200# 0.66fF
C2046 VN.n1809 a_400_38200# 1.01fF
C2047 VN.n1810 a_400_38200# 0.35fF
C2048 VN.n1811 a_400_38200# 0.35fF
C2049 VN.n1812 a_400_38200# 1.01fF
C2050 VN.n1813 a_400_38200# 1.19fF
C2051 VN.n1814 a_400_38200# 0.17fF
C2052 VN.n1815 a_400_38200# 5.41fF
C2053 VN.t209 a_400_38200# 0.03fF
C2054 VN.n1816 a_400_38200# 0.13fF
C2055 VN.n1817 a_400_38200# 0.16fF
C2056 VN.t360 a_400_38200# 0.03fF
C2057 VN.n1819 a_400_38200# 0.26fF
C2058 VN.n1820 a_400_38200# 1.00fF
C2059 VN.n1821 a_400_38200# 0.05fF
C2060 VN.n1822 a_400_38200# 2.05fF
C2061 VN.n1823 a_400_38200# 2.91fF
C2062 VN.t370 a_400_38200# 0.02fF
C2063 VN.n1824 a_400_38200# 0.26fF
C2064 VN.n1825 a_400_38200# 0.39fF
C2065 VN.n1826 a_400_38200# 0.66fF
C2066 VN.n1827 a_400_38200# 0.13fF
C2067 VN.t207 a_400_38200# 0.02fF
C2068 VN.n1828 a_400_38200# 0.15fF
C2069 VN.n1830 a_400_38200# 5.63fF
C2070 VN.t302 a_400_38200# 0.03fF
C2071 VN.n1831 a_400_38200# 0.13fF
C2072 VN.n1832 a_400_38200# 0.16fF
C2073 VN.t236 a_400_38200# 0.03fF
C2074 VN.n1834 a_400_38200# 0.26fF
C2075 VN.n1835 a_400_38200# 1.00fF
C2076 VN.n1836 a_400_38200# 0.05fF
C2077 VN.n1837 a_400_38200# 2.05fF
C2078 VN.n1838 a_400_38200# 2.91fF
C2079 VN.t248 a_400_38200# 0.02fF
C2080 VN.n1839 a_400_38200# 0.26fF
C2081 VN.n1840 a_400_38200# 0.39fF
C2082 VN.n1841 a_400_38200# 0.66fF
C2083 VN.n1842 a_400_38200# 0.13fF
C2084 VN.t78 a_400_38200# 0.02fF
C2085 VN.n1843 a_400_38200# 0.15fF
C2086 VN.n1845 a_400_38200# 2.05fF
C2087 VN.n1846 a_400_38200# 2.92fF
C2088 VN.t79 a_400_38200# 0.02fF
C2089 VN.n1847 a_400_38200# 0.26fF
C2090 VN.n1848 a_400_38200# 0.39fF
C2091 VN.n1849 a_400_38200# 0.66fF
C2092 VN.t46 a_400_38200# 0.02fF
C2093 VN.n1850 a_400_38200# 1.33fF
C2094 VN.n1851 a_400_38200# 0.46fF
C2095 VN.n1852 a_400_38200# 0.48fF
C2096 VN.n1853 a_400_38200# 0.40fF
C2097 VN.n1854 a_400_38200# 0.23fF
C2098 VN.n1855 a_400_38200# 0.27fF
C2099 VN.n1856 a_400_38200# 1.40fF
C2100 VN.n1857 a_400_38200# 0.39fF
C2101 VN.n1858 a_400_38200# 0.69fF
C2102 VN.n1859 a_400_38200# 1.26fF
C2103 VN.n1860 a_400_38200# 1.65fF
C2104 VN.n1861 a_400_38200# 0.65fF
C2105 VN.n1862 a_400_38200# 0.02fF
C2106 VN.n1863 a_400_38200# 1.06fF
C2107 VN.t45 a_400_38200# 9.89fF
C2108 VN.n1864 a_400_38200# 10.65fF
C2109 VN.n1866 a_400_38200# 0.41fF
C2110 VN.n1867 a_400_38200# 0.25fF
C2111 VN.n1868 a_400_38200# 3.08fF
C2112 VN.n1869 a_400_38200# 2.18fF
C2113 VN.n1870 a_400_38200# 4.45fF
C2114 VN.n1871 a_400_38200# 0.27fF
C2115 VN.n1872 a_400_38200# 0.01fF
C2116 VN.t260 a_400_38200# 0.02fF
C2117 VN.n1873 a_400_38200# 0.28fF
C2118 VN.t300 a_400_38200# 0.03fF
C2119 VN.n1874 a_400_38200# 1.04fF
C2120 VN.n1875 a_400_38200# 0.77fF
C2121 VN.n1876 a_400_38200# 0.85fF
C2122 VN.n1877 a_400_38200# 2.47fF
C2123 VN.n1878 a_400_38200# 2.05fF
C2124 VN.n1879 a_400_38200# 0.13fF
C2125 VN.t133 a_400_38200# 0.02fF
C2126 VN.n1880 a_400_38200# 0.15fF
C2127 VN.t291 a_400_38200# 0.02fF
C2128 VN.n1882 a_400_38200# 0.26fF
C2129 VN.n1883 a_400_38200# 0.39fF
C2130 VN.n1884 a_400_38200# 0.66fF
C2131 VN.n1885 a_400_38200# 1.51fF
C2132 VN.n1886 a_400_38200# 1.24fF
C2133 VN.n1887 a_400_38200# 0.38fF
C2134 VN.n1888 a_400_38200# 2.21fF
C2135 VN.t172 a_400_38200# 0.03fF
C2136 VN.n1889 a_400_38200# 0.26fF
C2137 VN.n1890 a_400_38200# 1.00fF
C2138 VN.n1891 a_400_38200# 0.05fF
C2139 VN.t154 a_400_38200# 0.03fF
C2140 VN.n1892 a_400_38200# 0.13fF
C2141 VN.n1893 a_400_38200# 0.16fF
C2142 VN.n1895 a_400_38200# 2.06fF
C2143 VN.n1896 a_400_38200# 2.05fF
C2144 VN.t160 a_400_38200# 0.02fF
C2145 VN.n1897 a_400_38200# 0.26fF
C2146 VN.n1898 a_400_38200# 0.39fF
C2147 VN.n1899 a_400_38200# 0.66fF
C2148 VN.n1900 a_400_38200# 0.13fF
C2149 VN.t367 a_400_38200# 0.02fF
C2150 VN.n1901 a_400_38200# 0.15fF
C2151 VN.n1903 a_400_38200# 1.26fF
C2152 VN.n1904 a_400_38200# 0.24fF
C2153 VN.n1905 a_400_38200# 2.06fF
C2154 VN.t34 a_400_38200# 0.03fF
C2155 VN.n1906 a_400_38200# 0.26fF
C2156 VN.n1907 a_400_38200# 1.00fF
C2157 VN.n1908 a_400_38200# 0.05fF
C2158 VN.t3 a_400_38200# 0.03fF
C2159 VN.n1909 a_400_38200# 0.13fF
C2160 VN.n1910 a_400_38200# 0.16fF
C2161 VN.n1912 a_400_38200# 9.61fF
C2162 VN.n1913 a_400_38200# 3.21fF
C2163 VN.n1914 a_400_38200# 2.05fF
C2164 VN.n1915 a_400_38200# 0.13fF
C2165 VN.t158 a_400_38200# 0.02fF
C2166 VN.n1916 a_400_38200# 0.15fF
C2167 VN.t334 a_400_38200# 0.02fF
C2168 VN.n1918 a_400_38200# 0.26fF
C2169 VN.n1919 a_400_38200# 0.39fF
C2170 VN.n1920 a_400_38200# 0.66fF
C2171 VN.n1921 a_400_38200# 1.19fF
C2172 VN.n1922 a_400_38200# 0.17fF
C2173 VN.n1923 a_400_38200# 2.29fF
C2174 VN.t193 a_400_38200# 0.03fF
C2175 VN.n1924 a_400_38200# 0.13fF
C2176 VN.n1925 a_400_38200# 0.16fF
C2177 VN.t229 a_400_38200# 0.03fF
C2178 VN.n1927 a_400_38200# 0.26fF
C2179 VN.n1928 a_400_38200# 1.00fF
C2180 VN.n1929 a_400_38200# 0.05fF
C2181 VN.n1930 a_400_38200# 2.05fF
C2182 VN.n1931 a_400_38200# 2.91fF
C2183 VN.t208 a_400_38200# 0.02fF
C2184 VN.n1932 a_400_38200# 0.26fF
C2185 VN.n1933 a_400_38200# 0.39fF
C2186 VN.n1934 a_400_38200# 0.66fF
C2187 VN.n1935 a_400_38200# 0.13fF
C2188 VN.t19 a_400_38200# 0.02fF
C2189 VN.n1936 a_400_38200# 0.15fF
C2190 VN.n1938 a_400_38200# 3.21fF
C2191 VN.n1939 a_400_38200# 2.51fF
C2192 VN.t65 a_400_38200# 0.03fF
C2193 VN.n1940 a_400_38200# 0.13fF
C2194 VN.n1941 a_400_38200# 0.16fF
C2195 VN.t103 a_400_38200# 0.03fF
C2196 VN.n1943 a_400_38200# 0.26fF
C2197 VN.n1944 a_400_38200# 1.00fF
C2198 VN.n1945 a_400_38200# 0.05fF
C2199 VN.n1946 a_400_38200# 0.13fF
C2200 VN.t166 a_400_38200# 0.02fF
C2201 VN.n1947 a_400_38200# 0.15fF
C2202 VN.t321 a_400_38200# 0.02fF
C2203 VN.n1949 a_400_38200# 0.26fF
C2204 VN.n1950 a_400_38200# 0.39fF
C2205 VN.n1951 a_400_38200# 0.66fF
C2206 VN.n1952 a_400_38200# 1.74fF
C2207 VN.n1953 a_400_38200# 0.15fF
C2208 VN.n1954 a_400_38200# 0.63fF
C2209 VN.n1955 a_400_38200# 0.58fF
C2210 VN.n1956 a_400_38200# 0.45fF
C2211 VN.n1957 a_400_38200# 0.27fF
C2212 VN.n1958 a_400_38200# 0.27fF
C2213 VN.n1959 a_400_38200# 0.74fF
C2214 VN.n1960 a_400_38200# 2.15fF
C2215 VN.t179 a_400_38200# 0.03fF
C2216 VN.n1961 a_400_38200# 0.13fF
C2217 VN.n1962 a_400_38200# 0.16fF
C2218 VN.t217 a_400_38200# 0.03fF
C2219 VN.n1964 a_400_38200# 0.26fF
C2220 VN.n1965 a_400_38200# 1.00fF
C2221 VN.n1966 a_400_38200# 0.05fF
C2222 VN.t2 a_400_38200# 21.51fF
C2223 VN.t339 a_400_38200# 0.03fF
C2224 VN.n1967 a_400_38200# 0.26fF
C2225 VN.n1968 a_400_38200# 1.00fF
C2226 VN.n1969 a_400_38200# 0.05fF
C2227 VN.t307 a_400_38200# 0.03fF
C2228 VN.n1970 a_400_38200# 0.13fF
C2229 VN.n1971 a_400_38200# 0.16fF
C2230 VN.n1973 a_400_38200# 0.13fF
C2231 VN.t275 a_400_38200# 0.02fF
C2232 VN.n1974 a_400_38200# 0.15fF
C2233 VN.n1976 a_400_38200# 5.64fF
C2234 VN.n1977 a_400_38200# 5.34fF
C2235 VN.t174 a_400_38200# 0.03fF
C2236 VN.n1978 a_400_38200# 0.13fF
C2237 VN.n1979 a_400_38200# 0.16fF
C2238 VN.t112 a_400_38200# 0.03fF
C2239 VN.n1981 a_400_38200# 0.26fF
C2240 VN.n1982 a_400_38200# 1.00fF
C2241 VN.n1983 a_400_38200# 0.05fF
C2242 VN.n1984 a_400_38200# 0.03fF
C2243 VN.n1985 a_400_38200# 0.13fF
C2244 VN.n1986 a_400_38200# 0.12fF
C2245 VN.n1987 a_400_38200# 0.39fF
C2246 VN.n1988 a_400_38200# 0.51fF
C2247 VN.n1989 a_400_38200# 1.24fF
C2248 VN.n1990 a_400_38200# 2.04fF
C2249 VN.n1991 a_400_38200# 0.13fF
C2250 VN.t320 a_400_38200# 0.02fF
C2251 VN.n1992 a_400_38200# 0.15fF
C2252 VN.t123 a_400_38200# 0.02fF
C2253 VN.n1994 a_400_38200# 0.26fF
C2254 VN.n1995 a_400_38200# 0.39fF
C2255 VN.n1996 a_400_38200# 0.66fF
C2256 VN.n1997 a_400_38200# 1.38fF
C2257 VN.n1998 a_400_38200# 2.60fF
C2258 VN.n1999 a_400_38200# 4.59fF
C2259 VN.t40 a_400_38200# 0.03fF
C2260 VN.n2000 a_400_38200# 0.13fF
C2261 VN.n2001 a_400_38200# 0.16fF
C2262 VN.t347 a_400_38200# 0.03fF
C2263 VN.n2003 a_400_38200# 0.26fF
C2264 VN.n2004 a_400_38200# 1.00fF
C2265 VN.n2005 a_400_38200# 0.05fF
C2266 VN.t39 a_400_38200# 21.10fF
C2267 VN.t310 a_400_38200# 0.03fF
C2268 VN.n2006 a_400_38200# 0.01fF
C2269 VN.n2007 a_400_38200# 0.28fF
C2270 VN.t224 a_400_38200# 0.03fF
C2271 VN.n2009 a_400_38200# 1.30fF
C2272 VN.n2010 a_400_38200# 0.05fF
C2273 VN.t361 a_400_38200# 0.02fF
C2274 VN.n2011 a_400_38200# 0.70fF
C2275 VN.n2012 a_400_38200# 0.66fF
C2276 VN.n2013 a_400_38200# 1.64fF
C2277 VN.n2014 a_400_38200# 0.02fF
C2278 VN.n2015 a_400_38200# 0.01fF
C2279 VN.n2016 a_400_38200# 0.01fF
C2280 VN.n2017 a_400_38200# 0.01fF
C2281 VN.n2018 a_400_38200# 0.02fF
C2282 VN.n2019 a_400_38200# 0.03fF
C2283 VN.n2020 a_400_38200# 0.03fF
C2284 VN.n2021 a_400_38200# 0.04fF
C2285 VN.n2022 a_400_38200# 0.18fF
C2286 VN.n2023 a_400_38200# 0.11fF
C2287 VN.n2024 a_400_38200# 0.18fF
C2288 VN.n2025 a_400_38200# 0.16fF
C2289 VN.n2026 a_400_38200# 0.30fF
C2290 VN.n2027 a_400_38200# 0.27fF
C2291 VN.n2028 a_400_38200# 5.12fF
C2292 VN.n2029 a_400_38200# 30.87fF
C2293 VN.n2030 a_400_38200# 28.96fF
C2294 fc2.n0 a_400_38200# 1.13fF
C2295 fc2.n1 a_400_38200# 0.87fF
C2296 fc2.n2 a_400_38200# 0.44fF
C2297 fc2.n3 a_400_38200# 0.15fF
C2298 fc2.t327 a_400_38200# 0.02fF
C2299 fc2.n4 a_400_38200# 1.14fF
C2300 fc2.n5 a_400_38200# 2.82fF
C2301 fc2.n6 a_400_38200# 0.01fF
C2302 fc2.t209 a_400_38200# 0.02fF
C2303 fc2.n7 a_400_38200# 0.32fF
C2304 fc2.n8 a_400_38200# 7.70fF
C2305 fc2.t278 a_400_38200# 0.02fF
C2306 fc2.n9 a_400_38200# 0.39fF
C2307 fc2.n10 a_400_38200# 62.63fF
C2308 fc2.n11 a_400_38200# 3.69fF
C2309 fc2.n12 a_400_38200# 2.70fF
C2310 fc2.n13 a_400_38200# 0.06fF
C2311 fc2.n14 a_400_38200# 0.17fF
C2312 fc2.n15 a_400_38200# 0.98fF
C2313 fc2.n16 a_400_38200# 1.63fF
C2314 fc2.t87 a_400_38200# 0.02fF
C2315 fc2.n17 a_400_38200# 0.78fF
C2316 fc2.t355 a_400_38200# 0.02fF
C2317 fc2.n18 a_400_38200# 0.78fF
C2318 fc2.n19 a_400_38200# 0.01fF
C2319 fc2.t156 a_400_38200# 0.02fF
C2320 fc2.n20 a_400_38200# 0.32fF
C2321 fc2.n21 a_400_38200# 3.95fF
C2322 fc2.n22 a_400_38200# 2.50fF
C2323 fc2.t328 a_400_38200# 0.02fF
C2324 fc2.n23 a_400_38200# 0.78fF
C2325 fc2.t58 a_400_38200# 0.02fF
C2326 fc2.n24 a_400_38200# 0.78fF
C2327 fc2.n25 a_400_38200# 2.39fF
C2328 fc2.n26 a_400_38200# 0.01fF
C2329 fc2.t222 a_400_38200# 0.02fF
C2330 fc2.n27 a_400_38200# 0.32fF
C2331 fc2.n28 a_400_38200# 3.65fF
C2332 fc2.n29 a_400_38200# 2.76fF
C2333 fc2.t300 a_400_38200# 0.02fF
C2334 fc2.n30 a_400_38200# 0.78fF
C2335 fc2.t15 a_400_38200# 0.02fF
C2336 fc2.n31 a_400_38200# 0.78fF
C2337 fc2.n32 a_400_38200# 2.82fF
C2338 fc2.n33 a_400_38200# 0.01fF
C2339 fc2.t100 a_400_38200# 0.02fF
C2340 fc2.n34 a_400_38200# 0.32fF
C2341 fc2.n35 a_400_38200# 4.26fF
C2342 fc2.n36 a_400_38200# 2.61fF
C2343 fc2.t173 a_400_38200# 0.02fF
C2344 fc2.n37 a_400_38200# 0.78fF
C2345 fc2.t269 a_400_38200# 0.02fF
C2346 fc2.n38 a_400_38200# 0.78fF
C2347 fc2.n39 a_400_38200# 1.96fF
C2348 fc2.n40 a_400_38200# 0.01fF
C2349 fc2.t340 a_400_38200# 0.02fF
C2350 fc2.n41 a_400_38200# 0.32fF
C2351 fc2.n42 a_400_38200# 4.26fF
C2352 fc2.n43 a_400_38200# 2.61fF
C2353 fc2.n44 a_400_38200# 1.96fF
C2354 fc2.t30 a_400_38200# 0.02fF
C2355 fc2.n45 a_400_38200# 0.78fF
C2356 fc2.n46 a_400_38200# 0.01fF
C2357 fc2.t86 a_400_38200# 0.02fF
C2358 fc2.n47 a_400_38200# 0.32fF
C2359 fc2.t289 a_400_38200# 0.02fF
C2360 fc2.n48 a_400_38200# 0.78fF
C2361 fc2.t40 a_400_38200# 0.02fF
C2362 fc2.n49 a_400_38200# 0.78fF
C2363 fc2.t146 a_400_38200# 0.02fF
C2364 fc2.n50 a_400_38200# 0.78fF
C2365 fc2.n51 a_400_38200# 3.65fF
C2366 fc2.n52 a_400_38200# 2.76fF
C2367 fc2.t14 a_400_38200# 53.44fF
C2368 fc2.n53 a_400_38200# 0.27fF
C2369 fc2.n54 a_400_38200# 0.15fF
C2370 fc2.n55 a_400_38200# 3.64fF
C2371 fc2.n56 a_400_38200# 0.82fF
C2372 fc2.n57 a_400_38200# 0.24fF
C2373 fc2.n58 a_400_38200# 1.41fF
C2374 fc2.n59 a_400_38200# 0.24fF
C2375 fc2.n60 a_400_38200# 1.41fF
C2376 fc2.n61 a_400_38200# 0.24fF
C2377 fc2.n62 a_400_38200# 1.41fF
C2378 fc2.n63 a_400_38200# 22.09fF
C2379 fc2.n64 a_400_38200# 12.40fF
C2380 fc2.n65 a_400_38200# 12.52fF
C2381 fc2.n66 a_400_38200# 11.42fF
C2382 fc2.n67 a_400_38200# 12.94fF
C2383 fc2.n68 a_400_38200# 11.42fF
C2384 fc2.n69 a_400_38200# 12.94fF
C2385 fc2.n70 a_400_38200# 11.42fF
C2386 fc2.n71 a_400_38200# 12.94fF
C2387 fc2.n72 a_400_38200# 11.91fF
C2388 fc2.n73 a_400_38200# 72.64fF
C2389 fc2.n74 a_400_38200# 368.26fF
C2390 fc2.n75 a_400_38200# 131.52fF
C2391 fc2.n76 a_400_38200# 0.09fF
C2392 fc2.n77 a_400_38200# 9.27fF
C2393 fc2.n78 a_400_38200# 2.95fF
C2394 fc2.n79 a_400_38200# 2.61fF
C2395 fc2.n80 a_400_38200# 7.90fF
C2396 fc2.n81 a_400_38200# 0.42fF
C2397 fc2.n82 a_400_38200# 2.09fF
C2398 fc2.n83 a_400_38200# 0.74fF
C2399 fc2.n84 a_400_38200# 0.15fF
C2400 fc2.n85 a_400_38200# 0.98fF
C2401 fc2.n86 a_400_38200# 0.24fF
C2402 fc2.n87 a_400_38200# 1.41fF
C2403 fc2.n88 a_400_38200# 0.24fF
C2404 fc2.n89 a_400_38200# 1.41fF
C2405 fc2.n90 a_400_38200# 0.24fF
C2406 fc2.n91 a_400_38200# 1.41fF
C2407 fc2.n92 a_400_38200# 22.65fF
C2408 fc2.n93 a_400_38200# 11.42fF
C2409 fc2.n94 a_400_38200# 12.94fF
C2410 fc2.n95 a_400_38200# 11.42fF
C2411 fc2.n96 a_400_38200# 12.94fF
C2412 fc2.n97 a_400_38200# 11.42fF
C2413 fc2.n98 a_400_38200# 12.94fF
C2414 fc2.n99 a_400_38200# 11.42fF
C2415 fc2.n100 a_400_38200# 12.94fF
C2416 fc2.n101 a_400_38200# 11.91fF
C2417 fc2.n102 a_400_38200# 72.64fF
C2418 fc2.n103 a_400_38200# 141.33fF
C2419 fc2.n104 a_400_38200# 368.23fF
C2420 fc2.n105 a_400_38200# 131.52fF
C2421 fc2.n106 a_400_38200# 3.72fF
C2422 fc2.n107 a_400_38200# 1.37fF
C2423 fc2.n108 a_400_38200# 0.25fF
C2424 fc2.n109 a_400_38200# 4.06fF
C2425 fc2.n110 a_400_38200# 0.08fF
C2426 fc2.n111 a_400_38200# 0.08fF
C2427 fc2.n112 a_400_38200# 0.30fF
C2428 fc2.n113 a_400_38200# 0.09fF
C2429 fc2.n114 a_400_38200# 0.18fF
C2430 fc2.n115 a_400_38200# 0.05fF
C2431 fc2.n116 a_400_38200# 0.02fF
C2432 fc2.n117 a_400_38200# 0.04fF
C2433 fc2.n118 a_400_38200# 0.20fF
C2434 fc2.n119 a_400_38200# 1.01fF
C2435 fc2.n120 a_400_38200# 0.02fF
C2436 fc2.n121 a_400_38200# 0.15fF
C2437 fc2.t44 a_400_38200# 0.02fF
C2438 fc2.n122 a_400_38200# 1.06fF
C2439 fc2.n123 a_400_38200# 0.03fF
C2440 fc2.n124 a_400_38200# 0.07fF
C2441 fc2.n125 a_400_38200# 0.05fF
C2442 fc2.n126 a_400_38200# 0.05fF
C2443 fc2.n127 a_400_38200# 0.64fF
C2444 fc2.n128 a_400_38200# 0.79fF
C2445 fc2.n129 a_400_38200# 1.01fF
C2446 fc2.n130 a_400_38200# 1.29fF
C2447 fc2.t8 a_400_38200# 7.96fF
C2448 fc2.n131 a_400_38200# 9.42fF
C2449 fc2.n133 a_400_38200# 0.33fF
C2450 fc2.n134 a_400_38200# 0.20fF
C2451 fc2.n135 a_400_38200# 3.05fF
C2452 fc2.n136 a_400_38200# 1.86fF
C2453 fc2.n137 a_400_38200# 0.03fF
C2454 fc2.n138 a_400_38200# 0.07fF
C2455 fc2.n139 a_400_38200# 0.24fF
C2456 fc2.n140 a_400_38200# 0.58fF
C2457 fc2.n141 a_400_38200# 0.44fF
C2458 fc2.n142 a_400_38200# 0.72fF
C2459 fc2.n143 a_400_38200# 0.74fF
C2460 fc2.n144 a_400_38200# 3.62fF
C2461 fc2.n145 a_400_38200# 0.22fF
C2462 fc2.n146 a_400_38200# 0.01fF
C2463 fc2.t252 a_400_38200# 0.02fF
C2464 fc2.n147 a_400_38200# 0.22fF
C2465 fc2.t208 a_400_38200# 0.02fF
C2466 fc2.n148 a_400_38200# 0.83fF
C2467 fc2.n149 a_400_38200# 0.62fF
C2468 fc2.n150 a_400_38200# 1.43fF
C2469 fc2.n151 a_400_38200# 0.51fF
C2470 fc2.n152 a_400_38200# 0.94fF
C2471 fc2.n153 a_400_38200# 0.18fF
C2472 fc2.n154 a_400_38200# 0.76fF
C2473 fc2.t290 a_400_38200# 0.02fF
C2474 fc2.n155 a_400_38200# 0.21fF
C2475 fc2.n156 a_400_38200# 0.31fF
C2476 fc2.n157 a_400_38200# 0.53fF
C2477 fc2.n158 a_400_38200# 0.10fF
C2478 fc2.t127 a_400_38200# 0.02fF
C2479 fc2.n159 a_400_38200# 0.12fF
C2480 fc2.n161 a_400_38200# 0.76fF
C2481 fc2.n162 a_400_38200# 0.44fF
C2482 fc2.n163 a_400_38200# 0.26fF
C2483 fc2.n164 a_400_38200# 0.70fF
C2484 fc2.n165 a_400_38200# 0.18fF
C2485 fc2.n166 a_400_38200# 1.49fF
C2486 fc2.t84 a_400_38200# 0.02fF
C2487 fc2.n167 a_400_38200# 0.21fF
C2488 fc2.n168 a_400_38200# 0.80fF
C2489 fc2.n169 a_400_38200# 0.04fF
C2490 fc2.t152 a_400_38200# 0.02fF
C2491 fc2.n170 a_400_38200# 0.10fF
C2492 fc2.n171 a_400_38200# 0.12fF
C2493 fc2.n173 a_400_38200# 7.70fF
C2494 fc2.n174 a_400_38200# 0.61fF
C2495 fc2.n175 a_400_38200# 0.25fF
C2496 fc2.n176 a_400_38200# 0.75fF
C2497 fc2.n177 a_400_38200# 0.18fF
C2498 fc2.n178 a_400_38200# 0.76fF
C2499 fc2.t230 a_400_38200# 0.02fF
C2500 fc2.n179 a_400_38200# 0.21fF
C2501 fc2.n180 a_400_38200# 0.31fF
C2502 fc2.n181 a_400_38200# 0.53fF
C2503 fc2.n182 a_400_38200# 0.10fF
C2504 fc2.t67 a_400_38200# 0.02fF
C2505 fc2.n183 a_400_38200# 0.12fF
C2506 fc2.n185 a_400_38200# 0.03fF
C2507 fc2.n186 a_400_38200# 0.01fF
C2508 fc2.n187 a_400_38200# 0.06fF
C2509 fc2.n188 a_400_38200# 0.24fF
C2510 fc2.n189 a_400_38200# 0.12fF
C2511 fc2.n190 a_400_38200# 0.27fF
C2512 fc2.n191 a_400_38200# 0.13fF
C2513 fc2.n192 a_400_38200# 0.06fF
C2514 fc2.n193 a_400_38200# 0.11fF
C2515 fc2.n194 a_400_38200# 0.05fF
C2516 fc2.n195 a_400_38200# 0.09fF
C2517 fc2.n196 a_400_38200# 0.03fF
C2518 fc2.n197 a_400_38200# 0.07fF
C2519 fc2.n198 a_400_38200# 0.32fF
C2520 fc2.n199 a_400_38200# 0.47fF
C2521 fc2.n200 a_400_38200# 0.29fF
C2522 fc2.n201 a_400_38200# 3.32fF
C2523 fc2.t97 a_400_38200# 0.02fF
C2524 fc2.n202 a_400_38200# 0.10fF
C2525 fc2.n203 a_400_38200# 0.12fF
C2526 fc2.t9 a_400_38200# 0.02fF
C2527 fc2.n205 a_400_38200# 0.21fF
C2528 fc2.n206 a_400_38200# 0.80fF
C2529 fc2.n207 a_400_38200# 0.04fF
C2530 fc2.n208 a_400_38200# 1.89fF
C2531 fc2.t110 a_400_38200# 0.02fF
C2532 fc2.n209 a_400_38200# 0.21fF
C2533 fc2.n210 a_400_38200# 0.31fF
C2534 fc2.n211 a_400_38200# 0.53fF
C2535 fc2.n212 a_400_38200# 0.10fF
C2536 fc2.t311 a_400_38200# 0.02fF
C2537 fc2.n213 a_400_38200# 0.12fF
C2538 fc2.n215 a_400_38200# 0.01fF
C2539 fc2.n216 a_400_38200# 0.03fF
C2540 fc2.n217 a_400_38200# 0.06fF
C2541 fc2.n218 a_400_38200# 0.24fF
C2542 fc2.n219 a_400_38200# 0.33fF
C2543 fc2.n220 a_400_38200# 0.13fF
C2544 fc2.n221 a_400_38200# 0.06fF
C2545 fc2.n222 a_400_38200# 0.11fF
C2546 fc2.n223 a_400_38200# 0.03fF
C2547 fc2.n224 a_400_38200# 0.07fF
C2548 fc2.n225 a_400_38200# 0.05fF
C2549 fc2.n226 a_400_38200# 0.09fF
C2550 fc2.n227 a_400_38200# 0.32fF
C2551 fc2.n228 a_400_38200# 0.47fF
C2552 fc2.n229 a_400_38200# 0.29fF
C2553 fc2.n230 a_400_38200# 1.59fF
C2554 fc2.n231 a_400_38200# 1.58fF
C2555 fc2.t338 a_400_38200# 0.02fF
C2556 fc2.n232 a_400_38200# 0.10fF
C2557 fc2.n233 a_400_38200# 0.12fF
C2558 fc2.t267 a_400_38200# 0.02fF
C2559 fc2.n235 a_400_38200# 0.21fF
C2560 fc2.n236 a_400_38200# 0.80fF
C2561 fc2.n237 a_400_38200# 0.04fF
C2562 fc2.n238 a_400_38200# 1.83fF
C2563 fc2.n239 a_400_38200# 0.58fF
C2564 fc2.n240 a_400_38200# 0.94fF
C2565 fc2.n241 a_400_38200# 0.18fF
C2566 fc2.n242 a_400_38200# 0.76fF
C2567 fc2.t347 a_400_38200# 0.02fF
C2568 fc2.n243 a_400_38200# 0.21fF
C2569 fc2.n244 a_400_38200# 0.31fF
C2570 fc2.n245 a_400_38200# 0.53fF
C2571 fc2.n246 a_400_38200# 0.10fF
C2572 fc2.t198 a_400_38200# 0.02fF
C2573 fc2.n247 a_400_38200# 0.12fF
C2574 fc2.n249 a_400_38200# 0.01fF
C2575 fc2.n250 a_400_38200# 0.03fF
C2576 fc2.n251 a_400_38200# 0.06fF
C2577 fc2.n252 a_400_38200# 0.24fF
C2578 fc2.n253 a_400_38200# 0.12fF
C2579 fc2.n254 a_400_38200# 0.27fF
C2580 fc2.n255 a_400_38200# 0.13fF
C2581 fc2.n256 a_400_38200# 0.06fF
C2582 fc2.n257 a_400_38200# 0.11fF
C2583 fc2.n258 a_400_38200# 0.03fF
C2584 fc2.n259 a_400_38200# 0.07fF
C2585 fc2.n260 a_400_38200# 0.05fF
C2586 fc2.n261 a_400_38200# 0.09fF
C2587 fc2.n262 a_400_38200# 0.32fF
C2588 fc2.n263 a_400_38200# 0.47fF
C2589 fc2.n264 a_400_38200# 0.29fF
C2590 fc2.n265 a_400_38200# 1.64fF
C2591 fc2.t206 a_400_38200# 0.02fF
C2592 fc2.n266 a_400_38200# 0.10fF
C2593 fc2.n267 a_400_38200# 0.12fF
C2594 fc2.t143 a_400_38200# 0.02fF
C2595 fc2.n269 a_400_38200# 0.21fF
C2596 fc2.n270 a_400_38200# 0.80fF
C2597 fc2.n271 a_400_38200# 0.04fF
C2598 fc2.n272 a_400_38200# 1.04fF
C2599 fc2.n273 a_400_38200# 0.12fF
C2600 fc2.n274 a_400_38200# 0.10fF
C2601 fc2.t191 a_400_38200# 0.02fF
C2602 fc2.n275 a_400_38200# 0.12fF
C2603 fc2.t360 a_400_38200# 0.02fF
C2604 fc2.n277 a_400_38200# 0.21fF
C2605 fc2.n278 a_400_38200# 0.31fF
C2606 fc2.n279 a_400_38200# 0.53fF
C2607 fc2.n280 a_400_38200# 1.94fF
C2608 fc2.n281 a_400_38200# 3.29fF
C2609 fc2.t218 a_400_38200# 0.02fF
C2610 fc2.n282 a_400_38200# 0.10fF
C2611 fc2.n283 a_400_38200# 0.12fF
C2612 fc2.t157 a_400_38200# 0.02fF
C2613 fc2.n285 a_400_38200# 0.21fF
C2614 fc2.n286 a_400_38200# 0.80fF
C2615 fc2.n287 a_400_38200# 0.04fF
C2616 fc2.t66 a_400_38200# 17.22fF
C2617 fc2.n288 a_400_38200# 0.10fF
C2618 fc2.t76 a_400_38200# 0.02fF
C2619 fc2.n289 a_400_38200# 0.12fF
C2620 fc2.n291 a_400_38200# 0.21fF
C2621 fc2.t25 a_400_38200# 0.02fF
C2622 fc2.n292 a_400_38200# 0.31fF
C2623 fc2.n293 a_400_38200# 0.32fF
C2624 fc2.n294 a_400_38200# 0.59fF
C2625 fc2.t82 a_400_38200# 0.02fF
C2626 fc2.n295 a_400_38200# 0.10fF
C2627 fc2.n296 a_400_38200# 0.12fF
C2628 fc2.n298 a_400_38200# 0.35fF
C2629 fc2.n299 a_400_38200# 0.21fF
C2630 fc2.t240 a_400_38200# 0.02fF
C2631 fc2.n300 a_400_38200# 0.31fF
C2632 fc2.n301 a_400_38200# 0.55fF
C2633 fc2.n302 a_400_38200# 0.35fF
C2634 fc2.n303 a_400_38200# 0.33fF
C2635 fc2.n304 a_400_38200# 0.13fF
C2636 fc2.n305 a_400_38200# 0.13fF
C2637 fc2.n306 a_400_38200# 0.05fF
C2638 fc2.n307 a_400_38200# 0.36fF
C2639 fc2.n308 a_400_38200# 0.49fF
C2640 fc2.n309 a_400_38200# 0.32fF
C2641 fc2.n310 a_400_38200# 0.10fF
C2642 fc2.n311 a_400_38200# 0.26fF
C2643 fc2.n312 a_400_38200# 0.82fF
C2644 fc2.n313 a_400_38200# 0.26fF
C2645 fc2.n314 a_400_38200# 0.52fF
C2646 fc2.n315 a_400_38200# 1.50fF
C2647 fc2.t243 a_400_38200# 0.02fF
C2648 fc2.n316 a_400_38200# 1.06fF
C2649 fc2.n317 a_400_38200# 0.46fF
C2650 fc2.n318 a_400_38200# 0.52fF
C2651 fc2.n319 a_400_38200# 0.46fF
C2652 fc2.n320 a_400_38200# 1.04fF
C2653 fc2.n321 a_400_38200# 0.12fF
C2654 fc2.n322 a_400_38200# 0.52fF
C2655 fc2.n323 a_400_38200# 0.10fF
C2656 fc2.t212 a_400_38200# 0.02fF
C2657 fc2.n324 a_400_38200# 0.12fF
C2658 fc2.t260 a_400_38200# 0.02fF
C2659 fc2.n326 a_400_38200# 0.21fF
C2660 fc2.n327 a_400_38200# 0.80fF
C2661 fc2.n328 a_400_38200# 0.04fF
C2662 fc2.t383 a_400_38200# 0.02fF
C2663 fc2.n329 a_400_38200# 0.21fF
C2664 fc2.n330 a_400_38200# 0.31fF
C2665 fc2.n331 a_400_38200# 0.53fF
C2666 fc2.n332 a_400_38200# 0.81fF
C2667 fc2.n333 a_400_38200# 0.88fF
C2668 fc2.n334 a_400_38200# 2.57fF
C2669 fc2.n335 a_400_38200# 3.37fF
C2670 fc2.t316 a_400_38200# 0.02fF
C2671 fc2.n336 a_400_38200# 0.10fF
C2672 fc2.n337 a_400_38200# 0.12fF
C2673 fc2.t125 a_400_38200# 0.02fF
C2674 fc2.n339 a_400_38200# 0.83fF
C2675 fc2.n340 a_400_38200# 0.62fF
C2676 fc2.n341 a_400_38200# 1.79fF
C2677 fc2.n342 a_400_38200# 0.05fF
C2678 fc2.n343 a_400_38200# 0.07fF
C2679 fc2.n344 a_400_38200# 1.14fF
C2680 fc2.n345 a_400_38200# 0.12fF
C2681 fc2.n346 a_400_38200# 0.05fF
C2682 fc2.n347 a_400_38200# 0.17fF
C2683 fc2.n348 a_400_38200# 0.06fF
C2684 fc2.n349 a_400_38200# 0.03fF
C2685 fc2.n350 a_400_38200# 0.10fF
C2686 fc2.n351 a_400_38200# 0.17fF
C2687 fc2.n352 a_400_38200# 0.68fF
C2688 fc2.t371 a_400_38200# 0.02fF
C2689 fc2.n353 a_400_38200# 0.21fF
C2690 fc2.n354 a_400_38200# 0.31fF
C2691 fc2.n355 a_400_38200# 0.53fF
C2692 fc2.n356 a_400_38200# 0.10fF
C2693 fc2.t202 a_400_38200# 0.02fF
C2694 fc2.n357 a_400_38200# 0.12fF
C2695 fc2.n359 a_400_38200# 0.01fF
C2696 fc2.n360 a_400_38200# 0.03fF
C2697 fc2.n361 a_400_38200# 0.06fF
C2698 fc2.n362 a_400_38200# 0.24fF
C2699 fc2.n363 a_400_38200# 0.05fF
C2700 fc2.n364 a_400_38200# 0.03fF
C2701 fc2.n365 a_400_38200# 0.33fF
C2702 fc2.n366 a_400_38200# 0.13fF
C2703 fc2.n367 a_400_38200# 0.06fF
C2704 fc2.n368 a_400_38200# 0.11fF
C2705 fc2.n369 a_400_38200# 0.03fF
C2706 fc2.n370 a_400_38200# 0.07fF
C2707 fc2.n371 a_400_38200# 0.03fF
C2708 fc2.n372 a_400_38200# 0.05fF
C2709 fc2.n373 a_400_38200# 0.05fF
C2710 fc2.n374 a_400_38200# 0.09fF
C2711 fc2.n375 a_400_38200# 0.32fF
C2712 fc2.n376 a_400_38200# 0.47fF
C2713 fc2.n377 a_400_38200# 0.29fF
C2714 fc2.n378 a_400_38200# 1.64fF
C2715 fc2.t250 a_400_38200# 0.02fF
C2716 fc2.n379 a_400_38200# 0.21fF
C2717 fc2.n380 a_400_38200# 0.80fF
C2718 fc2.n381 a_400_38200# 0.04fF
C2719 fc2.t323 a_400_38200# 0.02fF
C2720 fc2.n382 a_400_38200# 0.10fF
C2721 fc2.n383 a_400_38200# 0.12fF
C2722 fc2.n385 a_400_38200# 1.83fF
C2723 fc2.n386 a_400_38200# 2.55fF
C2724 fc2.t131 a_400_38200# 0.02fF
C2725 fc2.n387 a_400_38200# 0.21fF
C2726 fc2.n388 a_400_38200# 0.31fF
C2727 fc2.n389 a_400_38200# 0.53fF
C2728 fc2.n390 a_400_38200# 0.10fF
C2729 fc2.t331 a_400_38200# 0.02fF
C2730 fc2.n391 a_400_38200# 0.12fF
C2731 fc2.n393 a_400_38200# 0.01fF
C2732 fc2.n394 a_400_38200# 0.03fF
C2733 fc2.n395 a_400_38200# 0.06fF
C2734 fc2.n396 a_400_38200# 0.24fF
C2735 fc2.n397 a_400_38200# 0.05fF
C2736 fc2.n398 a_400_38200# 0.03fF
C2737 fc2.n399 a_400_38200# 0.33fF
C2738 fc2.n400 a_400_38200# 0.13fF
C2739 fc2.n401 a_400_38200# 0.06fF
C2740 fc2.n402 a_400_38200# 0.11fF
C2741 fc2.n403 a_400_38200# 0.03fF
C2742 fc2.n404 a_400_38200# 0.07fF
C2743 fc2.n405 a_400_38200# 0.03fF
C2744 fc2.n406 a_400_38200# 0.05fF
C2745 fc2.n407 a_400_38200# 0.05fF
C2746 fc2.n408 a_400_38200# 0.09fF
C2747 fc2.n409 a_400_38200# 0.32fF
C2748 fc2.n410 a_400_38200# 0.47fF
C2749 fc2.n411 a_400_38200# 0.29fF
C2750 fc2.n412 a_400_38200# 2.06fF
C2751 fc2.t377 a_400_38200# 0.02fF
C2752 fc2.n413 a_400_38200# 0.21fF
C2753 fc2.n414 a_400_38200# 0.80fF
C2754 fc2.n415 a_400_38200# 0.04fF
C2755 fc2.t63 a_400_38200# 0.02fF
C2756 fc2.n416 a_400_38200# 0.10fF
C2757 fc2.n417 a_400_38200# 0.12fF
C2758 fc2.n419 a_400_38200# 0.05fF
C2759 fc2.n420 a_400_38200# 0.07fF
C2760 fc2.n421 a_400_38200# 1.07fF
C2761 fc2.n422 a_400_38200# 0.12fF
C2762 fc2.n423 a_400_38200# 0.16fF
C2763 fc2.n424 a_400_38200# 0.05fF
C2764 fc2.n425 a_400_38200# 0.03fF
C2765 fc2.n426 a_400_38200# 0.10fF
C2766 fc2.n427 a_400_38200# 0.17fF
C2767 fc2.n428 a_400_38200# 0.69fF
C2768 fc2.t257 a_400_38200# 0.02fF
C2769 fc2.n429 a_400_38200# 0.21fF
C2770 fc2.n430 a_400_38200# 0.31fF
C2771 fc2.n431 a_400_38200# 0.53fF
C2772 fc2.n432 a_400_38200# 0.10fF
C2773 fc2.t91 a_400_38200# 0.02fF
C2774 fc2.n433 a_400_38200# 0.12fF
C2775 fc2.n435 a_400_38200# 0.03fF
C2776 fc2.n436 a_400_38200# 0.01fF
C2777 fc2.n437 a_400_38200# 0.06fF
C2778 fc2.n438 a_400_38200# 0.24fF
C2779 fc2.n439 a_400_38200# 0.33fF
C2780 fc2.n440 a_400_38200# 0.05fF
C2781 fc2.n441 a_400_38200# 0.03fF
C2782 fc2.n442 a_400_38200# 0.13fF
C2783 fc2.n443 a_400_38200# 0.06fF
C2784 fc2.n444 a_400_38200# 0.11fF
C2785 fc2.n445 a_400_38200# 0.03fF
C2786 fc2.n446 a_400_38200# 0.05fF
C2787 fc2.n447 a_400_38200# 0.05fF
C2788 fc2.n448 a_400_38200# 0.09fF
C2789 fc2.n449 a_400_38200# 0.03fF
C2790 fc2.n450 a_400_38200# 0.07fF
C2791 fc2.n451 a_400_38200# 0.32fF
C2792 fc2.n452 a_400_38200# 0.47fF
C2793 fc2.n453 a_400_38200# 0.29fF
C2794 fc2.n454 a_400_38200# 3.32fF
C2795 fc2.t135 a_400_38200# 0.02fF
C2796 fc2.n455 a_400_38200# 0.21fF
C2797 fc2.n456 a_400_38200# 0.80fF
C2798 fc2.n457 a_400_38200# 0.04fF
C2799 fc2.t186 a_400_38200# 0.02fF
C2800 fc2.n458 a_400_38200# 0.10fF
C2801 fc2.n459 a_400_38200# 0.12fF
C2802 fc2.n461 a_400_38200# 0.04fF
C2803 fc2.n462 a_400_38200# 0.05fF
C2804 fc2.n463 a_400_38200# 0.05fF
C2805 fc2.n464 a_400_38200# 0.03fF
C2806 fc2.n466 a_400_38200# 0.99fF
C2807 fc2.n467 a_400_38200# 0.22fF
C2808 fc2.n468 a_400_38200# 0.03fF
C2809 fc2.n469 a_400_38200# 0.01fF
C2810 fc2.n470 a_400_38200# 0.06fF
C2811 fc2.n471 a_400_38200# 0.62fF
C2812 fc2.t72 a_400_38200# 0.02fF
C2813 fc2.n472 a_400_38200# 0.21fF
C2814 fc2.n473 a_400_38200# 0.31fF
C2815 fc2.n474 a_400_38200# 0.53fF
C2816 fc2.n475 a_400_38200# 0.10fF
C2817 fc2.t270 a_400_38200# 0.02fF
C2818 fc2.n476 a_400_38200# 0.12fF
C2819 fc2.n478 a_400_38200# 0.01fF
C2820 fc2.n479 a_400_38200# 0.03fF
C2821 fc2.n480 a_400_38200# 0.06fF
C2822 fc2.n481 a_400_38200# 0.24fF
C2823 fc2.n482 a_400_38200# 0.05fF
C2824 fc2.n483 a_400_38200# 0.03fF
C2825 fc2.n484 a_400_38200# 0.32fF
C2826 fc2.n485 a_400_38200# 0.13fF
C2827 fc2.n486 a_400_38200# 0.06fF
C2828 fc2.n487 a_400_38200# 0.11fF
C2829 fc2.n488 a_400_38200# 0.03fF
C2830 fc2.n489 a_400_38200# 0.07fF
C2831 fc2.n490 a_400_38200# 0.03fF
C2832 fc2.n491 a_400_38200# 0.05fF
C2833 fc2.n492 a_400_38200# 0.05fF
C2834 fc2.n493 a_400_38200# 0.09fF
C2835 fc2.n494 a_400_38200# 0.32fF
C2836 fc2.n495 a_400_38200# 0.47fF
C2837 fc2.n496 a_400_38200# 0.29fF
C2838 fc2.n497 a_400_38200# 3.02fF
C2839 fc2.t318 a_400_38200# 0.02fF
C2840 fc2.n498 a_400_38200# 0.21fF
C2841 fc2.n499 a_400_38200# 0.80fF
C2842 fc2.n500 a_400_38200# 0.04fF
C2843 fc2.t373 a_400_38200# 0.02fF
C2844 fc2.n501 a_400_38200# 0.10fF
C2845 fc2.n502 a_400_38200# 0.12fF
C2846 fc2.n504 a_400_38200# 7.70fF
C2847 fc2.n505 a_400_38200# 2.05fF
C2848 fc2.n506 a_400_38200# 0.05fF
C2849 fc2.n507 a_400_38200# 0.07fF
C2850 fc2.n508 a_400_38200# 1.00fF
C2851 fc2.n509 a_400_38200# 0.12fF
C2852 fc2.n510 a_400_38200# 0.05fF
C2853 fc2.n511 a_400_38200# 0.17fF
C2854 fc2.n512 a_400_38200# 0.06fF
C2855 fc2.n513 a_400_38200# 0.03fF
C2856 fc2.n514 a_400_38200# 0.10fF
C2857 fc2.n515 a_400_38200# 0.17fF
C2858 fc2.n516 a_400_38200# 0.69fF
C2859 fc2.t141 a_400_38200# 0.02fF
C2860 fc2.n517 a_400_38200# 0.21fF
C2861 fc2.n518 a_400_38200# 0.31fF
C2862 fc2.n519 a_400_38200# 0.53fF
C2863 fc2.n520 a_400_38200# 0.10fF
C2864 fc2.t343 a_400_38200# 0.02fF
C2865 fc2.n521 a_400_38200# 0.12fF
C2866 fc2.n523 a_400_38200# 0.10fF
C2867 fc2.n524 a_400_38200# 0.04fF
C2868 fc2.n525 a_400_38200# 0.11fF
C2869 fc2.n526 a_400_38200# 0.07fF
C2870 fc2.n527 a_400_38200# 0.09fF
C2871 fc2.n528 a_400_38200# 0.12fF
C2872 fc2.n529 a_400_38200# 0.69fF
C2873 fc2.n530 a_400_38200# 0.11fF
C2874 fc2.n531 a_400_38200# 1.07fF
C2875 fc2.n532 a_400_38200# 0.13fF
C2876 fc2.n533 a_400_38200# 1.51fF
C2877 fc2.t245 a_400_38200# 0.02fF
C2878 fc2.n534 a_400_38200# 0.10fF
C2879 fc2.n535 a_400_38200# 0.12fF
C2880 fc2.t388 a_400_38200# 0.02fF
C2881 fc2.n537 a_400_38200# 0.21fF
C2882 fc2.n538 a_400_38200# 0.80fF
C2883 fc2.n539 a_400_38200# 0.04fF
C2884 fc2.t193 a_400_38200# 0.02fF
C2885 fc2.n540 a_400_38200# 0.01fF
C2886 fc2.n541 a_400_38200# 0.22fF
C2887 fc2.t62 a_400_38200# 17.21fF
C2888 fc2.n542 a_400_38200# 0.22fF
C2889 fc2.n543 a_400_38200# 1.23fF
C2890 fc2.n544 a_400_38200# 0.52fF
C2891 fc2.n545 a_400_38200# 0.15fF
C2892 fc2.n546 a_400_38200# 0.77fF
C2893 fc2.n547 a_400_38200# 0.52fF
C2894 fc2.n548 a_400_38200# 0.07fF
C2895 fc2.n549 a_400_38200# 1.89fF
C2896 fc2.n550 a_400_38200# 0.52fF
C2897 fc2.n551 a_400_38200# 0.19fF
C2898 fc2.n552 a_400_38200# 1.28fF
C2899 fc2.t43 a_400_38200# 7.96fF
C2900 fc2.n554 a_400_38200# 7.30fF
C2901 fc2.n556 a_400_38200# 1.22fF
C2902 fc2.n557 a_400_38200# 3.88fF
C2903 fc2.n558 a_400_38200# 1.81fF
C2904 fc2.n559 a_400_38200# 3.03fF
C2905 fc2.n560 a_400_38200# 0.28fF
C2906 fc2.n561 a_400_38200# 0.12fF
C2907 fc2.n562 a_400_38200# 0.18fF
C2908 fc2.n563 a_400_38200# 0.05fF
C2909 fc2.n564 a_400_38200# 0.04fF
C2910 fc2.n565 a_400_38200# 0.20fF
C2911 fc2.n566 a_400_38200# 1.01fF
C2912 fc2.n567 a_400_38200# 0.02fF
C2913 fc2.n568 a_400_38200# 1.68fF
C2914 fc2.n569 a_400_38200# 0.05fF
C2915 fc2.n570 a_400_38200# 0.06fF
C2916 fc2.n571 a_400_38200# 1.07fF
C2917 fc2.n572 a_400_38200# 0.12fF
C2918 fc2.n573 a_400_38200# 0.05fF
C2919 fc2.n574 a_400_38200# 0.16fF
C2920 fc2.n575 a_400_38200# 0.03fF
C2921 fc2.n576 a_400_38200# 0.08fF
C2922 fc2.n577 a_400_38200# 0.16fF
C2923 fc2.n578 a_400_38200# 0.71fF
C2924 fc2.t132 a_400_38200# 0.02fF
C2925 fc2.n579 a_400_38200# 0.21fF
C2926 fc2.n580 a_400_38200# 0.31fF
C2927 fc2.n581 a_400_38200# 0.53fF
C2928 fc2.n582 a_400_38200# 0.10fF
C2929 fc2.t332 a_400_38200# 0.02fF
C2930 fc2.n583 a_400_38200# 0.12fF
C2931 fc2.n585 a_400_38200# 0.01fF
C2932 fc2.n586 a_400_38200# 0.03fF
C2933 fc2.n587 a_400_38200# 0.06fF
C2934 fc2.n588 a_400_38200# 0.24fF
C2935 fc2.n589 a_400_38200# 0.05fF
C2936 fc2.n590 a_400_38200# 0.03fF
C2937 fc2.n591 a_400_38200# 0.33fF
C2938 fc2.n592 a_400_38200# 0.13fF
C2939 fc2.n593 a_400_38200# 0.06fF
C2940 fc2.n594 a_400_38200# 0.11fF
C2941 fc2.n595 a_400_38200# 0.03fF
C2942 fc2.n596 a_400_38200# 0.07fF
C2943 fc2.n597 a_400_38200# 0.03fF
C2944 fc2.n598 a_400_38200# 0.05fF
C2945 fc2.n599 a_400_38200# 0.05fF
C2946 fc2.n600 a_400_38200# 0.09fF
C2947 fc2.n601 a_400_38200# 0.32fF
C2948 fc2.n602 a_400_38200# 0.47fF
C2949 fc2.n603 a_400_38200# 0.29fF
C2950 fc2.n604 a_400_38200# 1.87fF
C2951 fc2.t378 a_400_38200# 0.02fF
C2952 fc2.n605 a_400_38200# 0.21fF
C2953 fc2.n606 a_400_38200# 0.80fF
C2954 fc2.n607 a_400_38200# 0.04fF
C2955 fc2.t231 a_400_38200# 0.02fF
C2956 fc2.n608 a_400_38200# 0.10fF
C2957 fc2.n609 a_400_38200# 0.12fF
C2958 fc2.n611 a_400_38200# 0.50fF
C2959 fc2.n612 a_400_38200# 0.94fF
C2960 fc2.n613 a_400_38200# 0.18fF
C2961 fc2.n614 a_400_38200# 0.76fF
C2962 fc2.t348 a_400_38200# 0.02fF
C2963 fc2.n615 a_400_38200# 0.21fF
C2964 fc2.n616 a_400_38200# 0.31fF
C2965 fc2.n617 a_400_38200# 0.53fF
C2966 fc2.t27 a_400_38200# 0.02fF
C2967 fc2.n618 a_400_38200# 1.06fF
C2968 fc2.n619 a_400_38200# 0.03fF
C2969 fc2.n620 a_400_38200# 0.07fF
C2970 fc2.n621 a_400_38200# 0.05fF
C2971 fc2.n622 a_400_38200# 0.05fF
C2972 fc2.n623 a_400_38200# 0.05fF
C2973 fc2.n624 a_400_38200# 0.64fF
C2974 fc2.n625 a_400_38200# 0.79fF
C2975 fc2.n626 a_400_38200# 1.01fF
C2976 fc2.n627 a_400_38200# 1.29fF
C2977 fc2.t2 a_400_38200# 7.96fF
C2978 fc2.n628 a_400_38200# 9.42fF
C2979 fc2.n630 a_400_38200# 0.33fF
C2980 fc2.n631 a_400_38200# 0.20fF
C2981 fc2.n632 a_400_38200# 3.05fF
C2982 fc2.n633 a_400_38200# 1.86fF
C2983 fc2.n634 a_400_38200# 0.03fF
C2984 fc2.n635 a_400_38200# 0.07fF
C2985 fc2.n636 a_400_38200# 0.24fF
C2986 fc2.n637 a_400_38200# 0.58fF
C2987 fc2.n638 a_400_38200# 0.44fF
C2988 fc2.n639 a_400_38200# 0.72fF
C2989 fc2.n640 a_400_38200# 0.74fF
C2990 fc2.n641 a_400_38200# 3.62fF
C2991 fc2.n642 a_400_38200# 0.22fF
C2992 fc2.n643 a_400_38200# 0.01fF
C2993 fc2.t239 a_400_38200# 0.02fF
C2994 fc2.n644 a_400_38200# 0.22fF
C2995 fc2.t199 a_400_38200# 0.02fF
C2996 fc2.n645 a_400_38200# 0.83fF
C2997 fc2.n646 a_400_38200# 0.62fF
C2998 fc2.n647 a_400_38200# 1.07fF
C2999 fc2.n648 a_400_38200# 0.25fF
C3000 fc2.n649 a_400_38200# 0.75fF
C3001 fc2.n650 a_400_38200# 0.18fF
C3002 fc2.n651 a_400_38200# 0.44fF
C3003 fc2.n652 a_400_38200# 0.79fF
C3004 fc2.t277 a_400_38200# 0.02fF
C3005 fc2.n653 a_400_38200# 0.21fF
C3006 fc2.n654 a_400_38200# 0.31fF
C3007 fc2.n655 a_400_38200# 0.53fF
C3008 fc2.n656 a_400_38200# 0.10fF
C3009 fc2.t114 a_400_38200# 0.02fF
C3010 fc2.n657 a_400_38200# 0.12fF
C3011 fc2.n659 a_400_38200# 0.01fF
C3012 fc2.n660 a_400_38200# 0.03fF
C3013 fc2.n661 a_400_38200# 0.06fF
C3014 fc2.n662 a_400_38200# 0.24fF
C3015 fc2.n663 a_400_38200# 0.33fF
C3016 fc2.n664 a_400_38200# 0.13fF
C3017 fc2.n665 a_400_38200# 0.06fF
C3018 fc2.n666 a_400_38200# 0.11fF
C3019 fc2.n667 a_400_38200# 0.03fF
C3020 fc2.n668 a_400_38200# 0.07fF
C3021 fc2.n669 a_400_38200# 0.05fF
C3022 fc2.n670 a_400_38200# 0.09fF
C3023 fc2.n671 a_400_38200# 0.32fF
C3024 fc2.n672 a_400_38200# 0.47fF
C3025 fc2.n673 a_400_38200# 0.29fF
C3026 fc2.n674 a_400_38200# 1.60fF
C3027 fc2.t74 a_400_38200# 0.02fF
C3028 fc2.n675 a_400_38200# 0.21fF
C3029 fc2.n676 a_400_38200# 0.80fF
C3030 fc2.n677 a_400_38200# 0.04fF
C3031 fc2.t140 a_400_38200# 0.02fF
C3032 fc2.n678 a_400_38200# 0.10fF
C3033 fc2.n679 a_400_38200# 0.12fF
C3034 fc2.n681 a_400_38200# 0.50fF
C3035 fc2.n682 a_400_38200# 0.94fF
C3036 fc2.n683 a_400_38200# 0.18fF
C3037 fc2.n684 a_400_38200# 0.76fF
C3038 fc2.t217 a_400_38200# 0.02fF
C3039 fc2.n685 a_400_38200# 0.21fF
C3040 fc2.n686 a_400_38200# 0.31fF
C3041 fc2.n687 a_400_38200# 0.53fF
C3042 fc2.n688 a_400_38200# 0.10fF
C3043 fc2.t53 a_400_38200# 0.02fF
C3044 fc2.n689 a_400_38200# 0.12fF
C3045 fc2.n691 a_400_38200# 0.76fF
C3046 fc2.n692 a_400_38200# 0.44fF
C3047 fc2.n693 a_400_38200# 1.07fF
C3048 fc2.n694 a_400_38200# 0.18fF
C3049 fc2.n695 a_400_38200# 3.23fF
C3050 fc2.t385 a_400_38200# 0.02fF
C3051 fc2.n696 a_400_38200# 0.21fF
C3052 fc2.n697 a_400_38200# 0.80fF
C3053 fc2.n698 a_400_38200# 0.04fF
C3054 fc2.t83 a_400_38200# 0.02fF
C3055 fc2.n699 a_400_38200# 0.10fF
C3056 fc2.n700 a_400_38200# 0.12fF
C3057 fc2.n702 a_400_38200# 7.70fF
C3058 fc2.n703 a_400_38200# 0.44fF
C3059 fc2.n704 a_400_38200# 0.25fF
C3060 fc2.n705 a_400_38200# 0.75fF
C3061 fc2.n706 a_400_38200# 0.18fF
C3062 fc2.n707 a_400_38200# 0.76fF
C3063 fc2.t337 a_400_38200# 0.02fF
C3064 fc2.n708 a_400_38200# 0.21fF
C3065 fc2.n709 a_400_38200# 0.31fF
C3066 fc2.n710 a_400_38200# 0.53fF
C3067 fc2.n711 a_400_38200# 0.10fF
C3068 fc2.t187 a_400_38200# 0.02fF
C3069 fc2.n712 a_400_38200# 0.12fF
C3070 fc2.n714 a_400_38200# 0.03fF
C3071 fc2.n715 a_400_38200# 0.01fF
C3072 fc2.n716 a_400_38200# 0.06fF
C3073 fc2.n717 a_400_38200# 0.24fF
C3074 fc2.n718 a_400_38200# 0.33fF
C3075 fc2.n719 a_400_38200# 0.13fF
C3076 fc2.n720 a_400_38200# 0.06fF
C3077 fc2.n721 a_400_38200# 0.11fF
C3078 fc2.n722 a_400_38200# 0.05fF
C3079 fc2.n723 a_400_38200# 0.09fF
C3080 fc2.n724 a_400_38200# 0.03fF
C3081 fc2.n725 a_400_38200# 0.07fF
C3082 fc2.n726 a_400_38200# 0.32fF
C3083 fc2.n727 a_400_38200# 0.47fF
C3084 fc2.n728 a_400_38200# 0.29fF
C3085 fc2.n729 a_400_38200# 3.32fF
C3086 fc2.t197 a_400_38200# 0.02fF
C3087 fc2.n730 a_400_38200# 0.10fF
C3088 fc2.n731 a_400_38200# 0.12fF
C3089 fc2.t133 a_400_38200# 0.02fF
C3090 fc2.n733 a_400_38200# 0.21fF
C3091 fc2.n734 a_400_38200# 0.80fF
C3092 fc2.n735 a_400_38200# 0.04fF
C3093 fc2.n736 a_400_38200# 1.71fF
C3094 fc2.n737 a_400_38200# 1.87fF
C3095 fc2.t226 a_400_38200# 0.02fF
C3096 fc2.n738 a_400_38200# 0.21fF
C3097 fc2.n739 a_400_38200# 0.31fF
C3098 fc2.n740 a_400_38200# 0.53fF
C3099 fc2.n741 a_400_38200# 0.10fF
C3100 fc2.t64 a_400_38200# 0.02fF
C3101 fc2.n742 a_400_38200# 0.12fF
C3102 fc2.n744 a_400_38200# 0.01fF
C3103 fc2.n745 a_400_38200# 0.03fF
C3104 fc2.n746 a_400_38200# 0.06fF
C3105 fc2.n747 a_400_38200# 0.24fF
C3106 fc2.n748 a_400_38200# 0.33fF
C3107 fc2.n749 a_400_38200# 0.13fF
C3108 fc2.n750 a_400_38200# 0.06fF
C3109 fc2.n751 a_400_38200# 0.11fF
C3110 fc2.n752 a_400_38200# 0.04fF
C3111 fc2.n753 a_400_38200# 0.08fF
C3112 fc2.n754 a_400_38200# 0.05fF
C3113 fc2.n755 a_400_38200# 0.09fF
C3114 fc2.n756 a_400_38200# 0.32fF
C3115 fc2.n757 a_400_38200# 0.47fF
C3116 fc2.n758 a_400_38200# 0.29fF
C3117 fc2.n759 a_400_38200# 1.78fF
C3118 fc2.t73 a_400_38200# 0.02fF
C3119 fc2.n760 a_400_38200# 0.10fF
C3120 fc2.n761 a_400_38200# 0.12fF
C3121 fc2.t3 a_400_38200# 0.02fF
C3122 fc2.n763 a_400_38200# 0.21fF
C3123 fc2.n764 a_400_38200# 0.80fF
C3124 fc2.n765 a_400_38200# 0.04fF
C3125 fc2.n766 a_400_38200# 1.04fF
C3126 fc2.n767 a_400_38200# 0.12fF
C3127 fc2.n768 a_400_38200# 0.10fF
C3128 fc2.t297 a_400_38200# 0.02fF
C3129 fc2.n769 a_400_38200# 0.12fF
C3130 fc2.t96 a_400_38200# 0.02fF
C3131 fc2.n771 a_400_38200# 0.21fF
C3132 fc2.n772 a_400_38200# 0.31fF
C3133 fc2.n773 a_400_38200# 0.53fF
C3134 fc2.n774 a_400_38200# 0.76fF
C3135 fc2.n775 a_400_38200# 0.50fF
C3136 fc2.n776 a_400_38200# 0.94fF
C3137 fc2.n777 a_400_38200# 0.18fF
C3138 fc2.n778 a_400_38200# 3.32fF
C3139 fc2.t325 a_400_38200# 0.02fF
C3140 fc2.n779 a_400_38200# 0.10fF
C3141 fc2.n780 a_400_38200# 0.12fF
C3142 fc2.t258 a_400_38200# 0.02fF
C3143 fc2.n782 a_400_38200# 0.21fF
C3144 fc2.n783 a_400_38200# 0.80fF
C3145 fc2.n784 a_400_38200# 0.04fF
C3146 fc2.t52 a_400_38200# 17.22fF
C3147 fc2.t144 a_400_38200# 0.02fF
C3148 fc2.n785 a_400_38200# 0.21fF
C3149 fc2.n786 a_400_38200# 0.80fF
C3150 fc2.n787 a_400_38200# 0.04fF
C3151 fc2.t207 a_400_38200# 0.02fF
C3152 fc2.n788 a_400_38200# 0.10fF
C3153 fc2.n789 a_400_38200# 0.12fF
C3154 fc2.n791 a_400_38200# 0.10fF
C3155 fc2.t180 a_400_38200# 0.02fF
C3156 fc2.n792 a_400_38200# 0.12fF
C3157 fc2.n794 a_400_38200# 0.01fF
C3158 fc2.n795 a_400_38200# 0.03fF
C3159 fc2.n796 a_400_38200# 0.06fF
C3160 fc2.n797 a_400_38200# 0.24fF
C3161 fc2.n798 a_400_38200# 0.33fF
C3162 fc2.n799 a_400_38200# 0.13fF
C3163 fc2.n800 a_400_38200# 0.06fF
C3164 fc2.n801 a_400_38200# 0.11fF
C3165 fc2.n802 a_400_38200# 0.03fF
C3166 fc2.n803 a_400_38200# 0.07fF
C3167 fc2.n804 a_400_38200# 0.05fF
C3168 fc2.n805 a_400_38200# 0.09fF
C3169 fc2.n806 a_400_38200# 0.32fF
C3170 fc2.n807 a_400_38200# 0.47fF
C3171 fc2.n808 a_400_38200# 0.29fF
C3172 fc2.n809 a_400_38200# 3.68fF
C3173 fc2.n810 a_400_38200# 1.75fF
C3174 fc2.n811 a_400_38200# 0.05fF
C3175 fc2.n812 a_400_38200# 0.07fF
C3176 fc2.n813 a_400_38200# 1.00fF
C3177 fc2.n814 a_400_38200# 0.12fF
C3178 fc2.n815 a_400_38200# 0.05fF
C3179 fc2.n816 a_400_38200# 0.17fF
C3180 fc2.n817 a_400_38200# 0.06fF
C3181 fc2.n818 a_400_38200# 0.03fF
C3182 fc2.n819 a_400_38200# 0.10fF
C3183 fc2.n820 a_400_38200# 0.17fF
C3184 fc2.n821 a_400_38200# 0.69fF
C3185 fc2.t372 a_400_38200# 0.02fF
C3186 fc2.n822 a_400_38200# 0.21fF
C3187 fc2.n823 a_400_38200# 0.31fF
C3188 fc2.n824 a_400_38200# 0.53fF
C3189 fc2.n825 a_400_38200# 0.10fF
C3190 fc2.t203 a_400_38200# 0.02fF
C3191 fc2.n826 a_400_38200# 0.12fF
C3192 fc2.n828 a_400_38200# 0.01fF
C3193 fc2.n829 a_400_38200# 0.03fF
C3194 fc2.n830 a_400_38200# 0.06fF
C3195 fc2.n831 a_400_38200# 0.24fF
C3196 fc2.n832 a_400_38200# 0.05fF
C3197 fc2.n833 a_400_38200# 0.03fF
C3198 fc2.n834 a_400_38200# 0.33fF
C3199 fc2.n835 a_400_38200# 0.13fF
C3200 fc2.n836 a_400_38200# 0.06fF
C3201 fc2.n837 a_400_38200# 0.11fF
C3202 fc2.n838 a_400_38200# 0.03fF
C3203 fc2.n839 a_400_38200# 0.07fF
C3204 fc2.n840 a_400_38200# 0.03fF
C3205 fc2.n841 a_400_38200# 0.05fF
C3206 fc2.n842 a_400_38200# 0.05fF
C3207 fc2.n843 a_400_38200# 0.09fF
C3208 fc2.n844 a_400_38200# 0.32fF
C3209 fc2.n845 a_400_38200# 0.47fF
C3210 fc2.n846 a_400_38200# 0.29fF
C3211 fc2.n847 a_400_38200# 1.53fF
C3212 fc2.t251 a_400_38200# 0.02fF
C3213 fc2.n848 a_400_38200# 0.21fF
C3214 fc2.n849 a_400_38200# 0.80fF
C3215 fc2.n850 a_400_38200# 0.04fF
C3216 fc2.t305 a_400_38200# 0.02fF
C3217 fc2.n851 a_400_38200# 0.10fF
C3218 fc2.n852 a_400_38200# 0.12fF
C3219 fc2.n854 a_400_38200# 1.81fF
C3220 fc2.n855 a_400_38200# 0.05fF
C3221 fc2.n856 a_400_38200# 0.07fF
C3222 fc2.n857 a_400_38200# 1.00fF
C3223 fc2.n858 a_400_38200# 0.12fF
C3224 fc2.n859 a_400_38200# 0.05fF
C3225 fc2.n860 a_400_38200# 0.17fF
C3226 fc2.n861 a_400_38200# 0.06fF
C3227 fc2.n862 a_400_38200# 0.03fF
C3228 fc2.n863 a_400_38200# 0.10fF
C3229 fc2.n864 a_400_38200# 0.17fF
C3230 fc2.n865 a_400_38200# 0.69fF
C3231 fc2.t244 a_400_38200# 0.02fF
C3232 fc2.n866 a_400_38200# 0.21fF
C3233 fc2.n867 a_400_38200# 0.31fF
C3234 fc2.n868 a_400_38200# 0.53fF
C3235 fc2.n869 a_400_38200# 0.10fF
C3236 fc2.t80 a_400_38200# 0.02fF
C3237 fc2.n870 a_400_38200# 0.12fF
C3238 fc2.n872 a_400_38200# 0.76fF
C3239 fc2.n873 a_400_38200# 0.44fF
C3240 fc2.n874 a_400_38200# 1.07fF
C3241 fc2.n875 a_400_38200# 0.18fF
C3242 fc2.n876 a_400_38200# 1.51fF
C3243 fc2.t126 a_400_38200# 0.02fF
C3244 fc2.n877 a_400_38200# 0.21fF
C3245 fc2.n878 a_400_38200# 0.80fF
C3246 fc2.n879 a_400_38200# 0.04fF
C3247 fc2.t176 a_400_38200# 0.02fF
C3248 fc2.n880 a_400_38200# 0.10fF
C3249 fc2.n881 a_400_38200# 0.12fF
C3250 fc2.n883 a_400_38200# 7.70fF
C3251 fc2.n884 a_400_38200# 0.04fF
C3252 fc2.n885 a_400_38200# 0.05fF
C3253 fc2.n886 a_400_38200# 0.05fF
C3254 fc2.n887 a_400_38200# 0.03fF
C3255 fc2.n888 a_400_38200# 1.06fF
C3256 fc2.n889 a_400_38200# 0.21fF
C3257 fc2.n890 a_400_38200# 0.10fF
C3258 fc2.n891 a_400_38200# 0.64fF
C3259 fc2.t60 a_400_38200# 0.02fF
C3260 fc2.n892 a_400_38200# 0.21fF
C3261 fc2.n893 a_400_38200# 0.31fF
C3262 fc2.n894 a_400_38200# 0.53fF
C3263 fc2.n895 a_400_38200# 0.10fF
C3264 fc2.t262 a_400_38200# 0.02fF
C3265 fc2.n896 a_400_38200# 0.12fF
C3266 fc2.n898 a_400_38200# 0.01fF
C3267 fc2.n899 a_400_38200# 0.03fF
C3268 fc2.n900 a_400_38200# 0.06fF
C3269 fc2.n901 a_400_38200# 0.24fF
C3270 fc2.n902 a_400_38200# 0.03fF
C3271 fc2.n903 a_400_38200# 0.32fF
C3272 fc2.n904 a_400_38200# 0.13fF
C3273 fc2.n905 a_400_38200# 0.06fF
C3274 fc2.n906 a_400_38200# 0.11fF
C3275 fc2.n907 a_400_38200# 0.03fF
C3276 fc2.n908 a_400_38200# 0.07fF
C3277 fc2.n909 a_400_38200# 0.03fF
C3278 fc2.n910 a_400_38200# 0.05fF
C3279 fc2.n911 a_400_38200# 0.05fF
C3280 fc2.n912 a_400_38200# 0.09fF
C3281 fc2.n913 a_400_38200# 0.32fF
C3282 fc2.n914 a_400_38200# 0.47fF
C3283 fc2.n915 a_400_38200# 0.29fF
C3284 fc2.n916 a_400_38200# 3.03fF
C3285 fc2.t361 a_400_38200# 0.02fF
C3286 fc2.n917 a_400_38200# 0.10fF
C3287 fc2.n918 a_400_38200# 0.12fF
C3288 fc2.t308 a_400_38200# 0.02fF
C3289 fc2.n920 a_400_38200# 0.21fF
C3290 fc2.n921 a_400_38200# 0.80fF
C3291 fc2.n922 a_400_38200# 0.04fF
C3292 fc2.n923 a_400_38200# 0.05fF
C3293 fc2.n924 a_400_38200# 0.07fF
C3294 fc2.n925 a_400_38200# 1.27fF
C3295 fc2.n926 a_400_38200# 0.12fF
C3296 fc2.n927 a_400_38200# 0.16fF
C3297 fc2.n928 a_400_38200# 0.05fF
C3298 fc2.n929 a_400_38200# 0.03fF
C3299 fc2.n930 a_400_38200# 0.10fF
C3300 fc2.n931 a_400_38200# 0.17fF
C3301 fc2.n932 a_400_38200# 0.68fF
C3302 fc2.t358 a_400_38200# 0.02fF
C3303 fc2.n933 a_400_38200# 0.21fF
C3304 fc2.n934 a_400_38200# 0.31fF
C3305 fc2.n935 a_400_38200# 0.53fF
C3306 fc2.n936 a_400_38200# 0.10fF
C3307 fc2.t190 a_400_38200# 0.02fF
C3308 fc2.n937 a_400_38200# 0.12fF
C3309 fc2.n939 a_400_38200# 0.03fF
C3310 fc2.n940 a_400_38200# 0.01fF
C3311 fc2.n941 a_400_38200# 0.06fF
C3312 fc2.n942 a_400_38200# 0.24fF
C3313 fc2.n943 a_400_38200# 0.33fF
C3314 fc2.n944 a_400_38200# 0.05fF
C3315 fc2.n945 a_400_38200# 0.03fF
C3316 fc2.n946 a_400_38200# 0.13fF
C3317 fc2.n947 a_400_38200# 0.06fF
C3318 fc2.n948 a_400_38200# 0.11fF
C3319 fc2.n949 a_400_38200# 0.03fF
C3320 fc2.n950 a_400_38200# 0.05fF
C3321 fc2.n951 a_400_38200# 0.05fF
C3322 fc2.n952 a_400_38200# 0.09fF
C3323 fc2.n953 a_400_38200# 0.03fF
C3324 fc2.n954 a_400_38200# 0.07fF
C3325 fc2.n955 a_400_38200# 0.32fF
C3326 fc2.n956 a_400_38200# 0.47fF
C3327 fc2.n957 a_400_38200# 0.29fF
C3328 fc2.n958 a_400_38200# 3.32fF
C3329 fc2.t312 a_400_38200# 0.02fF
C3330 fc2.n959 a_400_38200# 0.10fF
C3331 fc2.n960 a_400_38200# 0.12fF
C3332 fc2.t238 a_400_38200# 0.02fF
C3333 fc2.n962 a_400_38200# 0.21fF
C3334 fc2.n963 a_400_38200# 0.80fF
C3335 fc2.n964 a_400_38200# 0.04fF
C3336 fc2.n965 a_400_38200# 0.46fF
C3337 fc2.n966 a_400_38200# 0.52fF
C3338 fc2.n967 a_400_38200# 0.46fF
C3339 fc2.n968 a_400_38200# 1.04fF
C3340 fc2.n969 a_400_38200# 0.12fF
C3341 fc2.n970 a_400_38200# 0.52fF
C3342 fc2.n971 a_400_38200# 0.10fF
C3343 fc2.t321 a_400_38200# 0.02fF
C3344 fc2.n972 a_400_38200# 0.12fF
C3345 fc2.t121 a_400_38200# 0.02fF
C3346 fc2.n974 a_400_38200# 0.21fF
C3347 fc2.n975 a_400_38200# 0.31fF
C3348 fc2.n976 a_400_38200# 0.53fF
C3349 fc2.n977 a_400_38200# 0.05fF
C3350 fc2.n978 a_400_38200# 0.17fF
C3351 fc2.n979 a_400_38200# 0.06fF
C3352 fc2.n980 a_400_38200# 0.03fF
C3353 fc2.n981 a_400_38200# 0.10fF
C3354 fc2.n982 a_400_38200# 0.17fF
C3355 fc2.n983 a_400_38200# 0.69fF
C3356 fc2.n984 a_400_38200# 0.05fF
C3357 fc2.n985 a_400_38200# 0.07fF
C3358 fc2.n986 a_400_38200# 1.00fF
C3359 fc2.n987 a_400_38200# 0.12fF
C3360 fc2.n988 a_400_38200# 3.32fF
C3361 fc2.t48 a_400_38200# 0.02fF
C3362 fc2.n989 a_400_38200# 0.10fF
C3363 fc2.n990 a_400_38200# 0.12fF
C3364 fc2.t368 a_400_38200# 0.02fF
C3365 fc2.n992 a_400_38200# 0.21fF
C3366 fc2.n993 a_400_38200# 0.80fF
C3367 fc2.n994 a_400_38200# 0.04fF
C3368 fc2.t47 a_400_38200# 16.88fF
C3369 fc2.t183 a_400_38200# 0.02fF
C3370 fc2.n995 a_400_38200# 0.01fF
C3371 fc2.n996 a_400_38200# 0.22fF
C3372 fc2.t113 a_400_38200# 0.02fF
C3373 fc2.n998 a_400_38200# 1.04fF
C3374 fc2.n999 a_400_38200# 0.04fF
C3375 fc2.t229 a_400_38200# 0.02fF
C3376 fc2.n1000 a_400_38200# 0.56fF
C3377 fc2.n1001 a_400_38200# 0.53fF
C3378 fc2.n1002 a_400_38200# 0.52fF
C3379 fc2.n1003 a_400_38200# 0.15fF
C3380 fc2.n1004 a_400_38200# 0.77fF
C3381 fc2.n1005 a_400_38200# 0.52fF
C3382 fc2.n1006 a_400_38200# 0.07fF
C3383 fc2.n1007 a_400_38200# 1.89fF
C3384 fc2.n1008 a_400_38200# 0.52fF
C3385 fc2.n1009 a_400_38200# 0.19fF
C3386 fc2.n1010 a_400_38200# 1.28fF
C3387 fc2.t26 a_400_38200# 7.96fF
C3388 fc2.n1012 a_400_38200# 7.30fF
C3389 fc2.n1014 a_400_38200# 1.22fF
C3390 fc2.n1015 a_400_38200# 3.88fF
C3391 fc2.n1016 a_400_38200# 2.29fF
C3392 fc2.n1017 a_400_38200# 3.86fF
C3393 fc2.n1018 a_400_38200# 2.19fF
C3394 fc2.t111 a_400_38200# 0.02fF
C3395 fc2.n1019 a_400_38200# 0.56fF
C3396 fc2.n1020 a_400_38200# 0.53fF
C3397 fc2.n1021 a_400_38200# 2.57fF
C3398 fc2.n1022 a_400_38200# 1.36fF
C3399 fc2.n1023 a_400_38200# 0.79fF
C3400 fc2.n1024 a_400_38200# 0.03fF
C3401 fc2.n1025 a_400_38200# 0.05fF
C3402 fc2.n1026 a_400_38200# 0.05fF
C3403 fc2.n1027 a_400_38200# 0.07fF
C3404 fc2.n1028 a_400_38200# 0.15fF
C3405 fc2.n1029 a_400_38200# 0.05fF
C3406 fc2.n1030 a_400_38200# 0.03fF
C3407 fc2.n1031 a_400_38200# 0.07fF
C3408 fc2.n1032 a_400_38200# 0.24fF
C3409 fc2.n1033 a_400_38200# 0.58fF
C3410 fc2.n1034 a_400_38200# 0.44fF
C3411 fc2.t374 a_400_38200# 0.02fF
C3412 fc2.n1035 a_400_38200# 0.21fF
C3413 fc2.n1036 a_400_38200# 0.31fF
C3414 fc2.n1037 a_400_38200# 0.53fF
C3415 fc2.n1038 a_400_38200# 0.10fF
C3416 fc2.t249 a_400_38200# 0.02fF
C3417 fc2.n1039 a_400_38200# 0.12fF
C3418 fc2.n1041 a_400_38200# 0.01fF
C3419 fc2.n1042 a_400_38200# 0.03fF
C3420 fc2.n1043 a_400_38200# 0.06fF
C3421 fc2.n1044 a_400_38200# 0.26fF
C3422 fc2.n1045 a_400_38200# 0.09fF
C3423 fc2.n1046 a_400_38200# 0.08fF
C3424 fc2.n1047 a_400_38200# 0.10fF
C3425 fc2.n1048 a_400_38200# 0.06fF
C3426 fc2.n1049 a_400_38200# 0.04fF
C3427 fc2.n1050 a_400_38200# 0.04fF
C3428 fc2.n1051 a_400_38200# 0.06fF
C3429 fc2.n1052 a_400_38200# 0.03fF
C3430 fc2.n1053 a_400_38200# 0.05fF
C3431 fc2.n1054 a_400_38200# 0.15fF
C3432 fc2.n1055 a_400_38200# 0.13fF
C3433 fc2.n1056 a_400_38200# 0.11fF
C3434 fc2.n1057 a_400_38200# 0.50fF
C3435 fc2.n1058 a_400_38200# 0.03fF
C3436 fc2.n1059 a_400_38200# 0.22fF
C3437 fc2.n1060 a_400_38200# 0.09fF
C3438 fc2.n1061 a_400_38200# 0.11fF
C3439 fc2.n1062 a_400_38200# 0.09fF
C3440 fc2.n1063 a_400_38200# 1.55fF
C3441 fc2.t294 a_400_38200# 0.02fF
C3442 fc2.n1064 a_400_38200# 0.21fF
C3443 fc2.n1065 a_400_38200# 0.80fF
C3444 fc2.n1066 a_400_38200# 0.04fF
C3445 fc2.t150 a_400_38200# 0.02fF
C3446 fc2.n1067 a_400_38200# 0.10fF
C3447 fc2.n1068 a_400_38200# 0.12fF
C3448 fc2.n1070 a_400_38200# 0.26fF
C3449 fc2.n1071 a_400_38200# 0.14fF
C3450 fc2.n1072 a_400_38200# 0.90fF
C3451 fc2.t265 a_400_38200# 0.02fF
C3452 fc2.n1073 a_400_38200# 0.21fF
C3453 fc2.n1074 a_400_38200# 0.31fF
C3454 fc2.n1075 a_400_38200# 0.53fF
C3455 fc2.t322 a_400_38200# 0.02fF
C3456 fc2.n1076 a_400_38200# 1.06fF
C3457 fc2.n1077 a_400_38200# 0.03fF
C3458 fc2.n1078 a_400_38200# 0.07fF
C3459 fc2.n1079 a_400_38200# 0.03fF
C3460 fc2.n1080 a_400_38200# 0.06fF
C3461 fc2.n1081 a_400_38200# 0.05fF
C3462 fc2.n1082 a_400_38200# 0.06fF
C3463 fc2.n1083 a_400_38200# 0.64fF
C3464 fc2.n1084 a_400_38200# 0.79fF
C3465 fc2.n1085 a_400_38200# 1.01fF
C3466 fc2.n1086 a_400_38200# 1.29fF
C3467 fc2.t41 a_400_38200# 7.96fF
C3468 fc2.n1087 a_400_38200# 9.42fF
C3469 fc2.n1089 a_400_38200# 0.33fF
C3470 fc2.n1090 a_400_38200# 0.20fF
C3471 fc2.n1091 a_400_38200# 3.05fF
C3472 fc2.n1092 a_400_38200# 1.86fF
C3473 fc2.n1093 a_400_38200# 0.03fF
C3474 fc2.n1094 a_400_38200# 0.04fF
C3475 fc2.n1095 a_400_38200# 0.08fF
C3476 fc2.n1096 a_400_38200# 0.06fF
C3477 fc2.n1097 a_400_38200# 0.05fF
C3478 fc2.n1098 a_400_38200# 0.06fF
C3479 fc2.n1099 a_400_38200# 0.08fF
C3480 fc2.n1100 a_400_38200# 0.11fF
C3481 fc2.n1101 a_400_38200# 0.68fF
C3482 fc2.n1102 a_400_38200# 0.26fF
C3483 fc2.n1103 a_400_38200# 0.72fF
C3484 fc2.n1104 a_400_38200# 0.65fF
C3485 fc2.n1105 a_400_38200# 3.60fF
C3486 fc2.n1106 a_400_38200# 0.22fF
C3487 fc2.n1107 a_400_38200# 0.01fF
C3488 fc2.t158 a_400_38200# 0.02fF
C3489 fc2.n1108 a_400_38200# 0.22fF
C3490 fc2.t120 a_400_38200# 0.02fF
C3491 fc2.n1109 a_400_38200# 0.83fF
C3492 fc2.n1110 a_400_38200# 0.62fF
C3493 fc2.n1111 a_400_38200# 0.50fF
C3494 fc2.n1112 a_400_38200# 0.94fF
C3495 fc2.n1113 a_400_38200# 0.18fF
C3496 fc2.n1114 a_400_38200# 0.76fF
C3497 fc2.t254 a_400_38200# 0.02fF
C3498 fc2.n1115 a_400_38200# 0.21fF
C3499 fc2.n1116 a_400_38200# 0.31fF
C3500 fc2.n1117 a_400_38200# 0.53fF
C3501 fc2.n1118 a_400_38200# 0.10fF
C3502 fc2.t109 a_400_38200# 0.02fF
C3503 fc2.n1119 a_400_38200# 0.12fF
C3504 fc2.n1121 a_400_38200# 0.76fF
C3505 fc2.n1122 a_400_38200# 0.44fF
C3506 fc2.n1123 a_400_38200# 1.07fF
C3507 fc2.n1124 a_400_38200# 0.18fF
C3508 fc2.n1125 a_400_38200# 3.23fF
C3509 fc2.t42 a_400_38200# 0.02fF
C3510 fc2.n1126 a_400_38200# 0.21fF
C3511 fc2.n1127 a_400_38200# 0.80fF
C3512 fc2.n1128 a_400_38200# 0.04fF
C3513 fc2.t119 a_400_38200# 0.02fF
C3514 fc2.n1129 a_400_38200# 0.10fF
C3515 fc2.n1130 a_400_38200# 0.12fF
C3516 fc2.n1132 a_400_38200# 7.70fF
C3517 fc2.n1133 a_400_38200# 1.07fF
C3518 fc2.n1134 a_400_38200# 1.53fF
C3519 fc2.t192 a_400_38200# 0.02fF
C3520 fc2.n1135 a_400_38200# 0.21fF
C3521 fc2.n1136 a_400_38200# 0.31fF
C3522 fc2.n1137 a_400_38200# 0.53fF
C3523 fc2.n1138 a_400_38200# 0.10fF
C3524 fc2.t11 a_400_38200# 0.02fF
C3525 fc2.n1139 a_400_38200# 0.12fF
C3526 fc2.n1141 a_400_38200# 0.01fF
C3527 fc2.n1142 a_400_38200# 0.03fF
C3528 fc2.n1143 a_400_38200# 0.06fF
C3529 fc2.n1144 a_400_38200# 0.24fF
C3530 fc2.n1145 a_400_38200# 0.33fF
C3531 fc2.n1146 a_400_38200# 0.13fF
C3532 fc2.n1147 a_400_38200# 0.06fF
C3533 fc2.n1148 a_400_38200# 0.11fF
C3534 fc2.n1149 a_400_38200# 0.03fF
C3535 fc2.n1150 a_400_38200# 0.07fF
C3536 fc2.n1151 a_400_38200# 0.05fF
C3537 fc2.n1152 a_400_38200# 0.05fF
C3538 fc2.n1153 a_400_38200# 0.09fF
C3539 fc2.n1154 a_400_38200# 0.32fF
C3540 fc2.n1155 a_400_38200# 0.47fF
C3541 fc2.n1156 a_400_38200# 0.29fF
C3542 fc2.n1157 a_400_38200# 1.90fF
C3543 fc2.t55 a_400_38200# 0.02fF
C3544 fc2.n1158 a_400_38200# 0.10fF
C3545 fc2.n1159 a_400_38200# 0.12fF
C3546 fc2.t357 a_400_38200# 0.02fF
C3547 fc2.n1161 a_400_38200# 0.21fF
C3548 fc2.n1162 a_400_38200# 0.80fF
C3549 fc2.n1163 a_400_38200# 0.04fF
C3550 fc2.n1164 a_400_38200# 0.93fF
C3551 fc2.n1165 a_400_38200# 0.18fF
C3552 fc2.n1166 a_400_38200# 0.10fF
C3553 fc2.t346 a_400_38200# 0.02fF
C3554 fc2.n1167 a_400_38200# 0.12fF
C3555 fc2.t145 a_400_38200# 0.02fF
C3556 fc2.n1169 a_400_38200# 0.21fF
C3557 fc2.n1170 a_400_38200# 0.31fF
C3558 fc2.n1171 a_400_38200# 0.53fF
C3559 fc2.n1172 a_400_38200# 0.02fF
C3560 fc2.n1173 a_400_38200# 0.18fF
C3561 fc2.n1174 a_400_38200# 0.12fF
C3562 fc2.n1175 a_400_38200# 1.21fF
C3563 fc2.n1176 a_400_38200# 0.06fF
C3564 fc2.n1177 a_400_38200# 0.31fF
C3565 fc2.n1178 a_400_38200# 0.06fF
C3566 fc2.n1179 a_400_38200# 3.43fF
C3567 fc2.t354 a_400_38200# 0.02fF
C3568 fc2.n1180 a_400_38200# 0.10fF
C3569 fc2.n1181 a_400_38200# 0.12fF
C3570 fc2.t310 a_400_38200# 0.02fF
C3571 fc2.n1183 a_400_38200# 0.21fF
C3572 fc2.n1184 a_400_38200# 0.80fF
C3573 fc2.n1185 a_400_38200# 0.04fF
C3574 fc2.t10 a_400_38200# 17.22fF
C3575 fc2.t59 a_400_38200# 0.02fF
C3576 fc2.n1186 a_400_38200# 0.21fF
C3577 fc2.n1187 a_400_38200# 0.80fF
C3578 fc2.n1188 a_400_38200# 0.04fF
C3579 fc2.t130 a_400_38200# 0.02fF
C3580 fc2.n1189 a_400_38200# 0.10fF
C3581 fc2.n1190 a_400_38200# 0.12fF
C3582 fc2.n1192 a_400_38200# 0.10fF
C3583 fc2.t102 a_400_38200# 0.02fF
C3584 fc2.n1193 a_400_38200# 0.12fF
C3585 fc2.n1195 a_400_38200# 0.01fF
C3586 fc2.n1196 a_400_38200# 0.03fF
C3587 fc2.n1197 a_400_38200# 0.06fF
C3588 fc2.n1198 a_400_38200# 0.24fF
C3589 fc2.n1199 a_400_38200# 0.33fF
C3590 fc2.n1200 a_400_38200# 0.13fF
C3591 fc2.n1201 a_400_38200# 0.06fF
C3592 fc2.n1202 a_400_38200# 0.11fF
C3593 fc2.n1203 a_400_38200# 0.03fF
C3594 fc2.n1204 a_400_38200# 0.07fF
C3595 fc2.n1205 a_400_38200# 0.05fF
C3596 fc2.n1206 a_400_38200# 0.05fF
C3597 fc2.n1207 a_400_38200# 0.09fF
C3598 fc2.n1208 a_400_38200# 0.32fF
C3599 fc2.n1209 a_400_38200# 0.47fF
C3600 fc2.n1210 a_400_38200# 0.29fF
C3601 fc2.n1211 a_400_38200# 3.80fF
C3602 fc2.n1212 a_400_38200# 1.94fF
C3603 fc2.n1213 a_400_38200# 0.12fF
C3604 fc2.n1214 a_400_38200# 1.18fF
C3605 fc2.n1215 a_400_38200# 0.13fF
C3606 fc2.n1216 a_400_38200# 0.37fF
C3607 fc2.n1217 a_400_38200# 0.14fF
C3608 fc2.n1218 a_400_38200# 0.17fF
C3609 fc2.n1219 a_400_38200# 0.11fF
C3610 fc2.n1220 a_400_38200# 0.11fF
C3611 fc2.n1221 a_400_38200# 0.21fF
C3612 fc2.n1222 a_400_38200# 0.71fF
C3613 fc2.t246 a_400_38200# 0.02fF
C3614 fc2.n1223 a_400_38200# 0.21fF
C3615 fc2.n1224 a_400_38200# 0.31fF
C3616 fc2.n1225 a_400_38200# 0.53fF
C3617 fc2.n1226 a_400_38200# 0.10fF
C3618 fc2.t124 a_400_38200# 0.02fF
C3619 fc2.n1227 a_400_38200# 0.12fF
C3620 fc2.n1229 a_400_38200# 0.01fF
C3621 fc2.n1230 a_400_38200# 0.03fF
C3622 fc2.n1231 a_400_38200# 0.06fF
C3623 fc2.n1232 a_400_38200# 0.26fF
C3624 fc2.n1233 a_400_38200# 0.09fF
C3625 fc2.n1234 a_400_38200# 0.08fF
C3626 fc2.n1235 a_400_38200# 0.10fF
C3627 fc2.n1236 a_400_38200# 0.06fF
C3628 fc2.n1237 a_400_38200# 0.04fF
C3629 fc2.n1238 a_400_38200# 0.04fF
C3630 fc2.n1239 a_400_38200# 0.06fF
C3631 fc2.n1240 a_400_38200# 0.03fF
C3632 fc2.n1241 a_400_38200# 0.05fF
C3633 fc2.n1242 a_400_38200# 0.15fF
C3634 fc2.n1243 a_400_38200# 0.13fF
C3635 fc2.n1244 a_400_38200# 0.11fF
C3636 fc2.n1245 a_400_38200# 0.50fF
C3637 fc2.n1246 a_400_38200# 0.03fF
C3638 fc2.n1247 a_400_38200# 0.22fF
C3639 fc2.n1248 a_400_38200# 0.09fF
C3640 fc2.n1249 a_400_38200# 0.11fF
C3641 fc2.n1250 a_400_38200# 0.09fF
C3642 fc2.n1251 a_400_38200# 1.54fF
C3643 fc2.t166 a_400_38200# 0.02fF
C3644 fc2.n1252 a_400_38200# 0.21fF
C3645 fc2.n1253 a_400_38200# 0.80fF
C3646 fc2.n1254 a_400_38200# 0.04fF
C3647 fc2.t215 a_400_38200# 0.02fF
C3648 fc2.n1255 a_400_38200# 0.10fF
C3649 fc2.n1256 a_400_38200# 0.12fF
C3650 fc2.n1258 a_400_38200# 0.26fF
C3651 fc2.n1259 a_400_38200# 0.14fF
C3652 fc2.n1260 a_400_38200# 0.90fF
C3653 fc2.t138 a_400_38200# 0.02fF
C3654 fc2.n1261 a_400_38200# 0.21fF
C3655 fc2.n1262 a_400_38200# 0.31fF
C3656 fc2.n1263 a_400_38200# 0.53fF
C3657 fc2.t301 a_400_38200# 0.02fF
C3658 fc2.n1264 a_400_38200# 0.21fF
C3659 fc2.n1265 a_400_38200# 0.80fF
C3660 fc2.n1266 a_400_38200# 0.04fF
C3661 fc2.t370 a_400_38200# 0.02fF
C3662 fc2.n1267 a_400_38200# 0.10fF
C3663 fc2.n1268 a_400_38200# 0.12fF
C3664 fc2.n1270 a_400_38200# 0.10fF
C3665 fc2.t341 a_400_38200# 0.02fF
C3666 fc2.n1271 a_400_38200# 0.12fF
C3667 fc2.n1273 a_400_38200# 0.01fF
C3668 fc2.n1274 a_400_38200# 0.03fF
C3669 fc2.n1275 a_400_38200# 0.06fF
C3670 fc2.n1276 a_400_38200# 0.24fF
C3671 fc2.n1277 a_400_38200# 0.33fF
C3672 fc2.n1278 a_400_38200# 0.13fF
C3673 fc2.n1279 a_400_38200# 0.06fF
C3674 fc2.n1280 a_400_38200# 0.11fF
C3675 fc2.n1281 a_400_38200# 0.03fF
C3676 fc2.n1282 a_400_38200# 0.07fF
C3677 fc2.n1283 a_400_38200# 0.05fF
C3678 fc2.n1284 a_400_38200# 0.05fF
C3679 fc2.n1285 a_400_38200# 0.09fF
C3680 fc2.n1286 a_400_38200# 0.32fF
C3681 fc2.n1287 a_400_38200# 0.47fF
C3682 fc2.n1288 a_400_38200# 0.29fF
C3683 fc2.n1289 a_400_38200# 3.44fF
C3684 fc2.n1290 a_400_38200# 1.94fF
C3685 fc2.n1291 a_400_38200# 0.12fF
C3686 fc2.n1292 a_400_38200# 1.18fF
C3687 fc2.n1293 a_400_38200# 0.13fF
C3688 fc2.n1294 a_400_38200# 0.37fF
C3689 fc2.n1295 a_400_38200# 0.14fF
C3690 fc2.n1296 a_400_38200# 0.17fF
C3691 fc2.n1297 a_400_38200# 0.11fF
C3692 fc2.n1298 a_400_38200# 0.11fF
C3693 fc2.n1299 a_400_38200# 0.21fF
C3694 fc2.n1300 a_400_38200# 0.71fF
C3695 fc2.t122 a_400_38200# 0.02fF
C3696 fc2.n1301 a_400_38200# 0.21fF
C3697 fc2.n1302 a_400_38200# 0.31fF
C3698 fc2.n1303 a_400_38200# 0.53fF
C3699 fc2.n1304 a_400_38200# 0.10fF
C3700 fc2.t366 a_400_38200# 0.02fF
C3701 fc2.n1305 a_400_38200# 0.12fF
C3702 fc2.n1307 a_400_38200# 0.01fF
C3703 fc2.n1308 a_400_38200# 0.03fF
C3704 fc2.n1309 a_400_38200# 0.06fF
C3705 fc2.n1310 a_400_38200# 0.26fF
C3706 fc2.n1311 a_400_38200# 0.09fF
C3707 fc2.n1312 a_400_38200# 0.08fF
C3708 fc2.n1313 a_400_38200# 0.10fF
C3709 fc2.n1314 a_400_38200# 0.06fF
C3710 fc2.n1315 a_400_38200# 0.04fF
C3711 fc2.n1316 a_400_38200# 0.04fF
C3712 fc2.n1317 a_400_38200# 0.06fF
C3713 fc2.n1318 a_400_38200# 0.03fF
C3714 fc2.n1319 a_400_38200# 0.05fF
C3715 fc2.n1320 a_400_38200# 0.15fF
C3716 fc2.n1321 a_400_38200# 0.13fF
C3717 fc2.n1322 a_400_38200# 0.11fF
C3718 fc2.n1323 a_400_38200# 0.50fF
C3719 fc2.n1324 a_400_38200# 0.03fF
C3720 fc2.n1325 a_400_38200# 0.22fF
C3721 fc2.n1326 a_400_38200# 0.09fF
C3722 fc2.n1327 a_400_38200# 0.11fF
C3723 fc2.n1328 a_400_38200# 0.09fF
C3724 fc2.n1329 a_400_38200# 1.54fF
C3725 fc2.t32 a_400_38200# 0.02fF
C3726 fc2.n1330 a_400_38200# 0.21fF
C3727 fc2.n1331 a_400_38200# 0.80fF
C3728 fc2.n1332 a_400_38200# 0.04fF
C3729 fc2.t95 a_400_38200# 0.02fF
C3730 fc2.n1333 a_400_38200# 0.10fF
C3731 fc2.n1334 a_400_38200# 0.12fF
C3732 fc2.n1336 a_400_38200# 0.26fF
C3733 fc2.n1337 a_400_38200# 0.14fF
C3734 fc2.n1338 a_400_38200# 0.98fF
C3735 fc2.t381 a_400_38200# 0.02fF
C3736 fc2.n1339 a_400_38200# 0.21fF
C3737 fc2.n1340 a_400_38200# 0.31fF
C3738 fc2.n1341 a_400_38200# 0.53fF
C3739 fc2.t174 a_400_38200# 0.02fF
C3740 fc2.n1342 a_400_38200# 0.21fF
C3741 fc2.n1343 a_400_38200# 0.80fF
C3742 fc2.n1344 a_400_38200# 0.04fF
C3743 fc2.t242 a_400_38200# 0.02fF
C3744 fc2.n1345 a_400_38200# 0.10fF
C3745 fc2.n1346 a_400_38200# 0.12fF
C3746 fc2.n1348 a_400_38200# 0.10fF
C3747 fc2.t210 a_400_38200# 0.02fF
C3748 fc2.n1349 a_400_38200# 0.12fF
C3749 fc2.n1351 a_400_38200# 0.01fF
C3750 fc2.n1352 a_400_38200# 0.03fF
C3751 fc2.n1353 a_400_38200# 0.06fF
C3752 fc2.n1354 a_400_38200# 0.24fF
C3753 fc2.n1355 a_400_38200# 0.33fF
C3754 fc2.n1356 a_400_38200# 0.13fF
C3755 fc2.n1357 a_400_38200# 0.06fF
C3756 fc2.n1358 a_400_38200# 0.11fF
C3757 fc2.n1359 a_400_38200# 0.03fF
C3758 fc2.n1360 a_400_38200# 0.07fF
C3759 fc2.n1361 a_400_38200# 0.05fF
C3760 fc2.n1362 a_400_38200# 0.05fF
C3761 fc2.n1363 a_400_38200# 0.09fF
C3762 fc2.n1364 a_400_38200# 0.32fF
C3763 fc2.n1365 a_400_38200# 0.47fF
C3764 fc2.n1366 a_400_38200# 0.29fF
C3765 fc2.n1367 a_400_38200# 3.41fF
C3766 fc2.n1368 a_400_38200# 1.94fF
C3767 fc2.n1369 a_400_38200# 0.13fF
C3768 fc2.n1370 a_400_38200# 0.94fF
C3769 fc2.n1371 a_400_38200# 0.13fF
C3770 fc2.n1372 a_400_38200# 0.37fF
C3771 fc2.n1373 a_400_38200# 0.14fF
C3772 fc2.n1374 a_400_38200# 0.16fF
C3773 fc2.n1375 a_400_38200# 0.11fF
C3774 fc2.n1376 a_400_38200# 0.11fF
C3775 fc2.n1377 a_400_38200# 0.24fF
C3776 fc2.n1378 a_400_38200# 0.69fF
C3777 fc2.t363 a_400_38200# 0.02fF
C3778 fc2.n1379 a_400_38200# 0.21fF
C3779 fc2.n1380 a_400_38200# 0.31fF
C3780 fc2.n1381 a_400_38200# 0.53fF
C3781 fc2.n1382 a_400_38200# 0.10fF
C3782 fc2.t236 a_400_38200# 0.02fF
C3783 fc2.n1383 a_400_38200# 0.12fF
C3784 fc2.n1385 a_400_38200# 0.01fF
C3785 fc2.n1386 a_400_38200# 0.03fF
C3786 fc2.n1387 a_400_38200# 0.06fF
C3787 fc2.n1388 a_400_38200# 0.26fF
C3788 fc2.n1389 a_400_38200# 0.09fF
C3789 fc2.n1390 a_400_38200# 0.08fF
C3790 fc2.n1391 a_400_38200# 0.10fF
C3791 fc2.n1392 a_400_38200# 0.06fF
C3792 fc2.n1393 a_400_38200# 0.04fF
C3793 fc2.n1394 a_400_38200# 0.04fF
C3794 fc2.n1395 a_400_38200# 0.06fF
C3795 fc2.n1396 a_400_38200# 0.03fF
C3796 fc2.n1397 a_400_38200# 0.05fF
C3797 fc2.n1398 a_400_38200# 0.15fF
C3798 fc2.n1399 a_400_38200# 0.13fF
C3799 fc2.n1400 a_400_38200# 0.11fF
C3800 fc2.n1401 a_400_38200# 0.50fF
C3801 fc2.n1402 a_400_38200# 0.03fF
C3802 fc2.n1403 a_400_38200# 0.22fF
C3803 fc2.n1404 a_400_38200# 0.09fF
C3804 fc2.n1405 a_400_38200# 0.11fF
C3805 fc2.n1406 a_400_38200# 0.09fF
C3806 fc2.n1407 a_400_38200# 1.54fF
C3807 fc2.t282 a_400_38200# 0.02fF
C3808 fc2.n1408 a_400_38200# 0.21fF
C3809 fc2.n1409 a_400_38200# 0.80fF
C3810 fc2.n1410 a_400_38200# 0.04fF
C3811 fc2.t336 a_400_38200# 0.02fF
C3812 fc2.n1411 a_400_38200# 0.10fF
C3813 fc2.n1412 a_400_38200# 0.12fF
C3814 fc2.n1414 a_400_38200# 1.68fF
C3815 fc2.n1415 a_400_38200# 0.05fF
C3816 fc2.n1416 a_400_38200# 0.07fF
C3817 fc2.n1417 a_400_38200# 1.10fF
C3818 fc2.n1418 a_400_38200# 0.12fF
C3819 fc2.n1419 a_400_38200# 0.05fF
C3820 fc2.n1420 a_400_38200# 0.17fF
C3821 fc2.n1421 a_400_38200# 0.06fF
C3822 fc2.n1422 a_400_38200# 0.03fF
C3823 fc2.n1423 a_400_38200# 0.10fF
C3824 fc2.n1424 a_400_38200# 0.17fF
C3825 fc2.n1425 a_400_38200# 0.68fF
C3826 fc2.t232 a_400_38200# 0.02fF
C3827 fc2.n1426 a_400_38200# 0.21fF
C3828 fc2.n1427 a_400_38200# 0.31fF
C3829 fc2.n1428 a_400_38200# 0.53fF
C3830 fc2.n1429 a_400_38200# 0.10fF
C3831 fc2.t112 a_400_38200# 0.02fF
C3832 fc2.n1430 a_400_38200# 0.12fF
C3833 fc2.n1432 a_400_38200# 0.76fF
C3834 fc2.n1433 a_400_38200# 0.44fF
C3835 fc2.n1434 a_400_38200# 0.16fF
C3836 fc2.n1435 a_400_38200# 0.26fF
C3837 fc2.n1436 a_400_38200# 0.75fF
C3838 fc2.n1437 a_400_38200# 0.18fF
C3839 fc2.n1438 a_400_38200# 1.51fF
C3840 fc2.t155 a_400_38200# 0.02fF
C3841 fc2.n1439 a_400_38200# 0.21fF
C3842 fc2.n1440 a_400_38200# 0.80fF
C3843 fc2.n1441 a_400_38200# 0.04fF
C3844 fc2.t224 a_400_38200# 0.02fF
C3845 fc2.n1442 a_400_38200# 0.10fF
C3846 fc2.n1443 a_400_38200# 0.12fF
C3847 fc2.t21 a_400_38200# 8.91fF
C3848 fc2.n1445 a_400_38200# 7.70fF
C3849 fc2.n1446 a_400_38200# 0.12fF
C3850 fc2.n1447 a_400_38200# 0.06fF
C3851 fc2.n1448 a_400_38200# 0.03fF
C3852 fc2.n1449 a_400_38200# 0.04fF
C3853 fc2.n1450 a_400_38200# 0.29fF
C3854 fc2.n1451 a_400_38200# 0.04fF
C3855 fc2.n1452 a_400_38200# 0.05fF
C3856 fc2.n1453 a_400_38200# 0.07fF
C3857 fc2.n1454 a_400_38200# 0.05fF
C3858 fc2.n1455 a_400_38200# 0.05fF
C3859 fc2.n1456 a_400_38200# 0.05fF
C3860 fc2.n1457 a_400_38200# 0.06fF
C3861 fc2.n1458 a_400_38200# 0.12fF
C3862 fc2.n1459 a_400_38200# 0.10fF
C3863 fc2.n1460 a_400_38200# 0.10fF
C3864 fc2.n1461 a_400_38200# 0.02fF
C3865 fc2.n1462 a_400_38200# 0.32fF
C3866 fc2.n1463 a_400_38200# 0.40fF
C3867 fc2.n1464 a_400_38200# 0.22fF
C3868 fc2.n1465 a_400_38200# 0.11fF
C3869 fc2.n1466 a_400_38200# 0.25fF
C3870 fc2.n1467 a_400_38200# 0.03fF
C3871 fc2.t302 a_400_38200# 0.02fF
C3872 fc2.n1468 a_400_38200# 0.21fF
C3873 fc2.n1469 a_400_38200# 0.31fF
C3874 fc2.n1470 a_400_38200# 0.53fF
C3875 fc2.n1471 a_400_38200# 0.10fF
C3876 fc2.t177 a_400_38200# 0.02fF
C3877 fc2.n1472 a_400_38200# 0.12fF
C3878 fc2.n1474 a_400_38200# 0.02fF
C3879 fc2.n1475 a_400_38200# 0.03fF
C3880 fc2.n1476 a_400_38200# 0.07fF
C3881 fc2.n1477 a_400_38200# 0.07fF
C3882 fc2.n1478 a_400_38200# 0.15fF
C3883 fc2.n1479 a_400_38200# 0.03fF
C3884 fc2.n1480 a_400_38200# 0.05fF
C3885 fc2.n1481 a_400_38200# 0.05fF
C3886 fc2.n1482 a_400_38200# 0.05fF
C3887 fc2.n1483 a_400_38200# 0.25fF
C3888 fc2.n1484 a_400_38200# 0.55fF
C3889 fc2.n1485 a_400_38200# 0.01fF
C3890 fc2.n1486 a_400_38200# 0.09fF
C3891 fc2.n1487 a_400_38200# 0.30fF
C3892 fc2.n1488 a_400_38200# 0.03fF
C3893 fc2.n1489 a_400_38200# 0.10fF
C3894 fc2.n1490 a_400_38200# 0.05fF
C3895 fc2.n1491 a_400_38200# 0.15fF
C3896 fc2.n1492 a_400_38200# 0.18fF
C3897 fc2.n1493 a_400_38200# 0.26fF
C3898 fc2.n1494 a_400_38200# 3.12fF
C3899 fc2.t276 a_400_38200# 0.02fF
C3900 fc2.n1495 a_400_38200# 0.10fF
C3901 fc2.n1496 a_400_38200# 0.12fF
C3902 fc2.t219 a_400_38200# 0.02fF
C3903 fc2.n1498 a_400_38200# 0.21fF
C3904 fc2.n1499 a_400_38200# 0.80fF
C3905 fc2.n1500 a_400_38200# 0.04fF
C3906 fc2.t94 a_400_38200# 16.88fF
C3907 fc2.t7 a_400_38200# 0.02fF
C3908 fc2.n1501 a_400_38200# 1.04fF
C3909 fc2.n1502 a_400_38200# 0.04fF
C3910 fc2.t103 a_400_38200# 0.02fF
C3911 fc2.n1503 a_400_38200# 0.01fF
C3912 fc2.n1504 a_400_38200# 0.22fF
C3913 fc2.n1506 a_400_38200# 0.27fF
C3914 fc2.n1507 a_400_38200# 0.17fF
C3915 fc2.n1508 a_400_38200# 0.26fF
C3916 fc2.n1509 a_400_38200# 0.04fF
C3917 fc2.n1510 a_400_38200# 0.02fF
C3918 fc2.n1511 a_400_38200# 0.18fF
C3919 fc2.n1512 a_400_38200# 0.77fF
C3920 fc2.n1513 a_400_38200# 0.07fF
C3921 fc2.n1514 a_400_38200# 0.77fF
C3922 fc2.n1515 a_400_38200# 1.89fF
C3923 fc2.n1516 a_400_38200# 4.60fF
C3924 fc2.n1517 a_400_38200# 0.45fF
C3925 fc2.n1518 a_400_38200# 0.79fF
C3926 fc2.n1519 a_400_38200# 0.52fF
C3927 fc2.n1520 a_400_38200# 0.19fF
C3928 fc2.n1521 a_400_38200# 1.28fF
C3929 fc2.t6 a_400_38200# 7.96fF
C3930 fc2.n1523 a_400_38200# 7.30fF
C3931 fc2.n1525 a_400_38200# 1.22fF
C3932 fc2.n1526 a_400_38200# 0.18fF
C3933 fc2.n1527 a_400_38200# 5.12fF
C3934 fc2.n1528 a_400_38200# 1.20fF
C3935 fc2.n1529 a_400_38200# 0.09fF
C3936 fc2.n1530 a_400_38200# 1.61fF
C3937 fc2.n1531 a_400_38200# 1.85fF
C3938 fc2.n1532 a_400_38200# 0.52fF
C3939 fc2.n1533 a_400_38200# 0.15fF
C3940 fc2.n1534 a_400_38200# 0.52fF
C3941 fc2.n1535 a_400_38200# 0.07fF
C3942 fc2.n1536 a_400_38200# 1.89fF
C3943 fc2.n1537 a_400_38200# 0.52fF
C3944 fc2.n1538 a_400_38200# 0.19fF
C3945 fc2.n1539 a_400_38200# 1.28fF
C3946 fc2.t50 a_400_38200# 7.96fF
C3947 fc2.n1541 a_400_38200# 7.30fF
C3948 fc2.n1543 a_400_38200# 1.22fF
C3949 fc2.n1544 a_400_38200# 4.71fF
C3950 fc2.n1545 a_400_38200# 2.13fF
C3951 fc2.t188 a_400_38200# 0.02fF
C3952 fc2.n1546 a_400_38200# 0.56fF
C3953 fc2.n1547 a_400_38200# 0.53fF
C3954 fc2.n1548 a_400_38200# 1.68fF
C3955 fc2.n1549 a_400_38200# 0.05fF
C3956 fc2.n1550 a_400_38200# 0.06fF
C3957 fc2.n1551 a_400_38200# 1.08fF
C3958 fc2.n1552 a_400_38200# 0.12fF
C3959 fc2.n1553 a_400_38200# 0.05fF
C3960 fc2.n1554 a_400_38200# 0.16fF
C3961 fc2.n1555 a_400_38200# 0.03fF
C3962 fc2.n1556 a_400_38200# 0.08fF
C3963 fc2.n1557 a_400_38200# 0.16fF
C3964 fc2.n1558 a_400_38200# 0.71fF
C3965 fc2.t88 a_400_38200# 0.02fF
C3966 fc2.n1559 a_400_38200# 0.21fF
C3967 fc2.n1560 a_400_38200# 0.31fF
C3968 fc2.n1561 a_400_38200# 0.53fF
C3969 fc2.n1562 a_400_38200# 0.10fF
C3970 fc2.t291 a_400_38200# 0.02fF
C3971 fc2.n1563 a_400_38200# 0.12fF
C3972 fc2.n1565 a_400_38200# 0.01fF
C3973 fc2.n1566 a_400_38200# 0.03fF
C3974 fc2.n1567 a_400_38200# 0.06fF
C3975 fc2.n1568 a_400_38200# 0.24fF
C3976 fc2.n1569 a_400_38200# 0.05fF
C3977 fc2.n1570 a_400_38200# 0.03fF
C3978 fc2.n1571 a_400_38200# 0.33fF
C3979 fc2.n1572 a_400_38200# 0.13fF
C3980 fc2.n1573 a_400_38200# 0.06fF
C3981 fc2.n1574 a_400_38200# 0.11fF
C3982 fc2.n1575 a_400_38200# 0.03fF
C3983 fc2.n1576 a_400_38200# 0.07fF
C3984 fc2.n1577 a_400_38200# 0.03fF
C3985 fc2.n1578 a_400_38200# 0.05fF
C3986 fc2.n1579 a_400_38200# 0.05fF
C3987 fc2.n1580 a_400_38200# 0.09fF
C3988 fc2.n1581 a_400_38200# 0.32fF
C3989 fc2.n1582 a_400_38200# 0.47fF
C3990 fc2.n1583 a_400_38200# 0.29fF
C3991 fc2.n1584 a_400_38200# 1.87fF
C3992 fc2.t335 a_400_38200# 0.02fF
C3993 fc2.n1585 a_400_38200# 0.21fF
C3994 fc2.n1586 a_400_38200# 0.80fF
C3995 fc2.n1587 a_400_38200# 0.04fF
C3996 fc2.t189 a_400_38200# 0.02fF
C3997 fc2.n1588 a_400_38200# 0.10fF
C3998 fc2.n1589 a_400_38200# 0.12fF
C3999 fc2.n1591 a_400_38200# 0.25fF
C4000 fc2.n1592 a_400_38200# 0.75fF
C4001 fc2.n1593 a_400_38200# 0.18fF
C4002 fc2.n1594 a_400_38200# 0.42fF
C4003 fc2.n1595 a_400_38200# 0.79fF
C4004 fc2.t309 a_400_38200# 0.02fF
C4005 fc2.n1596 a_400_38200# 0.21fF
C4006 fc2.n1597 a_400_38200# 0.31fF
C4007 fc2.n1598 a_400_38200# 0.53fF
C4008 fc2.t106 a_400_38200# 0.02fF
C4009 fc2.n1599 a_400_38200# 0.21fF
C4010 fc2.n1600 a_400_38200# 0.80fF
C4011 fc2.n1601 a_400_38200# 0.04fF
C4012 fc2.t168 a_400_38200# 0.02fF
C4013 fc2.n1602 a_400_38200# 0.10fF
C4014 fc2.n1603 a_400_38200# 0.12fF
C4015 fc2.n1605 a_400_38200# 0.10fF
C4016 fc2.t139 a_400_38200# 0.02fF
C4017 fc2.n1606 a_400_38200# 0.12fF
C4018 fc2.n1608 a_400_38200# 0.01fF
C4019 fc2.n1609 a_400_38200# 0.03fF
C4020 fc2.n1610 a_400_38200# 0.06fF
C4021 fc2.n1611 a_400_38200# 0.24fF
C4022 fc2.n1612 a_400_38200# 0.33fF
C4023 fc2.n1613 a_400_38200# 0.13fF
C4024 fc2.n1614 a_400_38200# 0.06fF
C4025 fc2.n1615 a_400_38200# 0.11fF
C4026 fc2.n1616 a_400_38200# 0.03fF
C4027 fc2.n1617 a_400_38200# 0.07fF
C4028 fc2.n1618 a_400_38200# 0.05fF
C4029 fc2.n1619 a_400_38200# 0.09fF
C4030 fc2.n1620 a_400_38200# 0.32fF
C4031 fc2.n1621 a_400_38200# 0.47fF
C4032 fc2.n1622 a_400_38200# 0.29fF
C4033 fc2.n1623 a_400_38200# 3.69fF
C4034 fc2.n1624 a_400_38200# 1.75fF
C4035 fc2.n1625 a_400_38200# 0.05fF
C4036 fc2.n1626 a_400_38200# 0.06fF
C4037 fc2.n1627 a_400_38200# 1.08fF
C4038 fc2.n1628 a_400_38200# 0.12fF
C4039 fc2.n1629 a_400_38200# 0.05fF
C4040 fc2.n1630 a_400_38200# 0.16fF
C4041 fc2.n1631 a_400_38200# 0.03fF
C4042 fc2.n1632 a_400_38200# 0.08fF
C4043 fc2.n1633 a_400_38200# 0.16fF
C4044 fc2.n1634 a_400_38200# 0.71fF
C4045 fc2.t329 a_400_38200# 0.02fF
C4046 fc2.n1635 a_400_38200# 0.21fF
C4047 fc2.n1636 a_400_38200# 0.31fF
C4048 fc2.n1637 a_400_38200# 0.53fF
C4049 fc2.n1638 a_400_38200# 0.10fF
C4050 fc2.t163 a_400_38200# 0.02fF
C4051 fc2.n1639 a_400_38200# 0.12fF
C4052 fc2.n1641 a_400_38200# 0.01fF
C4053 fc2.n1642 a_400_38200# 0.03fF
C4054 fc2.n1643 a_400_38200# 0.06fF
C4055 fc2.n1644 a_400_38200# 0.24fF
C4056 fc2.n1645 a_400_38200# 0.05fF
C4057 fc2.n1646 a_400_38200# 0.03fF
C4058 fc2.n1647 a_400_38200# 0.33fF
C4059 fc2.n1648 a_400_38200# 0.13fF
C4060 fc2.n1649 a_400_38200# 0.06fF
C4061 fc2.n1650 a_400_38200# 0.11fF
C4062 fc2.n1651 a_400_38200# 0.03fF
C4063 fc2.n1652 a_400_38200# 0.07fF
C4064 fc2.n1653 a_400_38200# 0.03fF
C4065 fc2.n1654 a_400_38200# 0.05fF
C4066 fc2.n1655 a_400_38200# 0.05fF
C4067 fc2.n1656 a_400_38200# 0.09fF
C4068 fc2.n1657 a_400_38200# 0.32fF
C4069 fc2.n1658 a_400_38200# 0.47fF
C4070 fc2.n1659 a_400_38200# 0.29fF
C4071 fc2.n1660 a_400_38200# 1.54fF
C4072 fc2.t205 a_400_38200# 0.02fF
C4073 fc2.n1661 a_400_38200# 0.21fF
C4074 fc2.n1662 a_400_38200# 0.80fF
C4075 fc2.n1663 a_400_38200# 0.04fF
C4076 fc2.t261 a_400_38200# 0.02fF
C4077 fc2.n1664 a_400_38200# 0.10fF
C4078 fc2.n1665 a_400_38200# 0.12fF
C4079 fc2.n1667 a_400_38200# 0.50fF
C4080 fc2.n1668 a_400_38200# 0.94fF
C4081 fc2.n1669 a_400_38200# 0.18fF
C4082 fc2.n1670 a_400_38200# 0.76fF
C4083 fc2.t179 a_400_38200# 0.02fF
C4084 fc2.n1671 a_400_38200# 0.21fF
C4085 fc2.n1672 a_400_38200# 0.31fF
C4086 fc2.n1673 a_400_38200# 0.53fF
C4087 fc2.t365 a_400_38200# 0.02fF
C4088 fc2.n1674 a_400_38200# 1.06fF
C4089 fc2.n1675 a_400_38200# 0.03fF
C4090 fc2.n1676 a_400_38200# 0.07fF
C4091 fc2.n1677 a_400_38200# 0.03fF
C4092 fc2.n1678 a_400_38200# 0.05fF
C4093 fc2.n1679 a_400_38200# 0.05fF
C4094 fc2.n1680 a_400_38200# 0.05fF
C4095 fc2.n1681 a_400_38200# 0.64fF
C4096 fc2.n1682 a_400_38200# 0.79fF
C4097 fc2.n1683 a_400_38200# 1.01fF
C4098 fc2.n1684 a_400_38200# 1.29fF
C4099 fc2.t16 a_400_38200# 7.96fF
C4100 fc2.n1685 a_400_38200# 9.42fF
C4101 fc2.n1687 a_400_38200# 0.33fF
C4102 fc2.n1688 a_400_38200# 0.20fF
C4103 fc2.n1689 a_400_38200# 3.05fF
C4104 fc2.n1690 a_400_38200# 1.86fF
C4105 fc2.n1691 a_400_38200# 0.03fF
C4106 fc2.n1692 a_400_38200# 0.07fF
C4107 fc2.n1693 a_400_38200# 0.24fF
C4108 fc2.n1694 a_400_38200# 0.58fF
C4109 fc2.n1695 a_400_38200# 0.44fF
C4110 fc2.n1696 a_400_38200# 0.72fF
C4111 fc2.n1697 a_400_38200# 0.74fF
C4112 fc2.n1698 a_400_38200# 3.62fF
C4113 fc2.n1699 a_400_38200# 0.22fF
C4114 fc2.n1700 a_400_38200# 0.01fF
C4115 fc2.t196 a_400_38200# 0.02fF
C4116 fc2.n1701 a_400_38200# 0.22fF
C4117 fc2.t161 a_400_38200# 0.02fF
C4118 fc2.n1702 a_400_38200# 0.83fF
C4119 fc2.n1703 a_400_38200# 0.62fF
C4120 fc2.n1704 a_400_38200# 1.07fF
C4121 fc2.n1705 a_400_38200# 0.25fF
C4122 fc2.n1706 a_400_38200# 0.75fF
C4123 fc2.n1707 a_400_38200# 0.18fF
C4124 fc2.n1708 a_400_38200# 0.44fF
C4125 fc2.n1709 a_400_38200# 0.79fF
C4126 fc2.t235 a_400_38200# 0.02fF
C4127 fc2.n1710 a_400_38200# 0.21fF
C4128 fc2.n1711 a_400_38200# 0.31fF
C4129 fc2.n1712 a_400_38200# 0.53fF
C4130 fc2.n1713 a_400_38200# 0.10fF
C4131 fc2.t71 a_400_38200# 0.02fF
C4132 fc2.n1714 a_400_38200# 0.12fF
C4133 fc2.n1716 a_400_38200# 0.01fF
C4134 fc2.n1717 a_400_38200# 0.03fF
C4135 fc2.n1718 a_400_38200# 0.06fF
C4136 fc2.n1719 a_400_38200# 0.24fF
C4137 fc2.n1720 a_400_38200# 0.33fF
C4138 fc2.n1721 a_400_38200# 0.13fF
C4139 fc2.n1722 a_400_38200# 0.06fF
C4140 fc2.n1723 a_400_38200# 0.11fF
C4141 fc2.n1724 a_400_38200# 0.03fF
C4142 fc2.n1725 a_400_38200# 0.07fF
C4143 fc2.n1726 a_400_38200# 0.05fF
C4144 fc2.n1727 a_400_38200# 0.09fF
C4145 fc2.n1728 a_400_38200# 0.32fF
C4146 fc2.n1729 a_400_38200# 0.47fF
C4147 fc2.n1730 a_400_38200# 0.29fF
C4148 fc2.n1731 a_400_38200# 1.60fF
C4149 fc2.t17 a_400_38200# 0.02fF
C4150 fc2.n1732 a_400_38200# 0.21fF
C4151 fc2.n1733 a_400_38200# 0.80fF
C4152 fc2.n1734 a_400_38200# 0.04fF
C4153 fc2.t101 a_400_38200# 0.02fF
C4154 fc2.n1735 a_400_38200# 0.10fF
C4155 fc2.n1736 a_400_38200# 0.12fF
C4156 fc2.n1738 a_400_38200# 0.50fF
C4157 fc2.n1739 a_400_38200# 0.94fF
C4158 fc2.n1740 a_400_38200# 0.18fF
C4159 fc2.n1741 a_400_38200# 0.76fF
C4160 fc2.t51 a_400_38200# 0.02fF
C4161 fc2.n1742 a_400_38200# 0.21fF
C4162 fc2.n1743 a_400_38200# 0.31fF
C4163 fc2.n1744 a_400_38200# 0.53fF
C4164 fc2.n1745 a_400_38200# 0.10fF
C4165 fc2.t256 a_400_38200# 0.02fF
C4166 fc2.n1746 a_400_38200# 0.12fF
C4167 fc2.n1748 a_400_38200# 0.76fF
C4168 fc2.n1749 a_400_38200# 0.44fF
C4169 fc2.n1750 a_400_38200# 1.07fF
C4170 fc2.n1751 a_400_38200# 0.18fF
C4171 fc2.n1752 a_400_38200# 3.23fF
C4172 fc2.t211 a_400_38200# 0.02fF
C4173 fc2.n1753 a_400_38200# 0.21fF
C4174 fc2.n1754 a_400_38200# 0.80fF
C4175 fc2.n1755 a_400_38200# 0.04fF
C4176 fc2.t285 a_400_38200# 0.02fF
C4177 fc2.n1756 a_400_38200# 0.10fF
C4178 fc2.n1757 a_400_38200# 0.12fF
C4179 fc2.n1759 a_400_38200# 7.70fF
C4180 fc2.n1760 a_400_38200# 2.48fF
C4181 fc2.t185 a_400_38200# 0.02fF
C4182 fc2.n1761 a_400_38200# 0.21fF
C4183 fc2.n1762 a_400_38200# 0.31fF
C4184 fc2.n1763 a_400_38200# 0.53fF
C4185 fc2.n1764 a_400_38200# 0.10fF
C4186 fc2.t389 a_400_38200# 0.02fF
C4187 fc2.n1765 a_400_38200# 0.12fF
C4188 fc2.n1767 a_400_38200# 0.03fF
C4189 fc2.n1768 a_400_38200# 0.01fF
C4190 fc2.n1769 a_400_38200# 0.06fF
C4191 fc2.n1770 a_400_38200# 0.24fF
C4192 fc2.n1771 a_400_38200# 0.33fF
C4193 fc2.n1772 a_400_38200# 0.13fF
C4194 fc2.n1773 a_400_38200# 0.06fF
C4195 fc2.n1774 a_400_38200# 0.11fF
C4196 fc2.n1775 a_400_38200# 0.06fF
C4197 fc2.n1776 a_400_38200# 0.05fF
C4198 fc2.n1777 a_400_38200# 0.10fF
C4199 fc2.n1778 a_400_38200# 0.08fF
C4200 fc2.n1779 a_400_38200# 0.32fF
C4201 fc2.n1780 a_400_38200# 0.47fF
C4202 fc2.n1781 a_400_38200# 0.29fF
C4203 fc2.n1782 a_400_38200# 3.45fF
C4204 fc2.t13 a_400_38200# 0.02fF
C4205 fc2.n1783 a_400_38200# 0.10fF
C4206 fc2.n1784 a_400_38200# 0.12fF
C4207 fc2.t350 a_400_38200# 0.02fF
C4208 fc2.n1786 a_400_38200# 0.21fF
C4209 fc2.n1787 a_400_38200# 0.80fF
C4210 fc2.n1788 a_400_38200# 0.04fF
C4211 fc2.n1789 a_400_38200# 1.04fF
C4212 fc2.n1790 a_400_38200# 0.12fF
C4213 fc2.n1791 a_400_38200# 0.10fF
C4214 fc2.t147 a_400_38200# 0.02fF
C4215 fc2.n1792 a_400_38200# 0.12fF
C4216 fc2.t296 a_400_38200# 0.02fF
C4217 fc2.n1794 a_400_38200# 0.21fF
C4218 fc2.n1795 a_400_38200# 0.31fF
C4219 fc2.n1796 a_400_38200# 0.53fF
C4220 fc2.n1797 a_400_38200# 0.76fF
C4221 fc2.n1798 a_400_38200# 0.50fF
C4222 fc2.n1799 a_400_38200# 1.21fF
C4223 fc2.n1800 a_400_38200# 0.18fF
C4224 fc2.n1801 a_400_38200# 3.32fF
C4225 fc2.t160 a_400_38200# 0.02fF
C4226 fc2.n1802 a_400_38200# 0.10fF
C4227 fc2.n1803 a_400_38200# 0.12fF
C4228 fc2.t89 a_400_38200# 0.02fF
C4229 fc2.n1805 a_400_38200# 0.21fF
C4230 fc2.n1806 a_400_38200# 0.80fF
C4231 fc2.n1807 a_400_38200# 0.04fF
C4232 fc2.t12 a_400_38200# 17.22fF
C4233 fc2.t342 a_400_38200# 0.02fF
C4234 fc2.n1808 a_400_38200# 0.21fF
C4235 fc2.n1809 a_400_38200# 0.80fF
C4236 fc2.n1810 a_400_38200# 0.04fF
C4237 fc2.t33 a_400_38200# 0.02fF
C4238 fc2.n1811 a_400_38200# 0.10fF
C4239 fc2.n1812 a_400_38200# 0.12fF
C4240 fc2.n1814 a_400_38200# 0.10fF
C4241 fc2.t382 a_400_38200# 0.02fF
C4242 fc2.n1815 a_400_38200# 0.12fF
C4243 fc2.n1817 a_400_38200# 0.01fF
C4244 fc2.n1818 a_400_38200# 0.03fF
C4245 fc2.n1819 a_400_38200# 0.06fF
C4246 fc2.n1820 a_400_38200# 0.24fF
C4247 fc2.n1821 a_400_38200# 0.33fF
C4248 fc2.n1822 a_400_38200# 0.13fF
C4249 fc2.n1823 a_400_38200# 0.06fF
C4250 fc2.n1824 a_400_38200# 0.11fF
C4251 fc2.n1825 a_400_38200# 0.03fF
C4252 fc2.n1826 a_400_38200# 0.07fF
C4253 fc2.n1827 a_400_38200# 0.05fF
C4254 fc2.n1828 a_400_38200# 0.09fF
C4255 fc2.n1829 a_400_38200# 0.32fF
C4256 fc2.n1830 a_400_38200# 0.47fF
C4257 fc2.n1831 a_400_38200# 0.29fF
C4258 fc2.n1832 a_400_38200# 3.31fF
C4259 fc2.n1833 a_400_38200# 1.75fF
C4260 fc2.n1834 a_400_38200# 0.05fF
C4261 fc2.n1835 a_400_38200# 0.07fF
C4262 fc2.n1836 a_400_38200# 1.01fF
C4263 fc2.n1837 a_400_38200# 0.12fF
C4264 fc2.n1838 a_400_38200# 0.05fF
C4265 fc2.n1839 a_400_38200# 0.17fF
C4266 fc2.n1840 a_400_38200# 0.06fF
C4267 fc2.n1841 a_400_38200# 0.03fF
C4268 fc2.n1842 a_400_38200# 0.10fF
C4269 fc2.n1843 a_400_38200# 0.17fF
C4270 fc2.n1844 a_400_38200# 0.69fF
C4271 fc2.t201 a_400_38200# 0.02fF
C4272 fc2.n1845 a_400_38200# 0.21fF
C4273 fc2.n1846 a_400_38200# 0.31fF
C4274 fc2.n1847 a_400_38200# 0.53fF
C4275 fc2.n1848 a_400_38200# 0.10fF
C4276 fc2.t29 a_400_38200# 0.02fF
C4277 fc2.n1849 a_400_38200# 0.12fF
C4278 fc2.n1851 a_400_38200# 0.01fF
C4279 fc2.n1852 a_400_38200# 0.03fF
C4280 fc2.n1853 a_400_38200# 0.06fF
C4281 fc2.n1854 a_400_38200# 0.24fF
C4282 fc2.n1855 a_400_38200# 0.05fF
C4283 fc2.n1856 a_400_38200# 0.03fF
C4284 fc2.n1857 a_400_38200# 0.33fF
C4285 fc2.n1858 a_400_38200# 0.13fF
C4286 fc2.n1859 a_400_38200# 0.06fF
C4287 fc2.n1860 a_400_38200# 0.11fF
C4288 fc2.n1861 a_400_38200# 0.03fF
C4289 fc2.n1862 a_400_38200# 0.07fF
C4290 fc2.n1863 a_400_38200# 0.03fF
C4291 fc2.n1864 a_400_38200# 0.05fF
C4292 fc2.n1865 a_400_38200# 0.05fF
C4293 fc2.n1866 a_400_38200# 0.09fF
C4294 fc2.n1867 a_400_38200# 0.32fF
C4295 fc2.n1868 a_400_38200# 0.47fF
C4296 fc2.n1869 a_400_38200# 0.29fF
C4297 fc2.n1870 a_400_38200# 1.53fF
C4298 fc2.t81 a_400_38200# 0.02fF
C4299 fc2.n1871 a_400_38200# 0.21fF
C4300 fc2.n1872 a_400_38200# 0.80fF
C4301 fc2.n1873 a_400_38200# 0.04fF
C4302 fc2.t136 a_400_38200# 0.02fF
C4303 fc2.n1874 a_400_38200# 0.10fF
C4304 fc2.n1875 a_400_38200# 0.12fF
C4305 fc2.n1877 a_400_38200# 1.81fF
C4306 fc2.n1878 a_400_38200# 0.05fF
C4307 fc2.n1879 a_400_38200# 0.07fF
C4308 fc2.n1880 a_400_38200# 1.00fF
C4309 fc2.n1881 a_400_38200# 0.12fF
C4310 fc2.n1882 a_400_38200# 0.05fF
C4311 fc2.n1883 a_400_38200# 0.17fF
C4312 fc2.n1884 a_400_38200# 0.06fF
C4313 fc2.n1885 a_400_38200# 0.03fF
C4314 fc2.n1886 a_400_38200# 0.10fF
C4315 fc2.n1887 a_400_38200# 0.17fF
C4316 fc2.n1888 a_400_38200# 0.69fF
C4317 fc2.t78 a_400_38200# 0.02fF
C4318 fc2.n1889 a_400_38200# 0.21fF
C4319 fc2.n1890 a_400_38200# 0.31fF
C4320 fc2.n1891 a_400_38200# 0.53fF
C4321 fc2.n1892 a_400_38200# 0.10fF
C4322 fc2.t279 a_400_38200# 0.02fF
C4323 fc2.n1893 a_400_38200# 0.12fF
C4324 fc2.n1895 a_400_38200# 0.76fF
C4325 fc2.n1896 a_400_38200# 0.44fF
C4326 fc2.n1897 a_400_38200# 1.07fF
C4327 fc2.n1898 a_400_38200# 0.18fF
C4328 fc2.n1899 a_400_38200# 1.51fF
C4329 fc2.t324 a_400_38200# 0.02fF
C4330 fc2.n1900 a_400_38200# 0.21fF
C4331 fc2.n1901 a_400_38200# 0.80fF
C4332 fc2.n1902 a_400_38200# 0.04fF
C4333 fc2.t379 a_400_38200# 0.02fF
C4334 fc2.n1903 a_400_38200# 0.10fF
C4335 fc2.n1904 a_400_38200# 0.12fF
C4336 fc2.n1906 a_400_38200# 7.70fF
C4337 fc2.n1907 a_400_38200# 0.04fF
C4338 fc2.n1908 a_400_38200# 0.05fF
C4339 fc2.n1909 a_400_38200# 0.05fF
C4340 fc2.n1910 a_400_38200# 0.03fF
C4341 fc2.n1911 a_400_38200# 1.03fF
C4342 fc2.n1912 a_400_38200# 0.21fF
C4343 fc2.n1913 a_400_38200# 0.10fF
C4344 fc2.n1914 a_400_38200# 0.64fF
C4345 fc2.t387 a_400_38200# 0.02fF
C4346 fc2.n1915 a_400_38200# 0.21fF
C4347 fc2.n1916 a_400_38200# 0.31fF
C4348 fc2.n1917 a_400_38200# 0.53fF
C4349 fc2.n1918 a_400_38200# 0.10fF
C4350 fc2.t216 a_400_38200# 0.02fF
C4351 fc2.n1919 a_400_38200# 0.12fF
C4352 fc2.n1921 a_400_38200# 0.01fF
C4353 fc2.n1922 a_400_38200# 0.03fF
C4354 fc2.n1923 a_400_38200# 0.06fF
C4355 fc2.n1924 a_400_38200# 0.24fF
C4356 fc2.n1925 a_400_38200# 0.32fF
C4357 fc2.n1926 a_400_38200# 0.13fF
C4358 fc2.n1927 a_400_38200# 0.06fF
C4359 fc2.n1928 a_400_38200# 0.11fF
C4360 fc2.n1929 a_400_38200# 0.03fF
C4361 fc2.n1930 a_400_38200# 0.07fF
C4362 fc2.n1931 a_400_38200# 0.03fF
C4363 fc2.n1932 a_400_38200# 0.05fF
C4364 fc2.n1933 a_400_38200# 0.05fF
C4365 fc2.n1934 a_400_38200# 0.09fF
C4366 fc2.n1935 a_400_38200# 0.32fF
C4367 fc2.n1936 a_400_38200# 0.47fF
C4368 fc2.n1937 a_400_38200# 0.29fF
C4369 fc2.n1938 a_400_38200# 3.03fF
C4370 fc2.t319 a_400_38200# 0.02fF
C4371 fc2.n1939 a_400_38200# 0.10fF
C4372 fc2.n1940 a_400_38200# 0.12fF
C4373 fc2.t264 a_400_38200# 0.02fF
C4374 fc2.n1942 a_400_38200# 0.21fF
C4375 fc2.n1943 a_400_38200# 0.80fF
C4376 fc2.n1944 a_400_38200# 0.04fF
C4377 fc2.n1945 a_400_38200# 0.52fF
C4378 fc2.n1946 a_400_38200# 0.46fF
C4379 fc2.n1947 a_400_38200# 0.76fF
C4380 fc2.n1948 a_400_38200# 0.46fF
C4381 fc2.n1949 a_400_38200# 1.04fF
C4382 fc2.n1950 a_400_38200# 0.12fF
C4383 fc2.n1951 a_400_38200# 0.10fF
C4384 fc2.t151 a_400_38200# 0.02fF
C4385 fc2.n1952 a_400_38200# 0.12fF
C4386 fc2.t317 a_400_38200# 0.02fF
C4387 fc2.n1954 a_400_38200# 0.21fF
C4388 fc2.n1955 a_400_38200# 0.31fF
C4389 fc2.n1956 a_400_38200# 0.53fF
C4390 fc2.n1957 a_400_38200# 0.02fF
C4391 fc2.n1958 a_400_38200# 0.08fF
C4392 fc2.n1959 a_400_38200# 0.12fF
C4393 fc2.n1960 a_400_38200# 0.04fF
C4394 fc2.n1961 a_400_38200# 0.03fF
C4395 fc2.n1962 a_400_38200# 0.03fF
C4396 fc2.n1963 a_400_38200# 0.13fF
C4397 fc2.n1964 a_400_38200# 0.60fF
C4398 fc2.n1965 a_400_38200# 1.35fF
C4399 fc2.n1966 a_400_38200# 3.31fF
C4400 fc2.t266 a_400_38200# 0.02fF
C4401 fc2.n1967 a_400_38200# 0.10fF
C4402 fc2.n1968 a_400_38200# 0.12fF
C4403 fc2.t194 a_400_38200# 0.02fF
C4404 fc2.n1970 a_400_38200# 0.21fF
C4405 fc2.n1971 a_400_38200# 0.80fF
C4406 fc2.n1972 a_400_38200# 0.04fF
C4407 fc2.t28 a_400_38200# 16.88fF
C4408 fc2.t68 a_400_38200# 0.02fF
C4409 fc2.n1973 a_400_38200# 1.04fF
C4410 fc2.n1974 a_400_38200# 0.04fF
C4411 fc2.t142 a_400_38200# 0.02fF
C4412 fc2.n1975 a_400_38200# 0.01fF
C4413 fc2.n1976 a_400_38200# 0.22fF
C4414 fc2.n1978 a_400_38200# 0.04fF
C4415 fc2.n1979 a_400_38200# 0.18fF
C4416 fc2.n1980 a_400_38200# 0.11fF
C4417 fc2.n1981 a_400_38200# 0.10fF
C4418 fc2.n1982 a_400_38200# 0.82fF
C4419 fc2.n1983 a_400_38200# 0.05fF
C4420 fc2.n1984 a_400_38200# 0.16fF
C4421 fc2.n1985 a_400_38200# 0.08fF
C4422 fc2.n1986 a_400_38200# 1.57fF
C4423 fc2.n1987 a_400_38200# 1.85fF
C4424 fc2.n1988 a_400_38200# 2.13fF
C4425 fc2.t268 a_400_38200# 0.02fF
C4426 fc2.n1989 a_400_38200# 0.21fF
C4427 fc2.n1990 a_400_38200# 0.31fF
C4428 fc2.n1991 a_400_38200# 0.53fF
C4429 fc2.t79 a_400_38200# 0.02fF
C4430 fc2.n1992 a_400_38200# 1.06fF
C4431 fc2.n1993 a_400_38200# 0.03fF
C4432 fc2.n1994 a_400_38200# 0.07fF
C4433 fc2.n1995 a_400_38200# 0.05fF
C4434 fc2.n1996 a_400_38200# 0.05fF
C4435 fc2.n1997 a_400_38200# 0.64fF
C4436 fc2.n1998 a_400_38200# 0.79fF
C4437 fc2.n1999 a_400_38200# 1.01fF
C4438 fc2.n2000 a_400_38200# 1.29fF
C4439 fc2.t34 a_400_38200# 7.96fF
C4440 fc2.n2001 a_400_38200# 9.42fF
C4441 fc2.n2003 a_400_38200# 0.33fF
C4442 fc2.n2004 a_400_38200# 0.20fF
C4443 fc2.n2005 a_400_38200# 3.05fF
C4444 fc2.n2006 a_400_38200# 1.86fF
C4445 fc2.n2007 a_400_38200# 0.03fF
C4446 fc2.n2008 a_400_38200# 0.07fF
C4447 fc2.n2009 a_400_38200# 0.24fF
C4448 fc2.n2010 a_400_38200# 0.58fF
C4449 fc2.n2011 a_400_38200# 0.44fF
C4450 fc2.n2012 a_400_38200# 0.72fF
C4451 fc2.n2013 a_400_38200# 0.74fF
C4452 fc2.n2014 a_400_38200# 3.62fF
C4453 fc2.n2015 a_400_38200# 0.22fF
C4454 fc2.n2016 a_400_38200# 0.01fF
C4455 fc2.t281 a_400_38200# 0.02fF
C4456 fc2.n2017 a_400_38200# 0.22fF
C4457 fc2.t169 a_400_38200# 0.02fF
C4458 fc2.n2018 a_400_38200# 0.83fF
C4459 fc2.n2019 a_400_38200# 0.62fF
C4460 fc2.n2020 a_400_38200# 1.07fF
C4461 fc2.n2021 a_400_38200# 0.52fF
C4462 fc2.n2022 a_400_38200# 0.94fF
C4463 fc2.n2023 a_400_38200# 0.18fF
C4464 fc2.n2024 a_400_38200# 0.76fF
C4465 fc2.t320 a_400_38200# 0.02fF
C4466 fc2.n2025 a_400_38200# 0.21fF
C4467 fc2.n2026 a_400_38200# 0.31fF
C4468 fc2.n2027 a_400_38200# 0.53fF
C4469 fc2.n2028 a_400_38200# 0.10fF
C4470 fc2.t154 a_400_38200# 0.02fF
C4471 fc2.n2029 a_400_38200# 0.12fF
C4472 fc2.n2031 a_400_38200# 0.01fF
C4473 fc2.n2032 a_400_38200# 0.03fF
C4474 fc2.n2033 a_400_38200# 0.06fF
C4475 fc2.n2034 a_400_38200# 0.24fF
C4476 fc2.n2035 a_400_38200# 0.33fF
C4477 fc2.n2036 a_400_38200# 0.13fF
C4478 fc2.n2037 a_400_38200# 0.06fF
C4479 fc2.n2038 a_400_38200# 0.11fF
C4480 fc2.n2039 a_400_38200# 0.03fF
C4481 fc2.n2040 a_400_38200# 0.07fF
C4482 fc2.n2041 a_400_38200# 0.05fF
C4483 fc2.n2042 a_400_38200# 0.09fF
C4484 fc2.n2043 a_400_38200# 0.32fF
C4485 fc2.n2044 a_400_38200# 0.47fF
C4486 fc2.n2045 a_400_38200# 0.29fF
C4487 fc2.n2046 a_400_38200# 1.59fF
C4488 fc2.t35 a_400_38200# 0.02fF
C4489 fc2.n2047 a_400_38200# 0.21fF
C4490 fc2.n2048 a_400_38200# 0.80fF
C4491 fc2.n2049 a_400_38200# 0.04fF
C4492 fc2.t181 a_400_38200# 0.02fF
C4493 fc2.n2050 a_400_38200# 0.10fF
C4494 fc2.n2051 a_400_38200# 0.12fF
C4495 fc2.n2053 a_400_38200# 0.50fF
C4496 fc2.n2054 a_400_38200# 0.94fF
C4497 fc2.n2055 a_400_38200# 0.18fF
C4498 fc2.n2056 a_400_38200# 0.76fF
C4499 fc2.t1 a_400_38200# 0.02fF
C4500 fc2.n2057 a_400_38200# 0.21fF
C4501 fc2.n2058 a_400_38200# 0.31fF
C4502 fc2.n2059 a_400_38200# 0.53fF
C4503 fc2.n2060 a_400_38200# 0.10fF
C4504 fc2.t220 a_400_38200# 0.02fF
C4505 fc2.n2061 a_400_38200# 0.12fF
C4506 fc2.n2063 a_400_38200# 0.76fF
C4507 fc2.n2064 a_400_38200# 0.44fF
C4508 fc2.n2065 a_400_38200# 1.07fF
C4509 fc2.n2066 a_400_38200# 0.18fF
C4510 fc2.n2067 a_400_38200# 3.23fF
C4511 fc2.t116 a_400_38200# 0.02fF
C4512 fc2.n2068 a_400_38200# 0.21fF
C4513 fc2.n2069 a_400_38200# 0.80fF
C4514 fc2.n2070 a_400_38200# 0.04fF
C4515 fc2.t253 a_400_38200# 0.02fF
C4516 fc2.n2071 a_400_38200# 0.10fF
C4517 fc2.n2072 a_400_38200# 0.12fF
C4518 fc2.n2074 a_400_38200# 7.70fF
C4519 fc2.n2075 a_400_38200# 0.44fF
C4520 fc2.n2076 a_400_38200# 0.25fF
C4521 fc2.n2077 a_400_38200# 0.75fF
C4522 fc2.n2078 a_400_38200# 0.18fF
C4523 fc2.n2079 a_400_38200# 0.76fF
C4524 fc2.t137 a_400_38200# 0.02fF
C4525 fc2.n2080 a_400_38200# 0.21fF
C4526 fc2.n2081 a_400_38200# 0.31fF
C4527 fc2.n2082 a_400_38200# 0.53fF
C4528 fc2.n2083 a_400_38200# 0.10fF
C4529 fc2.t339 a_400_38200# 0.02fF
C4530 fc2.n2084 a_400_38200# 0.12fF
C4531 fc2.n2086 a_400_38200# 0.03fF
C4532 fc2.n2087 a_400_38200# 0.01fF
C4533 fc2.n2088 a_400_38200# 0.06fF
C4534 fc2.n2089 a_400_38200# 0.24fF
C4535 fc2.n2090 a_400_38200# 0.33fF
C4536 fc2.n2091 a_400_38200# 0.13fF
C4537 fc2.n2092 a_400_38200# 0.06fF
C4538 fc2.n2093 a_400_38200# 0.11fF
C4539 fc2.n2094 a_400_38200# 0.05fF
C4540 fc2.n2095 a_400_38200# 0.09fF
C4541 fc2.n2096 a_400_38200# 0.03fF
C4542 fc2.n2097 a_400_38200# 0.07fF
C4543 fc2.n2098 a_400_38200# 0.32fF
C4544 fc2.n2099 a_400_38200# 0.47fF
C4545 fc2.n2100 a_400_38200# 0.29fF
C4546 fc2.n2101 a_400_38200# 3.32fF
C4547 fc2.t369 a_400_38200# 0.02fF
C4548 fc2.n2102 a_400_38200# 0.10fF
C4549 fc2.n2103 a_400_38200# 0.12fF
C4550 fc2.t225 a_400_38200# 0.02fF
C4551 fc2.n2105 a_400_38200# 0.21fF
C4552 fc2.n2106 a_400_38200# 0.80fF
C4553 fc2.n2107 a_400_38200# 0.04fF
C4554 fc2.n2108 a_400_38200# 1.79fF
C4555 fc2.n2109 a_400_38200# 0.58fF
C4556 fc2.n2110 a_400_38200# 0.94fF
C4557 fc2.n2111 a_400_38200# 0.18fF
C4558 fc2.n2112 a_400_38200# 0.76fF
C4559 fc2.t380 a_400_38200# 0.02fF
C4560 fc2.n2113 a_400_38200# 0.21fF
C4561 fc2.n2114 a_400_38200# 0.31fF
C4562 fc2.n2115 a_400_38200# 0.53fF
C4563 fc2.n2116 a_400_38200# 0.10fF
C4564 fc2.t228 a_400_38200# 0.02fF
C4565 fc2.n2117 a_400_38200# 0.12fF
C4566 fc2.n2119 a_400_38200# 0.01fF
C4567 fc2.n2120 a_400_38200# 0.03fF
C4568 fc2.n2121 a_400_38200# 0.06fF
C4569 fc2.n2122 a_400_38200# 0.24fF
C4570 fc2.n2123 a_400_38200# 0.33fF
C4571 fc2.n2124 a_400_38200# 0.13fF
C4572 fc2.n2125 a_400_38200# 0.06fF
C4573 fc2.n2126 a_400_38200# 0.11fF
C4574 fc2.n2127 a_400_38200# 0.03fF
C4575 fc2.n2128 a_400_38200# 0.07fF
C4576 fc2.n2129 a_400_38200# 0.05fF
C4577 fc2.n2130 a_400_38200# 0.09fF
C4578 fc2.n2131 a_400_38200# 0.32fF
C4579 fc2.n2132 a_400_38200# 0.47fF
C4580 fc2.n2133 a_400_38200# 0.29fF
C4581 fc2.n2134 a_400_38200# 1.64fF
C4582 fc2.t241 a_400_38200# 0.02fF
C4583 fc2.n2135 a_400_38200# 0.10fF
C4584 fc2.n2136 a_400_38200# 0.12fF
C4585 fc2.t104 a_400_38200# 0.02fF
C4586 fc2.n2138 a_400_38200# 0.21fF
C4587 fc2.n2139 a_400_38200# 0.80fF
C4588 fc2.n2140 a_400_38200# 0.04fF
C4589 fc2.n2141 a_400_38200# 1.04fF
C4590 fc2.n2142 a_400_38200# 0.12fF
C4591 fc2.n2143 a_400_38200# 0.10fF
C4592 fc2.t99 a_400_38200# 0.02fF
C4593 fc2.n2144 a_400_38200# 0.12fF
C4594 fc2.t263 a_400_38200# 0.02fF
C4595 fc2.n2146 a_400_38200# 0.21fF
C4596 fc2.n2147 a_400_38200# 0.31fF
C4597 fc2.n2148 a_400_38200# 0.53fF
C4598 fc2.n2149 a_400_38200# 0.94fF
C4599 fc2.n2150 a_400_38200# 0.18fF
C4600 fc2.n2151 a_400_38200# 3.32fF
C4601 fc2.t128 a_400_38200# 0.02fF
C4602 fc2.n2152 a_400_38200# 0.10fF
C4603 fc2.n2153 a_400_38200# 0.12fF
C4604 fc2.t352 a_400_38200# 0.02fF
C4605 fc2.n2155 a_400_38200# 0.21fF
C4606 fc2.n2156 a_400_38200# 0.80fF
C4607 fc2.n2157 a_400_38200# 0.04fF
C4608 fc2.t98 a_400_38200# 17.22fF
C4609 fc2.t362 a_400_38200# 0.02fF
C4610 fc2.n2158 a_400_38200# 0.21fF
C4611 fc2.n2159 a_400_38200# 0.80fF
C4612 fc2.n2160 a_400_38200# 0.04fF
C4613 fc2.t118 a_400_38200# 0.02fF
C4614 fc2.n2161 a_400_38200# 0.10fF
C4615 fc2.n2162 a_400_38200# 0.12fF
C4616 fc2.n2164 a_400_38200# 0.10fF
C4617 fc2.t108 a_400_38200# 0.02fF
C4618 fc2.n2165 a_400_38200# 0.12fF
C4619 fc2.n2167 a_400_38200# 0.01fF
C4620 fc2.n2168 a_400_38200# 0.03fF
C4621 fc2.n2169 a_400_38200# 0.06fF
C4622 fc2.n2170 a_400_38200# 0.24fF
C4623 fc2.n2171 a_400_38200# 0.33fF
C4624 fc2.n2172 a_400_38200# 0.13fF
C4625 fc2.n2173 a_400_38200# 0.06fF
C4626 fc2.n2174 a_400_38200# 0.11fF
C4627 fc2.n2175 a_400_38200# 0.04fF
C4628 fc2.n2176 a_400_38200# 0.08fF
C4629 fc2.n2177 a_400_38200# 0.05fF
C4630 fc2.n2178 a_400_38200# 0.09fF
C4631 fc2.n2179 a_400_38200# 0.32fF
C4632 fc2.n2180 a_400_38200# 0.47fF
C4633 fc2.n2181 a_400_38200# 0.29fF
C4634 fc2.n2182 a_400_38200# 1.65fF
C4635 fc2.n2183 a_400_38200# 1.71fF
C4636 fc2.n2184 a_400_38200# 0.28fF
C4637 fc2.n2185 a_400_38200# 0.12fF
C4638 fc2.n2186 a_400_38200# 0.18fF
C4639 fc2.n2187 a_400_38200# 0.05fF
C4640 fc2.n2188 a_400_38200# 0.04fF
C4641 fc2.n2189 a_400_38200# 0.20fF
C4642 fc2.n2190 a_400_38200# 1.01fF
C4643 fc2.n2191 a_400_38200# 0.02fF
C4644 fc2.n2192 a_400_38200# 1.68fF
C4645 fc2.n2193 a_400_38200# 0.05fF
C4646 fc2.n2194 a_400_38200# 0.07fF
C4647 fc2.n2195 a_400_38200# 1.00fF
C4648 fc2.n2196 a_400_38200# 0.12fF
C4649 fc2.n2197 a_400_38200# 0.05fF
C4650 fc2.n2198 a_400_38200# 0.17fF
C4651 fc2.n2199 a_400_38200# 0.06fF
C4652 fc2.n2200 a_400_38200# 0.03fF
C4653 fc2.n2201 a_400_38200# 0.10fF
C4654 fc2.n2202 a_400_38200# 0.17fF
C4655 fc2.n2203 a_400_38200# 0.69fF
C4656 fc2.t171 a_400_38200# 0.02fF
C4657 fc2.n2204 a_400_38200# 0.21fF
C4658 fc2.n2205 a_400_38200# 0.31fF
C4659 fc2.n2206 a_400_38200# 0.53fF
C4660 fc2.n2207 a_400_38200# 0.10fF
C4661 fc2.t376 a_400_38200# 0.02fF
C4662 fc2.n2208 a_400_38200# 0.12fF
C4663 fc2.n2210 a_400_38200# 0.01fF
C4664 fc2.n2211 a_400_38200# 0.03fF
C4665 fc2.n2212 a_400_38200# 0.06fF
C4666 fc2.n2213 a_400_38200# 0.24fF
C4667 fc2.n2214 a_400_38200# 0.05fF
C4668 fc2.n2215 a_400_38200# 0.03fF
C4669 fc2.n2216 a_400_38200# 0.33fF
C4670 fc2.n2217 a_400_38200# 0.13fF
C4671 fc2.n2218 a_400_38200# 0.06fF
C4672 fc2.n2219 a_400_38200# 0.11fF
C4673 fc2.n2220 a_400_38200# 0.03fF
C4674 fc2.n2221 a_400_38200# 0.07fF
C4675 fc2.n2222 a_400_38200# 0.03fF
C4676 fc2.n2223 a_400_38200# 0.05fF
C4677 fc2.n2224 a_400_38200# 0.05fF
C4678 fc2.n2225 a_400_38200# 0.09fF
C4679 fc2.n2226 a_400_38200# 0.32fF
C4680 fc2.n2227 a_400_38200# 0.47fF
C4681 fc2.n2228 a_400_38200# 0.29fF
C4682 fc2.n2229 a_400_38200# 1.87fF
C4683 fc2.t46 a_400_38200# 0.02fF
C4684 fc2.n2230 a_400_38200# 0.21fF
C4685 fc2.n2231 a_400_38200# 0.80fF
C4686 fc2.n2232 a_400_38200# 0.04fF
C4687 fc2.t274 a_400_38200# 0.02fF
C4688 fc2.n2233 a_400_38200# 0.10fF
C4689 fc2.n2234 a_400_38200# 0.12fF
C4690 fc2.t293 a_400_38200# 0.02fF
C4691 fc2.n2236 a_400_38200# 0.21fF
C4692 fc2.n2237 a_400_38200# 0.80fF
C4693 fc2.n2238 a_400_38200# 0.04fF
C4694 fc2.n2239 a_400_38200# 1.81fF
C4695 fc2.n2240 a_400_38200# 0.05fF
C4696 fc2.n2241 a_400_38200# 0.07fF
C4697 fc2.n2242 a_400_38200# 1.00fF
C4698 fc2.n2243 a_400_38200# 0.12fF
C4699 fc2.n2244 a_400_38200# 0.05fF
C4700 fc2.n2245 a_400_38200# 0.17fF
C4701 fc2.n2246 a_400_38200# 0.06fF
C4702 fc2.n2247 a_400_38200# 0.03fF
C4703 fc2.n2248 a_400_38200# 0.10fF
C4704 fc2.n2249 a_400_38200# 0.17fF
C4705 fc2.n2250 a_400_38200# 0.69fF
C4706 fc2.t37 a_400_38200# 0.02fF
C4707 fc2.n2251 a_400_38200# 0.21fF
C4708 fc2.n2252 a_400_38200# 0.31fF
C4709 fc2.n2253 a_400_38200# 0.53fF
C4710 fc2.n2254 a_400_38200# 0.10fF
C4711 fc2.t248 a_400_38200# 0.02fF
C4712 fc2.n2255 a_400_38200# 0.12fF
C4713 fc2.n2257 a_400_38200# 0.76fF
C4714 fc2.n2258 a_400_38200# 0.44fF
C4715 fc2.n2259 a_400_38200# 1.07fF
C4716 fc2.n2260 a_400_38200# 0.18fF
C4717 fc2.n2261 a_400_38200# 1.51fF
C4718 fc2.t345 a_400_38200# 0.02fF
C4719 fc2.n2262 a_400_38200# 0.10fF
C4720 fc2.n2263 a_400_38200# 0.12fF
C4721 fc2.n2265 a_400_38200# 7.70fF
C4722 fc2.n2266 a_400_38200# 0.04fF
C4723 fc2.n2267 a_400_38200# 0.05fF
C4724 fc2.n2268 a_400_38200# 0.05fF
C4725 fc2.n2269 a_400_38200# 0.03fF
C4726 fc2.n2270 a_400_38200# 1.06fF
C4727 fc2.n2271 a_400_38200# 0.21fF
C4728 fc2.n2272 a_400_38200# 0.10fF
C4729 fc2.n2273 a_400_38200# 0.64fF
C4730 fc2.t105 a_400_38200# 0.02fF
C4731 fc2.n2274 a_400_38200# 0.21fF
C4732 fc2.n2275 a_400_38200# 0.31fF
C4733 fc2.n2276 a_400_38200# 0.53fF
C4734 fc2.t349 a_400_38200# 0.02fF
C4735 fc2.n2277 a_400_38200# 0.21fF
C4736 fc2.n2278 a_400_38200# 0.80fF
C4737 fc2.n2279 a_400_38200# 0.04fF
C4738 fc2.n2280 a_400_38200# 0.10fF
C4739 fc2.t304 a_400_38200# 0.02fF
C4740 fc2.n2281 a_400_38200# 0.12fF
C4741 fc2.n2283 a_400_38200# 0.01fF
C4742 fc2.n2284 a_400_38200# 0.03fF
C4743 fc2.n2285 a_400_38200# 0.06fF
C4744 fc2.n2286 a_400_38200# 0.24fF
C4745 fc2.n2287 a_400_38200# 0.05fF
C4746 fc2.n2288 a_400_38200# 0.03fF
C4747 fc2.n2289 a_400_38200# 0.32fF
C4748 fc2.n2290 a_400_38200# 0.13fF
C4749 fc2.n2291 a_400_38200# 0.06fF
C4750 fc2.n2292 a_400_38200# 0.11fF
C4751 fc2.n2293 a_400_38200# 0.03fF
C4752 fc2.n2294 a_400_38200# 0.07fF
C4753 fc2.n2295 a_400_38200# 0.03fF
C4754 fc2.n2296 a_400_38200# 0.05fF
C4755 fc2.n2297 a_400_38200# 0.05fF
C4756 fc2.n2298 a_400_38200# 0.09fF
C4757 fc2.n2299 a_400_38200# 0.32fF
C4758 fc2.n2300 a_400_38200# 0.47fF
C4759 fc2.n2301 a_400_38200# 0.29fF
C4760 fc2.n2302 a_400_38200# 3.03fF
C4761 fc2.t24 a_400_38200# 0.02fF
C4762 fc2.n2303 a_400_38200# 0.10fF
C4763 fc2.n2304 a_400_38200# 0.12fF
C4764 fc2.n2306 a_400_38200# 0.05fF
C4765 fc2.n2307 a_400_38200# 0.07fF
C4766 fc2.n2308 a_400_38200# 1.07fF
C4767 fc2.n2309 a_400_38200# 0.12fF
C4768 fc2.n2310 a_400_38200# 0.16fF
C4769 fc2.n2311 a_400_38200# 0.05fF
C4770 fc2.n2312 a_400_38200# 0.03fF
C4771 fc2.n2313 a_400_38200# 0.10fF
C4772 fc2.n2314 a_400_38200# 0.17fF
C4773 fc2.n2315 a_400_38200# 0.69fF
C4774 fc2.t162 a_400_38200# 0.02fF
C4775 fc2.n2316 a_400_38200# 0.21fF
C4776 fc2.n2317 a_400_38200# 0.31fF
C4777 fc2.n2318 a_400_38200# 0.53fF
C4778 fc2.n2319 a_400_38200# 0.10fF
C4779 fc2.t364 a_400_38200# 0.02fF
C4780 fc2.n2320 a_400_38200# 0.12fF
C4781 fc2.n2322 a_400_38200# 0.03fF
C4782 fc2.n2323 a_400_38200# 0.01fF
C4783 fc2.n2324 a_400_38200# 0.06fF
C4784 fc2.n2325 a_400_38200# 0.24fF
C4785 fc2.n2326 a_400_38200# 0.33fF
C4786 fc2.n2327 a_400_38200# 0.05fF
C4787 fc2.n2328 a_400_38200# 0.03fF
C4788 fc2.n2329 a_400_38200# 0.13fF
C4789 fc2.n2330 a_400_38200# 0.06fF
C4790 fc2.n2331 a_400_38200# 0.11fF
C4791 fc2.n2332 a_400_38200# 0.03fF
C4792 fc2.n2333 a_400_38200# 0.05fF
C4793 fc2.n2334 a_400_38200# 0.05fF
C4794 fc2.n2335 a_400_38200# 0.09fF
C4795 fc2.n2336 a_400_38200# 0.03fF
C4796 fc2.n2337 a_400_38200# 0.07fF
C4797 fc2.n2338 a_400_38200# 0.32fF
C4798 fc2.n2339 a_400_38200# 0.47fF
C4799 fc2.n2340 a_400_38200# 0.29fF
C4800 fc2.n2341 a_400_38200# 3.32fF
C4801 fc2.t93 a_400_38200# 0.02fF
C4802 fc2.n2342 a_400_38200# 0.10fF
C4803 fc2.n2343 a_400_38200# 0.12fF
C4804 fc2.t31 a_400_38200# 0.02fF
C4805 fc2.n2345 a_400_38200# 0.21fF
C4806 fc2.n2346 a_400_38200# 0.80fF
C4807 fc2.n2347 a_400_38200# 0.04fF
C4808 fc2.n2348 a_400_38200# 1.79fF
C4809 fc2.n2349 a_400_38200# 0.05fF
C4810 fc2.n2350 a_400_38200# 0.07fF
C4811 fc2.n2351 a_400_38200# 1.17fF
C4812 fc2.n2352 a_400_38200# 0.12fF
C4813 fc2.n2353 a_400_38200# 0.05fF
C4814 fc2.n2354 a_400_38200# 0.17fF
C4815 fc2.n2355 a_400_38200# 0.06fF
C4816 fc2.n2356 a_400_38200# 0.03fF
C4817 fc2.n2357 a_400_38200# 0.10fF
C4818 fc2.n2358 a_400_38200# 0.17fF
C4819 fc2.n2359 a_400_38200# 0.69fF
C4820 fc2.t18 a_400_38200# 0.02fF
C4821 fc2.n2360 a_400_38200# 0.21fF
C4822 fc2.n2361 a_400_38200# 0.31fF
C4823 fc2.n2362 a_400_38200# 0.53fF
C4824 fc2.n2363 a_400_38200# 0.10fF
C4825 fc2.t234 a_400_38200# 0.02fF
C4826 fc2.n2364 a_400_38200# 0.12fF
C4827 fc2.n2366 a_400_38200# 0.01fF
C4828 fc2.n2367 a_400_38200# 0.03fF
C4829 fc2.n2368 a_400_38200# 0.06fF
C4830 fc2.n2369 a_400_38200# 0.24fF
C4831 fc2.n2370 a_400_38200# 0.05fF
C4832 fc2.n2371 a_400_38200# 0.03fF
C4833 fc2.n2372 a_400_38200# 0.33fF
C4834 fc2.n2373 a_400_38200# 0.13fF
C4835 fc2.n2374 a_400_38200# 0.06fF
C4836 fc2.n2375 a_400_38200# 0.11fF
C4837 fc2.n2376 a_400_38200# 0.03fF
C4838 fc2.n2377 a_400_38200# 0.07fF
C4839 fc2.n2378 a_400_38200# 0.03fF
C4840 fc2.n2379 a_400_38200# 0.05fF
C4841 fc2.n2380 a_400_38200# 0.05fF
C4842 fc2.n2381 a_400_38200# 0.09fF
C4843 fc2.n2382 a_400_38200# 0.32fF
C4844 fc2.n2383 a_400_38200# 0.47fF
C4845 fc2.n2384 a_400_38200# 0.29fF
C4846 fc2.n2385 a_400_38200# 1.64fF
C4847 fc2.t351 a_400_38200# 0.02fF
C4848 fc2.n2386 a_400_38200# 0.10fF
C4849 fc2.n2387 a_400_38200# 0.12fF
C4850 fc2.t280 a_400_38200# 0.02fF
C4851 fc2.n2389 a_400_38200# 0.21fF
C4852 fc2.n2390 a_400_38200# 0.80fF
C4853 fc2.n2391 a_400_38200# 0.04fF
C4854 fc2.n2392 a_400_38200# 0.46fF
C4855 fc2.n2393 a_400_38200# 0.52fF
C4856 fc2.n2394 a_400_38200# 0.46fF
C4857 fc2.n2395 a_400_38200# 1.04fF
C4858 fc2.n2396 a_400_38200# 0.12fF
C4859 fc2.n2397 a_400_38200# 0.52fF
C4860 fc2.n2398 a_400_38200# 0.10fF
C4861 fc2.t123 a_400_38200# 0.02fF
C4862 fc2.n2399 a_400_38200# 0.12fF
C4863 fc2.t287 a_400_38200# 0.02fF
C4864 fc2.n2401 a_400_38200# 0.21fF
C4865 fc2.n2402 a_400_38200# 0.31fF
C4866 fc2.n2403 a_400_38200# 0.53fF
C4867 fc2.n2404 a_400_38200# 0.05fF
C4868 fc2.n2405 a_400_38200# 0.17fF
C4869 fc2.n2406 a_400_38200# 0.06fF
C4870 fc2.n2407 a_400_38200# 0.03fF
C4871 fc2.n2408 a_400_38200# 0.10fF
C4872 fc2.n2409 a_400_38200# 0.17fF
C4873 fc2.n2410 a_400_38200# 0.69fF
C4874 fc2.n2411 a_400_38200# 0.05fF
C4875 fc2.n2412 a_400_38200# 0.07fF
C4876 fc2.n2413 a_400_38200# 1.00fF
C4877 fc2.n2414 a_400_38200# 0.12fF
C4878 fc2.n2415 a_400_38200# 3.32fF
C4879 fc2.t214 a_400_38200# 0.02fF
C4880 fc2.n2416 a_400_38200# 0.10fF
C4881 fc2.n2417 a_400_38200# 0.12fF
C4882 fc2.t165 a_400_38200# 0.02fF
C4883 fc2.n2419 a_400_38200# 0.21fF
C4884 fc2.n2420 a_400_38200# 0.80fF
C4885 fc2.n2421 a_400_38200# 0.04fF
C4886 fc2.t23 a_400_38200# 16.88fF
C4887 fc2.t223 a_400_38200# 0.02fF
C4888 fc2.n2422 a_400_38200# 0.01fF
C4889 fc2.n2423 a_400_38200# 0.22fF
C4890 fc2.t153 a_400_38200# 0.02fF
C4891 fc2.n2425 a_400_38200# 1.04fF
C4892 fc2.n2426 a_400_38200# 0.04fF
C4893 fc2.t271 a_400_38200# 0.02fF
C4894 fc2.n2427 a_400_38200# 0.56fF
C4895 fc2.n2428 a_400_38200# 0.53fF
C4896 fc2.n2429 a_400_38200# 0.52fF
C4897 fc2.n2430 a_400_38200# 0.15fF
C4898 fc2.n2431 a_400_38200# 0.77fF
C4899 fc2.n2432 a_400_38200# 0.52fF
C4900 fc2.n2433 a_400_38200# 0.07fF
C4901 fc2.n2434 a_400_38200# 1.89fF
C4902 fc2.n2435 a_400_38200# 0.52fF
C4903 fc2.n2436 a_400_38200# 0.19fF
C4904 fc2.n2437 a_400_38200# 1.28fF
C4905 fc2.t0 a_400_38200# 7.96fF
C4906 fc2.n2439 a_400_38200# 7.30fF
C4907 fc2.n2441 a_400_38200# 1.22fF
C4908 fc2.n2442 a_400_38200# 3.88fF
C4909 fc2.n2443 a_400_38200# 2.29fF
C4910 fc2.n2444 a_400_38200# 3.86fF
C4911 fc2.n2445 a_400_38200# 0.30fF
C4912 fc2.n2446 a_400_38200# 0.09fF
C4913 fc2.n2447 a_400_38200# 0.18fF
C4914 fc2.n2448 a_400_38200# 0.05fF
C4915 fc2.n2449 a_400_38200# 0.02fF
C4916 fc2.n2450 a_400_38200# 0.04fF
C4917 fc2.n2451 a_400_38200# 0.20fF
C4918 fc2.n2452 a_400_38200# 1.01fF
C4919 fc2.n2453 a_400_38200# 0.02fF
C4920 fc2.n2454 a_400_38200# 7.70fF
C4921 fc2.n2455 a_400_38200# 0.53fF
C4922 fc2.n2456 a_400_38200# 1.00fF
C4923 fc2.n2457 a_400_38200# 0.23fF
C4924 fc2.n2458 a_400_38200# 0.74fF
C4925 fc2.t115 a_400_38200# 0.02fF
C4926 fc2.n2459 a_400_38200# 0.21fF
C4927 fc2.n2460 a_400_38200# 0.31fF
C4928 fc2.n2461 a_400_38200# 0.53fF
C4929 fc2.n2462 a_400_38200# 0.10fF
C4930 fc2.t315 a_400_38200# 0.02fF
C4931 fc2.n2463 a_400_38200# 0.12fF
C4932 fc2.n2465 a_400_38200# 0.11fF
C4933 fc2.n2466 a_400_38200# 0.64fF
C4934 fc2.n2467 a_400_38200# 0.05fF
C4935 fc2.n2468 a_400_38200# 0.03fF
C4936 fc2.n2470 a_400_38200# 1.07fF
C4937 fc2.n2471 a_400_38200# 0.21fF
C4938 fc2.n2472 a_400_38200# 3.25fF
C4939 fc2.t39 a_400_38200# 0.02fF
C4940 fc2.n2473 a_400_38200# 0.10fF
C4941 fc2.n2474 a_400_38200# 0.12fF
C4942 fc2.t359 a_400_38200# 0.02fF
C4943 fc2.n2476 a_400_38200# 0.21fF
C4944 fc2.n2477 a_400_38200# 0.80fF
C4945 fc2.n2478 a_400_38200# 0.04fF
C4946 fc2.n2479 a_400_38200# 2.19fF
C4947 fc2.n2480 a_400_38200# 2.41fF
C4948 fc2.t54 a_400_38200# 0.02fF
C4949 fc2.n2481 a_400_38200# 0.21fF
C4950 fc2.n2482 a_400_38200# 0.31fF
C4951 fc2.n2483 a_400_38200# 0.53fF
C4952 fc2.n2484 a_400_38200# 0.10fF
C4953 fc2.t259 a_400_38200# 0.02fF
C4954 fc2.n2485 a_400_38200# 0.12fF
C4955 fc2.n2487 a_400_38200# 0.10fF
C4956 fc2.n2488 a_400_38200# 0.26fF
C4957 fc2.n2489 a_400_38200# 0.12fF
C4958 fc2.n2490 a_400_38200# 0.27fF
C4959 fc2.n2491 a_400_38200# 0.05fF
C4960 fc2.n2492 a_400_38200# 0.05fF
C4961 fc2.n2493 a_400_38200# 0.03fF
C4962 fc2.n2494 a_400_38200# 0.13fF
C4963 fc2.n2495 a_400_38200# 0.13fF
C4964 fc2.n2496 a_400_38200# 0.03fF
C4965 fc2.n2497 a_400_38200# 0.05fF
C4966 fc2.n2498 a_400_38200# 0.05fF
C4967 fc2.n2499 a_400_38200# 0.06fF
C4968 fc2.n2500 a_400_38200# 0.05fF
C4969 fc2.n2501 a_400_38200# 0.03fF
C4970 fc2.n2502 a_400_38200# 0.04fF
C4971 fc2.n2503 a_400_38200# 0.07fF
C4972 fc2.n2504 a_400_38200# 0.15fF
C4973 fc2.n2505 a_400_38200# 0.52fF
C4974 fc2.n2506 a_400_38200# 0.32fF
C4975 fc2.n2507 a_400_38200# 3.82fF
C4976 fc2.t356 a_400_38200# 0.02fF
C4977 fc2.n2508 a_400_38200# 0.10fF
C4978 fc2.n2509 a_400_38200# 0.12fF
C4979 fc2.t303 a_400_38200# 0.02fF
C4980 fc2.n2511 a_400_38200# 0.21fF
C4981 fc2.n2512 a_400_38200# 0.80fF
C4982 fc2.n2513 a_400_38200# 0.04fF
C4983 fc2.n2514 a_400_38200# 0.05fF
C4984 fc2.n2515 a_400_38200# 0.05fF
C4985 fc2.n2516 a_400_38200# 0.03fF
C4986 fc2.n2517 a_400_38200# 0.12fF
C4987 fc2.n2518 a_400_38200# 0.27fF
C4988 fc2.n2519 a_400_38200# 0.13fF
C4989 fc2.n2520 a_400_38200# 0.13fF
C4990 fc2.n2521 a_400_38200# 0.03fF
C4991 fc2.n2522 a_400_38200# 0.07fF
C4992 fc2.n2523 a_400_38200# 0.03fF
C4993 fc2.n2524 a_400_38200# 0.05fF
C4994 fc2.n2525 a_400_38200# 0.05fF
C4995 fc2.n2526 a_400_38200# 0.09fF
C4996 fc2.n2527 a_400_38200# 0.32fF
C4997 fc2.n2528 a_400_38200# 0.49fF
C4998 fc2.n2529 a_400_38200# 0.32fF
C4999 fc2.n2530 a_400_38200# 0.10fF
C5000 fc2.n2531 a_400_38200# 0.26fF
C5001 fc2.n2532 a_400_38200# 1.76fF
C5002 fc2.n2533 a_400_38200# 0.10fF
C5003 fc2.t134 a_400_38200# 0.02fF
C5004 fc2.n2534 a_400_38200# 0.12fF
C5005 fc2.t298 a_400_38200# 0.02fF
C5006 fc2.n2536 a_400_38200# 0.21fF
C5007 fc2.n2537 a_400_38200# 0.31fF
C5008 fc2.n2538 a_400_38200# 0.53fF
C5009 fc2.n2539 a_400_38200# 2.67fF
C5010 fc2.n2540 a_400_38200# 1.99fF
C5011 fc2.t227 a_400_38200# 0.02fF
C5012 fc2.n2541 a_400_38200# 0.10fF
C5013 fc2.n2542 a_400_38200# 0.12fF
C5014 fc2.t175 a_400_38200# 0.02fF
C5015 fc2.n2544 a_400_38200# 0.21fF
C5016 fc2.n2545 a_400_38200# 0.80fF
C5017 fc2.n2546 a_400_38200# 0.04fF
C5018 fc2.n2547 a_400_38200# 2.53fF
C5019 fc2.t170 a_400_38200# 0.02fF
C5020 fc2.n2548 a_400_38200# 0.21fF
C5021 fc2.n2549 a_400_38200# 0.31fF
C5022 fc2.n2550 a_400_38200# 0.53fF
C5023 fc2.n2551 a_400_38200# 0.10fF
C5024 fc2.t375 a_400_38200# 0.02fF
C5025 fc2.n2552 a_400_38200# 0.12fF
C5026 fc2.n2554 a_400_38200# 0.10fF
C5027 fc2.n2555 a_400_38200# 0.26fF
C5028 fc2.n2556 a_400_38200# 0.12fF
C5029 fc2.n2557 a_400_38200# 0.27fF
C5030 fc2.n2558 a_400_38200# 0.05fF
C5031 fc2.n2559 a_400_38200# 0.05fF
C5032 fc2.n2560 a_400_38200# 0.03fF
C5033 fc2.n2561 a_400_38200# 0.13fF
C5034 fc2.n2562 a_400_38200# 0.13fF
C5035 fc2.n2563 a_400_38200# 0.03fF
C5036 fc2.n2564 a_400_38200# 0.04fF
C5037 fc2.n2565 a_400_38200# 0.07fF
C5038 fc2.n2566 a_400_38200# 0.03fF
C5039 fc2.n2567 a_400_38200# 0.05fF
C5040 fc2.n2568 a_400_38200# 0.05fF
C5041 fc2.n2569 a_400_38200# 0.06fF
C5042 fc2.n2570 a_400_38200# 0.05fF
C5043 fc2.n2571 a_400_38200# 0.15fF
C5044 fc2.n2572 a_400_38200# 0.52fF
C5045 fc2.n2573 a_400_38200# 0.32fF
C5046 fc2.n2574 a_400_38200# 1.69fF
C5047 fc2.n2575 a_400_38200# 2.00fF
C5048 fc2.t107 a_400_38200# 0.02fF
C5049 fc2.n2576 a_400_38200# 0.10fF
C5050 fc2.n2577 a_400_38200# 0.12fF
C5051 fc2.t45 a_400_38200# 0.02fF
C5052 fc2.n2579 a_400_38200# 0.21fF
C5053 fc2.n2580 a_400_38200# 0.80fF
C5054 fc2.n2581 a_400_38200# 0.04fF
C5055 fc2.t367 a_400_38200# 0.02fF
C5056 fc2.n2582 a_400_38200# 0.10fF
C5057 fc2.n2583 a_400_38200# 0.12fF
C5058 fc2.n2584 a_400_38200# 0.21fF
C5059 fc2.t292 a_400_38200# 0.02fF
C5060 fc2.n2585 a_400_38200# 0.31fF
C5061 fc2.n2586 a_400_38200# 0.32fF
C5062 fc2.n2587 a_400_38200# 0.59fF
C5063 fc2.n2588 a_400_38200# 0.05fF
C5064 fc2.n2589 a_400_38200# 0.05fF
C5065 fc2.n2590 a_400_38200# 0.03fF
C5066 fc2.n2591 a_400_38200# 0.12fF
C5067 fc2.n2592 a_400_38200# 0.27fF
C5068 fc2.n2593 a_400_38200# 0.13fF
C5069 fc2.n2594 a_400_38200# 0.13fF
C5070 fc2.n2595 a_400_38200# 0.03fF
C5071 fc2.n2596 a_400_38200# 0.07fF
C5072 fc2.n2597 a_400_38200# 0.03fF
C5073 fc2.n2598 a_400_38200# 0.05fF
C5074 fc2.n2599 a_400_38200# 0.05fF
C5075 fc2.n2600 a_400_38200# 0.09fF
C5076 fc2.n2601 a_400_38200# 0.32fF
C5077 fc2.n2602 a_400_38200# 0.49fF
C5078 fc2.n2603 a_400_38200# 0.32fF
C5079 fc2.n2604 a_400_38200# 0.10fF
C5080 fc2.n2605 a_400_38200# 0.26fF
C5081 fc2.n2606 a_400_38200# 1.76fF
C5082 fc2.n2607 a_400_38200# 2.79fF
C5083 fc2.n2608 a_400_38200# 0.90fF
C5084 fc2.n2609 a_400_38200# 0.21fF
C5085 fc2.t36 a_400_38200# 0.02fF
C5086 fc2.n2610 a_400_38200# 0.31fF
C5087 fc2.n2611 a_400_38200# 0.55fF
C5088 fc2.n2612 a_400_38200# 0.35fF
C5089 fc2.n2613 a_400_38200# 0.35fF
C5090 fc2.n2615 a_400_38200# 0.10fF
C5091 fc2.t247 a_400_38200# 0.02fF
C5092 fc2.n2616 a_400_38200# 0.12fF
C5093 fc2.t330 a_400_38200# 0.02fF
C5094 fc2.n2618 a_400_38200# 0.21fF
C5095 fc2.n2619 a_400_38200# 0.31fF
C5096 fc2.n2620 a_400_38200# 0.53fF
C5097 fc2.t184 a_400_38200# 0.02fF
C5098 fc2.n2621 a_400_38200# 0.21fF
C5099 fc2.n2622 a_400_38200# 0.81fF
C5100 fc2.n2623 a_400_38200# 0.03fF
C5101 fc2.n2624 a_400_38200# 0.04fF
C5102 fc2.n2625 a_400_38200# 0.07fF
C5103 fc2.n2626 a_400_38200# 0.06fF
C5104 fc2.n2627 a_400_38200# 0.28fF
C5105 fc2.n2628 a_400_38200# 0.55fF
C5106 fc2.n2629 a_400_38200# 1.42fF
C5107 fc2.n2630 a_400_38200# 1.84fF
C5108 fc2.t295 a_400_38200# 0.02fF
C5109 fc2.n2631 a_400_38200# 0.10fF
C5110 fc2.n2632 a_400_38200# 0.12fF
C5111 fc2.n2633 a_400_38200# 0.10fF
C5112 fc2.t284 a_400_38200# 0.02fF
C5113 fc2.n2634 a_400_38200# 0.12fF
C5114 fc2.t90 a_400_38200# 0.02fF
C5115 fc2.n2635 a_400_38200# 1.06fF
C5116 fc2.n2636 a_400_38200# 1.21fF
C5117 fc2.n2637 a_400_38200# 1.01fF
C5118 fc2.n2638 a_400_38200# 1.29fF
C5119 fc2.t69 a_400_38200# 7.96fF
C5120 fc2.n2639 a_400_38200# 0.74fF
C5121 fc2.n2640 a_400_38200# 9.42fF
C5122 fc2.n2642 a_400_38200# 0.33fF
C5123 fc2.n2643 a_400_38200# 0.20fF
C5124 fc2.n2644 a_400_38200# 3.17fF
C5125 fc2.n2645 a_400_38200# 2.26fF
C5126 fc2.n2646 a_400_38200# 0.03fF
C5127 fc2.n2647 a_400_38200# 0.07fF
C5128 fc2.n2648 a_400_38200# 0.05fF
C5129 fc2.n2649 a_400_38200# 0.04fF
C5130 fc2.n2650 a_400_38200# 0.64fF
C5131 fc2.n2651 a_400_38200# 1.86fF
C5132 fc2.n2652 a_400_38200# 3.79fF
C5133 fc2.n2653 a_400_38200# 0.22fF
C5134 fc2.n2654 a_400_38200# 0.01fF
C5135 fc2.t334 a_400_38200# 0.02fF
C5136 fc2.n2655 a_400_38200# 0.22fF
C5137 fc2.t255 a_400_38200# 0.02fF
C5138 fc2.n2656 a_400_38200# 0.83fF
C5139 fc2.n2657 a_400_38200# 0.62fF
C5140 fc2.n2658 a_400_38200# 7.70fF
C5141 fc2.n2659 a_400_38200# 1.95fF
C5142 fc2.t20 a_400_38200# 0.02fF
C5143 fc2.n2660 a_400_38200# 0.21fF
C5144 fc2.n2661 a_400_38200# 0.31fF
C5145 fc2.n2662 a_400_38200# 0.53fF
C5146 fc2.n2663 a_400_38200# 0.10fF
C5147 fc2.t275 a_400_38200# 0.02fF
C5148 fc2.n2664 a_400_38200# 0.12fF
C5149 fc2.n2666 a_400_38200# 0.06fF
C5150 fc2.n2667 a_400_38200# 0.28fF
C5151 fc2.n2668 a_400_38200# 0.03fF
C5152 fc2.n2669 a_400_38200# 0.04fF
C5153 fc2.n2670 a_400_38200# 0.07fF
C5154 fc2.n2671 a_400_38200# 0.62fF
C5155 fc2.n2672 a_400_38200# 1.42fF
C5156 fc2.n2673 a_400_38200# 1.54fF
C5157 fc2.t307 a_400_38200# 0.02fF
C5158 fc2.n2674 a_400_38200# 0.10fF
C5159 fc2.n2675 a_400_38200# 0.12fF
C5160 fc2.t195 a_400_38200# 0.02fF
C5161 fc2.n2677 a_400_38200# 0.21fF
C5162 fc2.n2678 a_400_38200# 0.80fF
C5163 fc2.n2679 a_400_38200# 0.04fF
C5164 fc2.n2680 a_400_38200# 0.03fF
C5165 fc2.n2681 a_400_38200# 0.04fF
C5166 fc2.n2682 a_400_38200# 0.07fF
C5167 fc2.n2683 a_400_38200# 0.06fF
C5168 fc2.n2684 a_400_38200# 0.28fF
C5169 fc2.n2685 a_400_38200# 0.55fF
C5170 fc2.n2686 a_400_38200# 1.42fF
C5171 fc2.n2687 a_400_38200# 1.85fF
C5172 fc2.n2688 a_400_38200# 0.10fF
C5173 fc2.t149 a_400_38200# 0.02fF
C5174 fc2.n2689 a_400_38200# 0.12fF
C5175 fc2.t272 a_400_38200# 0.02fF
C5176 fc2.n2691 a_400_38200# 0.21fF
C5177 fc2.n2692 a_400_38200# 0.31fF
C5178 fc2.n2693 a_400_38200# 0.53fF
C5179 fc2.n2694 a_400_38200# 3.50fF
C5180 fc2.t178 a_400_38200# 0.02fF
C5181 fc2.n2695 a_400_38200# 0.10fF
C5182 fc2.n2696 a_400_38200# 0.12fF
C5183 fc2.t70 a_400_38200# 0.02fF
C5184 fc2.n2698 a_400_38200# 0.21fF
C5185 fc2.n2699 a_400_38200# 0.80fF
C5186 fc2.n2700 a_400_38200# 0.04fF
C5187 fc2.n2701 a_400_38200# 0.72fF
C5188 fc2.n2702 a_400_38200# 0.03fF
C5189 fc2.n2703 a_400_38200# 0.04fF
C5190 fc2.n2704 a_400_38200# 0.07fF
C5191 fc2.n2705 a_400_38200# 0.06fF
C5192 fc2.n2706 a_400_38200# 0.05fF
C5193 fc2.n2707 a_400_38200# 0.15fF
C5194 fc2.n2708 a_400_38200# 0.52fF
C5195 fc2.n2709 a_400_38200# 0.82fF
C5196 fc2.n2710 a_400_38200# 0.36fF
C5197 fc2.n2711 a_400_38200# 2.01fF
C5198 fc2.n2712 a_400_38200# 0.10fF
C5199 fc2.t5 a_400_38200# 0.02fF
C5200 fc2.n2713 a_400_38200# 0.12fF
C5201 fc2.t148 a_400_38200# 0.02fF
C5202 fc2.n2715 a_400_38200# 0.21fF
C5203 fc2.n2716 a_400_38200# 0.31fF
C5204 fc2.n2717 a_400_38200# 0.53fF
C5205 fc2.n2718 a_400_38200# 3.24fF
C5206 fc2.t49 a_400_38200# 0.02fF
C5207 fc2.n2719 a_400_38200# 0.10fF
C5208 fc2.n2720 a_400_38200# 0.12fF
C5209 fc2.t313 a_400_38200# 0.02fF
C5210 fc2.n2722 a_400_38200# 0.21fF
C5211 fc2.n2723 a_400_38200# 0.80fF
C5212 fc2.n2724 a_400_38200# 0.04fF
C5213 fc2.n2725 a_400_38200# 1.78fF
C5214 fc2.t283 a_400_38200# 0.02fF
C5215 fc2.n2726 a_400_38200# 0.21fF
C5216 fc2.n2727 a_400_38200# 0.31fF
C5217 fc2.n2728 a_400_38200# 0.53fF
C5218 fc2.n2729 a_400_38200# 0.10fF
C5219 fc2.t159 a_400_38200# 0.02fF
C5220 fc2.n2730 a_400_38200# 0.12fF
C5221 fc2.n2732 a_400_38200# 0.36fF
C5222 fc2.n2733 a_400_38200# 0.72fF
C5223 fc2.n2734 a_400_38200# 0.05fF
C5224 fc2.n2735 a_400_38200# 0.08fF
C5225 fc2.n2736 a_400_38200# 0.08fF
C5226 fc2.n2737 a_400_38200# 0.36fF
C5227 fc2.n2738 a_400_38200# 0.49fF
C5228 fc2.n2739 a_400_38200# 0.82fF
C5229 fc2.n2740 a_400_38200# 3.54fF
C5230 fc2.t167 a_400_38200# 0.02fF
C5231 fc2.n2741 a_400_38200# 0.10fF
C5232 fc2.n2742 a_400_38200# 0.12fF
C5233 fc2.t77 a_400_38200# 0.02fF
C5234 fc2.n2744 a_400_38200# 0.21fF
C5235 fc2.n2745 a_400_38200# 0.80fF
C5236 fc2.n2746 a_400_38200# 0.04fF
C5237 fc2.n2747 a_400_38200# 0.21fF
C5238 fc2.t390 a_400_38200# 0.02fF
C5239 fc2.n2748 a_400_38200# 0.80fF
C5240 fc2.t4 a_400_38200# 20.79fF
C5241 fc2.t129 a_400_38200# 0.02fF
C5242 fc2.n2749 a_400_38200# 0.21fF
C5243 fc2.n2750 a_400_38200# 0.80fF
C5244 fc2.n2751 a_400_38200# 0.04fF
C5245 fc2.t233 a_400_38200# 0.02fF
C5246 fc2.n2752 a_400_38200# 0.10fF
C5247 fc2.n2753 a_400_38200# 0.12fF
C5248 fc2.n2755 a_400_38200# 0.10fF
C5249 fc2.t204 a_400_38200# 0.02fF
C5250 fc2.n2756 a_400_38200# 0.12fF
C5251 fc2.n2758 a_400_38200# 0.03fF
C5252 fc2.n2759 a_400_38200# 0.08fF
C5253 fc2.n2760 a_400_38200# 0.19fF
C5254 fc2.n2761 a_400_38200# 0.69fF
C5255 fc2.n2762 a_400_38200# 0.05fF
C5256 fc2.n2763 a_400_38200# 0.06fF
C5257 fc2.n2764 a_400_38200# 1.12fF
C5258 fc2.n2765 a_400_38200# 0.12fF
C5259 fc2.n2766 a_400_38200# 5.20fF
C5260 fc2.n2767 a_400_38200# 2.75fF
C5261 fc2.t182 a_400_38200# 0.02fF
C5262 fc2.n2768 a_400_38200# 0.21fF
C5263 fc2.n2769 a_400_38200# 0.31fF
C5264 fc2.n2770 a_400_38200# 0.53fF
C5265 fc2.n2771 a_400_38200# 0.10fF
C5266 fc2.t386 a_400_38200# 0.02fF
C5267 fc2.n2772 a_400_38200# 0.12fF
C5268 fc2.n2774 a_400_38200# 0.52fF
C5269 fc2.n2775 a_400_38200# 0.72fF
C5270 fc2.n2776 a_400_38200# 1.49fF
C5271 fc2.n2777 a_400_38200# 3.95fF
C5272 fc2.t288 a_400_38200# 0.02fF
C5273 fc2.n2778 a_400_38200# 0.10fF
C5274 fc2.n2779 a_400_38200# 0.12fF
C5275 fc2.t61 a_400_38200# 0.02fF
C5276 fc2.n2781 a_400_38200# 0.21fF
C5277 fc2.n2782 a_400_38200# 0.80fF
C5278 fc2.n2783 a_400_38200# 0.04fF
C5279 fc2.t38 a_400_38200# 16.88fF
C5280 fc2.t237 a_400_38200# 0.02fF
C5281 fc2.n2784 a_400_38200# 0.01fF
C5282 fc2.n2785 a_400_38200# 0.22fF
C5283 fc2.t164 a_400_38200# 0.02fF
C5284 fc2.n2787 a_400_38200# 1.04fF
C5285 fc2.n2788 a_400_38200# 0.04fF
C5286 fc2.t286 a_400_38200# 0.02fF
C5287 fc2.n2789 a_400_38200# 0.56fF
C5288 fc2.n2790 a_400_38200# 0.53fF
C5289 fc2.n2791 a_400_38200# 0.52fF
C5290 fc2.n2792 a_400_38200# 0.15fF
C5291 fc2.n2793 a_400_38200# 0.77fF
C5292 fc2.n2794 a_400_38200# 0.52fF
C5293 fc2.n2795 a_400_38200# 0.07fF
C5294 fc2.n2796 a_400_38200# 1.89fF
C5295 fc2.n2797 a_400_38200# 0.52fF
C5296 fc2.n2798 a_400_38200# 0.19fF
C5297 fc2.n2799 a_400_38200# 1.28fF
C5298 fc2.t19 a_400_38200# 7.96fF
C5299 fc2.n2801 a_400_38200# 7.30fF
C5300 fc2.n2803 a_400_38200# 1.22fF
C5301 fc2.n2804 a_400_38200# 3.88fF
C5302 fc2.n2805 a_400_38200# 2.28fF
C5303 fc2.n2806 a_400_38200# 3.93fF
C5304 fc2.n2807 a_400_38200# 135.03fF
C5305 fc2.n2808 a_400_38200# 2.19fF
C5306 fc2.t579 a_400_38200# -0.02fF
C5307 fc2.n2809 a_400_38200# 0.57fF
C5308 fc2.t562 a_400_38200# -0.02fF
C5309 fc2.n2810 a_400_38200# 0.21fF
C5310 fc2.t428 a_400_38200# -0.01fF
C5311 fc2.n2811 a_400_38200# 0.56fF
C5312 fc2.n2812 a_400_38200# 2.83fF
C5313 fc2.n2813 a_400_38200# 1.64fF
C5314 fc2.n2814 a_400_38200# 2.39fF
C5315 fc2.t589 a_400_38200# -0.06fF
C5316 fc2.n2815 a_400_38200# 0.62fF
C5317 fc2.t457 a_400_38200# -0.02fF
C5318 fc2.n2816 a_400_38200# 0.21fF
C5319 fc2.t570 a_400_38200# -0.02fF
C5320 fc2.n2818 a_400_38200# 0.21fF
C5321 fc2.t708 a_400_38200# -0.06fF
C5322 fc2.n2819 a_400_38200# 0.62fF
C5323 fc2.n2821 a_400_38200# 1.72fF
C5324 fc2.t643 a_400_38200# -0.06fF
C5325 fc2.n2822 a_400_38200# 0.26fF
C5326 fc2.t432 a_400_38200# 0.00fF
C5327 fc2.n2823 a_400_38200# 0.34fF
C5328 fc2.t706 a_400_38200# -0.00fF
C5329 fc2.n2824 a_400_38200# 0.34fF
C5330 fc2.n2825 a_400_38200# 12.20fF
C5331 fc2.n2826 a_400_38200# 1.96fF
C5332 fc2.t509 a_400_38200# -0.06fF
C5333 fc2.n2827 a_400_38200# 0.62fF
C5334 fc2.t455 a_400_38200# -0.02fF
C5335 fc2.n2828 a_400_38200# 0.21fF
C5336 fc2.t750 a_400_38200# -0.02fF
C5337 fc2.n2830 a_400_38200# 0.21fF
C5338 fc2.t677 a_400_38200# -0.06fF
C5339 fc2.n2831 a_400_38200# 0.62fF
C5340 fc2.n2833 a_400_38200# 2.39fF
C5341 fc2.n2834 a_400_38200# 2.28fF
C5342 fc2.n2835 a_400_38200# 1.61fF
C5343 fc2.n2836 a_400_38200# 2.34fF
C5344 fc2.t461 a_400_38200# -0.06fF
C5345 fc2.n2837 a_400_38200# 0.62fF
C5346 fc2.t581 a_400_38200# -0.02fF
C5347 fc2.n2838 a_400_38200# 0.21fF
C5348 fc2.t556 a_400_38200# -0.02fF
C5349 fc2.n2840 a_400_38200# 0.21fF
C5350 fc2.t595 a_400_38200# -0.06fF
C5351 fc2.n2841 a_400_38200# 0.62fF
C5352 fc2.n2843 a_400_38200# 2.38fF
C5353 fc2.n2844 a_400_38200# 2.30fF
C5354 fc2.n2845 a_400_38200# 1.61fF
C5355 fc2.t600 a_400_38200# -0.02fF
C5356 fc2.n2846 a_400_38200# 0.21fF
C5357 fc2.t425 a_400_38200# -0.06fF
C5358 fc2.n2847 a_400_38200# 0.62fF
C5359 fc2.t663 a_400_38200# -0.02fF
C5360 fc2.n2849 a_400_38200# 0.21fF
C5361 fc2.t737 a_400_38200# -0.06fF
C5362 fc2.n2850 a_400_38200# 0.62fF
C5363 fc2.n2852 a_400_38200# 2.11fF
C5364 fc2.n2853 a_400_38200# 1.87fF
C5365 fc2.n2854 a_400_38200# 2.29fF
C5366 fc2.n2855 a_400_38200# 1.61fF
C5367 fc2.n2856 a_400_38200# 2.39fF
C5368 fc2.t636 a_400_38200# -0.06fF
C5369 fc2.n2857 a_400_38200# 0.62fF
C5370 fc2.t634 a_400_38200# -0.02fF
C5371 fc2.n2858 a_400_38200# 0.21fF
C5372 fc2.t616 a_400_38200# -0.02fF
C5373 fc2.n2860 a_400_38200# 0.21fF
C5374 fc2.t749 a_400_38200# -0.06fF
C5375 fc2.n2861 a_400_38200# 0.62fF
C5376 fc2.n2863 a_400_38200# 1.87fF
C5377 fc2.n2864 a_400_38200# 2.30fF
C5378 fc2.n2865 a_400_38200# 1.61fF
C5379 fc2.t705 a_400_38200# -0.02fF
C5380 fc2.n2866 a_400_38200# 0.21fF
C5381 fc2.t700 a_400_38200# -0.06fF
C5382 fc2.n2867 a_400_38200# 0.62fF
C5383 fc2.t660 a_400_38200# -0.02fF
C5384 fc2.n2869 a_400_38200# 0.21fF
C5385 fc2.t690 a_400_38200# -0.06fF
C5386 fc2.n2870 a_400_38200# 0.62fF
C5387 fc2.n2872 a_400_38200# 2.39fF
C5388 fc2.n2873 a_400_38200# 1.87fF
C5389 fc2.n2874 a_400_38200# 2.29fF
C5390 fc2.n2875 a_400_38200# 1.61fF
C5391 fc2.n2876 a_400_38200# 2.39fF
C5392 fc2.t508 a_400_38200# -0.06fF
C5393 fc2.n2877 a_400_38200# 0.62fF
C5394 fc2.t622 a_400_38200# -0.02fF
C5395 fc2.n2878 a_400_38200# 0.21fF
C5396 fc2.t654 a_400_38200# -0.02fF
C5397 fc2.n2880 a_400_38200# 0.21fF
C5398 fc2.t667 a_400_38200# -0.06fF
C5399 fc2.n2881 a_400_38200# 0.62fF
C5400 fc2.n2883 a_400_38200# 1.87fF
C5401 fc2.n2884 a_400_38200# 2.30fF
C5402 fc2.n2885 a_400_38200# 1.61fF
C5403 fc2.t739 a_400_38200# -0.02fF
C5404 fc2.n2886 a_400_38200# 0.21fF
C5405 fc2.t631 a_400_38200# -0.06fF
C5406 fc2.n2887 a_400_38200# 0.62fF
C5407 fc2.t575 a_400_38200# -0.02fF
C5408 fc2.n2889 a_400_38200# 0.21fF
C5409 fc2.t671 a_400_38200# -0.06fF
C5410 fc2.n2890 a_400_38200# 0.62fF
C5411 fc2.n2892 a_400_38200# 2.39fF
C5412 fc2.n2893 a_400_38200# 1.87fF
C5413 fc2.n2894 a_400_38200# 2.29fF
C5414 fc2.n2895 a_400_38200# 2.31fF
C5415 fc2.n2896 a_400_38200# 1.70fF
C5416 fc2.n2897 a_400_38200# 1.39fF
C5417 fc2.n2898 a_400_38200# 2.09fF
C5418 fc2.n2899 a_400_38200# 2.19fF
C5419 fc2.t620 a_400_38200# -0.02fF
C5420 fc2.n2900 a_400_38200# 0.57fF
C5421 fc2.t630 a_400_38200# -0.02fF
C5422 fc2.n2901 a_400_38200# 0.21fF
C5423 fc2.t476 a_400_38200# -0.01fF
C5424 fc2.n2902 a_400_38200# 0.56fF
C5425 fc2.n2903 a_400_38200# 2.83fF
C5426 fc2.n2904 a_400_38200# 1.64fF
C5427 fc2.n2905 a_400_38200# 2.39fF
C5428 fc2.t639 a_400_38200# -0.06fF
C5429 fc2.n2906 a_400_38200# 0.62fF
C5430 fc2.t512 a_400_38200# -0.02fF
C5431 fc2.n2907 a_400_38200# 0.21fF
C5432 fc2.t718 a_400_38200# -0.02fF
C5433 fc2.n2909 a_400_38200# 0.21fF
C5434 fc2.t605 a_400_38200# -0.06fF
C5435 fc2.n2910 a_400_38200# 0.62fF
C5436 fc2.n2912 a_400_38200# 1.72fF
C5437 fc2.t741 a_400_38200# -0.06fF
C5438 fc2.n2913 a_400_38200# 0.26fF
C5439 fc2.t524 a_400_38200# 0.00fF
C5440 fc2.n2914 a_400_38200# 0.34fF
C5441 fc2.t613 a_400_38200# -0.00fF
C5442 fc2.n2915 a_400_38200# 0.34fF
C5443 fc2.n2916 a_400_38200# 12.20fF
C5444 fc2.n2917 a_400_38200# 1.96fF
C5445 fc2.t629 a_400_38200# -0.06fF
C5446 fc2.n2918 a_400_38200# 0.62fF
C5447 fc2.t527 a_400_38200# -0.02fF
C5448 fc2.n2919 a_400_38200# 0.21fF
C5449 fc2.t406 a_400_38200# -0.02fF
C5450 fc2.n2921 a_400_38200# 0.21fF
C5451 fc2.t462 a_400_38200# -0.06fF
C5452 fc2.n2922 a_400_38200# 0.62fF
C5453 fc2.n2924 a_400_38200# 2.39fF
C5454 fc2.n2925 a_400_38200# 2.28fF
C5455 fc2.n2926 a_400_38200# 1.61fF
C5456 fc2.n2927 a_400_38200# 2.34fF
C5457 fc2.t496 a_400_38200# -0.06fF
C5458 fc2.n2928 a_400_38200# 0.62fF
C5459 fc2.t724 a_400_38200# -0.02fF
C5460 fc2.n2929 a_400_38200# 0.21fF
C5461 fc2.t646 a_400_38200# -0.02fF
C5462 fc2.n2931 a_400_38200# 0.21fF
C5463 fc2.t430 a_400_38200# -0.06fF
C5464 fc2.n2932 a_400_38200# 0.62fF
C5465 fc2.n2934 a_400_38200# 2.38fF
C5466 fc2.n2935 a_400_38200# 2.30fF
C5467 fc2.n2936 a_400_38200# 1.61fF
C5468 fc2.t618 a_400_38200# -0.02fF
C5469 fc2.n2937 a_400_38200# 0.21fF
C5470 fc2.t664 a_400_38200# -0.06fF
C5471 fc2.n2938 a_400_38200# 0.62fF
C5472 fc2.t538 a_400_38200# -0.02fF
C5473 fc2.n2940 a_400_38200# 0.21fF
C5474 fc2.t624 a_400_38200# -0.06fF
C5475 fc2.n2941 a_400_38200# 0.62fF
C5476 fc2.n2943 a_400_38200# 2.11fF
C5477 fc2.n2944 a_400_38200# 1.87fF
C5478 fc2.n2945 a_400_38200# 2.29fF
C5479 fc2.n2946 a_400_38200# 2.31fF
C5480 fc2.n2947 a_400_38200# 1.70fF
C5481 fc2.n2948 a_400_38200# 1.39fF
C5482 fc2.n2949 a_400_38200# 2.09fF
C5483 fc2.n2950 a_400_38200# 1.59fF
C5484 fc2.n2951 a_400_38200# 2.49fF
C5485 fc2.t557 a_400_38200# -0.02fF
C5486 fc2.n2952 a_400_38200# 0.57fF
C5487 fc2.t415 a_400_38200# -0.02fF
C5488 fc2.n2953 a_400_38200# 0.21fF
C5489 fc2.t740 a_400_38200# -0.01fF
C5490 fc2.n2954 a_400_38200# 0.56fF
C5491 fc2.n2955 a_400_38200# 2.29fF
C5492 fc2.t523 a_400_38200# -0.06fF
C5493 fc2.n2956 a_400_38200# 0.26fF
C5494 fc2.t719 a_400_38200# 0.00fF
C5495 fc2.n2957 a_400_38200# 0.34fF
C5496 fc2.t715 a_400_38200# -0.00fF
C5497 fc2.n2958 a_400_38200# 0.34fF
C5498 fc2.n2959 a_400_38200# 11.12fF
C5499 fc2.n2960 a_400_38200# 2.54fF
C5500 fc2.n2961 a_400_38200# 138.87fF
C5501 fc2.n2962 a_400_38200# 2.83fF
C5502 fc2.t472 a_400_38200# -0.02fF
C5503 fc2.n2963 a_400_38200# 0.21fF
C5504 fc2.t642 a_400_38200# -0.01fF
C5505 fc2.n2964 a_400_38200# 0.56fF
C5506 fc2.t514 a_400_38200# -0.02fF
C5507 fc2.n2965 a_400_38200# 0.57fF
C5508 fc2.n2966 a_400_38200# 1.91fF
C5509 fc2.n2967 a_400_38200# 1.65fF
C5510 fc2.n2968 a_400_38200# 2.34fF
C5511 fc2.t720 a_400_38200# -0.06fF
C5512 fc2.n2969 a_400_38200# 0.62fF
C5513 fc2.t418 a_400_38200# -0.02fF
C5514 fc2.n2970 a_400_38200# 0.21fF
C5515 fc2.t488 a_400_38200# -0.02fF
C5516 fc2.n2972 a_400_38200# 0.21fF
C5517 fc2.t444 a_400_38200# -0.06fF
C5518 fc2.n2973 a_400_38200# 0.62fF
C5519 fc2.n2975 a_400_38200# 2.30fF
C5520 fc2.n2976 a_400_38200# 2.20fF
C5521 fc2.n2977 a_400_38200# 1.96fF
C5522 fc2.t445 a_400_38200# -0.06fF
C5523 fc2.n2978 a_400_38200# 0.62fF
C5524 fc2.t722 a_400_38200# -0.02fF
C5525 fc2.n2979 a_400_38200# 0.21fF
C5526 fc2.t714 a_400_38200# -0.02fF
C5527 fc2.n2981 a_400_38200# 0.21fF
C5528 fc2.t468 a_400_38200# -0.06fF
C5529 fc2.n2982 a_400_38200# 0.62fF
C5530 fc2.n2984 a_400_38200# 2.28fF
C5531 fc2.n2985 a_400_38200# 2.21fF
C5532 fc2.t693 a_400_38200# 0.00fF
C5533 fc2.t450 a_400_38200# -0.06fF
C5534 fc2.n2986 a_400_38200# 0.26fF
C5535 fc2.n2987 a_400_38200# 0.34fF
C5536 fc2.t467 a_400_38200# 0.00fF
C5537 fc2.n2988 a_400_38200# 0.34fF
C5538 fc2.n2989 a_400_38200# 11.39fF
C5539 fc2.n2990 a_400_38200# 2.07fF
C5540 fc2.n2991 a_400_38200# 1.71fF
C5541 fc2.n2992 a_400_38200# 2.26fF
C5542 fc2.n2993 a_400_38200# 2.19fF
C5543 fc2.t704 a_400_38200# -0.02fF
C5544 fc2.n2994 a_400_38200# 0.57fF
C5545 fc2.t601 a_400_38200# -0.02fF
C5546 fc2.n2995 a_400_38200# 0.21fF
C5547 fc2.t572 a_400_38200# -0.01fF
C5548 fc2.n2996 a_400_38200# 0.56fF
C5549 fc2.n2997 a_400_38200# 2.83fF
C5550 fc2.n2998 a_400_38200# 1.64fF
C5551 fc2.n2999 a_400_38200# 2.39fF
C5552 fc2.t563 a_400_38200# -0.06fF
C5553 fc2.n3000 a_400_38200# 0.62fF
C5554 fc2.t419 a_400_38200# -0.02fF
C5555 fc2.n3001 a_400_38200# 0.21fF
C5556 fc2.t437 a_400_38200# -0.02fF
C5557 fc2.n3003 a_400_38200# 0.21fF
C5558 fc2.t492 a_400_38200# -0.06fF
C5559 fc2.n3004 a_400_38200# 0.62fF
C5560 fc2.n3006 a_400_38200# 1.72fF
C5561 fc2.t531 a_400_38200# -0.06fF
C5562 fc2.n3007 a_400_38200# 0.26fF
C5563 fc2.t471 a_400_38200# 0.00fF
C5564 fc2.n3008 a_400_38200# 0.34fF
C5565 fc2.t443 a_400_38200# -0.00fF
C5566 fc2.n3009 a_400_38200# 0.34fF
C5567 fc2.n3010 a_400_38200# 12.20fF
C5568 fc2.n3011 a_400_38200# 1.96fF
C5569 fc2.t483 a_400_38200# -0.06fF
C5570 fc2.n3012 a_400_38200# 0.62fF
C5571 fc2.t522 a_400_38200# -0.02fF
C5572 fc2.n3013 a_400_38200# 0.21fF
C5573 fc2.t626 a_400_38200# -0.02fF
C5574 fc2.n3015 a_400_38200# 0.21fF
C5575 fc2.t482 a_400_38200# -0.06fF
C5576 fc2.n3016 a_400_38200# 0.62fF
C5577 fc2.n3018 a_400_38200# 2.39fF
C5578 fc2.n3019 a_400_38200# 2.28fF
C5579 fc2.n3020 a_400_38200# 1.61fF
C5580 fc2.n3021 a_400_38200# 2.34fF
C5581 fc2.t426 a_400_38200# -0.06fF
C5582 fc2.n3022 a_400_38200# 0.62fF
C5583 fc2.t695 a_400_38200# -0.02fF
C5584 fc2.n3023 a_400_38200# 0.21fF
C5585 fc2.t497 a_400_38200# -0.02fF
C5586 fc2.n3025 a_400_38200# 0.21fF
C5587 fc2.t421 a_400_38200# -0.06fF
C5588 fc2.n3026 a_400_38200# 0.62fF
C5589 fc2.n3028 a_400_38200# 2.38fF
C5590 fc2.n3029 a_400_38200# 2.30fF
C5591 fc2.n3030 a_400_38200# 1.61fF
C5592 fc2.t438 a_400_38200# -0.02fF
C5593 fc2.n3031 a_400_38200# 0.21fF
C5594 fc2.t578 a_400_38200# -0.06fF
C5595 fc2.n3032 a_400_38200# 0.62fF
C5596 fc2.t685 a_400_38200# -0.02fF
C5597 fc2.n3034 a_400_38200# 0.21fF
C5598 fc2.t552 a_400_38200# -0.06fF
C5599 fc2.n3035 a_400_38200# 0.62fF
C5600 fc2.n3037 a_400_38200# 2.11fF
C5601 fc2.n3038 a_400_38200# 1.87fF
C5602 fc2.n3039 a_400_38200# 2.29fF
C5603 fc2.n3040 a_400_38200# 1.61fF
C5604 fc2.n3041 a_400_38200# 2.39fF
C5605 fc2.t498 a_400_38200# -0.06fF
C5606 fc2.n3042 a_400_38200# 0.62fF
C5607 fc2.t507 a_400_38200# -0.02fF
C5608 fc2.n3043 a_400_38200# 0.21fF
C5609 fc2.t707 a_400_38200# -0.02fF
C5610 fc2.n3045 a_400_38200# 0.21fF
C5611 fc2.t478 a_400_38200# -0.06fF
C5612 fc2.n3046 a_400_38200# 0.62fF
C5613 fc2.n3048 a_400_38200# 1.87fF
C5614 fc2.n3049 a_400_38200# 2.30fF
C5615 fc2.n3050 a_400_38200# 1.61fF
C5616 fc2.t573 a_400_38200# -0.02fF
C5617 fc2.n3051 a_400_38200# 0.21fF
C5618 fc2.t717 a_400_38200# -0.06fF
C5619 fc2.n3052 a_400_38200# 0.62fF
C5620 fc2.t623 a_400_38200# -0.02fF
C5621 fc2.n3054 a_400_38200# 0.21fF
C5622 fc2.t500 a_400_38200# -0.06fF
C5623 fc2.n3055 a_400_38200# 0.62fF
C5624 fc2.n3057 a_400_38200# 2.39fF
C5625 fc2.n3058 a_400_38200# 1.87fF
C5626 fc2.n3059 a_400_38200# 2.29fF
C5627 fc2.n3060 a_400_38200# 2.31fF
C5628 fc2.n3061 a_400_38200# 1.70fF
C5629 fc2.n3062 a_400_38200# 1.39fF
C5630 fc2.n3063 a_400_38200# 2.09fF
C5631 fc2.n3064 a_400_38200# 2.19fF
C5632 fc2.t394 a_400_38200# -0.02fF
C5633 fc2.n3065 a_400_38200# 0.57fF
C5634 fc2.t611 a_400_38200# -0.02fF
C5635 fc2.n3066 a_400_38200# 0.21fF
C5636 fc2.t526 a_400_38200# -0.01fF
C5637 fc2.n3067 a_400_38200# 0.56fF
C5638 fc2.n3068 a_400_38200# 2.83fF
C5639 fc2.n3069 a_400_38200# 1.64fF
C5640 fc2.n3070 a_400_38200# 2.39fF
C5641 fc2.t583 a_400_38200# -0.06fF
C5642 fc2.n3071 a_400_38200# 0.62fF
C5643 fc2.t423 a_400_38200# -0.02fF
C5644 fc2.n3072 a_400_38200# 0.21fF
C5645 fc2.t439 a_400_38200# -0.02fF
C5646 fc2.n3074 a_400_38200# 0.21fF
C5647 fc2.t672 a_400_38200# -0.06fF
C5648 fc2.n3075 a_400_38200# 0.62fF
C5649 fc2.n3077 a_400_38200# 1.72fF
C5650 fc2.t410 a_400_38200# -0.06fF
C5651 fc2.n3078 a_400_38200# 0.26fF
C5652 fc2.t547 a_400_38200# 0.00fF
C5653 fc2.n3079 a_400_38200# 0.34fF
C5654 fc2.t619 a_400_38200# -0.00fF
C5655 fc2.n3080 a_400_38200# 0.34fF
C5656 fc2.n3081 a_400_38200# 12.20fF
C5657 fc2.n3082 a_400_38200# 1.96fF
C5658 fc2.t540 a_400_38200# -0.06fF
C5659 fc2.n3083 a_400_38200# 0.62fF
C5660 fc2.t621 a_400_38200# -0.02fF
C5661 fc2.n3084 a_400_38200# 0.21fF
C5662 fc2.t680 a_400_38200# -0.02fF
C5663 fc2.n3086 a_400_38200# 0.21fF
C5664 fc2.t398 a_400_38200# -0.06fF
C5665 fc2.n3087 a_400_38200# 0.62fF
C5666 fc2.n3089 a_400_38200# 2.39fF
C5667 fc2.n3090 a_400_38200# 2.28fF
C5668 fc2.n3091 a_400_38200# 1.61fF
C5669 fc2.n3092 a_400_38200# 2.34fF
C5670 fc2.t548 a_400_38200# -0.06fF
C5671 fc2.n3093 a_400_38200# 0.62fF
C5672 fc2.t503 a_400_38200# -0.02fF
C5673 fc2.n3094 a_400_38200# 0.21fF
C5674 fc2.t559 a_400_38200# -0.02fF
C5675 fc2.n3096 a_400_38200# 0.21fF
C5676 fc2.t662 a_400_38200# -0.06fF
C5677 fc2.n3097 a_400_38200# 0.62fF
C5678 fc2.n3099 a_400_38200# 2.38fF
C5679 fc2.n3100 a_400_38200# 2.30fF
C5680 fc2.n3101 a_400_38200# 1.61fF
C5681 fc2.t659 a_400_38200# -0.02fF
C5682 fc2.n3102 a_400_38200# 0.21fF
C5683 fc2.t678 a_400_38200# -0.06fF
C5684 fc2.n3103 a_400_38200# 0.62fF
C5685 fc2.t473 a_400_38200# -0.02fF
C5686 fc2.n3105 a_400_38200# 0.21fF
C5687 fc2.t454 a_400_38200# -0.06fF
C5688 fc2.n3106 a_400_38200# 0.62fF
C5689 fc2.n3108 a_400_38200# 2.11fF
C5690 fc2.n3109 a_400_38200# 1.87fF
C5691 fc2.n3110 a_400_38200# 2.29fF
C5692 fc2.n3111 a_400_38200# 1.61fF
C5693 fc2.n3112 a_400_38200# 2.39fF
C5694 fc2.t549 a_400_38200# -0.06fF
C5695 fc2.n3113 a_400_38200# 0.62fF
C5696 fc2.t701 a_400_38200# -0.02fF
C5697 fc2.n3114 a_400_38200# 0.21fF
C5698 fc2.t734 a_400_38200# -0.02fF
C5699 fc2.n3116 a_400_38200# 0.21fF
C5700 fc2.t692 a_400_38200# -0.06fF
C5701 fc2.n3117 a_400_38200# 0.62fF
C5702 fc2.n3119 a_400_38200# 1.87fF
C5703 fc2.n3120 a_400_38200# 2.30fF
C5704 fc2.n3121 a_400_38200# 1.61fF
C5705 fc2.t747 a_400_38200# -0.02fF
C5706 fc2.n3122 a_400_38200# 0.21fF
C5707 fc2.t743 a_400_38200# -0.06fF
C5708 fc2.n3123 a_400_38200# 0.62fF
C5709 fc2.t480 a_400_38200# -0.02fF
C5710 fc2.n3125 a_400_38200# 0.21fF
C5711 fc2.t564 a_400_38200# -0.06fF
C5712 fc2.n3126 a_400_38200# 0.62fF
C5713 fc2.n3128 a_400_38200# 2.39fF
C5714 fc2.n3129 a_400_38200# 1.87fF
C5715 fc2.n3130 a_400_38200# 2.29fF
C5716 fc2.n3131 a_400_38200# 1.61fF
C5717 fc2.n3132 a_400_38200# 2.39fF
C5718 fc2.t520 a_400_38200# -0.06fF
C5719 fc2.n3133 a_400_38200# 0.62fF
C5720 fc2.t752 a_400_38200# -0.02fF
C5721 fc2.n3134 a_400_38200# 0.21fF
C5722 fc2.t417 a_400_38200# -0.02fF
C5723 fc2.n3136 a_400_38200# 0.21fF
C5724 fc2.t744 a_400_38200# -0.06fF
C5725 fc2.n3137 a_400_38200# 0.62fF
C5726 fc2.n3139 a_400_38200# 1.87fF
C5727 fc2.n3140 a_400_38200# 2.30fF
C5728 fc2.n3141 a_400_38200# 1.61fF
C5729 fc2.t459 a_400_38200# -0.02fF
C5730 fc2.n3142 a_400_38200# 0.21fF
C5731 fc2.t712 a_400_38200# -0.06fF
C5732 fc2.n3143 a_400_38200# 0.62fF
C5733 fc2.t447 a_400_38200# -0.02fF
C5734 fc2.n3145 a_400_38200# 0.21fF
C5735 fc2.t584 a_400_38200# -0.06fF
C5736 fc2.n3146 a_400_38200# 0.62fF
C5737 fc2.n3148 a_400_38200# 2.39fF
C5738 fc2.n3149 a_400_38200# 1.87fF
C5739 fc2.n3150 a_400_38200# 2.29fF
C5740 fc2.n3151 a_400_38200# 1.61fF
C5741 fc2.n3152 a_400_38200# 2.39fF
C5742 fc2.t491 a_400_38200# -0.06fF
C5743 fc2.n3153 a_400_38200# 0.62fF
C5744 fc2.t607 a_400_38200# -0.02fF
C5745 fc2.n3154 a_400_38200# 0.21fF
C5746 fc2.t723 a_400_38200# -0.02fF
C5747 fc2.n3156 a_400_38200# 0.21fF
C5748 fc2.t698 a_400_38200# -0.06fF
C5749 fc2.n3157 a_400_38200# 0.62fF
C5750 fc2.n3159 a_400_38200# 1.87fF
C5751 fc2.n3160 a_400_38200# 2.30fF
C5752 fc2.n3161 a_400_38200# 1.61fF
C5753 fc2.t554 a_400_38200# -0.02fF
C5754 fc2.n3162 a_400_38200# 0.21fF
C5755 fc2.t610 a_400_38200# -0.06fF
C5756 fc2.n3163 a_400_38200# 0.62fF
C5757 fc2.t580 a_400_38200# -0.02fF
C5758 fc2.n3165 a_400_38200# 0.21fF
C5759 fc2.t635 a_400_38200# -0.06fF
C5760 fc2.n3166 a_400_38200# 0.62fF
C5761 fc2.n3168 a_400_38200# 2.39fF
C5762 fc2.n3169 a_400_38200# 1.87fF
C5763 fc2.n3170 a_400_38200# 2.29fF
C5764 fc2.n3171 a_400_38200# 2.31fF
C5765 fc2.n3172 a_400_38200# 1.70fF
C5766 fc2.n3173 a_400_38200# 1.39fF
C5767 fc2.n3174 a_400_38200# 2.09fF
C5768 fc2.n3175 a_400_38200# 0.27fF
C5769 fc2.n3176 a_400_38200# 0.20fF
C5770 fc2.t745 a_400_38200# -0.00fF
C5771 fc2.t682 a_400_38200# -0.01fF
C5772 fc2.n3177 a_400_38200# 0.74fF
C5773 fc2.n3178 a_400_38200# 3.12fF
C5774 fc2.t558 a_400_38200# -0.02fF
C5775 fc2.t555 a_400_38200# 0.00fF
C5776 fc2.n3179 a_400_38200# 0.54fF
C5777 fc2.n3180 a_400_38200# 9.58fF
C5778 fc2.n3181 a_400_38200# 1.74fF
C5779 fc2.t568 a_400_38200# -0.02fF
C5780 fc2.n3182 a_400_38200# 0.21fF
C5781 fc2.t716 a_400_38200# -0.06fF
C5782 fc2.n3183 a_400_38200# 0.62fF
C5783 fc2.t529 a_400_38200# -0.02fF
C5784 fc2.n3185 a_400_38200# 0.21fF
C5785 fc2.t506 a_400_38200# -0.06fF
C5786 fc2.n3186 a_400_38200# 0.62fF
C5787 fc2.n3188 a_400_38200# 2.14fF
C5788 fc2.n3189 a_400_38200# 2.19fF
C5789 fc2.n3190 a_400_38200# 1.61fF
C5790 fc2.t416 a_400_38200# -0.02fF
C5791 fc2.n3191 a_400_38200# 0.21fF
C5792 fc2.t485 a_400_38200# -0.06fF
C5793 fc2.n3192 a_400_38200# 0.62fF
C5794 fc2.t458 a_400_38200# -0.02fF
C5795 fc2.n3194 a_400_38200# 0.21fF
C5796 fc2.t590 a_400_38200# -0.06fF
C5797 fc2.n3195 a_400_38200# 0.62fF
C5798 fc2.n3197 a_400_38200# 2.02fF
C5799 fc2.n3198 a_400_38200# 2.54fF
C5800 fc2.n3199 a_400_38200# 2.11fF
C5801 fc2.n3200 a_400_38200# 2.30fF
C5802 fc2.n3201 a_400_38200# 1.61fF
C5803 fc2.t699 a_400_38200# -0.02fF
C5804 fc2.n3202 a_400_38200# 0.21fF
C5805 fc2.t486 a_400_38200# -0.06fF
C5806 fc2.n3203 a_400_38200# 0.62fF
C5807 fc2.t501 a_400_38200# -0.02fF
C5808 fc2.n3205 a_400_38200# 0.21fF
C5809 fc2.t542 a_400_38200# -0.06fF
C5810 fc2.n3206 a_400_38200# 0.62fF
C5811 fc2.n3208 a_400_38200# 2.09fF
C5812 fc2.n3209 a_400_38200# 1.87fF
C5813 fc2.n3210 a_400_38200# 2.30fF
C5814 fc2.n3211 a_400_38200# 1.61fF
C5815 fc2.t675 a_400_38200# -0.02fF
C5816 fc2.n3212 a_400_38200# 0.21fF
C5817 fc2.t596 a_400_38200# -0.06fF
C5818 fc2.n3213 a_400_38200# 0.62fF
C5819 fc2.t442 a_400_38200# -0.02fF
C5820 fc2.n3215 a_400_38200# 0.21fF
C5821 fc2.t628 a_400_38200# -0.06fF
C5822 fc2.n3216 a_400_38200# 0.62fF
C5823 fc2.n3218 a_400_38200# 2.39fF
C5824 fc2.n3219 a_400_38200# 1.87fF
C5825 fc2.n3220 a_400_38200# 2.30fF
C5826 fc2.n3221 a_400_38200# 1.61fF
C5827 fc2.t713 a_400_38200# -0.02fF
C5828 fc2.n3222 a_400_38200# 0.21fF
C5829 fc2.t434 a_400_38200# -0.06fF
C5830 fc2.n3223 a_400_38200# 0.62fF
C5831 fc2.t736 a_400_38200# -0.02fF
C5832 fc2.n3225 a_400_38200# 0.21fF
C5833 fc2.t640 a_400_38200# -0.06fF
C5834 fc2.n3226 a_400_38200# 0.62fF
C5835 fc2.n3228 a_400_38200# 2.39fF
C5836 fc2.n3229 a_400_38200# 1.87fF
C5837 fc2.n3230 a_400_38200# 2.30fF
C5838 fc2.n3231 a_400_38200# 1.61fF
C5839 fc2.t644 a_400_38200# -0.02fF
C5840 fc2.n3232 a_400_38200# 0.21fF
C5841 fc2.t391 a_400_38200# -0.06fF
C5842 fc2.n3233 a_400_38200# 0.62fF
C5843 fc2.t574 a_400_38200# -0.02fF
C5844 fc2.n3235 a_400_38200# 0.21fF
C5845 fc2.t511 a_400_38200# -0.06fF
C5846 fc2.n3236 a_400_38200# 0.62fF
C5847 fc2.n3238 a_400_38200# 2.39fF
C5848 fc2.n3239 a_400_38200# 1.87fF
C5849 fc2.n3240 a_400_38200# 2.30fF
C5850 fc2.n3241 a_400_38200# 1.61fF
C5851 fc2.t545 a_400_38200# -0.02fF
C5852 fc2.n3242 a_400_38200# 0.21fF
C5853 fc2.t397 a_400_38200# -0.06fF
C5854 fc2.n3243 a_400_38200# 0.62fF
C5855 fc2.t615 a_400_38200# -0.02fF
C5856 fc2.n3245 a_400_38200# 0.21fF
C5857 fc2.t627 a_400_38200# -0.06fF
C5858 fc2.n3246 a_400_38200# 0.62fF
C5859 fc2.n3248 a_400_38200# 2.39fF
C5860 fc2.n3249 a_400_38200# 1.87fF
C5861 fc2.n3250 a_400_38200# 2.30fF
C5862 fc2.n3251 a_400_38200# 1.61fF
C5863 fc2.t691 a_400_38200# -0.02fF
C5864 fc2.n3252 a_400_38200# 0.21fF
C5865 fc2.t598 a_400_38200# -0.06fF
C5866 fc2.n3253 a_400_38200# 0.62fF
C5867 fc2.t694 a_400_38200# -0.02fF
C5868 fc2.n3255 a_400_38200# 0.21fF
C5869 fc2.t449 a_400_38200# -0.06fF
C5870 fc2.n3256 a_400_38200# 0.62fF
C5871 fc2.n3258 a_400_38200# 2.39fF
C5872 fc2.n3259 a_400_38200# 1.87fF
C5873 fc2.n3260 a_400_38200# 2.30fF
C5874 fc2.n3261 a_400_38200# 1.61fF
C5875 fc2.t436 a_400_38200# -0.02fF
C5876 fc2.n3262 a_400_38200# 0.21fF
C5877 fc2.t687 a_400_38200# -0.06fF
C5878 fc2.n3263 a_400_38200# 0.62fF
C5879 fc2.t499 a_400_38200# -0.02fF
C5880 fc2.n3265 a_400_38200# 0.21fF
C5881 fc2.t647 a_400_38200# -0.06fF
C5882 fc2.n3266 a_400_38200# 0.62fF
C5883 fc2.n3268 a_400_38200# 2.39fF
C5884 fc2.n3269 a_400_38200# 1.87fF
C5885 fc2.n3270 a_400_38200# 2.30fF
C5886 fc2.n3271 a_400_38200# 1.61fF
C5887 fc2.t477 a_400_38200# -0.02fF
C5888 fc2.n3272 a_400_38200# 0.21fF
C5889 fc2.t729 a_400_38200# -0.06fF
C5890 fc2.n3273 a_400_38200# 0.62fF
C5891 fc2.t532 a_400_38200# -0.02fF
C5892 fc2.n3275 a_400_38200# 0.21fF
C5893 fc2.t676 a_400_38200# -0.06fF
C5894 fc2.n3276 a_400_38200# 0.62fF
C5895 fc2.n3278 a_400_38200# 2.39fF
C5896 fc2.n3279 a_400_38200# 1.87fF
C5897 fc2.n3280 a_400_38200# 2.30fF
C5898 fc2.n3281 a_400_38200# 1.61fF
C5899 fc2.t725 a_400_38200# -0.02fF
C5900 fc2.n3282 a_400_38200# 0.21fF
C5901 fc2.t632 a_400_38200# -0.06fF
C5902 fc2.n3283 a_400_38200# 0.62fF
C5903 fc2.t727 a_400_38200# -0.02fF
C5904 fc2.n3285 a_400_38200# 0.21fF
C5905 fc2.t440 a_400_38200# -0.06fF
C5906 fc2.n3286 a_400_38200# 0.62fF
C5907 fc2.n3288 a_400_38200# 2.39fF
C5908 fc2.n3289 a_400_38200# 1.87fF
C5909 fc2.n3290 a_400_38200# 2.30fF
C5910 fc2.n3291 a_400_38200# 1.57fF
C5911 fc2.t565 a_400_38200# -0.02fF
C5912 fc2.n3292 a_400_38200# 0.21fF
C5913 fc2.t517 a_400_38200# -0.06fF
C5914 fc2.n3293 a_400_38200# 0.62fF
C5915 fc2.t502 a_400_38200# -0.02fF
C5916 fc2.n3295 a_400_38200# 0.21fF
C5917 fc2.t481 a_400_38200# -0.06fF
C5918 fc2.n3296 a_400_38200# 0.62fF
C5919 fc2.n3298 a_400_38200# 2.36fF
C5920 fc2.n3299 a_400_38200# 1.87fF
C5921 fc2.n3300 a_400_38200# 2.13fF
C5922 fc2.n3301 a_400_38200# 1.15fF
C5923 fc2.n3302 a_400_38200# 3.12fF
C5924 fc2.n3303 a_400_38200# 0.83fF
C5925 fc2.n3304 a_400_38200# 2.74fF
C5926 fc2.n3305 a_400_38200# 0.02fF
C5927 fc2.n3306 a_400_38200# 0.21fF
C5928 fc2.n3307 a_400_38200# 1.47fF
C5929 fc2.n3308 a_400_38200# 134.70fF
C5930 fc2.n3309 a_400_38200# 40.87fF
C5931 fc2.n3310 a_400_38200# 24.84fF
C5932 fc2.n3311 a_400_38200# 24.84fF
C5933 fc2.n3312 a_400_38200# 24.84fF
C5934 fc2.n3313 a_400_38200# 24.84fF
C5935 fc2.t22 a_400_38200# 0.02fF
C5936 fc2.n3314 a_400_38200# 1.14fF
C5937 fc2.n3315 a_400_38200# 0.16fF
C5938 fc2.n3316 a_400_38200# 24.10fF
C5939 fc2.n3317 a_400_38200# 13.94fF
C5940 fc2.n3318 a_400_38200# 13.51fF
C5941 fc2.n3319 a_400_38200# 10.63fF
C5942 fc2.n3320 a_400_38200# 25.07fF
C5943 fc2.n3321 a_400_38200# 3.48fF
C5944 fc2.n3322 a_400_38200# 10.76fF
C5945 fc2.n3323 a_400_38200# 13.59fF
C5946 fc2.n3324 a_400_38200# 10.76fF
C5947 fc2.n3325 a_400_38200# 13.59fF
C5948 fc2.n3326 a_400_38200# 10.76fF
C5949 fc2.n3327 a_400_38200# 25.09fF
C5950 fc2.n3328 a_400_38200# 3.46fF
C5951 fc2.n3329 a_400_38200# 25.44fF
C5952 fc2.n3330 a_400_38200# 3.78fF
C5953 fc2.n3331 a_400_38200# 3.78fF
C5954 fc2.n3332 a_400_38200# 3.99fF
C5955 fc2.n3333 a_400_38200# 3.78fF
C5956 fc2.n3334 a_400_38200# 3.78fF
C5957 fc2.n3335 a_400_38200# 40.47fF
C5958 fc2.n3336 a_400_38200# 3.79fF
C5959 fc2.n3337 a_400_38200# 3.03fF
C5960 fc2.n3338 a_400_38200# 0.16fF
C5961 fc2.n3339 a_400_38200# 8.14fF
C5962 fc2.n3340 a_400_38200# 0.22fF
C5963 fc2.t117 a_400_38200# 0.02fF
C5964 fc2.n3341 a_400_38200# 0.38fF
C5965 fc2.n3342 a_400_38200# 0.35fF
C5966 fc2.n3343 a_400_38200# 0.17fF
C5967 fc2.n3344 a_400_38200# 0.18fF
C5968 fc2.n3345 a_400_38200# 0.06fF
C5969 fc2.n3346 a_400_38200# 0.09fF
C5970 fc2.n3347 a_400_38200# 0.10fF
C5971 fc2.n3348 a_400_38200# 0.16fF
C5972 fc2.n3349 a_400_38200# 0.78fF
C5973 fc2.t65 a_400_38200# 0.02fF
C5974 fc2.n3350 a_400_38200# 0.78fF
C5975 fc2.t75 a_400_38200# 0.02fF
C5976 fc2.n3351 a_400_38200# 0.78fF
C5977 fc2.n3352 a_400_38200# 2.09fF
C5978 fc2.n3353 a_400_38200# 0.33fF
C5979 fc2.n3354 a_400_38200# 13.59fF
C5980 fc2.n3355 a_400_38200# 13.49fF
C5981 fc2.n3356 a_400_38200# 0.88fF
C5982 fc2.n3357 a_400_38200# 79.24fF
C5983 fc2.n3358 a_400_38200# 24.56fF
C5984 fc2.n3359 a_400_38200# 1.04fF
C5985 fc2.n3360 a_400_38200# 2.88fF
C5986 fc2.n3361 a_400_38200# 0.11fF
C5987 fc2.n3362 a_400_38200# 1.05fF
C5988 fc2.t333 a_400_38200# 0.02fF
C5989 fc2.n3363 a_400_38200# 0.01fF
C5990 fc2.n3364 a_400_38200# 0.32fF
C5991 fc2.n3365 a_400_38200# 1.75fF
C5992 fc2.t172 a_400_38200# 0.02fF
C5993 fc2.n3366 a_400_38200# 0.78fF
C5994 fc2.t200 a_400_38200# 0.02fF
C5995 fc2.n3367 a_400_38200# 0.78fF
C5996 fc2.n3368 a_400_38200# 2.09fF
C5997 fc2.n3369 a_400_38200# 0.33fF
C5998 fc2.n3370 a_400_38200# 13.59fF
C5999 fc2.n3371 a_400_38200# 10.76fF
C6000 fc2.n3372 a_400_38200# 0.88fF
C6001 fc2.n3373 a_400_38200# 24.48fF
C6002 fc2.n3374 a_400_38200# 1.32fF
C6003 fc2.n3375 a_400_38200# 2.44fF
C6004 fc2.n3376 a_400_38200# 0.11fF
C6005 fc2.n3377 a_400_38200# 1.05fF
C6006 fc2.t92 a_400_38200# 0.02fF
C6007 fc2.n3378 a_400_38200# 0.01fF
C6008 fc2.n3379 a_400_38200# 0.32fF
C6009 fc2.n3380 a_400_38200# 1.75fF
C6010 fc2.t299 a_400_38200# 0.02fF
C6011 fc2.n3381 a_400_38200# 0.78fF
C6012 fc2.t326 a_400_38200# 0.02fF
C6013 fc2.n3382 a_400_38200# 0.78fF
C6014 fc2.n3383 a_400_38200# 2.09fF
C6015 fc2.n3384 a_400_38200# 0.33fF
C6016 fc2.n3385 a_400_38200# 0.88fF
C6017 fc2.n3386 a_400_38200# 1.32fF
C6018 fc2.n3387 a_400_38200# 2.44fF
C6019 fc2.n3388 a_400_38200# 0.11fF
C6020 fc2.n3389 a_400_38200# 1.05fF
C6021 fc2.t213 a_400_38200# 0.02fF
C6022 fc2.n3390 a_400_38200# 0.01fF
C6023 fc2.n3391 a_400_38200# 0.32fF
C6024 fc2.n3392 a_400_38200# 1.01fF
C6025 fc2.n3393 a_400_38200# 0.01fF
C6026 fc2.n3394 a_400_38200# 0.28fF
C6027 fc2.t57 a_400_38200# 0.02fF
C6028 fc2.n3395 a_400_38200# 0.78fF
C6029 fc2.t85 a_400_38200# 0.02fF
C6030 fc2.n3396 a_400_38200# 0.78fF
C6031 fc2.n3397 a_400_38200# 2.09fF
C6032 fc2.n3398 a_400_38200# 0.33fF
C6033 fc2.n3399 a_400_38200# 0.88fF
C6034 fc2.n3400 a_400_38200# 0.08fF
C6035 fc2.n3402 a_400_38200# 0.42fF
C6036 fc2.n3403 a_400_38200# 1.27fF
C6037 fc2.n3404 a_400_38200# 2.06fF
C6038 fc2.n3405 a_400_38200# 0.11fF
C6039 fc2.n3406 a_400_38200# 1.05fF
C6040 fc2.t344 a_400_38200# 0.02fF
C6041 fc2.n3407 a_400_38200# 0.01fF
C6042 fc2.n3408 a_400_38200# 0.32fF
C6043 fc2.n3409 a_400_38200# 0.08fF
C6044 fc2.n3411 a_400_38200# 0.28fF
C6045 fc2.n3412 a_400_38200# 0.88fF
C6046 fc2.n3413 a_400_38200# 0.32fF
C6047 fc2.n3414 a_400_38200# 0.88fF
C6048 fc2.n3415 a_400_38200# 2.77fF
C6049 fc2.n3416 a_400_38200# 0.11fF
C6050 fc2.n3417 a_400_38200# 1.05fF
C6051 fc2.t353 a_400_38200# 0.02fF
C6052 fc2.n3418 a_400_38200# 0.78fF
C6053 fc2.t384 a_400_38200# 0.02fF
C6054 fc2.n3419 a_400_38200# 0.78fF
C6055 fc2.n3420 a_400_38200# 2.13fF
C6056 fc2.n3421 a_400_38200# 0.01fF
C6057 fc2.n3422 a_400_38200# 0.15fF
C6058 fc2.n3423 a_400_38200# 1.05fF
C6059 fc2.t273 a_400_38200# 0.02fF
C6060 fc2.n3424 a_400_38200# 0.01fF
C6061 fc2.n3425 a_400_38200# 0.32fF
C6062 fc2.n3426 a_400_38200# 0.49fF
C6063 fc2.n3427 a_400_38200# 0.63fF
C6064 fc2.n3428 a_400_38200# 0.78fF
C6065 fc2.n3429 a_400_38200# 0.35fF
C6066 fc2.n3430 a_400_38200# 0.17fF
C6067 fc2.n3431 a_400_38200# 0.09fF
C6068 fc2.n3432 a_400_38200# 0.10fF
C6069 fc2.n3433 a_400_38200# 0.16fF
C6070 fc2.n3434 a_400_38200# 1.37fF
C6071 fc2.n3435 a_400_38200# 2.85fF
C6072 fc2.n3436 a_400_38200# 79.14fF
C6073 fc2.n3437 a_400_38200# 1.04fF
C6074 fc2.n3438 a_400_38200# 0.78fF
C6075 fc2.t306 a_400_38200# 0.02fF
C6076 fc2.n3439 a_400_38200# 0.78fF
C6077 fc2.t314 a_400_38200# 0.02fF
C6078 fc2.n3440 a_400_38200# 0.78fF
C6079 fc2.t221 a_400_38200# 0.02fF
C6080 fc2.n3441 a_400_38200# 0.01fF
C6081 fc2.n3442 a_400_38200# 0.32fF
C6082 fc2.t56 a_400_38200# 38.43fF
C6083 fc2.n3443 a_400_38200# 2.05fF
C6084 fc2.n3444 a_400_38200# 79.46fF
C6085 fc2.n3445 a_400_38200# 307.24fF
C6086 fc2.n3446 a_400_38200# 0.05fF
C6087 fc2.n3447 a_400_38200# 0.10fF
C6088 fc2.n3448 a_400_38200# 0.03fF
C6089 fc2.n3449 a_400_38200# 0.04fF
C6090 fc2.n3450 a_400_38200# 0.68fF
C6091 fc2.n3451 a_400_38200# 0.25fF
C6092 fc2.n3452 a_400_38200# 0.08fF
C6093 fc2.n3453 a_400_38200# 0.10fF
C6094 fc2.n3454 a_400_38200# 0.11fF
C6095 fc2.n3455 a_400_38200# 0.46fF
C6096 fc2.n3456 a_400_38200# 0.05fF
C6097 fc2.n3457 a_400_38200# 0.24fF
C6098 fc2.n3458 a_400_38200# 2.12fF
C6099 fc2.t661 a_400_38200# -0.02fF
C6100 fc2.n3459 a_400_38200# 0.57fF
C6101 fc2.t587 a_400_38200# -0.02fF
C6102 fc2.n3460 a_400_38200# 0.21fF
C6103 fc2.t742 a_400_38200# -0.01fF
C6104 fc2.n3461 a_400_38200# 0.56fF
C6105 fc2.n3462 a_400_38200# 0.25fF
C6106 fc2.n3463 a_400_38200# 2.12fF
C6107 fc2.n3464 a_400_38200# 4.09fF
C6108 fc2.n3465 a_400_38200# 0.05fF
C6109 fc2.n3466 a_400_38200# 0.46fF
C6110 fc2.n3467 a_400_38200# 1.19fF
C6111 fc2.n3468 a_400_38200# 1.72fF
C6112 fc2.t537 a_400_38200# -0.02fF
C6113 fc2.n3469 a_400_38200# 0.21fF
C6114 fc2.t721 a_400_38200# -0.06fF
C6115 fc2.n3470 a_400_38200# 0.62fF
C6116 fc2.t609 a_400_38200# -0.02fF
C6117 fc2.n3472 a_400_38200# 0.21fF
C6118 fc2.t656 a_400_38200# -0.06fF
C6119 fc2.n3473 a_400_38200# 0.62fF
C6120 fc2.n3475 a_400_38200# 1.20fF
C6121 fc2.n3476 a_400_38200# 1.75fF
C6122 fc2.n3477 a_400_38200# 1.80fF
C6123 fc2.n3478 a_400_38200# 1.83fF
C6124 fc2.n3479 a_400_38200# 2.30fF
C6125 fc2.t474 a_400_38200# -0.02fF
C6126 fc2.n3480 a_400_38200# 0.21fF
C6127 fc2.t637 a_400_38200# -0.06fF
C6128 fc2.n3481 a_400_38200# 0.62fF
C6129 fc2.t731 a_400_38200# -0.02fF
C6130 fc2.n3483 a_400_38200# 0.21fF
C6131 fc2.t528 a_400_38200# -0.06fF
C6132 fc2.n3484 a_400_38200# 0.62fF
C6133 fc2.n3486 a_400_38200# 2.59fF
C6134 fc2.n3487 a_400_38200# 1.69fF
C6135 fc2.n3488 a_400_38200# 1.77fF
C6136 fc2.n3489 a_400_38200# 2.30fF
C6137 fc2.t681 a_400_38200# -0.02fF
C6138 fc2.n3490 a_400_38200# 0.21fF
C6139 fc2.t604 a_400_38200# -0.06fF
C6140 fc2.n3491 a_400_38200# 0.62fF
C6141 fc2.t400 a_400_38200# -0.02fF
C6142 fc2.n3493 a_400_38200# 0.21fF
C6143 fc2.t504 a_400_38200# -0.06fF
C6144 fc2.n3494 a_400_38200# 0.62fF
C6145 fc2.n3496 a_400_38200# 2.39fF
C6146 fc2.n3497 a_400_38200# 1.69fF
C6147 fc2.n3498 a_400_38200# 1.77fF
C6148 fc2.n3499 a_400_38200# 2.30fF
C6149 fc2.t470 a_400_38200# -0.02fF
C6150 fc2.n3500 a_400_38200# 0.21fF
C6151 fc2.t582 a_400_38200# -0.06fF
C6152 fc2.n3501 a_400_38200# 0.62fF
C6153 fc2.t606 a_400_38200# -0.02fF
C6154 fc2.n3503 a_400_38200# 0.21fF
C6155 fc2.t585 a_400_38200# -0.06fF
C6156 fc2.n3504 a_400_38200# 0.62fF
C6157 fc2.n3506 a_400_38200# 2.39fF
C6158 fc2.n3507 a_400_38200# 1.69fF
C6159 fc2.n3508 a_400_38200# 1.77fF
C6160 fc2.n3509 a_400_38200# 2.30fF
C6161 fc2.t401 a_400_38200# -0.02fF
C6162 fc2.n3510 a_400_38200# 0.21fF
C6163 fc2.t539 a_400_38200# -0.06fF
C6164 fc2.n3511 a_400_38200# 0.62fF
C6165 fc2.t489 a_400_38200# -0.02fF
C6166 fc2.n3513 a_400_38200# 0.21fF
C6167 fc2.t551 a_400_38200# -0.06fF
C6168 fc2.n3514 a_400_38200# 0.62fF
C6169 fc2.n3516 a_400_38200# 2.39fF
C6170 fc2.n3517 a_400_38200# 1.69fF
C6171 fc2.n3518 a_400_38200# 1.77fF
C6172 fc2.n3519 a_400_38200# 2.30fF
C6173 fc2.t469 a_400_38200# -0.02fF
C6174 fc2.n3520 a_400_38200# 0.21fF
C6175 fc2.t414 a_400_38200# -0.06fF
C6176 fc2.n3521 a_400_38200# 0.62fF
C6177 fc2.t567 a_400_38200# -0.02fF
C6178 fc2.n3523 a_400_38200# 0.21fF
C6179 fc2.t571 a_400_38200# -0.06fF
C6180 fc2.n3524 a_400_38200# 0.62fF
C6181 fc2.n3526 a_400_38200# 2.39fF
C6182 fc2.n3527 a_400_38200# 1.69fF
C6183 fc2.n3528 a_400_38200# 1.77fF
C6184 fc2.n3529 a_400_38200# 2.30fF
C6185 fc2.t413 a_400_38200# -0.02fF
C6186 fc2.n3530 a_400_38200# 0.21fF
C6187 fc2.t688 a_400_38200# -0.06fF
C6188 fc2.n3531 a_400_38200# 0.62fF
C6189 fc2.t746 a_400_38200# -0.02fF
C6190 fc2.n3533 a_400_38200# 0.21fF
C6191 fc2.t452 a_400_38200# -0.06fF
C6192 fc2.n3534 a_400_38200# 0.62fF
C6193 fc2.n3536 a_400_38200# 2.39fF
C6194 fc2.n3537 a_400_38200# 1.69fF
C6195 fc2.n3538 a_400_38200# 1.77fF
C6196 fc2.n3539 a_400_38200# 2.30fF
C6197 fc2.t466 a_400_38200# -0.02fF
C6198 fc2.n3540 a_400_38200# 0.21fF
C6199 fc2.t453 a_400_38200# -0.06fF
C6200 fc2.n3541 a_400_38200# 0.62fF
C6201 fc2.t429 a_400_38200# -0.02fF
C6202 fc2.n3543 a_400_38200# 0.21fF
C6203 fc2.t411 a_400_38200# -0.06fF
C6204 fc2.n3544 a_400_38200# 0.62fF
C6205 fc2.n3546 a_400_38200# 2.39fF
C6206 fc2.n3547 a_400_38200# 1.69fF
C6207 fc2.n3548 a_400_38200# 1.77fF
C6208 fc2.n3549 a_400_38200# 2.30fF
C6209 fc2.t543 a_400_38200# -0.02fF
C6210 fc2.n3550 a_400_38200# 0.21fF
C6211 fc2.t553 a_400_38200# -0.06fF
C6212 fc2.n3551 a_400_38200# 0.62fF
C6213 fc2.t521 a_400_38200# -0.02fF
C6214 fc2.n3553 a_400_38200# 0.21fF
C6215 fc2.t495 a_400_38200# -0.06fF
C6216 fc2.n3554 a_400_38200# 0.62fF
C6217 fc2.n3556 a_400_38200# 2.39fF
C6218 fc2.n3557 a_400_38200# 1.69fF
C6219 fc2.n3558 a_400_38200# 1.77fF
C6220 fc2.n3559 a_400_38200# 1.20fF
C6221 fc2.n3560 a_400_38200# 1.97fF
C6222 fc2.t617 a_400_38200# -0.02fF
C6223 fc2.n3561 a_400_38200# 0.21fF
C6224 fc2.t518 a_400_38200# -0.06fF
C6225 fc2.n3562 a_400_38200# 0.62fF
C6226 fc2.t703 a_400_38200# -0.02fF
C6227 fc2.n3564 a_400_38200# 0.21fF
C6228 fc2.t405 a_400_38200# -0.06fF
C6229 fc2.n3565 a_400_38200# 0.62fF
C6230 fc2.n3567 a_400_38200# 2.49fF
C6231 fc2.n3568 a_400_38200# 1.69fF
C6232 fc2.n3569 a_400_38200# 1.72fF
C6233 fc2.n3570 a_400_38200# 1.01fF
C6234 fc2.t633 a_400_38200# -0.06fF
C6235 fc2.n3571 a_400_38200# 0.26fF
C6236 fc2.t686 a_400_38200# 0.00fF
C6237 fc2.n3572 a_400_38200# 0.34fF
C6238 fc2.t487 a_400_38200# -0.00fF
C6239 fc2.n3573 a_400_38200# 0.34fF
C6240 fc2.n3574 a_400_38200# 0.03fF
C6241 fc2.n3575 a_400_38200# 0.04fF
C6242 fc2.n3576 a_400_38200# 0.68fF
C6243 fc2.n3577 a_400_38200# 0.25fF
C6244 fc2.n3578 a_400_38200# 0.08fF
C6245 fc2.n3579 a_400_38200# 0.11fF
C6246 fc2.n3580 a_400_38200# 0.84fF
C6247 fc2.n3581 a_400_38200# 1.91fF
C6248 fc2.n3582 a_400_38200# 0.05fF
C6249 fc2.n3583 a_400_38200# 0.36fF
C6250 fc2.n3584 a_400_38200# 0.38fF
C6251 fc2.n3585 a_400_38200# 0.74fF
C6252 fc2.n3586 a_400_38200# 0.05fF
C6253 fc2.n3587 a_400_38200# 0.10fF
C6254 fc2.n3588 a_400_38200# 0.03fF
C6255 fc2.n3589 a_400_38200# 0.04fF
C6256 fc2.n3590 a_400_38200# 0.68fF
C6257 fc2.n3591 a_400_38200# 0.25fF
C6258 fc2.n3592 a_400_38200# 0.08fF
C6259 fc2.n3593 a_400_38200# 0.10fF
C6260 fc2.n3594 a_400_38200# 0.11fF
C6261 fc2.n3595 a_400_38200# 0.46fF
C6262 fc2.n3596 a_400_38200# 0.05fF
C6263 fc2.n3597 a_400_38200# 0.24fF
C6264 fc2.n3598 a_400_38200# 2.12fF
C6265 fc2.t424 a_400_38200# -0.02fF
C6266 fc2.n3599 a_400_38200# 0.57fF
C6267 fc2.t683 a_400_38200# -0.02fF
C6268 fc2.n3600 a_400_38200# 0.21fF
C6269 fc2.t464 a_400_38200# -0.01fF
C6270 fc2.n3601 a_400_38200# 0.56fF
C6271 fc2.n3602 a_400_38200# 0.25fF
C6272 fc2.n3603 a_400_38200# 2.12fF
C6273 fc2.n3604 a_400_38200# 4.09fF
C6274 fc2.n3605 a_400_38200# 0.05fF
C6275 fc2.n3606 a_400_38200# 0.46fF
C6276 fc2.n3607 a_400_38200# 1.19fF
C6277 fc2.n3608 a_400_38200# 1.72fF
C6278 fc2.t597 a_400_38200# -0.02fF
C6279 fc2.n3609 a_400_38200# 0.21fF
C6280 fc2.t666 a_400_38200# -0.06fF
C6281 fc2.n3610 a_400_38200# 0.62fF
C6282 fc2.t655 a_400_38200# -0.02fF
C6283 fc2.n3612 a_400_38200# 0.21fF
C6284 fc2.t402 a_400_38200# -0.06fF
C6285 fc2.n3613 a_400_38200# 0.62fF
C6286 fc2.n3615 a_400_38200# 1.20fF
C6287 fc2.n3616 a_400_38200# 1.75fF
C6288 fc2.n3617 a_400_38200# 1.80fF
C6289 fc2.n3618 a_400_38200# 1.83fF
C6290 fc2.n3619 a_400_38200# 2.30fF
C6291 fc2.t396 a_400_38200# -0.02fF
C6292 fc2.n3620 a_400_38200# 0.21fF
C6293 fc2.t702 a_400_38200# -0.06fF
C6294 fc2.n3621 a_400_38200# 0.62fF
C6295 fc2.t550 a_400_38200# -0.02fF
C6296 fc2.n3623 a_400_38200# 0.21fF
C6297 fc2.t460 a_400_38200# -0.06fF
C6298 fc2.n3624 a_400_38200# 0.62fF
C6299 fc2.n3626 a_400_38200# 2.59fF
C6300 fc2.n3627 a_400_38200# 1.69fF
C6301 fc2.n3628 a_400_38200# 1.77fF
C6302 fc2.n3629 a_400_38200# 2.30fF
C6303 fc2.t479 a_400_38200# -0.02fF
C6304 fc2.n3630 a_400_38200# 0.21fF
C6305 fc2.t566 a_400_38200# -0.06fF
C6306 fc2.n3631 a_400_38200# 0.62fF
C6307 fc2.t673 a_400_38200# -0.02fF
C6308 fc2.n3633 a_400_38200# 0.21fF
C6309 fc2.t403 a_400_38200# -0.06fF
C6310 fc2.n3634 a_400_38200# 0.62fF
C6311 fc2.n3636 a_400_38200# 2.39fF
C6312 fc2.n3637 a_400_38200# 1.69fF
C6313 fc2.n3638 a_400_38200# 1.77fF
C6314 fc2.n3639 a_400_38200# 2.30fF
C6315 fc2.t638 a_400_38200# -0.02fF
C6316 fc2.n3640 a_400_38200# 0.21fF
C6317 fc2.t412 a_400_38200# -0.06fF
C6318 fc2.n3641 a_400_38200# 0.62fF
C6319 fc2.t544 a_400_38200# -0.02fF
C6320 fc2.n3643 a_400_38200# 0.21fF
C6321 fc2.t435 a_400_38200# -0.06fF
C6322 fc2.n3644 a_400_38200# 0.62fF
C6323 fc2.n3646 a_400_38200# 2.39fF
C6324 fc2.n3647 a_400_38200# 1.69fF
C6325 fc2.n3648 a_400_38200# 1.77fF
C6326 fc2.n3649 a_400_38200# 2.30fF
C6327 fc2.t561 a_400_38200# -0.02fF
C6328 fc2.n3650 a_400_38200# 0.21fF
C6329 fc2.t586 a_400_38200# -0.06fF
C6330 fc2.n3651 a_400_38200# 0.62fF
C6331 fc2.t404 a_400_38200# -0.02fF
C6332 fc2.n3653 a_400_38200# 0.21fF
C6333 fc2.t733 a_400_38200# -0.06fF
C6334 fc2.n3654 a_400_38200# 0.62fF
C6335 fc2.n3656 a_400_38200# 2.39fF
C6336 fc2.n3657 a_400_38200# 1.69fF
C6337 fc2.n3658 a_400_38200# 1.77fF
C6338 fc2.n3659 a_400_38200# 1.20fF
C6339 fc2.n3660 a_400_38200# 1.97fF
C6340 fc2.t433 a_400_38200# -0.02fF
C6341 fc2.n3661 a_400_38200# 0.21fF
C6342 fc2.t649 a_400_38200# -0.06fF
C6343 fc2.n3662 a_400_38200# 0.62fF
C6344 fc2.t456 a_400_38200# -0.02fF
C6345 fc2.n3664 a_400_38200# 0.21fF
C6346 fc2.t451 a_400_38200# -0.06fF
C6347 fc2.n3665 a_400_38200# 0.62fF
C6348 fc2.n3667 a_400_38200# 2.49fF
C6349 fc2.n3668 a_400_38200# 1.69fF
C6350 fc2.n3669 a_400_38200# 1.72fF
C6351 fc2.n3670 a_400_38200# 1.01fF
C6352 fc2.t748 a_400_38200# -0.06fF
C6353 fc2.n3671 a_400_38200# 0.26fF
C6354 fc2.t625 a_400_38200# 0.00fF
C6355 fc2.n3672 a_400_38200# 0.34fF
C6356 fc2.t603 a_400_38200# -0.00fF
C6357 fc2.n3673 a_400_38200# 0.34fF
C6358 fc2.n3674 a_400_38200# 0.03fF
C6359 fc2.n3675 a_400_38200# 0.04fF
C6360 fc2.n3676 a_400_38200# 0.68fF
C6361 fc2.n3677 a_400_38200# 0.25fF
C6362 fc2.n3678 a_400_38200# 0.08fF
C6363 fc2.n3679 a_400_38200# 0.11fF
C6364 fc2.n3680 a_400_38200# 0.84fF
C6365 fc2.n3681 a_400_38200# 1.91fF
C6366 fc2.n3682 a_400_38200# 0.05fF
C6367 fc2.n3683 a_400_38200# 0.36fF
C6368 fc2.n3684 a_400_38200# 0.38fF
C6369 fc2.n3685 a_400_38200# 0.74fF
C6370 fc2.n3686 a_400_38200# 0.05fF
C6371 fc2.n3687 a_400_38200# 2.70fF
C6372 fc2.t751 a_400_38200# -0.06fF
C6373 fc2.n3688 a_400_38200# 0.62fF
C6374 fc2.t602 a_400_38200# -0.02fF
C6375 fc2.n3689 a_400_38200# 0.21fF
C6376 fc2.t510 a_400_38200# -0.02fF
C6377 fc2.n3691 a_400_38200# 0.21fF
C6378 fc2.t653 a_400_38200# -0.06fF
C6379 fc2.n3692 a_400_38200# 0.62fF
C6380 fc2.n3694 a_400_38200# 1.20fF
C6381 fc2.n3695 a_400_38200# 1.96fF
C6382 fc2.n3696 a_400_38200# 1.69fF
C6383 fc2.n3697 a_400_38200# 0.05fF
C6384 fc2.n3698 a_400_38200# 0.46fF
C6385 fc2.n3699 a_400_38200# 1.19fF
C6386 fc2.n3700 a_400_38200# 1.73fF
C6387 fc2.t652 a_400_38200# -0.02fF
C6388 fc2.n3701 a_400_38200# 0.21fF
C6389 fc2.t668 a_400_38200# -0.06fF
C6390 fc2.n3702 a_400_38200# 0.62fF
C6391 fc2.t599 a_400_38200# -0.02fF
C6392 fc2.n3704 a_400_38200# 0.21fF
C6393 fc2.t463 a_400_38200# -0.06fF
C6394 fc2.n3705 a_400_38200# 0.62fF
C6395 fc2.n3707 a_400_38200# 1.75fF
C6396 fc2.n3708 a_400_38200# 1.80fF
C6397 fc2.n3709 a_400_38200# 0.25fF
C6398 fc2.n3710 a_400_38200# 2.12fF
C6399 fc2.t431 a_400_38200# -0.02fF
C6400 fc2.n3711 a_400_38200# 0.21fF
C6401 fc2.t730 a_400_38200# -0.01fF
C6402 fc2.n3712 a_400_38200# 0.56fF
C6403 fc2.t657 a_400_38200# -0.02fF
C6404 fc2.n3713 a_400_38200# 0.57fF
C6405 fc2.n3714 a_400_38200# 0.24fF
C6406 fc2.n3715 a_400_38200# 2.12fF
C6407 fc2.n3716 a_400_38200# 1.20fF
C6408 fc2.n3717 a_400_38200# 0.46fF
C6409 fc2.n3718 a_400_38200# 0.05fF
C6410 fc2.n3719 a_400_38200# 4.09fF
C6411 fc2.n3720 a_400_38200# 1.83fF
C6412 fc2.n3721 a_400_38200# 1.72fF
C6413 fc2.n3722 a_400_38200# 1.01fF
C6414 fc2.n3723 a_400_38200# 0.10fF
C6415 fc2.n3724 a_400_38200# 0.03fF
C6416 fc2.n3725 a_400_38200# 0.04fF
C6417 fc2.n3726 a_400_38200# 0.68fF
C6418 fc2.n3727 a_400_38200# 0.25fF
C6419 fc2.n3728 a_400_38200# 0.08fF
C6420 fc2.n3729 a_400_38200# 0.10fF
C6421 fc2.n3730 a_400_38200# 0.11fF
C6422 fc2.t593 a_400_38200# -0.06fF
C6423 fc2.n3731 a_400_38200# 0.26fF
C6424 fc2.t588 a_400_38200# 0.00fF
C6425 fc2.n3732 a_400_38200# 0.34fF
C6426 fc2.t689 a_400_38200# -0.00fF
C6427 fc2.n3733 a_400_38200# 0.34fF
C6428 fc2.n3734 a_400_38200# 0.03fF
C6429 fc2.n3735 a_400_38200# 0.04fF
C6430 fc2.n3736 a_400_38200# 0.68fF
C6431 fc2.n3737 a_400_38200# 0.25fF
C6432 fc2.n3738 a_400_38200# 0.08fF
C6433 fc2.n3739 a_400_38200# 0.11fF
C6434 fc2.n3740 a_400_38200# 0.84fF
C6435 fc2.n3741 a_400_38200# 1.91fF
C6436 fc2.n3742 a_400_38200# 0.05fF
C6437 fc2.n3743 a_400_38200# 0.36fF
C6438 fc2.n3744 a_400_38200# 0.38fF
C6439 fc2.n3745 a_400_38200# 0.74fF
C6440 fc2.n3746 a_400_38200# 0.12fF
C6441 fc2.n3747 a_400_38200# 1.88fF
C6442 fc2.t446 a_400_38200# -0.02fF
C6443 fc2.n3748 a_400_38200# 0.21fF
C6444 fc2.t422 a_400_38200# -0.01fF
C6445 fc2.n3749 a_400_38200# 0.56fF
C6446 fc2.t515 a_400_38200# -0.02fF
C6447 fc2.n3750 a_400_38200# 0.57fF
C6448 fc2.n3751 a_400_38200# 0.38fF
C6449 fc2.n3752 a_400_38200# 1.88fF
C6450 fc2.n3753 a_400_38200# 0.05fF
C6451 fc2.n3754 a_400_38200# 0.05fF
C6452 fc2.n3755 a_400_38200# 4.22fF
C6453 fc2.n3756 a_400_38200# 0.05fF
C6454 fc2.n3757 a_400_38200# 0.05fF
C6455 fc2.n3758 a_400_38200# 0.38fF
C6456 fc2.n3759 a_400_38200# 0.27fF
C6457 fc2.n3760 a_400_38200# 0.21fF
C6458 fc2.n3761 a_400_38200# 0.09fF
C6459 fc2.n3762 a_400_38200# 1.19fF
C6460 fc2.n3763 a_400_38200# 0.33fF
C6461 fc2.n3764 a_400_38200# 3.90fF
C6462 fc2.n3765 a_400_38200# 0.23fF
C6463 fc2.t490 a_400_38200# -0.06fF
C6464 fc2.n3766 a_400_38200# 0.26fF
C6465 fc2.t648 a_400_38200# 0.00fF
C6466 fc2.n3767 a_400_38200# 0.34fF
C6467 fc2.t493 a_400_38200# -0.00fF
C6468 fc2.n3768 a_400_38200# 0.34fF
C6469 fc2.n3769 a_400_38200# 0.27fF
C6470 fc2.n3770 a_400_38200# 0.21fF
C6471 fc2.n3771 a_400_38200# 0.08fF
C6472 fc2.n3772 a_400_38200# 1.20fF
C6473 fc2.n3773 a_400_38200# 0.30fF
C6474 fc2.n3774 a_400_38200# 3.90fF
C6475 fc2.n3775 a_400_38200# 0.24fF
C6476 fc2.n3776 a_400_38200# 0.13fF
C6477 fc2.n3777 a_400_38200# 1.92fF
C6478 fc2.n3778 a_400_38200# 3.43fF
C6479 fc2.n3779 a_400_38200# 21.84fF
C6480 fc2.n3780 a_400_38200# 0.41fF
C6481 fc2.n3781 a_400_38200# 13.20fF
C6482 fc2.n3782 a_400_38200# 0.10fF
C6483 fc2.n3783 a_400_38200# 0.25fF
C6484 fc2.n3784 a_400_38200# 0.24fF
C6485 fc2.n3785 a_400_38200# 2.12fF
C6486 fc2.t641 a_400_38200# -0.02fF
C6487 fc2.n3786 a_400_38200# 0.57fF
C6488 fc2.t541 a_400_38200# -0.02fF
C6489 fc2.n3787 a_400_38200# 0.21fF
C6490 fc2.t409 a_400_38200# -0.01fF
C6491 fc2.n3788 a_400_38200# 0.56fF
C6492 fc2.n3789 a_400_38200# 2.12fF
C6493 fc2.n3790 a_400_38200# 4.75fF
C6494 fc2.n3791 a_400_38200# 0.05fF
C6495 fc2.n3792 a_400_38200# 0.46fF
C6496 fc2.n3793 a_400_38200# 1.19fF
C6497 fc2.n3794 a_400_38200# 1.63fF
C6498 fc2.t726 a_400_38200# -0.02fF
C6499 fc2.n3795 a_400_38200# 0.21fF
C6500 fc2.t732 a_400_38200# -0.06fF
C6501 fc2.n3796 a_400_38200# 0.62fF
C6502 fc2.t399 a_400_38200# -0.02fF
C6503 fc2.n3798 a_400_38200# 0.21fF
C6504 fc2.t728 a_400_38200# -0.06fF
C6505 fc2.n3799 a_400_38200# 0.62fF
C6506 fc2.n3801 a_400_38200# 0.05fF
C6507 fc2.n3802 a_400_38200# 0.46fF
C6508 fc2.n3803 a_400_38200# 1.20fF
C6509 fc2.n3804 a_400_38200# 1.75fF
C6510 fc2.n3805 a_400_38200# 1.98fF
C6511 fc2.n3806 a_400_38200# 1.72fF
C6512 fc2.n3807 a_400_38200# 1.61fF
C6513 fc2.t735 a_400_38200# -0.02fF
C6514 fc2.n3808 a_400_38200# 0.21fF
C6515 fc2.t684 a_400_38200# -0.06fF
C6516 fc2.n3809 a_400_38200# 0.62fF
C6517 fc2.t612 a_400_38200# -0.02fF
C6518 fc2.n3811 a_400_38200# 0.21fF
C6519 fc2.t530 a_400_38200# -0.06fF
C6520 fc2.n3812 a_400_38200# 0.62fF
C6521 fc2.n3814 a_400_38200# 2.59fF
C6522 fc2.n3815 a_400_38200# 1.87fF
C6523 fc2.n3816 a_400_38200# 2.30fF
C6524 fc2.n3817 a_400_38200# 1.61fF
C6525 fc2.t591 a_400_38200# -0.02fF
C6526 fc2.n3818 a_400_38200# 0.21fF
C6527 fc2.t614 a_400_38200# -0.06fF
C6528 fc2.n3819 a_400_38200# 0.62fF
C6529 fc2.t665 a_400_38200# -0.02fF
C6530 fc2.n3821 a_400_38200# 0.21fF
C6531 fc2.t408 a_400_38200# -0.06fF
C6532 fc2.n3822 a_400_38200# 0.62fF
C6533 fc2.n3824 a_400_38200# 2.39fF
C6534 fc2.n3825 a_400_38200# 1.87fF
C6535 fc2.n3826 a_400_38200# 2.30fF
C6536 fc2.n3827 a_400_38200# 1.61fF
C6537 fc2.t407 a_400_38200# -0.02fF
C6538 fc2.n3828 a_400_38200# 0.21fF
C6539 fc2.t645 a_400_38200# -0.06fF
C6540 fc2.n3829 a_400_38200# 0.62fF
C6541 fc2.t651 a_400_38200# -0.02fF
C6542 fc2.n3831 a_400_38200# 0.21fF
C6543 fc2.t650 a_400_38200# -0.06fF
C6544 fc2.n3832 a_400_38200# 0.62fF
C6545 fc2.n3834 a_400_38200# 2.49fF
C6546 fc2.n3835 a_400_38200# 1.87fF
C6547 fc2.n3836 a_400_38200# 1.97fF
C6548 fc2.n3837 a_400_38200# 1.20fF
C6549 fc2.n3838 a_400_38200# 0.03fF
C6550 fc2.n3839 a_400_38200# 0.04fF
C6551 fc2.n3840 a_400_38200# 0.24fF
C6552 fc2.n3841 a_400_38200# 1.41fF
C6553 fc2.n3842 a_400_38200# 0.68fF
C6554 fc2.n3843 a_400_38200# 0.25fF
C6555 fc2.n3844 a_400_38200# 0.08fF
C6556 fc2.n3845 a_400_38200# 0.10fF
C6557 fc2.n3846 a_400_38200# 0.11fF
C6558 fc2.t577 a_400_38200# -0.06fF
C6559 fc2.n3847 a_400_38200# 0.26fF
C6560 fc2.t709 a_400_38200# 0.00fF
C6561 fc2.n3848 a_400_38200# 0.34fF
C6562 fc2.t395 a_400_38200# -0.00fF
C6563 fc2.n3849 a_400_38200# 0.34fF
C6564 fc2.n3850 a_400_38200# 0.03fF
C6565 fc2.n3851 a_400_38200# 0.04fF
C6566 fc2.n3852 a_400_38200# 0.24fF
C6567 fc2.n3853 a_400_38200# 1.41fF
C6568 fc2.n3854 a_400_38200# 0.68fF
C6569 fc2.n3855 a_400_38200# 0.25fF
C6570 fc2.n3856 a_400_38200# 0.08fF
C6571 fc2.n3857 a_400_38200# 0.11fF
C6572 fc2.n3858 a_400_38200# 0.84fF
C6573 fc2.n3859 a_400_38200# 1.92fF
C6574 fc2.n3860 a_400_38200# 1.61fF
C6575 fc2.n3861 a_400_38200# 21.40fF
C6576 fc2.n3862 a_400_38200# 14.33fF
C6577 fc2.n3863 a_400_38200# 0.41fF
C6578 fc2.n3864 a_400_38200# 13.20fF
C6579 fc2.n3865 a_400_38200# 0.10fF
C6580 fc2.n3866 a_400_38200# 0.25fF
C6581 fc2.n3867 a_400_38200# 0.24fF
C6582 fc2.n3868 a_400_38200# 2.12fF
C6583 fc2.t427 a_400_38200# -0.02fF
C6584 fc2.n3869 a_400_38200# 0.57fF
C6585 fc2.t393 a_400_38200# -0.02fF
C6586 fc2.n3870 a_400_38200# 0.21fF
C6587 fc2.t536 a_400_38200# -0.01fF
C6588 fc2.n3871 a_400_38200# 0.56fF
C6589 fc2.n3872 a_400_38200# 2.12fF
C6590 fc2.n3873 a_400_38200# 4.75fF
C6591 fc2.n3874 a_400_38200# 0.05fF
C6592 fc2.n3875 a_400_38200# 0.46fF
C6593 fc2.n3876 a_400_38200# 1.19fF
C6594 fc2.n3877 a_400_38200# 1.63fF
C6595 fc2.t513 a_400_38200# -0.02fF
C6596 fc2.n3878 a_400_38200# 0.21fF
C6597 fc2.t475 a_400_38200# -0.06fF
C6598 fc2.n3879 a_400_38200# 0.62fF
C6599 fc2.t441 a_400_38200# -0.02fF
C6600 fc2.n3881 a_400_38200# 0.21fF
C6601 fc2.t465 a_400_38200# -0.06fF
C6602 fc2.n3882 a_400_38200# 0.62fF
C6603 fc2.n3884 a_400_38200# 0.05fF
C6604 fc2.n3885 a_400_38200# 0.46fF
C6605 fc2.n3886 a_400_38200# 1.20fF
C6606 fc2.n3887 a_400_38200# 1.75fF
C6607 fc2.n3888 a_400_38200# 1.98fF
C6608 fc2.n3889 a_400_38200# 1.72fF
C6609 fc2.n3890 a_400_38200# 1.61fF
C6610 fc2.t569 a_400_38200# -0.02fF
C6611 fc2.n3891 a_400_38200# 0.21fF
C6612 fc2.t546 a_400_38200# -0.06fF
C6613 fc2.n3892 a_400_38200# 0.62fF
C6614 fc2.t592 a_400_38200# -0.02fF
C6615 fc2.n3894 a_400_38200# 0.21fF
C6616 fc2.t535 a_400_38200# -0.06fF
C6617 fc2.n3895 a_400_38200# 0.62fF
C6618 fc2.n3897 a_400_38200# 2.59fF
C6619 fc2.n3898 a_400_38200# 1.87fF
C6620 fc2.n3899 a_400_38200# 2.30fF
C6621 fc2.n3900 a_400_38200# 1.61fF
C6622 fc2.t484 a_400_38200# -0.02fF
C6623 fc2.n3901 a_400_38200# 0.21fF
C6624 fc2.t658 a_400_38200# -0.06fF
C6625 fc2.n3902 a_400_38200# 0.62fF
C6626 fc2.t534 a_400_38200# -0.02fF
C6627 fc2.n3904 a_400_38200# 0.21fF
C6628 fc2.t711 a_400_38200# -0.06fF
C6629 fc2.n3905 a_400_38200# 0.62fF
C6630 fc2.n3907 a_400_38200# 2.39fF
C6631 fc2.n3908 a_400_38200# 1.87fF
C6632 fc2.n3909 a_400_38200# 2.30fF
C6633 fc2.n3910 a_400_38200# 1.61fF
C6634 fc2.t505 a_400_38200# -0.02fF
C6635 fc2.n3911 a_400_38200# 0.21fF
C6636 fc2.t608 a_400_38200# -0.06fF
C6637 fc2.n3912 a_400_38200# 0.62fF
C6638 fc2.t448 a_400_38200# -0.02fF
C6639 fc2.n3914 a_400_38200# 0.21fF
C6640 fc2.t533 a_400_38200# -0.06fF
C6641 fc2.n3915 a_400_38200# 0.62fF
C6642 fc2.n3917 a_400_38200# 2.39fF
C6643 fc2.n3918 a_400_38200# 1.87fF
C6644 fc2.n3919 a_400_38200# 2.30fF
C6645 fc2.n3920 a_400_38200# 1.61fF
C6646 fc2.t710 a_400_38200# -0.02fF
C6647 fc2.n3921 a_400_38200# 0.21fF
C6648 fc2.t392 a_400_38200# -0.06fF
C6649 fc2.n3922 a_400_38200# 0.62fF
C6650 fc2.t674 a_400_38200# -0.02fF
C6651 fc2.n3924 a_400_38200# 0.21fF
C6652 fc2.t697 a_400_38200# -0.06fF
C6653 fc2.n3925 a_400_38200# 0.62fF
C6654 fc2.n3927 a_400_38200# 2.39fF
C6655 fc2.n3928 a_400_38200# 1.87fF
C6656 fc2.n3929 a_400_38200# 2.30fF
C6657 fc2.n3930 a_400_38200# 1.61fF
C6658 fc2.t519 a_400_38200# -0.02fF
C6659 fc2.n3931 a_400_38200# 0.21fF
C6660 fc2.t754 a_400_38200# -0.06fF
C6661 fc2.n3932 a_400_38200# 0.62fF
C6662 fc2.t420 a_400_38200# -0.02fF
C6663 fc2.n3934 a_400_38200# 0.21fF
C6664 fc2.t494 a_400_38200# -0.06fF
C6665 fc2.n3935 a_400_38200# 0.62fF
C6666 fc2.n3937 a_400_38200# 2.39fF
C6667 fc2.n3938 a_400_38200# 1.87fF
C6668 fc2.n3939 a_400_38200# 2.30fF
C6669 fc2.n3940 a_400_38200# 1.61fF
C6670 fc2.t696 a_400_38200# -0.02fF
C6671 fc2.n3941 a_400_38200# 0.21fF
C6672 fc2.t560 a_400_38200# -0.06fF
C6673 fc2.n3942 a_400_38200# 0.62fF
C6674 fc2.t516 a_400_38200# -0.02fF
C6675 fc2.n3944 a_400_38200# 0.21fF
C6676 fc2.t753 a_400_38200# -0.06fF
C6677 fc2.n3945 a_400_38200# 0.62fF
C6678 fc2.n3947 a_400_38200# 2.39fF
C6679 fc2.n3948 a_400_38200# 1.87fF
C6680 fc2.n3949 a_400_38200# 2.30fF
C6681 fc2.n3950 a_400_38200# 1.61fF
C6682 fc2.t670 a_400_38200# -0.02fF
C6683 fc2.n3951 a_400_38200# 0.21fF
C6684 fc2.t669 a_400_38200# -0.06fF
C6685 fc2.n3952 a_400_38200# 0.62fF
C6686 fc2.t594 a_400_38200# -0.02fF
C6687 fc2.n3954 a_400_38200# 0.21fF
C6688 fc2.t576 a_400_38200# -0.06fF
C6689 fc2.n3955 a_400_38200# 0.62fF
C6690 fc2.n3957 a_400_38200# 2.49fF
C6691 fc2.n3958 a_400_38200# 1.87fF
C6692 fc2.n3959 a_400_38200# 1.97fF
C6693 fc2.n3960 a_400_38200# 1.20fF
C6694 fc2.n3961 a_400_38200# 0.03fF
C6695 fc2.n3962 a_400_38200# 0.04fF
C6696 fc2.n3963 a_400_38200# 0.24fF
C6697 fc2.n3964 a_400_38200# 1.41fF
C6698 fc2.n3965 a_400_38200# 0.68fF
C6699 fc2.n3966 a_400_38200# 0.25fF
C6700 fc2.n3967 a_400_38200# 0.08fF
C6701 fc2.n3968 a_400_38200# 0.10fF
C6702 fc2.n3969 a_400_38200# 0.11fF
C6703 fc2.t738 a_400_38200# -0.06fF
C6704 fc2.n3970 a_400_38200# 0.26fF
C6705 fc2.t525 a_400_38200# 0.00fF
C6706 fc2.n3971 a_400_38200# 0.34fF
C6707 fc2.t679 a_400_38200# -0.00fF
C6708 fc2.n3972 a_400_38200# 0.34fF
C6709 fc2.n3973 a_400_38200# 0.03fF
C6710 fc2.n3974 a_400_38200# 0.04fF
C6711 fc2.n3975 a_400_38200# 0.24fF
C6712 fc2.n3976 a_400_38200# 1.41fF
C6713 fc2.n3977 a_400_38200# 0.68fF
C6714 fc2.n3978 a_400_38200# 0.25fF
C6715 fc2.n3979 a_400_38200# 0.08fF
C6716 fc2.n3980 a_400_38200# 0.11fF
C6717 fc2.n3981 a_400_38200# 0.84fF
C6718 fc2.n3982 a_400_38200# 1.92fF
C6719 fc2.n3983 a_400_38200# 1.61fF
C6720 fc2.n3984 a_400_38200# 21.40fF
C6721 fc2.n3985 a_400_38200# 14.33fF
C6722 fc2.n3986 a_400_38200# 0.41fF
C6723 fc2.n3987 a_400_38200# 10.72fF
C6724 fc2.n3988 a_400_38200# 11.73fF
C6725 fc2.n3989 a_400_38200# 0.14fF
C6726 fc2.n3990 a_400_38200# 0.95fF
C6727 fc2.n3991 a_400_38200# 58.52fF
C6728 VP.n0 a_400_38200# 2.73fF
C6729 VP.n1 a_400_38200# 0.35fF
C6730 VP.n2 a_400_38200# 0.97fF
C6731 VP.n3 a_400_38200# 1.07fF
C6732 VP.n4 a_400_38200# 1.05fF
C6733 VP.n5 a_400_38200# 0.09fF
C6734 VP.n6 a_400_38200# 0.27fF
C6735 VP.n7 a_400_38200# 1.03fF
C6736 VP.n8 a_400_38200# 0.15fF
C6737 VP.n9 a_400_38200# 0.90fF
C6738 VP.n10 a_400_38200# 0.08fF
C6739 VP.n11 a_400_38200# 0.27fF
C6740 VP.n12 a_400_38200# 1.01fF
C6741 VP.n13 a_400_38200# 1.63fF
C6742 VP.n14 a_400_38200# 0.97fF
C6743 VP.n15 a_400_38200# 0.01fF
C6744 VP.n16 a_400_38200# 0.16fF
C6745 VP.n17 a_400_38200# 1.00fF
C6746 VP.n18 a_400_38200# 1.01fF
C6747 VP.n19 a_400_38200# 2.15fF
C6748 VP.n20 a_400_38200# 0.09fF
C6749 VP.n21 a_400_38200# 0.27fF
C6750 VP.n22 a_400_38200# 0.97fF
C6751 VP.n23 a_400_38200# 0.16fF
C6752 VP.n24 a_400_38200# 1.00fF
C6753 VP.n25 a_400_38200# 0.12fF
C6754 VP.n26 a_400_38200# 1.47fF
C6755 VP.n27 a_400_38200# 0.27fF
C6756 VP.n28 a_400_38200# 1.01fF
C6757 VP.n29 a_400_38200# 2.15fF
C6758 VP.n30 a_400_38200# 0.09fF
C6759 VP.n31 a_400_38200# 0.27fF
C6760 VP.n32 a_400_38200# 0.97fF
C6761 VP.n33 a_400_38200# 0.16fF
C6762 VP.n34 a_400_38200# 1.00fF
C6763 VP.n35 a_400_38200# 0.12fF
C6764 VP.n36 a_400_38200# 1.47fF
C6765 VP.n37 a_400_38200# 0.27fF
C6766 VP.n38 a_400_38200# 1.01fF
C6767 VP.n39 a_400_38200# 1.65fF
C6768 VP.n40 a_400_38200# 0.09fF
C6769 VP.n41 a_400_38200# 0.27fF
C6770 VP.n42 a_400_38200# 0.97fF
C6771 VP.n43 a_400_38200# 0.16fF
C6772 VP.n44 a_400_38200# 1.00fF
C6773 VP.n45 a_400_38200# 0.08fF
C6774 VP.n46 a_400_38200# 0.27fF
C6775 VP.n47 a_400_38200# 0.97fF
C6776 VP.n48 a_400_38200# 0.01fF
C6777 VP.n49 a_400_38200# 0.16fF
C6778 VP.n50 a_400_38200# 1.00fF
C6779 VP.n51 a_400_38200# 0.09fF
C6780 VP.n52 a_400_38200# 0.27fF
C6781 VP.n53 a_400_38200# 0.97fF
C6782 VP.n54 a_400_38200# 0.16fF
C6783 VP.n55 a_400_38200# 1.00fF
C6784 VP.n56 a_400_38200# 0.08fF
C6785 VP.n57 a_400_38200# 0.27fF
C6786 VP.n58 a_400_38200# 1.01fF
C6787 VP.n59 a_400_38200# 1.65fF
C6788 VP.n60 a_400_38200# 0.97fF
C6789 VP.n61 a_400_38200# 0.01fF
C6790 VP.n62 a_400_38200# 0.16fF
C6791 VP.n63 a_400_38200# 1.00fF
C6792 VP.n64 a_400_38200# 1.01fF
C6793 VP.n65 a_400_38200# 1.65fF
C6794 VP.n66 a_400_38200# 0.09fF
C6795 VP.n67 a_400_38200# 0.27fF
C6796 VP.n68 a_400_38200# 0.97fF
C6797 VP.n69 a_400_38200# 0.16fF
C6798 VP.n70 a_400_38200# 1.00fF
C6799 VP.n71 a_400_38200# 0.08fF
C6800 VP.n72 a_400_38200# 0.27fF
C6801 VP.n73 a_400_38200# 0.97fF
C6802 VP.n74 a_400_38200# 0.01fF
C6803 VP.n75 a_400_38200# 0.16fF
C6804 VP.n76 a_400_38200# 1.00fF
C6805 VP.n77 a_400_38200# 0.09fF
C6806 VP.n78 a_400_38200# 0.27fF
C6807 VP.n79 a_400_38200# 0.97fF
C6808 VP.n80 a_400_38200# 0.16fF
C6809 VP.n81 a_400_38200# 1.00fF
C6810 VP.n82 a_400_38200# 0.08fF
C6811 VP.n83 a_400_38200# 0.27fF
C6812 VP.n84 a_400_38200# 1.01fF
C6813 VP.n85 a_400_38200# 1.65fF
C6814 VP.n86 a_400_38200# 0.97fF
C6815 VP.n87 a_400_38200# 0.01fF
C6816 VP.n88 a_400_38200# 0.16fF
C6817 VP.n89 a_400_38200# 1.00fF
C6818 VP.n90 a_400_38200# 1.01fF
C6819 VP.n91 a_400_38200# 1.65fF
C6820 VP.n92 a_400_38200# 0.09fF
C6821 VP.n93 a_400_38200# 0.27fF
C6822 VP.n94 a_400_38200# 0.97fF
C6823 VP.n95 a_400_38200# 0.16fF
C6824 VP.n96 a_400_38200# 1.00fF
C6825 VP.n97 a_400_38200# 0.08fF
C6826 VP.n98 a_400_38200# 0.27fF
C6827 VP.n99 a_400_38200# 0.97fF
C6828 VP.n100 a_400_38200# 0.01fF
C6829 VP.n101 a_400_38200# 0.16fF
C6830 VP.n102 a_400_38200# 1.00fF
C6831 VP.n103 a_400_38200# 0.09fF
C6832 VP.n104 a_400_38200# 0.27fF
C6833 VP.n105 a_400_38200# 0.97fF
C6834 VP.n106 a_400_38200# 0.16fF
C6835 VP.n107 a_400_38200# 1.00fF
C6836 VP.n108 a_400_38200# 0.08fF
C6837 VP.n109 a_400_38200# 0.27fF
C6838 VP.n110 a_400_38200# 1.01fF
C6839 VP.n111 a_400_38200# 1.65fF
C6840 VP.n112 a_400_38200# 0.97fF
C6841 VP.n113 a_400_38200# 0.01fF
C6842 VP.n114 a_400_38200# 0.16fF
C6843 VP.n115 a_400_38200# 1.00fF
C6844 VP.n116 a_400_38200# 0.09fF
C6845 VP.n117 a_400_38200# 0.27fF
C6846 VP.n118 a_400_38200# 0.97fF
C6847 VP.n119 a_400_38200# 0.16fF
C6848 VP.n120 a_400_38200# 1.00fF
C6849 VP.n121 a_400_38200# 0.08fF
C6850 VP.n122 a_400_38200# 0.27fF
C6851 VP.n123 a_400_38200# 1.01fF
C6852 VP.n124 a_400_38200# 1.65fF
C6853 VP.n125 a_400_38200# 0.97fF
C6854 VP.n126 a_400_38200# 0.01fF
C6855 VP.n127 a_400_38200# 0.16fF
C6856 VP.n128 a_400_38200# 1.00fF
C6857 VP.t833 a_400_38200# 0.02fF
C6858 VP.n129 a_400_38200# 0.44fF
C6859 VP.n130 a_400_38200# 0.99fF
C6860 VP.n131 a_400_38200# 2.15fF
C6861 VP.n132 a_400_38200# 0.35fF
C6862 VP.n133 a_400_38200# 0.97fF
C6863 VP.n134 a_400_38200# 0.30fF
C6864 VP.n135 a_400_38200# 1.06fF
C6865 VP.n136 a_400_38200# 0.12fF
C6866 VP.n137 a_400_38200# 1.47fF
C6867 VP.n138 a_400_38200# 0.27fF
C6868 VP.t564 a_400_38200# 0.02fF
C6869 VP.n139 a_400_38200# 0.89fF
C6870 VP.t604 a_400_38200# 0.02fF
C6871 VP.n140 a_400_38200# 0.89fF
C6872 VP.t275 a_400_38200# 0.02fF
C6873 VP.n141 a_400_38200# 0.02fF
C6874 VP.n142 a_400_38200# 0.37fF
C6875 VP.n143 a_400_38200# 0.10fF
C6876 VP.n144 a_400_38200# 1.30fF
C6877 VP.n145 a_400_38200# 0.33fF
C6878 VP.t818 a_400_38200# 0.02fF
C6879 VP.n146 a_400_38200# 0.89fF
C6880 VP.t138 a_400_38200# 0.02fF
C6881 VP.n147 a_400_38200# 0.89fF
C6882 VP.n148 a_400_38200# 0.03fF
C6883 VP.n149 a_400_38200# 0.03fF
C6884 VP.n150 a_400_38200# 0.04fF
C6885 VP.n151 a_400_38200# 0.47fF
C6886 VP.n152 a_400_38200# 0.11fF
C6887 VP.n153 a_400_38200# 0.11fF
C6888 VP.n154 a_400_38200# 0.05fF
C6889 VP.n155 a_400_38200# 0.08fF
C6890 VP.n156 a_400_38200# 0.10fF
C6891 VP.n157 a_400_38200# 0.09fF
C6892 VP.n158 a_400_38200# 0.28fF
C6893 VP.n159 a_400_38200# 1.28fF
C6894 VP.n161 a_400_38200# 1.45fF
C6895 VP.n162 a_400_38200# 0.39fF
C6896 VP.n163 a_400_38200# 1.76fF
C6897 VP.n164 a_400_38200# 0.52fF
C6898 VP.n165 a_400_38200# 2.08fF
C6899 VP.n166 a_400_38200# 1.76fF
C6900 VP.n167 a_400_38200# 0.52fF
C6901 VP.n168 a_400_38200# 2.08fF
C6902 VP.n169 a_400_38200# 1.76fF
C6903 VP.n170 a_400_38200# 0.52fF
C6904 VP.n171 a_400_38200# 2.08fF
C6905 VP.n172 a_400_38200# 1.76fF
C6906 VP.n173 a_400_38200# 0.52fF
C6907 VP.n174 a_400_38200# 2.08fF
C6908 VP.n175 a_400_38200# 1.76fF
C6909 VP.n176 a_400_38200# 0.52fF
C6910 VP.n177 a_400_38200# 2.08fF
C6911 VP.n178 a_400_38200# 1.76fF
C6912 VP.n179 a_400_38200# 0.52fF
C6913 VP.n180 a_400_38200# 2.08fF
C6914 VP.n181 a_400_38200# 1.76fF
C6915 VP.n182 a_400_38200# 0.52fF
C6916 VP.n183 a_400_38200# 2.08fF
C6917 VP.n184 a_400_38200# 1.76fF
C6918 VP.n185 a_400_38200# 0.52fF
C6919 VP.n186 a_400_38200# 2.08fF
C6920 VP.n187 a_400_38200# 1.76fF
C6921 VP.n188 a_400_38200# 0.52fF
C6922 VP.n189 a_400_38200# 2.08fF
C6923 VP.n190 a_400_38200# 1.76fF
C6924 VP.n191 a_400_38200# 0.52fF
C6925 VP.n192 a_400_38200# 2.08fF
C6926 VP.n193 a_400_38200# 1.79fF
C6927 VP.n194 a_400_38200# 0.52fF
C6928 VP.n195 a_400_38200# 2.28fF
C6929 VP.n196 a_400_38200# 71.87fF
C6930 VP.n197 a_400_38200# 1.05fF
C6931 VP.n198 a_400_38200# 3.98fF
C6932 VP.n199 a_400_38200# 1.48fF
C6933 VP.t529 a_400_38200# 0.02fF
C6934 VP.n200 a_400_38200# 0.02fF
C6935 VP.n201 a_400_38200# 0.37fF
C6936 VP.n202 a_400_38200# 15.28fF
C6937 VP.t418 a_400_38200# 0.02fF
C6938 VP.n203 a_400_38200# 0.89fF
C6939 VP.t70 a_400_38200# 0.02fF
C6940 VP.n204 a_400_38200# 0.02fF
C6941 VP.n205 a_400_38200# 0.37fF
C6942 VP.t382 a_400_38200# 0.02fF
C6943 VP.n206 a_400_38200# 0.89fF
C6944 VP.t1273 a_400_38200# 0.02fF
C6945 VP.n207 a_400_38200# 0.89fF
C6946 VP.t952 a_400_38200# 0.02fF
C6947 VP.n208 a_400_38200# 0.02fF
C6948 VP.n209 a_400_38200# 0.37fF
C6949 VP.t1238 a_400_38200# 0.02fF
C6950 VP.n210 a_400_38200# 0.89fF
C6951 VP.t827 a_400_38200# 0.02fF
C6952 VP.n211 a_400_38200# 0.89fF
C6953 VP.t1201 a_400_38200# 0.02fF
C6954 VP.n212 a_400_38200# 0.02fF
C6955 VP.n213 a_400_38200# 0.37fF
C6956 VP.t179 a_400_38200# 0.02fF
C6957 VP.n214 a_400_38200# 0.89fF
C6958 VP.t1127 a_400_38200# 0.02fF
C6959 VP.n215 a_400_38200# 0.89fF
C6960 VP.t753 a_400_38200# 0.02fF
C6961 VP.n216 a_400_38200# 0.02fF
C6962 VP.n217 a_400_38200# 0.37fF
C6963 VP.t1031 a_400_38200# 0.02fF
C6964 VP.n218 a_400_38200# 0.89fF
C6965 VP.t679 a_400_38200# 0.02fF
C6966 VP.n219 a_400_38200# 0.89fF
C6967 VP.t298 a_400_38200# 0.02fF
C6968 VP.n220 a_400_38200# 0.02fF
C6969 VP.n221 a_400_38200# 0.37fF
C6970 VP.t583 a_400_38200# 0.02fF
C6971 VP.n222 a_400_38200# 0.89fF
C6972 VP.t235 a_400_38200# 0.02fF
C6973 VP.n223 a_400_38200# 0.89fF
C6974 VP.t1146 a_400_38200# 0.02fF
C6975 VP.n224 a_400_38200# 0.02fF
C6976 VP.n225 a_400_38200# 0.37fF
C6977 VP.t117 a_400_38200# 0.02fF
C6978 VP.n226 a_400_38200# 0.89fF
C6979 VP.t1090 a_400_38200# 0.02fF
C6980 VP.n227 a_400_38200# 0.89fF
C6981 VP.t699 a_400_38200# 0.02fF
C6982 VP.n228 a_400_38200# 0.02fF
C6983 VP.n229 a_400_38200# 0.37fF
C6984 VP.t988 a_400_38200# 0.02fF
C6985 VP.n230 a_400_38200# 0.89fF
C6986 VP.t648 a_400_38200# 0.02fF
C6987 VP.n231 a_400_38200# 0.89fF
C6988 VP.t254 a_400_38200# 0.02fF
C6989 VP.n232 a_400_38200# 0.02fF
C6990 VP.n233 a_400_38200# 0.37fF
C6991 VP.t542 a_400_38200# 0.02fF
C6992 VP.n234 a_400_38200# 0.89fF
C6993 VP.t202 a_400_38200# 0.02fF
C6994 VP.n235 a_400_38200# 0.89fF
C6995 VP.t1108 a_400_38200# 0.02fF
C6996 VP.n236 a_400_38200# 0.02fF
C6997 VP.n237 a_400_38200# 0.37fF
C6998 VP.t149 a_400_38200# 0.02fF
C6999 VP.n238 a_400_38200# 0.89fF
C7000 VP.t1053 a_400_38200# 0.02fF
C7001 VP.n239 a_400_38200# 0.89fF
C7002 VP.t723 a_400_38200# 0.02fF
C7003 VP.n240 a_400_38200# 0.02fF
C7004 VP.n241 a_400_38200# 0.37fF
C7005 VP.t1007 a_400_38200# 0.02fF
C7006 VP.n242 a_400_38200# 0.89fF
C7007 VP.t116 a_400_38200# 113.64fF
C7008 VP.t546 a_400_38200# 0.02fF
C7009 VP.n243 a_400_38200# 1.30fF
C7010 VP.n244 a_400_38200# 0.25fF
C7011 VP.n245 a_400_38200# 0.35fF
C7012 VP.n246 a_400_38200# 0.97fF
C7013 VP.n247 a_400_38200# 0.32fF
C7014 VP.n248 a_400_38200# 1.07fF
C7015 VP.n249 a_400_38200# 5.03fF
C7016 VP.n250 a_400_38200# 0.10fF
C7017 VP.n251 a_400_38200# 0.17fF
C7018 VP.n252 a_400_38200# 0.10fF
C7019 VP.n253 a_400_38200# 0.13fF
C7020 VP.n254 a_400_38200# 0.37fF
C7021 VP.n255 a_400_38200# 0.08fF
C7022 VP.n256 a_400_38200# 0.09fF
C7023 VP.n257 a_400_38200# 0.20fF
C7024 VP.n258 a_400_38200# 0.01fF
C7025 VP.n259 a_400_38200# 0.21fF
C7026 VP.n260 a_400_38200# 0.24fF
C7027 VP.n261 a_400_38200# 0.04fF
C7028 VP.n262 a_400_38200# 0.02fF
C7029 VP.n263 a_400_38200# 0.06fF
C7030 VP.n264 a_400_38200# 0.69fF
C7031 VP.n265 a_400_38200# 0.10fF
C7032 VP.n266 a_400_38200# 0.12fF
C7033 VP.t992 a_400_38200# 0.02fF
C7034 VP.n267 a_400_38200# 0.14fF
C7035 VP.n269 a_400_38200# 1.92fF
C7036 VP.t321 a_400_38200# 0.02fF
C7037 VP.n270 a_400_38200# 0.24fF
C7038 VP.n271 a_400_38200# 0.35fF
C7039 VP.n272 a_400_38200# 0.60fF
C7040 VP.n273 a_400_38200# 0.12fF
C7041 VP.t1175 a_400_38200# 0.02fF
C7042 VP.n274 a_400_38200# 0.14fF
C7043 VP.n276 a_400_38200# 0.04fF
C7044 VP.n277 a_400_38200# 0.02fF
C7045 VP.n278 a_400_38200# 0.06fF
C7046 VP.n279 a_400_38200# 0.30fF
C7047 VP.n280 a_400_38200# 0.10fF
C7048 VP.n281 a_400_38200# 0.28fF
C7049 VP.n282 a_400_38200# 0.15fF
C7050 VP.n283 a_400_38200# 0.08fF
C7051 VP.n284 a_400_38200# 0.14fF
C7052 VP.n285 a_400_38200# 1.39fF
C7053 VP.n286 a_400_38200# 0.34fF
C7054 VP.n287 a_400_38200# 2.18fF
C7055 VP.t1338 a_400_38200# 0.02fF
C7056 VP.n288 a_400_38200# 0.24fF
C7057 VP.n289 a_400_38200# 0.91fF
C7058 VP.n290 a_400_38200# 0.05fF
C7059 VP.t281 a_400_38200# 0.02fF
C7060 VP.n291 a_400_38200# 0.12fF
C7061 VP.n292 a_400_38200# 0.14fF
C7062 VP.n294 a_400_38200# 1.84fF
C7063 VP.n295 a_400_38200# 0.12fF
C7064 VP.t724 a_400_38200# 0.02fF
C7065 VP.n296 a_400_38200# 0.14fF
C7066 VP.t1163 a_400_38200# 0.02fF
C7067 VP.n298 a_400_38200# 0.24fF
C7068 VP.n299 a_400_38200# 0.35fF
C7069 VP.n300 a_400_38200# 0.60fF
C7070 VP.n301 a_400_38200# 0.17fF
C7071 VP.n302 a_400_38200# 1.38fF
C7072 VP.n303 a_400_38200# 0.36fF
C7073 VP.n304 a_400_38200# 0.12fF
C7074 VP.n305 a_400_38200# 0.03fF
C7075 VP.n306 a_400_38200# 0.02fF
C7076 VP.n307 a_400_38200# 0.04fF
C7077 VP.n308 a_400_38200# 0.02fF
C7078 VP.n309 a_400_38200# 0.09fF
C7079 VP.n310 a_400_38200# 0.03fF
C7080 VP.n311 a_400_38200# 0.12fF
C7081 VP.n312 a_400_38200# 0.09fF
C7082 VP.n313 a_400_38200# 2.30fF
C7083 VP.t888 a_400_38200# 0.02fF
C7084 VP.n314 a_400_38200# 0.24fF
C7085 VP.n315 a_400_38200# 0.91fF
C7086 VP.n316 a_400_38200# 0.05fF
C7087 VP.t1135 a_400_38200# 0.02fF
C7088 VP.n317 a_400_38200# 0.12fF
C7089 VP.n318 a_400_38200# 0.14fF
C7090 VP.n320 a_400_38200# 0.84fF
C7091 VP.n321 a_400_38200# 0.13fF
C7092 VP.n322 a_400_38200# 16.85fF
C7093 VP.n323 a_400_38200# 3.35fF
C7094 VP.n325 a_400_38200# 20.92fF
C7095 VP.n327 a_400_38200# 2.44fF
C7096 VP.n328 a_400_38200# 1.35fF
C7097 VP.n329 a_400_38200# 0.48fF
C7098 VP.n330 a_400_38200# 0.88fF
C7099 VP.n331 a_400_38200# 0.60fF
C7100 VP.n332 a_400_38200# 2.33fF
C7101 VP.n333 a_400_38200# 0.84fF
C7102 VP.n334 a_400_38200# 0.02fF
C7103 VP.n335 a_400_38200# 0.76fF
C7104 VP.n336 a_400_38200# 0.96fF
C7105 VP.t69 a_400_38200# 15.72fF
C7106 VP.n337 a_400_38200# 15.42fF
C7107 VP.n339 a_400_38200# 0.38fF
C7108 VP.n340 a_400_38200# 3.60fF
C7109 VP.n341 a_400_38200# 1.80fF
C7110 VP.t94 a_400_38200# 0.02fF
C7111 VP.n342 a_400_38200# 0.64fF
C7112 VP.n343 a_400_38200# 0.60fF
C7113 VP.n344 a_400_38200# 2.20fF
C7114 VP.n345 a_400_38200# 4.74fF
C7115 VP.t1130 a_400_38200# 0.02fF
C7116 VP.n346 a_400_38200# 1.19fF
C7117 VP.n347 a_400_38200# 0.05fF
C7118 VP.t58 a_400_38200# 0.02fF
C7119 VP.n348 a_400_38200# 0.01fF
C7120 VP.n349 a_400_38200# 0.26fF
C7121 VP.n351 a_400_38200# 15.28fF
C7122 VP.n352 a_400_38200# 0.10fF
C7123 VP.n353 a_400_38200# 0.17fF
C7124 VP.n354 a_400_38200# 0.10fF
C7125 VP.n355 a_400_38200# 0.13fF
C7126 VP.n356 a_400_38200# 0.37fF
C7127 VP.n357 a_400_38200# 0.08fF
C7128 VP.n358 a_400_38200# 0.09fF
C7129 VP.n359 a_400_38200# 0.20fF
C7130 VP.n360 a_400_38200# 0.01fF
C7131 VP.n361 a_400_38200# 0.21fF
C7132 VP.n362 a_400_38200# 0.24fF
C7133 VP.n363 a_400_38200# 0.04fF
C7134 VP.n364 a_400_38200# 0.02fF
C7135 VP.n365 a_400_38200# 0.06fF
C7136 VP.n366 a_400_38200# 0.69fF
C7137 VP.n367 a_400_38200# 0.10fF
C7138 VP.n368 a_400_38200# 1.92fF
C7139 VP.n369 a_400_38200# 0.12fF
C7140 VP.t545 a_400_38200# 0.02fF
C7141 VP.n370 a_400_38200# 0.14fF
C7142 VP.t982 a_400_38200# 0.02fF
C7143 VP.n372 a_400_38200# 0.24fF
C7144 VP.n373 a_400_38200# 0.35fF
C7145 VP.n374 a_400_38200# 0.60fF
C7146 VP.n375 a_400_38200# 0.27fF
C7147 VP.n376 a_400_38200# 0.03fF
C7148 VP.n377 a_400_38200# 0.05fF
C7149 VP.n378 a_400_38200# 0.06fF
C7150 VP.n379 a_400_38200# 0.15fF
C7151 VP.n380 a_400_38200# 0.12fF
C7152 VP.n381 a_400_38200# 0.04fF
C7153 VP.n382 a_400_38200# 0.03fF
C7154 VP.n383 a_400_38200# 0.07fF
C7155 VP.n384 a_400_38200# 0.09fF
C7156 VP.n385 a_400_38200# 0.24fF
C7157 VP.n386 a_400_38200# 0.03fF
C7158 VP.n387 a_400_38200# 0.05fF
C7159 VP.n388 a_400_38200# 0.05fF
C7160 VP.n389 a_400_38200# 0.04fF
C7161 VP.n390 a_400_38200# 0.66fF
C7162 VP.n391 a_400_38200# 0.97fF
C7163 VP.n392 a_400_38200# 1.90fF
C7164 VP.t959 a_400_38200# 0.02fF
C7165 VP.n393 a_400_38200# 0.12fF
C7166 VP.n394 a_400_38200# 0.14fF
C7167 VP.t694 a_400_38200# 0.02fF
C7168 VP.n396 a_400_38200# 0.24fF
C7169 VP.n397 a_400_38200# 0.91fF
C7170 VP.n398 a_400_38200# 0.05fF
C7171 VP.n399 a_400_38200# 0.10fF
C7172 VP.n400 a_400_38200# 0.17fF
C7173 VP.n401 a_400_38200# 0.10fF
C7174 VP.n402 a_400_38200# 0.13fF
C7175 VP.n403 a_400_38200# 0.37fF
C7176 VP.n404 a_400_38200# 0.08fF
C7177 VP.n405 a_400_38200# 0.09fF
C7178 VP.n406 a_400_38200# 0.20fF
C7179 VP.n407 a_400_38200# 0.01fF
C7180 VP.n408 a_400_38200# 0.21fF
C7181 VP.n409 a_400_38200# 0.24fF
C7182 VP.n410 a_400_38200# 0.04fF
C7183 VP.n411 a_400_38200# 0.02fF
C7184 VP.n412 a_400_38200# 0.06fF
C7185 VP.n413 a_400_38200# 0.69fF
C7186 VP.n414 a_400_38200# 0.10fF
C7187 VP.n415 a_400_38200# 1.92fF
C7188 VP.n416 a_400_38200# 0.12fF
C7189 VP.t68 a_400_38200# 0.02fF
C7190 VP.n417 a_400_38200# 0.14fF
C7191 VP.t534 a_400_38200# 0.02fF
C7192 VP.n419 a_400_38200# 0.24fF
C7193 VP.n420 a_400_38200# 0.35fF
C7194 VP.n421 a_400_38200# 0.60fF
C7195 VP.n422 a_400_38200# 0.27fF
C7196 VP.n423 a_400_38200# 0.03fF
C7197 VP.n424 a_400_38200# 0.05fF
C7198 VP.n425 a_400_38200# 0.06fF
C7199 VP.n426 a_400_38200# 0.15fF
C7200 VP.n427 a_400_38200# 0.12fF
C7201 VP.n428 a_400_38200# 0.04fF
C7202 VP.n429 a_400_38200# 0.03fF
C7203 VP.n430 a_400_38200# 0.07fF
C7204 VP.n431 a_400_38200# 0.09fF
C7205 VP.n432 a_400_38200# 0.24fF
C7206 VP.n433 a_400_38200# 0.03fF
C7207 VP.n434 a_400_38200# 0.05fF
C7208 VP.n435 a_400_38200# 0.05fF
C7209 VP.n436 a_400_38200# 0.04fF
C7210 VP.n437 a_400_38200# 0.66fF
C7211 VP.n438 a_400_38200# 0.97fF
C7212 VP.n439 a_400_38200# 1.90fF
C7213 VP.t512 a_400_38200# 0.02fF
C7214 VP.n440 a_400_38200# 0.12fF
C7215 VP.n441 a_400_38200# 0.14fF
C7216 VP.t249 a_400_38200# 0.02fF
C7217 VP.n443 a_400_38200# 0.24fF
C7218 VP.n444 a_400_38200# 0.91fF
C7219 VP.n445 a_400_38200# 0.05fF
C7220 VP.n446 a_400_38200# 0.10fF
C7221 VP.n447 a_400_38200# 0.17fF
C7222 VP.n448 a_400_38200# 0.10fF
C7223 VP.n449 a_400_38200# 0.13fF
C7224 VP.n450 a_400_38200# 0.37fF
C7225 VP.n451 a_400_38200# 0.08fF
C7226 VP.n452 a_400_38200# 0.09fF
C7227 VP.n453 a_400_38200# 0.20fF
C7228 VP.n454 a_400_38200# 0.01fF
C7229 VP.n455 a_400_38200# 0.21fF
C7230 VP.n456 a_400_38200# 0.24fF
C7231 VP.n457 a_400_38200# 0.04fF
C7232 VP.n458 a_400_38200# 0.02fF
C7233 VP.n459 a_400_38200# 0.06fF
C7234 VP.n460 a_400_38200# 0.69fF
C7235 VP.n461 a_400_38200# 0.10fF
C7236 VP.n462 a_400_38200# 1.92fF
C7237 VP.n463 a_400_38200# 0.12fF
C7238 VP.t410 a_400_38200# 0.02fF
C7239 VP.n464 a_400_38200# 0.14fF
C7240 VP.t792 a_400_38200# 0.02fF
C7241 VP.n466 a_400_38200# 0.24fF
C7242 VP.n467 a_400_38200# 0.35fF
C7243 VP.n468 a_400_38200# 0.60fF
C7244 VP.n469 a_400_38200# 0.27fF
C7245 VP.n470 a_400_38200# 0.03fF
C7246 VP.n471 a_400_38200# 0.05fF
C7247 VP.n472 a_400_38200# 0.06fF
C7248 VP.n473 a_400_38200# 0.15fF
C7249 VP.n474 a_400_38200# 0.12fF
C7250 VP.n475 a_400_38200# 0.04fF
C7251 VP.n476 a_400_38200# 0.03fF
C7252 VP.n477 a_400_38200# 0.07fF
C7253 VP.n478 a_400_38200# 0.09fF
C7254 VP.n479 a_400_38200# 0.24fF
C7255 VP.n480 a_400_38200# 0.03fF
C7256 VP.n481 a_400_38200# 0.05fF
C7257 VP.n482 a_400_38200# 0.05fF
C7258 VP.n483 a_400_38200# 0.04fF
C7259 VP.n484 a_400_38200# 0.66fF
C7260 VP.n485 a_400_38200# 0.97fF
C7261 VP.n486 a_400_38200# 1.90fF
C7262 VP.t761 a_400_38200# 0.02fF
C7263 VP.n487 a_400_38200# 0.12fF
C7264 VP.n488 a_400_38200# 0.14fF
C7265 VP.t506 a_400_38200# 0.02fF
C7266 VP.n490 a_400_38200# 0.24fF
C7267 VP.n491 a_400_38200# 0.91fF
C7268 VP.n492 a_400_38200# 0.05fF
C7269 VP.n493 a_400_38200# 0.10fF
C7270 VP.n494 a_400_38200# 0.17fF
C7271 VP.n495 a_400_38200# 0.10fF
C7272 VP.n496 a_400_38200# 0.13fF
C7273 VP.n497 a_400_38200# 0.37fF
C7274 VP.n498 a_400_38200# 0.08fF
C7275 VP.n499 a_400_38200# 0.09fF
C7276 VP.n500 a_400_38200# 0.20fF
C7277 VP.n501 a_400_38200# 0.01fF
C7278 VP.n502 a_400_38200# 0.21fF
C7279 VP.n503 a_400_38200# 0.24fF
C7280 VP.n504 a_400_38200# 0.04fF
C7281 VP.n505 a_400_38200# 0.02fF
C7282 VP.n506 a_400_38200# 0.06fF
C7283 VP.n507 a_400_38200# 0.69fF
C7284 VP.n508 a_400_38200# 0.10fF
C7285 VP.n509 a_400_38200# 1.92fF
C7286 VP.n510 a_400_38200# 0.12fF
C7287 VP.t1264 a_400_38200# 0.02fF
C7288 VP.n511 a_400_38200# 0.14fF
C7289 VP.t401 a_400_38200# 0.02fF
C7290 VP.n513 a_400_38200# 0.24fF
C7291 VP.n514 a_400_38200# 0.35fF
C7292 VP.n515 a_400_38200# 0.60fF
C7293 VP.n516 a_400_38200# 0.27fF
C7294 VP.n517 a_400_38200# 0.03fF
C7295 VP.n518 a_400_38200# 0.05fF
C7296 VP.n519 a_400_38200# 0.06fF
C7297 VP.n520 a_400_38200# 0.15fF
C7298 VP.n521 a_400_38200# 0.12fF
C7299 VP.n522 a_400_38200# 0.04fF
C7300 VP.n523 a_400_38200# 0.03fF
C7301 VP.n524 a_400_38200# 0.07fF
C7302 VP.n525 a_400_38200# 0.09fF
C7303 VP.n526 a_400_38200# 0.24fF
C7304 VP.n527 a_400_38200# 0.03fF
C7305 VP.n528 a_400_38200# 0.05fF
C7306 VP.n529 a_400_38200# 0.05fF
C7307 VP.n530 a_400_38200# 0.04fF
C7308 VP.n531 a_400_38200# 0.66fF
C7309 VP.n532 a_400_38200# 0.97fF
C7310 VP.n533 a_400_38200# 1.90fF
C7311 VP.t308 a_400_38200# 0.02fF
C7312 VP.n534 a_400_38200# 0.12fF
C7313 VP.n535 a_400_38200# 0.14fF
C7314 VP.t96 a_400_38200# 0.02fF
C7315 VP.n537 a_400_38200# 0.24fF
C7316 VP.n538 a_400_38200# 0.91fF
C7317 VP.n539 a_400_38200# 0.05fF
C7318 VP.n540 a_400_38200# 0.10fF
C7319 VP.n541 a_400_38200# 0.17fF
C7320 VP.n542 a_400_38200# 0.10fF
C7321 VP.n543 a_400_38200# 0.13fF
C7322 VP.n544 a_400_38200# 0.37fF
C7323 VP.n545 a_400_38200# 0.08fF
C7324 VP.n546 a_400_38200# 0.09fF
C7325 VP.n547 a_400_38200# 0.20fF
C7326 VP.n548 a_400_38200# 0.01fF
C7327 VP.n549 a_400_38200# 0.21fF
C7328 VP.n550 a_400_38200# 0.24fF
C7329 VP.n551 a_400_38200# 0.04fF
C7330 VP.n552 a_400_38200# 0.02fF
C7331 VP.n553 a_400_38200# 0.06fF
C7332 VP.n554 a_400_38200# 0.69fF
C7333 VP.n555 a_400_38200# 0.10fF
C7334 VP.n556 a_400_38200# 1.92fF
C7335 VP.n557 a_400_38200# 0.12fF
C7336 VP.t821 a_400_38200# 0.02fF
C7337 VP.n558 a_400_38200# 0.14fF
C7338 VP.t1258 a_400_38200# 0.02fF
C7339 VP.n560 a_400_38200# 0.24fF
C7340 VP.n561 a_400_38200# 0.35fF
C7341 VP.n562 a_400_38200# 0.60fF
C7342 VP.n563 a_400_38200# 0.27fF
C7343 VP.n564 a_400_38200# 0.03fF
C7344 VP.n565 a_400_38200# 0.05fF
C7345 VP.n566 a_400_38200# 0.06fF
C7346 VP.n567 a_400_38200# 0.15fF
C7347 VP.n568 a_400_38200# 0.12fF
C7348 VP.n569 a_400_38200# 0.04fF
C7349 VP.n570 a_400_38200# 0.03fF
C7350 VP.n571 a_400_38200# 0.07fF
C7351 VP.n572 a_400_38200# 0.09fF
C7352 VP.n573 a_400_38200# 0.24fF
C7353 VP.n574 a_400_38200# 0.03fF
C7354 VP.n575 a_400_38200# 0.05fF
C7355 VP.n576 a_400_38200# 0.05fF
C7356 VP.n577 a_400_38200# 0.04fF
C7357 VP.n578 a_400_38200# 0.66fF
C7358 VP.n579 a_400_38200# 0.97fF
C7359 VP.n580 a_400_38200# 1.90fF
C7360 VP.t1155 a_400_38200# 0.02fF
C7361 VP.n581 a_400_38200# 0.12fF
C7362 VP.n582 a_400_38200# 0.14fF
C7363 VP.t973 a_400_38200# 0.02fF
C7364 VP.n584 a_400_38200# 0.24fF
C7365 VP.n585 a_400_38200# 0.91fF
C7366 VP.n586 a_400_38200# 0.05fF
C7367 VP.n587 a_400_38200# 0.10fF
C7368 VP.n588 a_400_38200# 0.17fF
C7369 VP.n589 a_400_38200# 0.10fF
C7370 VP.n590 a_400_38200# 0.13fF
C7371 VP.n591 a_400_38200# 0.37fF
C7372 VP.n592 a_400_38200# 0.08fF
C7373 VP.n593 a_400_38200# 0.09fF
C7374 VP.n594 a_400_38200# 0.20fF
C7375 VP.n595 a_400_38200# 0.01fF
C7376 VP.n596 a_400_38200# 0.21fF
C7377 VP.n597 a_400_38200# 0.24fF
C7378 VP.n598 a_400_38200# 0.04fF
C7379 VP.n599 a_400_38200# 0.02fF
C7380 VP.n600 a_400_38200# 0.06fF
C7381 VP.n601 a_400_38200# 0.69fF
C7382 VP.n602 a_400_38200# 0.10fF
C7383 VP.n603 a_400_38200# 1.92fF
C7384 VP.n604 a_400_38200# 0.12fF
C7385 VP.t370 a_400_38200# 0.02fF
C7386 VP.n605 a_400_38200# 0.14fF
C7387 VP.t814 a_400_38200# 0.02fF
C7388 VP.n607 a_400_38200# 0.24fF
C7389 VP.n608 a_400_38200# 0.35fF
C7390 VP.n609 a_400_38200# 0.60fF
C7391 VP.n610 a_400_38200# 0.03fF
C7392 VP.n611 a_400_38200# 0.07fF
C7393 VP.n612 a_400_38200# 0.09fF
C7394 VP.n613 a_400_38200# 0.24fF
C7395 VP.n614 a_400_38200# 0.03fF
C7396 VP.n615 a_400_38200# 0.05fF
C7397 VP.n616 a_400_38200# 0.05fF
C7398 VP.n617 a_400_38200# 0.04fF
C7399 VP.n618 a_400_38200# 0.82fF
C7400 VP.n619 a_400_38200# 1.66fF
C7401 VP.n620 a_400_38200# 2.04fF
C7402 VP.t706 a_400_38200# 0.02fF
C7403 VP.n621 a_400_38200# 0.12fF
C7404 VP.n622 a_400_38200# 0.14fF
C7405 VP.t524 a_400_38200# 0.02fF
C7406 VP.n624 a_400_38200# 0.24fF
C7407 VP.n625 a_400_38200# 0.91fF
C7408 VP.n626 a_400_38200# 0.05fF
C7409 VP.n627 a_400_38200# 0.10fF
C7410 VP.n628 a_400_38200# 0.17fF
C7411 VP.n629 a_400_38200# 0.10fF
C7412 VP.n630 a_400_38200# 0.13fF
C7413 VP.n631 a_400_38200# 0.37fF
C7414 VP.n632 a_400_38200# 0.08fF
C7415 VP.n633 a_400_38200# 0.09fF
C7416 VP.n634 a_400_38200# 0.20fF
C7417 VP.n635 a_400_38200# 0.01fF
C7418 VP.n636 a_400_38200# 0.21fF
C7419 VP.n637 a_400_38200# 0.24fF
C7420 VP.n638 a_400_38200# 0.04fF
C7421 VP.n639 a_400_38200# 0.02fF
C7422 VP.n640 a_400_38200# 0.06fF
C7423 VP.n641 a_400_38200# 0.69fF
C7424 VP.n642 a_400_38200# 0.10fF
C7425 VP.n643 a_400_38200# 1.92fF
C7426 VP.n644 a_400_38200# 0.12fF
C7427 VP.t1225 a_400_38200# 0.02fF
C7428 VP.n645 a_400_38200# 0.14fF
C7429 VP.t363 a_400_38200# 0.02fF
C7430 VP.n647 a_400_38200# 0.24fF
C7431 VP.n648 a_400_38200# 0.35fF
C7432 VP.n649 a_400_38200# 0.60fF
C7433 VP.n650 a_400_38200# 2.21fF
C7434 VP.t262 a_400_38200# 0.02fF
C7435 VP.n651 a_400_38200# 0.12fF
C7436 VP.n652 a_400_38200# 0.14fF
C7437 VP.t46 a_400_38200# 0.02fF
C7438 VP.n654 a_400_38200# 0.24fF
C7439 VP.n655 a_400_38200# 0.91fF
C7440 VP.n656 a_400_38200# 0.05fF
C7441 VP.n657 a_400_38200# 0.10fF
C7442 VP.n658 a_400_38200# 0.17fF
C7443 VP.n659 a_400_38200# 0.10fF
C7444 VP.n660 a_400_38200# 0.13fF
C7445 VP.n661 a_400_38200# 0.37fF
C7446 VP.n662 a_400_38200# 0.08fF
C7447 VP.n663 a_400_38200# 0.09fF
C7448 VP.n664 a_400_38200# 0.20fF
C7449 VP.n665 a_400_38200# 0.01fF
C7450 VP.n666 a_400_38200# 0.21fF
C7451 VP.n667 a_400_38200# 0.24fF
C7452 VP.n668 a_400_38200# 0.04fF
C7453 VP.n669 a_400_38200# 0.02fF
C7454 VP.n670 a_400_38200# 0.06fF
C7455 VP.n671 a_400_38200# 0.69fF
C7456 VP.n672 a_400_38200# 0.10fF
C7457 VP.n673 a_400_38200# 1.92fF
C7458 VP.n674 a_400_38200# 0.12fF
C7459 VP.t780 a_400_38200# 0.02fF
C7460 VP.n675 a_400_38200# 0.14fF
C7461 VP.t1217 a_400_38200# 0.02fF
C7462 VP.n677 a_400_38200# 0.24fF
C7463 VP.n678 a_400_38200# 0.35fF
C7464 VP.n679 a_400_38200# 0.60fF
C7465 VP.n680 a_400_38200# 1.00fF
C7466 VP.n681 a_400_38200# 2.39fF
C7467 VP.n682 a_400_38200# 2.21fF
C7468 VP.t1117 a_400_38200# 0.02fF
C7469 VP.n683 a_400_38200# 0.12fF
C7470 VP.n684 a_400_38200# 0.14fF
C7471 VP.t935 a_400_38200# 0.02fF
C7472 VP.n686 a_400_38200# 0.24fF
C7473 VP.n687 a_400_38200# 0.91fF
C7474 VP.n688 a_400_38200# 0.05fF
C7475 VP.n689 a_400_38200# 0.10fF
C7476 VP.n690 a_400_38200# 0.17fF
C7477 VP.n691 a_400_38200# 0.10fF
C7478 VP.n692 a_400_38200# 0.13fF
C7479 VP.n693 a_400_38200# 0.37fF
C7480 VP.n694 a_400_38200# 0.08fF
C7481 VP.n695 a_400_38200# 0.09fF
C7482 VP.n696 a_400_38200# 0.20fF
C7483 VP.n697 a_400_38200# 0.01fF
C7484 VP.n698 a_400_38200# 0.21fF
C7485 VP.n699 a_400_38200# 0.24fF
C7486 VP.n700 a_400_38200# 0.04fF
C7487 VP.n701 a_400_38200# 0.02fF
C7488 VP.n702 a_400_38200# 0.06fF
C7489 VP.n703 a_400_38200# 0.69fF
C7490 VP.n704 a_400_38200# 0.10fF
C7491 VP.n705 a_400_38200# 1.92fF
C7492 VP.n706 a_400_38200# 0.12fF
C7493 VP.t331 a_400_38200# 0.02fF
C7494 VP.n707 a_400_38200# 0.14fF
C7495 VP.t772 a_400_38200# 0.02fF
C7496 VP.n709 a_400_38200# 0.24fF
C7497 VP.n710 a_400_38200# 0.35fF
C7498 VP.n711 a_400_38200# 0.60fF
C7499 VP.n712 a_400_38200# 0.03fF
C7500 VP.n713 a_400_38200# 0.07fF
C7501 VP.n714 a_400_38200# 0.09fF
C7502 VP.n715 a_400_38200# 0.24fF
C7503 VP.n716 a_400_38200# 0.03fF
C7504 VP.n717 a_400_38200# 0.05fF
C7505 VP.n718 a_400_38200# 0.05fF
C7506 VP.n719 a_400_38200# 0.04fF
C7507 VP.n720 a_400_38200# 0.89fF
C7508 VP.n721 a_400_38200# 1.18fF
C7509 VP.n722 a_400_38200# 2.07fF
C7510 VP.t733 a_400_38200# 0.02fF
C7511 VP.n723 a_400_38200# 0.12fF
C7512 VP.n724 a_400_38200# 0.14fF
C7513 VP.t489 a_400_38200# 0.02fF
C7514 VP.n726 a_400_38200# 0.24fF
C7515 VP.n727 a_400_38200# 0.91fF
C7516 VP.n728 a_400_38200# 0.05fF
C7517 VP.t57 a_400_38200# 34.79fF
C7518 VP.t78 a_400_38200# 0.02fF
C7519 VP.n729 a_400_38200# 0.12fF
C7520 VP.n730 a_400_38200# 0.14fF
C7521 VP.t1144 a_400_38200# 0.02fF
C7522 VP.n732 a_400_38200# 0.24fF
C7523 VP.n733 a_400_38200# 0.91fF
C7524 VP.n734 a_400_38200# 0.05fF
C7525 VP.t107 a_400_38200# 0.02fF
C7526 VP.n735 a_400_38200# 0.24fF
C7527 VP.n736 a_400_38200# 0.35fF
C7528 VP.n737 a_400_38200# 0.60fF
C7529 VP.n738 a_400_38200# 0.03fF
C7530 VP.n739 a_400_38200# 0.03fF
C7531 VP.n740 a_400_38200# 0.07fF
C7532 VP.n741 a_400_38200# 0.09fF
C7533 VP.n742 a_400_38200# 0.24fF
C7534 VP.n743 a_400_38200# 0.03fF
C7535 VP.n744 a_400_38200# 0.05fF
C7536 VP.n745 a_400_38200# 0.05fF
C7537 VP.n746 a_400_38200# 0.04fF
C7538 VP.n747 a_400_38200# 0.29fF
C7539 VP.n748 a_400_38200# 0.62fF
C7540 VP.n749 a_400_38200# 0.02fF
C7541 VP.n750 a_400_38200# 0.10fF
C7542 VP.n751 a_400_38200# 0.36fF
C7543 VP.n752 a_400_38200# 0.04fF
C7544 VP.n753 a_400_38200# 0.06fF
C7545 VP.n754 a_400_38200# 0.05fF
C7546 VP.n755 a_400_38200# 0.18fF
C7547 VP.n756 a_400_38200# 0.21fF
C7548 VP.n757 a_400_38200# 0.30fF
C7549 VP.n758 a_400_38200# 1.74fF
C7550 VP.n759 a_400_38200# 1.96fF
C7551 VP.n760 a_400_38200# 1.04fF
C7552 VP.n761 a_400_38200# 0.05fF
C7553 VP.n762 a_400_38200# 0.03fF
C7554 VP.n763 a_400_38200# 0.06fF
C7555 VP.n764 a_400_38200# 0.06fF
C7556 VP.n765 a_400_38200# 0.06fF
C7557 VP.n766 a_400_38200# 0.07fF
C7558 VP.n767 a_400_38200# 0.03fF
C7559 VP.n768 a_400_38200# 0.05fF
C7560 VP.n769 a_400_38200# 0.07fF
C7561 VP.n770 a_400_38200# 0.19fF
C7562 VP.n771 a_400_38200# 0.60fF
C7563 VP.n772 a_400_38200# 0.76fF
C7564 VP.n773 a_400_38200# 0.40fF
C7565 VP.n774 a_400_38200# 0.03fF
C7566 VP.n775 a_400_38200# 0.01fF
C7567 VP.t975 a_400_38200# 0.02fF
C7568 VP.n776 a_400_38200# 0.25fF
C7569 VP.t843 a_400_38200# 0.02fF
C7570 VP.n777 a_400_38200# 0.95fF
C7571 VP.n778 a_400_38200# 0.70fF
C7572 VP.n779 a_400_38200# 1.93fF
C7573 VP.n780 a_400_38200# 1.01fF
C7574 VP.n781 a_400_38200# 2.77fF
C7575 VP.n782 a_400_38200# 2.27fF
C7576 VP.t446 a_400_38200# 0.02fF
C7577 VP.n783 a_400_38200# 0.24fF
C7578 VP.n784 a_400_38200# 0.35fF
C7579 VP.n785 a_400_38200# 0.60fF
C7580 VP.t1199 a_400_38200# 0.02fF
C7581 VP.n786 a_400_38200# 0.12fF
C7582 VP.n787 a_400_38200# 0.14fF
C7583 VP.n789 a_400_38200# 0.12fF
C7584 VP.t1152 a_400_38200# 0.02fF
C7585 VP.n790 a_400_38200# 0.14fF
C7586 VP.n792 a_400_38200# 0.04fF
C7587 VP.n793 a_400_38200# 0.02fF
C7588 VP.n794 a_400_38200# 0.06fF
C7589 VP.n795 a_400_38200# 0.30fF
C7590 VP.n796 a_400_38200# 0.10fF
C7591 VP.n797 a_400_38200# 0.28fF
C7592 VP.n798 a_400_38200# 0.06fF
C7593 VP.n799 a_400_38200# 0.06fF
C7594 VP.n800 a_400_38200# 0.03fF
C7595 VP.n801 a_400_38200# 0.15fF
C7596 VP.n802 a_400_38200# 0.08fF
C7597 VP.n803 a_400_38200# 0.14fF
C7598 VP.n804 a_400_38200# 0.03fF
C7599 VP.n805 a_400_38200# 0.06fF
C7600 VP.n806 a_400_38200# 0.06fF
C7601 VP.n807 a_400_38200# 0.06fF
C7602 VP.n808 a_400_38200# 0.06fF
C7603 VP.n809 a_400_38200# 0.03fF
C7604 VP.n810 a_400_38200# 0.05fF
C7605 VP.n811 a_400_38200# 0.07fF
C7606 VP.n812 a_400_38200# 0.19fF
C7607 VP.n813 a_400_38200# 0.59fF
C7608 VP.n814 a_400_38200# 0.34fF
C7609 VP.n815 a_400_38200# 1.88fF
C7610 VP.t1017 a_400_38200# 0.02fF
C7611 VP.n816 a_400_38200# 0.24fF
C7612 VP.n817 a_400_38200# 0.91fF
C7613 VP.n818 a_400_38200# 0.05fF
C7614 VP.t572 a_400_38200# 0.02fF
C7615 VP.n819 a_400_38200# 0.24fF
C7616 VP.n820 a_400_38200# 0.91fF
C7617 VP.n821 a_400_38200# 0.05fF
C7618 VP.n822 a_400_38200# 0.19fF
C7619 VP.n823 a_400_38200# 0.10fF
C7620 VP.n824 a_400_38200# 0.10fF
C7621 VP.n825 a_400_38200# 0.18fF
C7622 VP.n826 a_400_38200# 0.09fF
C7623 VP.n827 a_400_38200# 0.04fF
C7624 VP.n828 a_400_38200# 0.03fF
C7625 VP.n829 a_400_38200# 0.03fF
C7626 VP.n830 a_400_38200# 0.08fF
C7627 VP.n831 a_400_38200# 0.26fF
C7628 VP.n832 a_400_38200# 1.07fF
C7629 VP.n833 a_400_38200# 0.06fF
C7630 VP.n834 a_400_38200# 0.44fF
C7631 VP.n835 a_400_38200# 0.13fF
C7632 VP.n836 a_400_38200# 0.02fF
C7633 VP.n837 a_400_38200# 1.81fF
C7634 VP.n838 a_400_38200# 0.12fF
C7635 VP.t704 a_400_38200# 0.02fF
C7636 VP.n839 a_400_38200# 0.14fF
C7637 VP.t1300 a_400_38200# 0.02fF
C7638 VP.n841 a_400_38200# 0.24fF
C7639 VP.n842 a_400_38200# 0.35fF
C7640 VP.n843 a_400_38200# 0.60fF
C7641 VP.n844 a_400_38200# 0.81fF
C7642 VP.n845 a_400_38200# 2.99fF
C7643 VP.n846 a_400_38200# 2.06fF
C7644 VP.n847 a_400_38200# 1.98fF
C7645 VP.t750 a_400_38200# 0.02fF
C7646 VP.n848 a_400_38200# 0.12fF
C7647 VP.n849 a_400_38200# 0.14fF
C7648 VP.n851 a_400_38200# 1.73fF
C7649 VP.n852 a_400_38200# 0.12fF
C7650 VP.n853 a_400_38200# 0.11fF
C7651 VP.n854 a_400_38200# 0.94fF
C7652 VP.n855 a_400_38200# 0.25fF
C7653 VP.n856 a_400_38200# 0.19fF
C7654 VP.n857 a_400_38200# 0.09fF
C7655 VP.n858 a_400_38200# 0.18fF
C7656 VP.n859 a_400_38200# 0.09fF
C7657 VP.n860 a_400_38200# 0.08fF
C7658 VP.n861 a_400_38200# 0.39fF
C7659 VP.n862 a_400_38200# 0.24fF
C7660 VP.n863 a_400_38200# 0.13fF
C7661 VP.n864 a_400_38200# 0.02fF
C7662 VP.n865 a_400_38200# 2.05fF
C7663 VP.n866 a_400_38200# 0.12fF
C7664 VP.t961 a_400_38200# 0.02fF
C7665 VP.n867 a_400_38200# 0.14fF
C7666 VP.t242 a_400_38200# 0.02fF
C7667 VP.n869 a_400_38200# 0.24fF
C7668 VP.n870 a_400_38200# 0.35fF
C7669 VP.n871 a_400_38200# 0.60fF
C7670 VP.n872 a_400_38200# 2.75fF
C7671 VP.n873 a_400_38200# 1.98fF
C7672 VP.t830 a_400_38200# 0.02fF
C7673 VP.n874 a_400_38200# 0.24fF
C7674 VP.n875 a_400_38200# 0.91fF
C7675 VP.n876 a_400_38200# 0.05fF
C7676 VP.t296 a_400_38200# 0.02fF
C7677 VP.n877 a_400_38200# 0.12fF
C7678 VP.n878 a_400_38200# 0.14fF
C7679 VP.n880 a_400_38200# 15.28fF
C7680 VP.n881 a_400_38200# 0.10fF
C7681 VP.n882 a_400_38200# 0.06fF
C7682 VP.n883 a_400_38200# 0.06fF
C7683 VP.n884 a_400_38200# 0.28fF
C7684 VP.n885 a_400_38200# 0.03fF
C7685 VP.n886 a_400_38200# 0.15fF
C7686 VP.n887 a_400_38200# 0.08fF
C7687 VP.n888 a_400_38200# 0.14fF
C7688 VP.n889 a_400_38200# 0.03fF
C7689 VP.n890 a_400_38200# 0.06fF
C7690 VP.n891 a_400_38200# 0.06fF
C7691 VP.n892 a_400_38200# 0.06fF
C7692 VP.n893 a_400_38200# 0.06fF
C7693 VP.n894 a_400_38200# 0.03fF
C7694 VP.n895 a_400_38200# 0.05fF
C7695 VP.n896 a_400_38200# 0.07fF
C7696 VP.n897 a_400_38200# 0.19fF
C7697 VP.n898 a_400_38200# 0.59fF
C7698 VP.n899 a_400_38200# 0.34fF
C7699 VP.n900 a_400_38200# 0.04fF
C7700 VP.n901 a_400_38200# 0.02fF
C7701 VP.n902 a_400_38200# 0.06fF
C7702 VP.n903 a_400_38200# 0.30fF
C7703 VP.n904 a_400_38200# 1.93fF
C7704 VP.n905 a_400_38200# 0.12fF
C7705 VP.t527 a_400_38200# 0.02fF
C7706 VP.n906 a_400_38200# 0.14fF
C7707 VP.t1109 a_400_38200# 0.02fF
C7708 VP.n908 a_400_38200# 0.24fF
C7709 VP.n909 a_400_38200# 0.35fF
C7710 VP.n910 a_400_38200# 0.60fF
C7711 VP.n911 a_400_38200# 0.07fF
C7712 VP.n912 a_400_38200# 0.72fF
C7713 VP.n913 a_400_38200# 0.20fF
C7714 VP.n914 a_400_38200# 0.19fF
C7715 VP.n915 a_400_38200# 0.10fF
C7716 VP.n916 a_400_38200# 0.11fF
C7717 VP.n917 a_400_38200# 0.09fF
C7718 VP.n918 a_400_38200# 0.16fF
C7719 VP.n919 a_400_38200# 0.11fF
C7720 VP.n920 a_400_38200# 0.36fF
C7721 VP.n921 a_400_38200# 1.05fF
C7722 VP.n922 a_400_38200# 0.15fF
C7723 VP.n924 a_400_38200# 1.72fF
C7724 VP.t563 a_400_38200# 0.02fF
C7725 VP.n925 a_400_38200# 0.12fF
C7726 VP.n926 a_400_38200# 0.14fF
C7727 VP.t391 a_400_38200# 0.02fF
C7728 VP.n928 a_400_38200# 0.24fF
C7729 VP.n929 a_400_38200# 0.91fF
C7730 VP.n930 a_400_38200# 0.05fF
C7731 VP.n931 a_400_38200# 0.10fF
C7732 VP.n932 a_400_38200# 0.06fF
C7733 VP.n933 a_400_38200# 0.06fF
C7734 VP.n934 a_400_38200# 0.28fF
C7735 VP.n935 a_400_38200# 0.03fF
C7736 VP.n936 a_400_38200# 0.15fF
C7737 VP.n937 a_400_38200# 0.08fF
C7738 VP.n938 a_400_38200# 0.14fF
C7739 VP.n939 a_400_38200# 0.03fF
C7740 VP.n940 a_400_38200# 0.06fF
C7741 VP.n941 a_400_38200# 0.06fF
C7742 VP.n942 a_400_38200# 0.06fF
C7743 VP.n943 a_400_38200# 0.06fF
C7744 VP.n944 a_400_38200# 0.03fF
C7745 VP.n945 a_400_38200# 0.05fF
C7746 VP.n946 a_400_38200# 0.07fF
C7747 VP.n947 a_400_38200# 0.19fF
C7748 VP.n948 a_400_38200# 0.59fF
C7749 VP.n949 a_400_38200# 0.34fF
C7750 VP.n950 a_400_38200# 0.04fF
C7751 VP.n951 a_400_38200# 0.02fF
C7752 VP.n952 a_400_38200# 0.06fF
C7753 VP.n953 a_400_38200# 0.30fF
C7754 VP.n954 a_400_38200# 1.93fF
C7755 VP.n955 a_400_38200# 0.12fF
C7756 VP.t50 a_400_38200# 0.02fF
C7757 VP.n956 a_400_38200# 0.14fF
C7758 VP.t667 a_400_38200# 0.02fF
C7759 VP.n958 a_400_38200# 0.24fF
C7760 VP.n959 a_400_38200# 0.35fF
C7761 VP.n960 a_400_38200# 0.60fF
C7762 VP.n961 a_400_38200# 0.07fF
C7763 VP.n962 a_400_38200# 0.72fF
C7764 VP.n963 a_400_38200# 0.20fF
C7765 VP.n964 a_400_38200# 0.19fF
C7766 VP.n965 a_400_38200# 0.10fF
C7767 VP.n966 a_400_38200# 0.11fF
C7768 VP.n967 a_400_38200# 0.09fF
C7769 VP.n968 a_400_38200# 0.16fF
C7770 VP.n969 a_400_38200# 0.11fF
C7771 VP.n970 a_400_38200# 0.36fF
C7772 VP.n971 a_400_38200# 1.05fF
C7773 VP.n972 a_400_38200# 0.15fF
C7774 VP.n974 a_400_38200# 1.72fF
C7775 VP.t93 a_400_38200# 0.02fF
C7776 VP.n975 a_400_38200# 0.12fF
C7777 VP.n976 a_400_38200# 0.14fF
C7778 VP.t1248 a_400_38200# 0.02fF
C7779 VP.n978 a_400_38200# 0.24fF
C7780 VP.n979 a_400_38200# 0.91fF
C7781 VP.n980 a_400_38200# 0.05fF
C7782 VP.n981 a_400_38200# 0.10fF
C7783 VP.n982 a_400_38200# 0.28fF
C7784 VP.n983 a_400_38200# 0.06fF
C7785 VP.n984 a_400_38200# 0.06fF
C7786 VP.n985 a_400_38200# 0.03fF
C7787 VP.n986 a_400_38200# 0.15fF
C7788 VP.n987 a_400_38200# 0.08fF
C7789 VP.n988 a_400_38200# 0.14fF
C7790 VP.n989 a_400_38200# 0.03fF
C7791 VP.n990 a_400_38200# 0.06fF
C7792 VP.n991 a_400_38200# 0.06fF
C7793 VP.n992 a_400_38200# 0.06fF
C7794 VP.n993 a_400_38200# 0.06fF
C7795 VP.n994 a_400_38200# 0.03fF
C7796 VP.n995 a_400_38200# 0.05fF
C7797 VP.n996 a_400_38200# 0.07fF
C7798 VP.n997 a_400_38200# 0.19fF
C7799 VP.n998 a_400_38200# 0.59fF
C7800 VP.n999 a_400_38200# 0.34fF
C7801 VP.n1000 a_400_38200# 0.04fF
C7802 VP.n1001 a_400_38200# 0.02fF
C7803 VP.n1002 a_400_38200# 0.06fF
C7804 VP.n1003 a_400_38200# 0.30fF
C7805 VP.n1004 a_400_38200# 1.93fF
C7806 VP.n1005 a_400_38200# 0.12fF
C7807 VP.t334 a_400_38200# 0.02fF
C7808 VP.n1006 a_400_38200# 0.14fF
C7809 VP.t921 a_400_38200# 0.02fF
C7810 VP.n1008 a_400_38200# 0.24fF
C7811 VP.n1009 a_400_38200# 0.35fF
C7812 VP.n1010 a_400_38200# 0.60fF
C7813 VP.n1011 a_400_38200# 0.07fF
C7814 VP.n1012 a_400_38200# 0.72fF
C7815 VP.n1013 a_400_38200# 0.20fF
C7816 VP.n1014 a_400_38200# 0.19fF
C7817 VP.n1015 a_400_38200# 0.10fF
C7818 VP.n1016 a_400_38200# 0.11fF
C7819 VP.n1017 a_400_38200# 0.09fF
C7820 VP.n1018 a_400_38200# 0.16fF
C7821 VP.n1019 a_400_38200# 0.11fF
C7822 VP.n1020 a_400_38200# 0.36fF
C7823 VP.n1021 a_400_38200# 1.05fF
C7824 VP.n1022 a_400_38200# 0.15fF
C7825 VP.n1024 a_400_38200# 1.72fF
C7826 VP.t969 a_400_38200# 0.02fF
C7827 VP.n1025 a_400_38200# 0.12fF
C7828 VP.n1026 a_400_38200# 0.14fF
C7829 VP.t194 a_400_38200# 0.02fF
C7830 VP.n1028 a_400_38200# 0.24fF
C7831 VP.n1029 a_400_38200# 0.91fF
C7832 VP.n1030 a_400_38200# 0.05fF
C7833 VP.n1031 a_400_38200# 0.10fF
C7834 VP.n1032 a_400_38200# 0.28fF
C7835 VP.n1033 a_400_38200# 0.06fF
C7836 VP.n1034 a_400_38200# 0.06fF
C7837 VP.n1035 a_400_38200# 0.03fF
C7838 VP.n1036 a_400_38200# 0.15fF
C7839 VP.n1037 a_400_38200# 0.08fF
C7840 VP.n1038 a_400_38200# 0.14fF
C7841 VP.n1039 a_400_38200# 0.03fF
C7842 VP.n1040 a_400_38200# 0.06fF
C7843 VP.n1041 a_400_38200# 0.06fF
C7844 VP.n1042 a_400_38200# 0.06fF
C7845 VP.n1043 a_400_38200# 0.06fF
C7846 VP.n1044 a_400_38200# 0.03fF
C7847 VP.n1045 a_400_38200# 0.05fF
C7848 VP.n1046 a_400_38200# 0.07fF
C7849 VP.n1047 a_400_38200# 0.19fF
C7850 VP.n1048 a_400_38200# 0.59fF
C7851 VP.n1049 a_400_38200# 0.34fF
C7852 VP.n1050 a_400_38200# 0.04fF
C7853 VP.n1051 a_400_38200# 0.02fF
C7854 VP.n1052 a_400_38200# 0.06fF
C7855 VP.n1053 a_400_38200# 0.30fF
C7856 VP.n1054 a_400_38200# 1.93fF
C7857 VP.n1055 a_400_38200# 0.12fF
C7858 VP.t1180 a_400_38200# 0.02fF
C7859 VP.n1056 a_400_38200# 0.14fF
C7860 VP.t472 a_400_38200# 0.02fF
C7861 VP.n1058 a_400_38200# 0.24fF
C7862 VP.n1059 a_400_38200# 0.35fF
C7863 VP.n1060 a_400_38200# 0.60fF
C7864 VP.n1061 a_400_38200# 0.07fF
C7865 VP.n1062 a_400_38200# 0.72fF
C7866 VP.n1063 a_400_38200# 0.20fF
C7867 VP.n1064 a_400_38200# 0.19fF
C7868 VP.n1065 a_400_38200# 0.10fF
C7869 VP.n1066 a_400_38200# 0.11fF
C7870 VP.n1067 a_400_38200# 0.09fF
C7871 VP.n1068 a_400_38200# 0.16fF
C7872 VP.n1069 a_400_38200# 0.11fF
C7873 VP.n1070 a_400_38200# 0.36fF
C7874 VP.n1071 a_400_38200# 1.05fF
C7875 VP.n1072 a_400_38200# 0.15fF
C7876 VP.n1074 a_400_38200# 1.72fF
C7877 VP.t1282 a_400_38200# 0.02fF
C7878 VP.n1075 a_400_38200# 0.12fF
C7879 VP.n1076 a_400_38200# 0.14fF
C7880 VP.t1048 a_400_38200# 0.02fF
C7881 VP.n1078 a_400_38200# 0.24fF
C7882 VP.n1079 a_400_38200# 0.91fF
C7883 VP.n1080 a_400_38200# 0.05fF
C7884 VP.n1081 a_400_38200# 0.10fF
C7885 VP.n1082 a_400_38200# 0.06fF
C7886 VP.n1083 a_400_38200# 0.06fF
C7887 VP.n1084 a_400_38200# 0.28fF
C7888 VP.n1085 a_400_38200# 0.03fF
C7889 VP.n1086 a_400_38200# 0.15fF
C7890 VP.n1087 a_400_38200# 0.08fF
C7891 VP.n1088 a_400_38200# 0.14fF
C7892 VP.n1089 a_400_38200# 0.03fF
C7893 VP.n1090 a_400_38200# 0.06fF
C7894 VP.n1091 a_400_38200# 0.06fF
C7895 VP.n1092 a_400_38200# 0.06fF
C7896 VP.n1093 a_400_38200# 0.06fF
C7897 VP.n1094 a_400_38200# 0.03fF
C7898 VP.n1095 a_400_38200# 0.05fF
C7899 VP.n1096 a_400_38200# 0.07fF
C7900 VP.n1097 a_400_38200# 0.19fF
C7901 VP.n1098 a_400_38200# 0.59fF
C7902 VP.n1099 a_400_38200# 0.34fF
C7903 VP.n1100 a_400_38200# 0.04fF
C7904 VP.n1101 a_400_38200# 0.02fF
C7905 VP.n1102 a_400_38200# 0.06fF
C7906 VP.n1103 a_400_38200# 0.30fF
C7907 VP.n1104 a_400_38200# 1.93fF
C7908 VP.n1105 a_400_38200# 0.12fF
C7909 VP.t728 a_400_38200# 0.02fF
C7910 VP.n1106 a_400_38200# 0.14fF
C7911 VP.t1320 a_400_38200# 0.02fF
C7912 VP.n1108 a_400_38200# 0.24fF
C7913 VP.n1109 a_400_38200# 0.35fF
C7914 VP.n1110 a_400_38200# 0.60fF
C7915 VP.n1111 a_400_38200# 0.07fF
C7916 VP.n1112 a_400_38200# 0.72fF
C7917 VP.n1113 a_400_38200# 0.20fF
C7918 VP.n1114 a_400_38200# 0.19fF
C7919 VP.n1115 a_400_38200# 0.10fF
C7920 VP.n1116 a_400_38200# 0.11fF
C7921 VP.n1117 a_400_38200# 0.09fF
C7922 VP.n1118 a_400_38200# 0.16fF
C7923 VP.n1119 a_400_38200# 0.11fF
C7924 VP.n1120 a_400_38200# 0.36fF
C7925 VP.n1121 a_400_38200# 1.05fF
C7926 VP.n1122 a_400_38200# 0.15fF
C7927 VP.n1124 a_400_38200# 1.72fF
C7928 VP.t837 a_400_38200# 0.02fF
C7929 VP.n1125 a_400_38200# 0.12fF
C7930 VP.n1126 a_400_38200# 0.14fF
C7931 VP.t598 a_400_38200# 0.02fF
C7932 VP.n1128 a_400_38200# 0.24fF
C7933 VP.n1129 a_400_38200# 0.91fF
C7934 VP.n1130 a_400_38200# 0.05fF
C7935 VP.n1131 a_400_38200# 0.10fF
C7936 VP.n1132 a_400_38200# 0.06fF
C7937 VP.n1133 a_400_38200# 0.06fF
C7938 VP.n1134 a_400_38200# 0.28fF
C7939 VP.n1135 a_400_38200# 0.03fF
C7940 VP.n1136 a_400_38200# 0.15fF
C7941 VP.n1137 a_400_38200# 0.08fF
C7942 VP.n1138 a_400_38200# 0.14fF
C7943 VP.n1139 a_400_38200# 0.03fF
C7944 VP.n1140 a_400_38200# 0.06fF
C7945 VP.n1141 a_400_38200# 0.06fF
C7946 VP.n1142 a_400_38200# 0.06fF
C7947 VP.n1143 a_400_38200# 0.06fF
C7948 VP.n1144 a_400_38200# 0.03fF
C7949 VP.n1145 a_400_38200# 0.05fF
C7950 VP.n1146 a_400_38200# 0.07fF
C7951 VP.n1147 a_400_38200# 0.19fF
C7952 VP.n1148 a_400_38200# 0.59fF
C7953 VP.n1149 a_400_38200# 0.34fF
C7954 VP.n1150 a_400_38200# 0.04fF
C7955 VP.n1151 a_400_38200# 0.02fF
C7956 VP.n1152 a_400_38200# 0.06fF
C7957 VP.n1153 a_400_38200# 0.30fF
C7958 VP.n1154 a_400_38200# 1.93fF
C7959 VP.n1155 a_400_38200# 0.12fF
C7960 VP.t278 a_400_38200# 0.02fF
C7961 VP.n1156 a_400_38200# 0.14fF
C7962 VP.t870 a_400_38200# 0.02fF
C7963 VP.n1158 a_400_38200# 0.24fF
C7964 VP.n1159 a_400_38200# 0.35fF
C7965 VP.n1160 a_400_38200# 0.60fF
C7966 VP.n1161 a_400_38200# 2.99fF
C7967 VP.n1162 a_400_38200# 1.88fF
C7968 VP.t386 a_400_38200# 0.02fF
C7969 VP.n1163 a_400_38200# 0.12fF
C7970 VP.n1164 a_400_38200# 0.14fF
C7971 VP.t130 a_400_38200# 0.02fF
C7972 VP.n1166 a_400_38200# 0.24fF
C7973 VP.n1167 a_400_38200# 0.91fF
C7974 VP.n1168 a_400_38200# 0.05fF
C7975 VP.n1169 a_400_38200# 0.10fF
C7976 VP.n1170 a_400_38200# 0.28fF
C7977 VP.n1171 a_400_38200# 0.06fF
C7978 VP.n1172 a_400_38200# 0.06fF
C7979 VP.n1173 a_400_38200# 0.03fF
C7980 VP.n1174 a_400_38200# 0.15fF
C7981 VP.n1175 a_400_38200# 0.08fF
C7982 VP.n1176 a_400_38200# 0.14fF
C7983 VP.n1177 a_400_38200# 0.03fF
C7984 VP.n1178 a_400_38200# 0.06fF
C7985 VP.n1179 a_400_38200# 0.06fF
C7986 VP.n1180 a_400_38200# 0.06fF
C7987 VP.n1181 a_400_38200# 0.06fF
C7988 VP.n1182 a_400_38200# 0.03fF
C7989 VP.n1183 a_400_38200# 0.05fF
C7990 VP.n1184 a_400_38200# 0.07fF
C7991 VP.n1185 a_400_38200# 0.19fF
C7992 VP.n1186 a_400_38200# 0.59fF
C7993 VP.n1187 a_400_38200# 0.34fF
C7994 VP.n1188 a_400_38200# 0.04fF
C7995 VP.n1189 a_400_38200# 0.02fF
C7996 VP.n1190 a_400_38200# 0.06fF
C7997 VP.n1191 a_400_38200# 0.30fF
C7998 VP.n1192 a_400_38200# 1.93fF
C7999 VP.n1193 a_400_38200# 0.12fF
C8000 VP.t1132 a_400_38200# 0.02fF
C8001 VP.n1194 a_400_38200# 0.14fF
C8002 VP.t424 a_400_38200# 0.02fF
C8003 VP.n1196 a_400_38200# 0.24fF
C8004 VP.n1197 a_400_38200# 0.35fF
C8005 VP.n1198 a_400_38200# 0.60fF
C8006 VP.n1199 a_400_38200# 1.00fF
C8007 VP.n1200 a_400_38200# 2.77fF
C8008 VP.n1201 a_400_38200# 2.25fF
C8009 VP.n1202 a_400_38200# 1.88fF
C8010 VP.t1242 a_400_38200# 0.02fF
C8011 VP.n1203 a_400_38200# 0.12fF
C8012 VP.n1204 a_400_38200# 0.14fF
C8013 VP.t997 a_400_38200# 0.02fF
C8014 VP.n1206 a_400_38200# 0.24fF
C8015 VP.n1207 a_400_38200# 0.91fF
C8016 VP.n1208 a_400_38200# 0.05fF
C8017 VP.n1209 a_400_38200# 0.10fF
C8018 VP.n1210 a_400_38200# 0.28fF
C8019 VP.n1211 a_400_38200# 0.06fF
C8020 VP.n1212 a_400_38200# 0.06fF
C8021 VP.n1213 a_400_38200# 0.03fF
C8022 VP.n1214 a_400_38200# 0.15fF
C8023 VP.n1215 a_400_38200# 0.08fF
C8024 VP.n1216 a_400_38200# 0.14fF
C8025 VP.n1217 a_400_38200# 0.03fF
C8026 VP.n1218 a_400_38200# 0.06fF
C8027 VP.n1219 a_400_38200# 0.06fF
C8028 VP.n1220 a_400_38200# 0.06fF
C8029 VP.n1221 a_400_38200# 0.06fF
C8030 VP.n1222 a_400_38200# 0.03fF
C8031 VP.n1223 a_400_38200# 0.05fF
C8032 VP.n1224 a_400_38200# 0.07fF
C8033 VP.n1225 a_400_38200# 0.19fF
C8034 VP.n1226 a_400_38200# 0.59fF
C8035 VP.n1227 a_400_38200# 0.34fF
C8036 VP.n1228 a_400_38200# 0.04fF
C8037 VP.n1229 a_400_38200# 0.02fF
C8038 VP.n1230 a_400_38200# 0.06fF
C8039 VP.n1231 a_400_38200# 0.30fF
C8040 VP.n1232 a_400_38200# 1.93fF
C8041 VP.n1233 a_400_38200# 0.12fF
C8042 VP.t685 a_400_38200# 0.02fF
C8043 VP.n1234 a_400_38200# 0.14fF
C8044 VP.t1278 a_400_38200# 0.02fF
C8045 VP.n1236 a_400_38200# 0.24fF
C8046 VP.n1237 a_400_38200# 0.35fF
C8047 VP.n1238 a_400_38200# 0.60fF
C8048 VP.n1239 a_400_38200# 0.72fF
C8049 VP.n1240 a_400_38200# 1.24fF
C8050 VP.n1241 a_400_38200# 0.54fF
C8051 VP.n1242 a_400_38200# 0.22fF
C8052 VP.n1243 a_400_38200# 1.73fF
C8053 VP.t797 a_400_38200# 0.02fF
C8054 VP.n1244 a_400_38200# 0.12fF
C8055 VP.n1245 a_400_38200# 0.14fF
C8056 VP.t552 a_400_38200# 0.02fF
C8057 VP.n1247 a_400_38200# 0.24fF
C8058 VP.n1248 a_400_38200# 0.91fF
C8059 VP.n1249 a_400_38200# 0.05fF
C8060 VP.n1250 a_400_38200# 0.10fF
C8061 VP.n1251 a_400_38200# 0.28fF
C8062 VP.n1252 a_400_38200# 0.06fF
C8063 VP.n1253 a_400_38200# 0.06fF
C8064 VP.n1254 a_400_38200# 0.03fF
C8065 VP.n1255 a_400_38200# 0.15fF
C8066 VP.n1256 a_400_38200# 0.08fF
C8067 VP.n1257 a_400_38200# 0.14fF
C8068 VP.n1258 a_400_38200# 0.03fF
C8069 VP.n1259 a_400_38200# 0.06fF
C8070 VP.n1260 a_400_38200# 0.06fF
C8071 VP.n1261 a_400_38200# 0.06fF
C8072 VP.n1262 a_400_38200# 0.06fF
C8073 VP.n1263 a_400_38200# 0.03fF
C8074 VP.n1264 a_400_38200# 0.05fF
C8075 VP.n1265 a_400_38200# 0.07fF
C8076 VP.n1266 a_400_38200# 0.19fF
C8077 VP.n1267 a_400_38200# 0.59fF
C8078 VP.n1268 a_400_38200# 0.34fF
C8079 VP.n1269 a_400_38200# 0.04fF
C8080 VP.n1270 a_400_38200# 0.02fF
C8081 VP.n1271 a_400_38200# 0.06fF
C8082 VP.n1272 a_400_38200# 0.30fF
C8083 VP.n1273 a_400_38200# 1.93fF
C8084 VP.n1274 a_400_38200# 0.12fF
C8085 VP.t305 a_400_38200# 0.02fF
C8086 VP.n1275 a_400_38200# 0.14fF
C8087 VP.t834 a_400_38200# 0.02fF
C8088 VP.n1277 a_400_38200# 0.24fF
C8089 VP.n1278 a_400_38200# 0.35fF
C8090 VP.n1279 a_400_38200# 0.60fF
C8091 VP.n1280 a_400_38200# 0.86fF
C8092 VP.n1281 a_400_38200# 1.97fF
C8093 VP.n1282 a_400_38200# 0.54fF
C8094 VP.n1283 a_400_38200# 0.21fF
C8095 VP.n1284 a_400_38200# 1.73fF
C8096 VP.t349 a_400_38200# 0.02fF
C8097 VP.n1285 a_400_38200# 0.12fF
C8098 VP.n1286 a_400_38200# 0.14fF
C8099 VP.t81 a_400_38200# 0.02fF
C8100 VP.n1288 a_400_38200# 0.24fF
C8101 VP.n1289 a_400_38200# 0.91fF
C8102 VP.n1290 a_400_38200# 0.05fF
C8103 VP.t49 a_400_38200# 35.17fF
C8104 VP.t256 a_400_38200# 0.02fF
C8105 VP.n1291 a_400_38200# 1.21fF
C8106 VP.n1292 a_400_38200# 0.25fF
C8107 VP.n1293 a_400_38200# 0.52fF
C8108 VP.n1294 a_400_38200# 10.38fF
C8109 VP.n1295 a_400_38200# 38.02fF
C8110 VP.n1296 a_400_38200# 38.02fF
C8111 VP.n1297 a_400_38200# 0.76fF
C8112 VP.n1298 a_400_38200# 0.27fF
C8113 VP.n1299 a_400_38200# 0.59fF
C8114 VP.n1300 a_400_38200# 0.10fF
C8115 VP.n1301 a_400_38200# 3.02fF
C8116 VP.t45 a_400_38200# 15.72fF
C8117 VP.n1302 a_400_38200# 1.15fF
C8118 VP.n1304 a_400_38200# 13.70fF
C8119 VP.n1306 a_400_38200# 1.99fF
C8120 VP.n1307 a_400_38200# 4.39fF
C8121 VP.n1308 a_400_38200# 0.03fF
C8122 VP.n1309 a_400_38200# 0.05fF
C8123 VP.n1310 a_400_38200# 0.07fF
C8124 VP.n1311 a_400_38200# 0.10fF
C8125 VP.n1312 a_400_38200# 0.04fF
C8126 VP.n1313 a_400_38200# 0.07fF
C8127 VP.n1314 a_400_38200# 0.06fF
C8128 VP.n1315 a_400_38200# 0.06fF
C8129 VP.n1316 a_400_38200# 0.07fF
C8130 VP.n1317 a_400_38200# 0.57fF
C8131 VP.n1318 a_400_38200# 1.88fF
C8132 VP.n1319 a_400_38200# 0.92fF
C8133 VP.n1320 a_400_38200# 2.63fF
C8134 VP.n1321 a_400_38200# 0.10fF
C8135 VP.n1322 a_400_38200# 0.28fF
C8136 VP.n1323 a_400_38200# 0.15fF
C8137 VP.n1324 a_400_38200# 0.08fF
C8138 VP.n1325 a_400_38200# 0.14fF
C8139 VP.n1326 a_400_38200# 0.06fF
C8140 VP.n1327 a_400_38200# 0.06fF
C8141 VP.n1328 a_400_38200# 0.03fF
C8142 VP.n1329 a_400_38200# 0.05fF
C8143 VP.n1330 a_400_38200# 0.07fF
C8144 VP.n1331 a_400_38200# 0.19fF
C8145 VP.n1332 a_400_38200# 0.59fF
C8146 VP.n1333 a_400_38200# 0.34fF
C8147 VP.n1334 a_400_38200# 0.04fF
C8148 VP.n1335 a_400_38200# 0.02fF
C8149 VP.n1336 a_400_38200# 0.06fF
C8150 VP.n1337 a_400_38200# 0.30fF
C8151 VP.n1338 a_400_38200# 0.12fF
C8152 VP.t1134 a_400_38200# 0.02fF
C8153 VP.n1339 a_400_38200# 0.14fF
C8154 VP.n1341 a_400_38200# 1.93fF
C8155 VP.t1065 a_400_38200# 0.02fF
C8156 VP.n1342 a_400_38200# 0.24fF
C8157 VP.n1343 a_400_38200# 0.35fF
C8158 VP.n1344 a_400_38200# 0.60fF
C8159 VP.n1345 a_400_38200# 0.12fF
C8160 VP.t478 a_400_38200# 0.02fF
C8161 VP.n1346 a_400_38200# 0.14fF
C8162 VP.n1348 a_400_38200# 0.04fF
C8163 VP.n1349 a_400_38200# 0.02fF
C8164 VP.n1350 a_400_38200# 0.06fF
C8165 VP.n1351 a_400_38200# 0.30fF
C8166 VP.n1352 a_400_38200# 0.10fF
C8167 VP.n1353 a_400_38200# 0.28fF
C8168 VP.n1354 a_400_38200# 0.15fF
C8169 VP.n1355 a_400_38200# 0.08fF
C8170 VP.n1356 a_400_38200# 0.14fF
C8171 VP.n1357 a_400_38200# 0.06fF
C8172 VP.n1358 a_400_38200# 0.06fF
C8173 VP.n1359 a_400_38200# 0.03fF
C8174 VP.n1360 a_400_38200# 0.05fF
C8175 VP.n1361 a_400_38200# 0.07fF
C8176 VP.n1362 a_400_38200# 0.19fF
C8177 VP.n1363 a_400_38200# 0.59fF
C8178 VP.n1364 a_400_38200# 0.34fF
C8179 VP.n1365 a_400_38200# 2.18fF
C8180 VP.t637 a_400_38200# 0.02fF
C8181 VP.n1366 a_400_38200# 0.24fF
C8182 VP.n1367 a_400_38200# 0.91fF
C8183 VP.n1368 a_400_38200# 0.05fF
C8184 VP.t884 a_400_38200# 0.02fF
C8185 VP.n1369 a_400_38200# 0.12fF
C8186 VP.n1370 a_400_38200# 0.14fF
C8187 VP.n1372 a_400_38200# 0.10fF
C8188 VP.n1373 a_400_38200# 0.10fF
C8189 VP.n1374 a_400_38200# 0.18fF
C8190 VP.n1375 a_400_38200# 0.09fF
C8191 VP.n1376 a_400_38200# 0.04fF
C8192 VP.n1377 a_400_38200# 0.26fF
C8193 VP.n1378 a_400_38200# 1.17fF
C8194 VP.n1379 a_400_38200# 0.06fF
C8195 VP.n1380 a_400_38200# 0.44fF
C8196 VP.n1381 a_400_38200# 0.13fF
C8197 VP.n1382 a_400_38200# 0.02fF
C8198 VP.n1383 a_400_38200# 1.81fF
C8199 VP.n1384 a_400_38200# 0.12fF
C8200 VP.t1325 a_400_38200# 0.02fF
C8201 VP.n1385 a_400_38200# 0.14fF
C8202 VP.t619 a_400_38200# 0.02fF
C8203 VP.n1387 a_400_38200# 0.24fF
C8204 VP.n1388 a_400_38200# 0.35fF
C8205 VP.n1389 a_400_38200# 0.60fF
C8206 VP.n1390 a_400_38200# 2.28fF
C8207 VP.t184 a_400_38200# 0.02fF
C8208 VP.n1391 a_400_38200# 0.24fF
C8209 VP.n1392 a_400_38200# 0.91fF
C8210 VP.n1393 a_400_38200# 0.05fF
C8211 VP.t435 a_400_38200# 0.02fF
C8212 VP.n1394 a_400_38200# 0.12fF
C8213 VP.n1395 a_400_38200# 0.14fF
C8214 VP.n1397 a_400_38200# 0.06fF
C8215 VP.n1398 a_400_38200# 0.11fF
C8216 VP.n1399 a_400_38200# 0.03fF
C8217 VP.n1400 a_400_38200# 0.09fF
C8218 VP.n1401 a_400_38200# 0.05fF
C8219 VP.n1402 a_400_38200# 0.11fF
C8220 VP.n1403 a_400_38200# 0.09fF
C8221 VP.n1404 a_400_38200# 0.09fF
C8222 VP.n1405 a_400_38200# 0.02fF
C8223 VP.n1406 a_400_38200# 0.46fF
C8224 VP.n1407 a_400_38200# 1.81fF
C8225 VP.n1408 a_400_38200# 0.12fF
C8226 VP.t874 a_400_38200# 0.02fF
C8227 VP.n1409 a_400_38200# 0.14fF
C8228 VP.t155 a_400_38200# 0.02fF
C8229 VP.n1411 a_400_38200# 0.24fF
C8230 VP.n1412 a_400_38200# 0.35fF
C8231 VP.n1413 a_400_38200# 0.60fF
C8232 VP.n1414 a_400_38200# 2.43fF
C8233 VP.t1035 a_400_38200# 0.02fF
C8234 VP.n1415 a_400_38200# 0.24fF
C8235 VP.n1416 a_400_38200# 0.91fF
C8236 VP.n1417 a_400_38200# 0.05fF
C8237 VP.t1290 a_400_38200# 0.02fF
C8238 VP.n1418 a_400_38200# 0.12fF
C8239 VP.n1419 a_400_38200# 0.14fF
C8240 VP.n1421 a_400_38200# 2.32fF
C8241 VP.n1422 a_400_38200# 1.29fF
C8242 VP.n1423 a_400_38200# 0.11fF
C8243 VP.n1424 a_400_38200# 0.86fF
C8244 VP.n1425 a_400_38200# 0.12fF
C8245 VP.n1426 a_400_38200# 0.03fF
C8246 VP.n1427 a_400_38200# 0.88fF
C8247 VP.n1428 a_400_38200# 0.48fF
C8248 VP.n1429 a_400_38200# 0.88fF
C8249 VP.n1430 a_400_38200# 0.60fF
C8250 VP.n1431 a_400_38200# 2.33fF
C8251 VP.n1432 a_400_38200# 0.59fF
C8252 VP.n1433 a_400_38200# 0.02fF
C8253 VP.n1434 a_400_38200# 0.96fF
C8254 VP.t80 a_400_38200# 15.72fF
C8255 VP.n1435 a_400_38200# 15.42fF
C8256 VP.n1437 a_400_38200# 0.38fF
C8257 VP.n1438 a_400_38200# 3.61fF
C8258 VP.n1439 a_400_38200# 1.90fF
C8259 VP.t412 a_400_38200# 0.02fF
C8260 VP.n1440 a_400_38200# 0.64fF
C8261 VP.n1441 a_400_38200# 0.60fF
C8262 VP.n1442 a_400_38200# 2.11fF
C8263 VP.t1283 a_400_38200# 0.02fF
C8264 VP.n1443 a_400_38200# 1.19fF
C8265 VP.n1444 a_400_38200# 0.05fF
C8266 VP.t234 a_400_38200# 0.02fF
C8267 VP.n1445 a_400_38200# 0.01fF
C8268 VP.n1446 a_400_38200# 0.26fF
C8269 VP.n1448 a_400_38200# 15.28fF
C8270 VP.n1449 a_400_38200# 0.10fF
C8271 VP.n1450 a_400_38200# 0.28fF
C8272 VP.n1451 a_400_38200# 0.15fF
C8273 VP.n1452 a_400_38200# 0.08fF
C8274 VP.n1453 a_400_38200# 0.14fF
C8275 VP.n1454 a_400_38200# 0.06fF
C8276 VP.n1455 a_400_38200# 0.06fF
C8277 VP.n1456 a_400_38200# 0.03fF
C8278 VP.n1457 a_400_38200# 0.05fF
C8279 VP.n1458 a_400_38200# 0.07fF
C8280 VP.n1459 a_400_38200# 0.19fF
C8281 VP.n1460 a_400_38200# 0.59fF
C8282 VP.n1461 a_400_38200# 0.34fF
C8283 VP.n1462 a_400_38200# 0.04fF
C8284 VP.n1463 a_400_38200# 0.02fF
C8285 VP.n1464 a_400_38200# 0.06fF
C8286 VP.n1465 a_400_38200# 0.30fF
C8287 VP.n1466 a_400_38200# 1.93fF
C8288 VP.n1467 a_400_38200# 0.12fF
C8289 VP.t686 a_400_38200# 0.02fF
C8290 VP.n1468 a_400_38200# 0.14fF
C8291 VP.t1281 a_400_38200# 0.02fF
C8292 VP.n1470 a_400_38200# 0.24fF
C8293 VP.n1471 a_400_38200# 0.35fF
C8294 VP.n1472 a_400_38200# 0.60fF
C8295 VP.n1473 a_400_38200# 0.07fF
C8296 VP.n1474 a_400_38200# 0.72fF
C8297 VP.n1475 a_400_38200# 0.09fF
C8298 VP.n1476 a_400_38200# 0.16fF
C8299 VP.n1477 a_400_38200# 0.98fF
C8300 VP.n1478 a_400_38200# 0.15fF
C8301 VP.n1480 a_400_38200# 1.72fF
C8302 VP.t1101 a_400_38200# 0.02fF
C8303 VP.n1481 a_400_38200# 0.12fF
C8304 VP.n1482 a_400_38200# 0.14fF
C8305 VP.t851 a_400_38200# 0.02fF
C8306 VP.n1484 a_400_38200# 0.24fF
C8307 VP.n1485 a_400_38200# 0.91fF
C8308 VP.n1486 a_400_38200# 0.05fF
C8309 VP.n1487 a_400_38200# 0.10fF
C8310 VP.n1488 a_400_38200# 0.28fF
C8311 VP.n1489 a_400_38200# 0.15fF
C8312 VP.n1490 a_400_38200# 0.08fF
C8313 VP.n1491 a_400_38200# 0.14fF
C8314 VP.n1492 a_400_38200# 0.06fF
C8315 VP.n1493 a_400_38200# 0.06fF
C8316 VP.n1494 a_400_38200# 0.03fF
C8317 VP.n1495 a_400_38200# 0.05fF
C8318 VP.n1496 a_400_38200# 0.07fF
C8319 VP.n1497 a_400_38200# 0.19fF
C8320 VP.n1498 a_400_38200# 0.59fF
C8321 VP.n1499 a_400_38200# 0.34fF
C8322 VP.n1500 a_400_38200# 0.04fF
C8323 VP.n1501 a_400_38200# 0.02fF
C8324 VP.n1502 a_400_38200# 0.06fF
C8325 VP.n1503 a_400_38200# 0.30fF
C8326 VP.n1504 a_400_38200# 1.93fF
C8327 VP.n1505 a_400_38200# 0.12fF
C8328 VP.t240 a_400_38200# 0.02fF
C8329 VP.n1506 a_400_38200# 0.14fF
C8330 VP.t836 a_400_38200# 0.02fF
C8331 VP.n1508 a_400_38200# 0.24fF
C8332 VP.n1509 a_400_38200# 0.35fF
C8333 VP.n1510 a_400_38200# 0.60fF
C8334 VP.n1511 a_400_38200# 0.07fF
C8335 VP.n1512 a_400_38200# 0.72fF
C8336 VP.n1513 a_400_38200# 0.09fF
C8337 VP.n1514 a_400_38200# 0.16fF
C8338 VP.n1515 a_400_38200# 0.98fF
C8339 VP.n1516 a_400_38200# 0.15fF
C8340 VP.n1518 a_400_38200# 1.72fF
C8341 VP.t659 a_400_38200# 0.02fF
C8342 VP.n1519 a_400_38200# 0.12fF
C8343 VP.n1520 a_400_38200# 0.14fF
C8344 VP.t402 a_400_38200# 0.02fF
C8345 VP.n1522 a_400_38200# 0.24fF
C8346 VP.n1523 a_400_38200# 0.91fF
C8347 VP.n1524 a_400_38200# 0.05fF
C8348 VP.n1525 a_400_38200# 0.10fF
C8349 VP.n1526 a_400_38200# 0.28fF
C8350 VP.n1527 a_400_38200# 0.15fF
C8351 VP.n1528 a_400_38200# 0.08fF
C8352 VP.n1529 a_400_38200# 0.14fF
C8353 VP.n1530 a_400_38200# 0.06fF
C8354 VP.n1531 a_400_38200# 0.06fF
C8355 VP.n1532 a_400_38200# 0.03fF
C8356 VP.n1533 a_400_38200# 0.05fF
C8357 VP.n1534 a_400_38200# 0.07fF
C8358 VP.n1535 a_400_38200# 0.19fF
C8359 VP.n1536 a_400_38200# 0.59fF
C8360 VP.n1537 a_400_38200# 0.34fF
C8361 VP.n1538 a_400_38200# 0.04fF
C8362 VP.n1539 a_400_38200# 0.02fF
C8363 VP.n1540 a_400_38200# 0.06fF
C8364 VP.n1541 a_400_38200# 0.30fF
C8365 VP.n1542 a_400_38200# 1.93fF
C8366 VP.n1543 a_400_38200# 0.12fF
C8367 VP.t555 a_400_38200# 0.02fF
C8368 VP.n1544 a_400_38200# 0.14fF
C8369 VP.t1081 a_400_38200# 0.02fF
C8370 VP.n1546 a_400_38200# 0.24fF
C8371 VP.n1547 a_400_38200# 0.35fF
C8372 VP.n1548 a_400_38200# 0.60fF
C8373 VP.n1549 a_400_38200# 0.07fF
C8374 VP.n1550 a_400_38200# 0.72fF
C8375 VP.n1551 a_400_38200# 0.09fF
C8376 VP.n1552 a_400_38200# 0.16fF
C8377 VP.n1553 a_400_38200# 0.98fF
C8378 VP.n1554 a_400_38200# 0.15fF
C8379 VP.n1556 a_400_38200# 1.72fF
C8380 VP.t910 a_400_38200# 0.02fF
C8381 VP.n1557 a_400_38200# 0.12fF
C8382 VP.n1558 a_400_38200# 0.14fF
C8383 VP.t653 a_400_38200# 0.02fF
C8384 VP.n1560 a_400_38200# 0.24fF
C8385 VP.n1561 a_400_38200# 0.91fF
C8386 VP.n1562 a_400_38200# 0.05fF
C8387 VP.n1563 a_400_38200# 0.10fF
C8388 VP.n1564 a_400_38200# 0.28fF
C8389 VP.n1565 a_400_38200# 0.15fF
C8390 VP.n1566 a_400_38200# 0.08fF
C8391 VP.n1567 a_400_38200# 0.14fF
C8392 VP.n1568 a_400_38200# 0.06fF
C8393 VP.n1569 a_400_38200# 0.06fF
C8394 VP.n1570 a_400_38200# 0.03fF
C8395 VP.n1571 a_400_38200# 0.05fF
C8396 VP.n1572 a_400_38200# 0.07fF
C8397 VP.n1573 a_400_38200# 0.19fF
C8398 VP.n1574 a_400_38200# 0.59fF
C8399 VP.n1575 a_400_38200# 0.34fF
C8400 VP.n1576 a_400_38200# 0.04fF
C8401 VP.n1577 a_400_38200# 0.02fF
C8402 VP.n1578 a_400_38200# 0.06fF
C8403 VP.n1579 a_400_38200# 0.30fF
C8404 VP.n1580 a_400_38200# 1.93fF
C8405 VP.n1581 a_400_38200# 0.12fF
C8406 VP.t85 a_400_38200# 0.02fF
C8407 VP.n1582 a_400_38200# 0.14fF
C8408 VP.t688 a_400_38200# 0.02fF
C8409 VP.n1584 a_400_38200# 0.24fF
C8410 VP.n1585 a_400_38200# 0.35fF
C8411 VP.n1586 a_400_38200# 0.60fF
C8412 VP.n1587 a_400_38200# 0.07fF
C8413 VP.n1588 a_400_38200# 0.72fF
C8414 VP.n1589 a_400_38200# 0.09fF
C8415 VP.n1590 a_400_38200# 0.16fF
C8416 VP.n1591 a_400_38200# 0.98fF
C8417 VP.n1592 a_400_38200# 0.15fF
C8418 VP.n1594 a_400_38200# 1.72fF
C8419 VP.t460 a_400_38200# 0.02fF
C8420 VP.n1595 a_400_38200# 0.12fF
C8421 VP.n1596 a_400_38200# 0.14fF
C8422 VP.t260 a_400_38200# 0.02fF
C8423 VP.n1598 a_400_38200# 0.24fF
C8424 VP.n1599 a_400_38200# 0.91fF
C8425 VP.n1600 a_400_38200# 0.05fF
C8426 VP.n1601 a_400_38200# 0.10fF
C8427 VP.n1602 a_400_38200# 0.28fF
C8428 VP.n1603 a_400_38200# 0.15fF
C8429 VP.n1604 a_400_38200# 0.08fF
C8430 VP.n1605 a_400_38200# 0.14fF
C8431 VP.n1606 a_400_38200# 0.06fF
C8432 VP.n1607 a_400_38200# 0.06fF
C8433 VP.n1608 a_400_38200# 0.03fF
C8434 VP.n1609 a_400_38200# 0.05fF
C8435 VP.n1610 a_400_38200# 0.07fF
C8436 VP.n1611 a_400_38200# 0.19fF
C8437 VP.n1612 a_400_38200# 0.59fF
C8438 VP.n1613 a_400_38200# 0.34fF
C8439 VP.n1614 a_400_38200# 0.04fF
C8440 VP.n1615 a_400_38200# 0.02fF
C8441 VP.n1616 a_400_38200# 0.06fF
C8442 VP.n1617 a_400_38200# 0.30fF
C8443 VP.n1618 a_400_38200# 1.93fF
C8444 VP.n1619 a_400_38200# 0.12fF
C8445 VP.t964 a_400_38200# 0.02fF
C8446 VP.n1620 a_400_38200# 0.14fF
C8447 VP.t244 a_400_38200# 0.02fF
C8448 VP.n1622 a_400_38200# 0.24fF
C8449 VP.n1623 a_400_38200# 0.35fF
C8450 VP.n1624 a_400_38200# 0.60fF
C8451 VP.n1625 a_400_38200# 2.59fF
C8452 VP.n1626 a_400_38200# 2.20fF
C8453 VP.t1309 a_400_38200# 0.02fF
C8454 VP.n1627 a_400_38200# 0.12fF
C8455 VP.n1628 a_400_38200# 0.14fF
C8456 VP.t1115 a_400_38200# 0.02fF
C8457 VP.n1630 a_400_38200# 0.24fF
C8458 VP.n1631 a_400_38200# 0.91fF
C8459 VP.n1632 a_400_38200# 0.05fF
C8460 VP.n1633 a_400_38200# 0.10fF
C8461 VP.n1634 a_400_38200# 0.28fF
C8462 VP.n1635 a_400_38200# 0.15fF
C8463 VP.n1636 a_400_38200# 0.08fF
C8464 VP.n1637 a_400_38200# 0.14fF
C8465 VP.n1638 a_400_38200# 0.06fF
C8466 VP.n1639 a_400_38200# 0.06fF
C8467 VP.n1640 a_400_38200# 0.03fF
C8468 VP.n1641 a_400_38200# 0.05fF
C8469 VP.n1642 a_400_38200# 0.07fF
C8470 VP.n1643 a_400_38200# 0.19fF
C8471 VP.n1644 a_400_38200# 0.59fF
C8472 VP.n1645 a_400_38200# 0.34fF
C8473 VP.n1646 a_400_38200# 0.04fF
C8474 VP.n1647 a_400_38200# 0.02fF
C8475 VP.n1648 a_400_38200# 0.06fF
C8476 VP.n1649 a_400_38200# 0.30fF
C8477 VP.n1650 a_400_38200# 1.93fF
C8478 VP.n1651 a_400_38200# 0.12fF
C8479 VP.t516 a_400_38200# 0.02fF
C8480 VP.n1652 a_400_38200# 0.14fF
C8481 VP.t1098 a_400_38200# 0.02fF
C8482 VP.n1654 a_400_38200# 0.24fF
C8483 VP.n1655 a_400_38200# 0.35fF
C8484 VP.n1656 a_400_38200# 0.60fF
C8485 VP.n1657 a_400_38200# 2.59fF
C8486 VP.n1658 a_400_38200# 2.20fF
C8487 VP.t862 a_400_38200# 0.02fF
C8488 VP.n1659 a_400_38200# 0.12fF
C8489 VP.n1660 a_400_38200# 0.14fF
C8490 VP.t671 a_400_38200# 0.02fF
C8491 VP.n1662 a_400_38200# 0.24fF
C8492 VP.n1663 a_400_38200# 0.91fF
C8493 VP.n1664 a_400_38200# 0.05fF
C8494 VP.n1665 a_400_38200# 0.10fF
C8495 VP.n1666 a_400_38200# 0.28fF
C8496 VP.n1667 a_400_38200# 0.15fF
C8497 VP.n1668 a_400_38200# 0.08fF
C8498 VP.n1669 a_400_38200# 0.14fF
C8499 VP.n1670 a_400_38200# 0.06fF
C8500 VP.n1671 a_400_38200# 0.06fF
C8501 VP.n1672 a_400_38200# 0.03fF
C8502 VP.n1673 a_400_38200# 0.05fF
C8503 VP.n1674 a_400_38200# 0.07fF
C8504 VP.n1675 a_400_38200# 0.19fF
C8505 VP.n1676 a_400_38200# 0.59fF
C8506 VP.n1677 a_400_38200# 0.34fF
C8507 VP.n1678 a_400_38200# 0.04fF
C8508 VP.n1679 a_400_38200# 0.02fF
C8509 VP.n1680 a_400_38200# 0.06fF
C8510 VP.n1681 a_400_38200# 0.30fF
C8511 VP.n1682 a_400_38200# 1.93fF
C8512 VP.n1683 a_400_38200# 0.12fF
C8513 VP.t35 a_400_38200# 0.02fF
C8514 VP.n1684 a_400_38200# 0.14fF
C8515 VP.t656 a_400_38200# 0.02fF
C8516 VP.n1686 a_400_38200# 0.24fF
C8517 VP.n1687 a_400_38200# 0.35fF
C8518 VP.n1688 a_400_38200# 0.60fF
C8519 VP.n1689 a_400_38200# 2.47fF
C8520 VP.n1690 a_400_38200# 2.20fF
C8521 VP.t415 a_400_38200# 0.02fF
C8522 VP.n1691 a_400_38200# 0.12fF
C8523 VP.n1692 a_400_38200# 0.14fF
C8524 VP.t224 a_400_38200# 0.02fF
C8525 VP.n1694 a_400_38200# 0.24fF
C8526 VP.n1695 a_400_38200# 0.91fF
C8527 VP.n1696 a_400_38200# 0.05fF
C8528 VP.n1697 a_400_38200# 0.10fF
C8529 VP.n1698 a_400_38200# 0.28fF
C8530 VP.n1699 a_400_38200# 0.15fF
C8531 VP.n1700 a_400_38200# 0.08fF
C8532 VP.n1701 a_400_38200# 0.14fF
C8533 VP.n1702 a_400_38200# 0.06fF
C8534 VP.n1703 a_400_38200# 0.06fF
C8535 VP.n1704 a_400_38200# 0.03fF
C8536 VP.n1705 a_400_38200# 0.05fF
C8537 VP.n1706 a_400_38200# 0.07fF
C8538 VP.n1707 a_400_38200# 0.19fF
C8539 VP.n1708 a_400_38200# 0.59fF
C8540 VP.n1709 a_400_38200# 0.34fF
C8541 VP.n1710 a_400_38200# 0.04fF
C8542 VP.n1711 a_400_38200# 0.02fF
C8543 VP.n1712 a_400_38200# 0.06fF
C8544 VP.n1713 a_400_38200# 0.30fF
C8545 VP.n1714 a_400_38200# 1.93fF
C8546 VP.n1715 a_400_38200# 0.12fF
C8547 VP.t926 a_400_38200# 0.02fF
C8548 VP.n1716 a_400_38200# 0.14fF
C8549 VP.t210 a_400_38200# 0.02fF
C8550 VP.n1718 a_400_38200# 0.24fF
C8551 VP.n1719 a_400_38200# 0.35fF
C8552 VP.n1720 a_400_38200# 0.60fF
C8553 VP.n1721 a_400_38200# 1.30fF
C8554 VP.n1722 a_400_38200# 1.01fF
C8555 VP.n1723 a_400_38200# 1.71fF
C8556 VP.t1272 a_400_38200# 0.02fF
C8557 VP.n1724 a_400_38200# 0.12fF
C8558 VP.n1725 a_400_38200# 0.14fF
C8559 VP.t1079 a_400_38200# 0.02fF
C8560 VP.n1727 a_400_38200# 0.24fF
C8561 VP.n1728 a_400_38200# 0.91fF
C8562 VP.n1729 a_400_38200# 0.05fF
C8563 VP.t34 a_400_38200# 34.79fF
C8564 VP.t246 a_400_38200# 0.02fF
C8565 VP.n1730 a_400_38200# 0.12fF
C8566 VP.n1731 a_400_38200# 0.14fF
C8567 VP.t1298 a_400_38200# 0.02fF
C8568 VP.n1733 a_400_38200# 0.24fF
C8569 VP.n1734 a_400_38200# 0.91fF
C8570 VP.n1735 a_400_38200# 0.05fF
C8571 VP.t427 a_400_38200# 0.02fF
C8572 VP.n1736 a_400_38200# 0.24fF
C8573 VP.n1737 a_400_38200# 0.35fF
C8574 VP.n1738 a_400_38200# 0.60fF
C8575 VP.n1739 a_400_38200# 0.04fF
C8576 VP.n1740 a_400_38200# 0.08fF
C8577 VP.n1741 a_400_38200# 0.72fF
C8578 VP.n1742 a_400_38200# 0.09fF
C8579 VP.n1743 a_400_38200# 0.00fF
C8580 VP.n1744 a_400_38200# 0.98fF
C8581 VP.n1745 a_400_38200# 0.19fF
C8582 VP.n1747 a_400_38200# 1.72fF
C8583 VP.n1748 a_400_38200# 1.96fF
C8584 VP.n1749 a_400_38200# 1.04fF
C8585 VP.n1750 a_400_38200# 0.05fF
C8586 VP.n1751 a_400_38200# 0.03fF
C8587 VP.n1752 a_400_38200# 0.06fF
C8588 VP.n1753 a_400_38200# 0.06fF
C8589 VP.n1754 a_400_38200# 0.06fF
C8590 VP.n1755 a_400_38200# 0.07fF
C8591 VP.n1756 a_400_38200# 0.03fF
C8592 VP.n1757 a_400_38200# 0.05fF
C8593 VP.n1758 a_400_38200# 0.07fF
C8594 VP.n1759 a_400_38200# 0.19fF
C8595 VP.n1760 a_400_38200# 0.60fF
C8596 VP.n1761 a_400_38200# 0.76fF
C8597 VP.n1762 a_400_38200# 0.40fF
C8598 VP.n1763 a_400_38200# 0.03fF
C8599 VP.n1764 a_400_38200# 0.01fF
C8600 VP.t1118 a_400_38200# 0.02fF
C8601 VP.n1765 a_400_38200# 0.25fF
C8602 VP.t985 a_400_38200# 0.02fF
C8603 VP.n1766 a_400_38200# 0.95fF
C8604 VP.n1767 a_400_38200# 0.70fF
C8605 VP.n1768 a_400_38200# 1.93fF
C8606 VP.n1769 a_400_38200# 1.80fF
C8607 VP.n1770 a_400_38200# 2.77fF
C8608 VP.n1771 a_400_38200# 0.83fF
C8609 VP.t976 a_400_38200# 0.02fF
C8610 VP.n1772 a_400_38200# 0.24fF
C8611 VP.n1773 a_400_38200# 0.35fF
C8612 VP.n1774 a_400_38200# 0.60fF
C8613 VP.n1775 a_400_38200# 0.12fF
C8614 VP.t457 a_400_38200# 0.02fF
C8615 VP.n1776 a_400_38200# 0.14fF
C8616 VP.n1778 a_400_38200# 0.04fF
C8617 VP.n1779 a_400_38200# 0.02fF
C8618 VP.n1780 a_400_38200# 0.06fF
C8619 VP.n1781 a_400_38200# 0.30fF
C8620 VP.n1782 a_400_38200# 0.10fF
C8621 VP.n1783 a_400_38200# 0.06fF
C8622 VP.n1784 a_400_38200# 0.06fF
C8623 VP.n1785 a_400_38200# 0.28fF
C8624 VP.n1786 a_400_38200# 0.03fF
C8625 VP.n1787 a_400_38200# 0.15fF
C8626 VP.n1788 a_400_38200# 0.08fF
C8627 VP.n1789 a_400_38200# 0.14fF
C8628 VP.n1790 a_400_38200# 0.03fF
C8629 VP.n1791 a_400_38200# 0.06fF
C8630 VP.n1792 a_400_38200# 0.06fF
C8631 VP.n1793 a_400_38200# 0.06fF
C8632 VP.n1794 a_400_38200# 0.06fF
C8633 VP.n1795 a_400_38200# 0.03fF
C8634 VP.n1796 a_400_38200# 0.05fF
C8635 VP.n1797 a_400_38200# 0.07fF
C8636 VP.n1798 a_400_38200# 0.19fF
C8637 VP.n1799 a_400_38200# 0.59fF
C8638 VP.n1800 a_400_38200# 0.34fF
C8639 VP.n1801 a_400_38200# 1.88fF
C8640 VP.t248 a_400_38200# 0.02fF
C8641 VP.n1802 a_400_38200# 0.24fF
C8642 VP.n1803 a_400_38200# 0.91fF
C8643 VP.n1804 a_400_38200# 0.05fF
C8644 VP.t495 a_400_38200# 0.02fF
C8645 VP.n1805 a_400_38200# 0.12fF
C8646 VP.n1806 a_400_38200# 0.14fF
C8647 VP.n1808 a_400_38200# 0.19fF
C8648 VP.n1809 a_400_38200# 0.10fF
C8649 VP.n1810 a_400_38200# 0.10fF
C8650 VP.n1811 a_400_38200# 0.18fF
C8651 VP.n1812 a_400_38200# 0.09fF
C8652 VP.n1813 a_400_38200# 0.04fF
C8653 VP.n1814 a_400_38200# 0.19fF
C8654 VP.n1815 a_400_38200# 0.26fF
C8655 VP.n1816 a_400_38200# 1.17fF
C8656 VP.n1817 a_400_38200# 0.06fF
C8657 VP.n1818 a_400_38200# 0.44fF
C8658 VP.n1819 a_400_38200# 0.13fF
C8659 VP.n1820 a_400_38200# 0.02fF
C8660 VP.n1821 a_400_38200# 1.81fF
C8661 VP.n1822 a_400_38200# 0.12fF
C8662 VP.t1307 a_400_38200# 0.02fF
C8663 VP.n1823 a_400_38200# 0.14fF
C8664 VP.t594 a_400_38200# 0.02fF
C8665 VP.n1825 a_400_38200# 0.24fF
C8666 VP.n1826 a_400_38200# 0.35fF
C8667 VP.n1827 a_400_38200# 0.60fF
C8668 VP.n1828 a_400_38200# 3.18fF
C8669 VP.n1829 a_400_38200# 2.06fF
C8670 VP.n1830 a_400_38200# 1.98fF
C8671 VP.t1166 a_400_38200# 0.02fF
C8672 VP.n1831 a_400_38200# 0.24fF
C8673 VP.n1832 a_400_38200# 0.91fF
C8674 VP.n1833 a_400_38200# 0.05fF
C8675 VP.t1346 a_400_38200# 0.02fF
C8676 VP.n1834 a_400_38200# 0.12fF
C8677 VP.n1835 a_400_38200# 0.14fF
C8678 VP.n1837 a_400_38200# 0.19fF
C8679 VP.n1838 a_400_38200# 0.03fF
C8680 VP.n1839 a_400_38200# 0.24fF
C8681 VP.n1840 a_400_38200# 0.99fF
C8682 VP.n1841 a_400_38200# 0.12fF
C8683 VP.n1842 a_400_38200# 0.19fF
C8684 VP.n1843 a_400_38200# 0.09fF
C8685 VP.n1844 a_400_38200# 0.18fF
C8686 VP.n1845 a_400_38200# 0.09fF
C8687 VP.n1846 a_400_38200# 0.08fF
C8688 VP.n1847 a_400_38200# 0.39fF
C8689 VP.n1848 a_400_38200# 0.24fF
C8690 VP.n1849 a_400_38200# 0.13fF
C8691 VP.n1850 a_400_38200# 0.02fF
C8692 VP.n1851 a_400_38200# 1.81fF
C8693 VP.n1852 a_400_38200# 0.12fF
C8694 VP.t860 a_400_38200# 0.02fF
C8695 VP.n1853 a_400_38200# 0.14fF
C8696 VP.t128 a_400_38200# 0.02fF
C8697 VP.n1855 a_400_38200# 0.24fF
C8698 VP.n1856 a_400_38200# 0.35fF
C8699 VP.n1857 a_400_38200# 0.60fF
C8700 VP.n1858 a_400_38200# 2.96fF
C8701 VP.n1859 a_400_38200# 2.27fF
C8702 VP.n1860 a_400_38200# 1.98fF
C8703 VP.t715 a_400_38200# 0.02fF
C8704 VP.n1861 a_400_38200# 0.24fF
C8705 VP.n1862 a_400_38200# 0.91fF
C8706 VP.n1863 a_400_38200# 0.05fF
C8707 VP.t899 a_400_38200# 0.02fF
C8708 VP.n1864 a_400_38200# 0.12fF
C8709 VP.n1865 a_400_38200# 0.14fF
C8710 VP.n1867 a_400_38200# 15.28fF
C8711 VP.n1868 a_400_38200# 0.10fF
C8712 VP.n1869 a_400_38200# 0.06fF
C8713 VP.n1870 a_400_38200# 0.06fF
C8714 VP.n1871 a_400_38200# 0.28fF
C8715 VP.n1872 a_400_38200# 0.03fF
C8716 VP.n1873 a_400_38200# 0.15fF
C8717 VP.n1874 a_400_38200# 0.08fF
C8718 VP.n1875 a_400_38200# 0.14fF
C8719 VP.n1876 a_400_38200# 0.03fF
C8720 VP.n1877 a_400_38200# 0.06fF
C8721 VP.n1878 a_400_38200# 0.06fF
C8722 VP.n1879 a_400_38200# 0.06fF
C8723 VP.n1880 a_400_38200# 0.06fF
C8724 VP.n1881 a_400_38200# 0.03fF
C8725 VP.n1882 a_400_38200# 0.05fF
C8726 VP.n1883 a_400_38200# 0.07fF
C8727 VP.n1884 a_400_38200# 0.19fF
C8728 VP.n1885 a_400_38200# 0.59fF
C8729 VP.n1886 a_400_38200# 0.34fF
C8730 VP.n1887 a_400_38200# 0.04fF
C8731 VP.n1888 a_400_38200# 0.02fF
C8732 VP.n1889 a_400_38200# 0.06fF
C8733 VP.n1890 a_400_38200# 0.30fF
C8734 VP.n1891 a_400_38200# 1.93fF
C8735 VP.n1892 a_400_38200# 0.12fF
C8736 VP.t673 a_400_38200# 0.02fF
C8737 VP.n1893 a_400_38200# 0.14fF
C8738 VP.t1265 a_400_38200# 0.02fF
C8739 VP.n1895 a_400_38200# 0.24fF
C8740 VP.n1896 a_400_38200# 0.35fF
C8741 VP.n1897 a_400_38200# 0.60fF
C8742 VP.n1898 a_400_38200# 0.07fF
C8743 VP.n1899 a_400_38200# 0.72fF
C8744 VP.n1900 a_400_38200# 0.20fF
C8745 VP.n1901 a_400_38200# 0.19fF
C8746 VP.n1902 a_400_38200# 0.10fF
C8747 VP.n1903 a_400_38200# 0.11fF
C8748 VP.n1904 a_400_38200# 0.09fF
C8749 VP.n1905 a_400_38200# 0.16fF
C8750 VP.n1906 a_400_38200# 0.10fF
C8751 VP.n1907 a_400_38200# 0.11fF
C8752 VP.n1908 a_400_38200# 0.19fF
C8753 VP.n1909 a_400_38200# 0.20fF
C8754 VP.n1910 a_400_38200# 0.98fF
C8755 VP.n1911 a_400_38200# 0.15fF
C8756 VP.n1913 a_400_38200# 1.72fF
C8757 VP.t703 a_400_38200# 0.02fF
C8758 VP.n1914 a_400_38200# 0.12fF
C8759 VP.n1915 a_400_38200# 0.14fF
C8760 VP.t537 a_400_38200# 0.02fF
C8761 VP.n1917 a_400_38200# 0.24fF
C8762 VP.n1918 a_400_38200# 0.91fF
C8763 VP.n1919 a_400_38200# 0.05fF
C8764 VP.n1920 a_400_38200# 0.10fF
C8765 VP.n1921 a_400_38200# 0.28fF
C8766 VP.n1922 a_400_38200# 0.06fF
C8767 VP.n1923 a_400_38200# 0.06fF
C8768 VP.n1924 a_400_38200# 0.03fF
C8769 VP.n1925 a_400_38200# 0.15fF
C8770 VP.n1926 a_400_38200# 0.08fF
C8771 VP.n1927 a_400_38200# 0.14fF
C8772 VP.n1928 a_400_38200# 0.03fF
C8773 VP.n1929 a_400_38200# 0.06fF
C8774 VP.n1930 a_400_38200# 0.06fF
C8775 VP.n1931 a_400_38200# 0.06fF
C8776 VP.n1932 a_400_38200# 0.06fF
C8777 VP.n1933 a_400_38200# 0.03fF
C8778 VP.n1934 a_400_38200# 0.05fF
C8779 VP.n1935 a_400_38200# 0.07fF
C8780 VP.n1936 a_400_38200# 0.19fF
C8781 VP.n1937 a_400_38200# 0.59fF
C8782 VP.n1938 a_400_38200# 0.34fF
C8783 VP.n1939 a_400_38200# 0.04fF
C8784 VP.n1940 a_400_38200# 0.02fF
C8785 VP.n1941 a_400_38200# 0.06fF
C8786 VP.n1942 a_400_38200# 0.30fF
C8787 VP.n1943 a_400_38200# 1.93fF
C8788 VP.n1944 a_400_38200# 0.12fF
C8789 VP.t227 a_400_38200# 0.02fF
C8790 VP.n1945 a_400_38200# 0.14fF
C8791 VP.t820 a_400_38200# 0.02fF
C8792 VP.n1947 a_400_38200# 0.24fF
C8793 VP.n1948 a_400_38200# 0.35fF
C8794 VP.n1949 a_400_38200# 0.60fF
C8795 VP.n1950 a_400_38200# 0.07fF
C8796 VP.n1951 a_400_38200# 0.72fF
C8797 VP.n1952 a_400_38200# 0.20fF
C8798 VP.n1953 a_400_38200# 0.19fF
C8799 VP.n1954 a_400_38200# 0.10fF
C8800 VP.n1955 a_400_38200# 0.11fF
C8801 VP.n1956 a_400_38200# 0.09fF
C8802 VP.n1957 a_400_38200# 0.16fF
C8803 VP.n1958 a_400_38200# 0.10fF
C8804 VP.n1959 a_400_38200# 0.11fF
C8805 VP.n1960 a_400_38200# 0.19fF
C8806 VP.n1961 a_400_38200# 0.20fF
C8807 VP.n1962 a_400_38200# 0.98fF
C8808 VP.n1963 a_400_38200# 0.15fF
C8809 VP.n1965 a_400_38200# 1.72fF
C8810 VP.t259 a_400_38200# 0.02fF
C8811 VP.n1966 a_400_38200# 0.12fF
C8812 VP.n1967 a_400_38200# 0.14fF
C8813 VP.t61 a_400_38200# 0.02fF
C8814 VP.n1969 a_400_38200# 0.24fF
C8815 VP.n1970 a_400_38200# 0.91fF
C8816 VP.n1971 a_400_38200# 0.05fF
C8817 VP.n1972 a_400_38200# 0.10fF
C8818 VP.n1973 a_400_38200# 0.06fF
C8819 VP.n1974 a_400_38200# 0.06fF
C8820 VP.n1975 a_400_38200# 0.28fF
C8821 VP.n1976 a_400_38200# 0.03fF
C8822 VP.n1977 a_400_38200# 0.15fF
C8823 VP.n1978 a_400_38200# 0.08fF
C8824 VP.n1979 a_400_38200# 0.14fF
C8825 VP.n1980 a_400_38200# 0.03fF
C8826 VP.n1981 a_400_38200# 0.06fF
C8827 VP.n1982 a_400_38200# 0.06fF
C8828 VP.n1983 a_400_38200# 0.06fF
C8829 VP.n1984 a_400_38200# 0.06fF
C8830 VP.n1985 a_400_38200# 0.03fF
C8831 VP.n1986 a_400_38200# 0.05fF
C8832 VP.n1987 a_400_38200# 0.07fF
C8833 VP.n1988 a_400_38200# 0.19fF
C8834 VP.n1989 a_400_38200# 0.59fF
C8835 VP.n1990 a_400_38200# 0.34fF
C8836 VP.n1991 a_400_38200# 0.04fF
C8837 VP.n1992 a_400_38200# 0.02fF
C8838 VP.n1993 a_400_38200# 0.06fF
C8839 VP.n1994 a_400_38200# 0.30fF
C8840 VP.n1995 a_400_38200# 1.93fF
C8841 VP.n1996 a_400_38200# 0.12fF
C8842 VP.t480 a_400_38200# 0.02fF
C8843 VP.n1997 a_400_38200# 0.14fF
C8844 VP.t1066 a_400_38200# 0.02fF
C8845 VP.n1999 a_400_38200# 0.24fF
C8846 VP.n2000 a_400_38200# 0.35fF
C8847 VP.n2001 a_400_38200# 0.60fF
C8848 VP.n2002 a_400_38200# 0.07fF
C8849 VP.n2003 a_400_38200# 0.72fF
C8850 VP.n2004 a_400_38200# 0.20fF
C8851 VP.n2005 a_400_38200# 0.19fF
C8852 VP.n2006 a_400_38200# 0.10fF
C8853 VP.n2007 a_400_38200# 0.11fF
C8854 VP.n2008 a_400_38200# 0.09fF
C8855 VP.n2009 a_400_38200# 0.16fF
C8856 VP.n2010 a_400_38200# 0.10fF
C8857 VP.n2011 a_400_38200# 0.11fF
C8858 VP.n2012 a_400_38200# 0.19fF
C8859 VP.n2013 a_400_38200# 0.20fF
C8860 VP.n2014 a_400_38200# 0.98fF
C8861 VP.n2015 a_400_38200# 0.15fF
C8862 VP.n2017 a_400_38200# 1.72fF
C8863 VP.t1112 a_400_38200# 0.02fF
C8864 VP.n2018 a_400_38200# 0.12fF
C8865 VP.n2019 a_400_38200# 0.14fF
C8866 VP.t347 a_400_38200# 0.02fF
C8867 VP.n2021 a_400_38200# 0.24fF
C8868 VP.n2022 a_400_38200# 0.91fF
C8869 VP.n2023 a_400_38200# 0.05fF
C8870 VP.n2024 a_400_38200# 0.10fF
C8871 VP.n2025 a_400_38200# 0.06fF
C8872 VP.n2026 a_400_38200# 0.06fF
C8873 VP.n2027 a_400_38200# 0.28fF
C8874 VP.n2028 a_400_38200# 0.03fF
C8875 VP.n2029 a_400_38200# 0.15fF
C8876 VP.n2030 a_400_38200# 0.08fF
C8877 VP.n2031 a_400_38200# 0.14fF
C8878 VP.n2032 a_400_38200# 0.03fF
C8879 VP.n2033 a_400_38200# 0.06fF
C8880 VP.n2034 a_400_38200# 0.06fF
C8881 VP.n2035 a_400_38200# 0.06fF
C8882 VP.n2036 a_400_38200# 0.06fF
C8883 VP.n2037 a_400_38200# 0.03fF
C8884 VP.n2038 a_400_38200# 0.05fF
C8885 VP.n2039 a_400_38200# 0.07fF
C8886 VP.n2040 a_400_38200# 0.19fF
C8887 VP.n2041 a_400_38200# 0.59fF
C8888 VP.n2042 a_400_38200# 0.34fF
C8889 VP.n2043 a_400_38200# 0.04fF
C8890 VP.n2044 a_400_38200# 0.02fF
C8891 VP.n2045 a_400_38200# 0.06fF
C8892 VP.n2046 a_400_38200# 0.30fF
C8893 VP.n2047 a_400_38200# 1.93fF
C8894 VP.n2048 a_400_38200# 0.12fF
C8895 VP.t1330 a_400_38200# 0.02fF
C8896 VP.n2049 a_400_38200# 0.14fF
C8897 VP.t620 a_400_38200# 0.02fF
C8898 VP.n2051 a_400_38200# 0.24fF
C8899 VP.n2052 a_400_38200# 0.35fF
C8900 VP.n2053 a_400_38200# 0.60fF
C8901 VP.n2054 a_400_38200# 0.07fF
C8902 VP.n2055 a_400_38200# 0.72fF
C8903 VP.n2056 a_400_38200# 0.20fF
C8904 VP.n2057 a_400_38200# 0.19fF
C8905 VP.n2058 a_400_38200# 0.10fF
C8906 VP.n2059 a_400_38200# 0.11fF
C8907 VP.n2060 a_400_38200# 0.09fF
C8908 VP.n2061 a_400_38200# 0.16fF
C8909 VP.n2062 a_400_38200# 0.10fF
C8910 VP.n2063 a_400_38200# 0.11fF
C8911 VP.n2064 a_400_38200# 0.19fF
C8912 VP.n2065 a_400_38200# 0.20fF
C8913 VP.n2066 a_400_38200# 0.98fF
C8914 VP.n2067 a_400_38200# 0.15fF
C8915 VP.n2069 a_400_38200# 1.72fF
C8916 VP.t102 a_400_38200# 0.02fF
C8917 VP.n2070 a_400_38200# 0.12fF
C8918 VP.n2071 a_400_38200# 0.14fF
C8919 VP.t1196 a_400_38200# 0.02fF
C8920 VP.n2073 a_400_38200# 0.24fF
C8921 VP.n2074 a_400_38200# 0.91fF
C8922 VP.n2075 a_400_38200# 0.05fF
C8923 VP.n2076 a_400_38200# 0.10fF
C8924 VP.n2077 a_400_38200# 0.28fF
C8925 VP.n2078 a_400_38200# 0.06fF
C8926 VP.n2079 a_400_38200# 0.06fF
C8927 VP.n2080 a_400_38200# 0.03fF
C8928 VP.n2081 a_400_38200# 0.15fF
C8929 VP.n2082 a_400_38200# 0.08fF
C8930 VP.n2083 a_400_38200# 0.14fF
C8931 VP.n2084 a_400_38200# 0.03fF
C8932 VP.n2085 a_400_38200# 0.06fF
C8933 VP.n2086 a_400_38200# 0.06fF
C8934 VP.n2087 a_400_38200# 0.06fF
C8935 VP.n2088 a_400_38200# 0.06fF
C8936 VP.n2089 a_400_38200# 0.03fF
C8937 VP.n2090 a_400_38200# 0.05fF
C8938 VP.n2091 a_400_38200# 0.07fF
C8939 VP.n2092 a_400_38200# 0.19fF
C8940 VP.n2093 a_400_38200# 0.59fF
C8941 VP.n2094 a_400_38200# 0.34fF
C8942 VP.n2095 a_400_38200# 0.04fF
C8943 VP.n2096 a_400_38200# 0.02fF
C8944 VP.n2097 a_400_38200# 0.06fF
C8945 VP.n2098 a_400_38200# 0.30fF
C8946 VP.n2099 a_400_38200# 1.93fF
C8947 VP.n2100 a_400_38200# 0.12fF
C8948 VP.t878 a_400_38200# 0.02fF
C8949 VP.n2101 a_400_38200# 0.14fF
C8950 VP.t161 a_400_38200# 0.02fF
C8951 VP.n2103 a_400_38200# 0.24fF
C8952 VP.n2104 a_400_38200# 0.35fF
C8953 VP.n2105 a_400_38200# 0.60fF
C8954 VP.n2106 a_400_38200# 0.72fF
C8955 VP.n2107 a_400_38200# 1.24fF
C8956 VP.n2108 a_400_38200# 0.54fF
C8957 VP.n2109 a_400_38200# 0.22fF
C8958 VP.n2110 a_400_38200# 1.73fF
C8959 VP.t978 a_400_38200# 0.02fF
C8960 VP.n2111 a_400_38200# 0.12fF
C8961 VP.n2112 a_400_38200# 0.14fF
C8962 VP.t743 a_400_38200# 0.02fF
C8963 VP.n2114 a_400_38200# 0.24fF
C8964 VP.n2115 a_400_38200# 0.91fF
C8965 VP.n2116 a_400_38200# 0.05fF
C8966 VP.n2117 a_400_38200# 0.10fF
C8967 VP.n2118 a_400_38200# 0.06fF
C8968 VP.n2119 a_400_38200# 0.06fF
C8969 VP.n2120 a_400_38200# 0.28fF
C8970 VP.n2121 a_400_38200# 0.03fF
C8971 VP.n2122 a_400_38200# 0.15fF
C8972 VP.n2123 a_400_38200# 0.08fF
C8973 VP.n2124 a_400_38200# 0.14fF
C8974 VP.n2125 a_400_38200# 0.03fF
C8975 VP.n2126 a_400_38200# 0.06fF
C8976 VP.n2127 a_400_38200# 0.06fF
C8977 VP.n2128 a_400_38200# 0.06fF
C8978 VP.n2129 a_400_38200# 0.06fF
C8979 VP.n2130 a_400_38200# 0.03fF
C8980 VP.n2131 a_400_38200# 0.05fF
C8981 VP.n2132 a_400_38200# 0.07fF
C8982 VP.n2133 a_400_38200# 0.19fF
C8983 VP.n2134 a_400_38200# 0.59fF
C8984 VP.n2135 a_400_38200# 0.34fF
C8985 VP.n2136 a_400_38200# 0.04fF
C8986 VP.n2137 a_400_38200# 0.02fF
C8987 VP.n2138 a_400_38200# 0.06fF
C8988 VP.n2139 a_400_38200# 0.30fF
C8989 VP.n2140 a_400_38200# 1.93fF
C8990 VP.n2141 a_400_38200# 0.12fF
C8991 VP.t430 a_400_38200# 0.02fF
C8992 VP.n2142 a_400_38200# 0.14fF
C8993 VP.t1012 a_400_38200# 0.02fF
C8994 VP.n2144 a_400_38200# 0.24fF
C8995 VP.n2145 a_400_38200# 0.35fF
C8996 VP.n2146 a_400_38200# 0.60fF
C8997 VP.n2147 a_400_38200# 0.72fF
C8998 VP.n2148 a_400_38200# 1.24fF
C8999 VP.n2149 a_400_38200# 0.54fF
C9000 VP.n2150 a_400_38200# 0.22fF
C9001 VP.n2151 a_400_38200# 1.73fF
C9002 VP.t532 a_400_38200# 0.02fF
C9003 VP.n2152 a_400_38200# 0.12fF
C9004 VP.n2153 a_400_38200# 0.14fF
C9005 VP.t290 a_400_38200# 0.02fF
C9006 VP.n2155 a_400_38200# 0.24fF
C9007 VP.n2156 a_400_38200# 0.91fF
C9008 VP.n2157 a_400_38200# 0.05fF
C9009 VP.n2158 a_400_38200# 0.10fF
C9010 VP.n2159 a_400_38200# 0.06fF
C9011 VP.n2160 a_400_38200# 0.06fF
C9012 VP.n2161 a_400_38200# 0.28fF
C9013 VP.n2162 a_400_38200# 0.03fF
C9014 VP.n2163 a_400_38200# 0.15fF
C9015 VP.n2164 a_400_38200# 0.08fF
C9016 VP.n2165 a_400_38200# 0.14fF
C9017 VP.n2166 a_400_38200# 0.03fF
C9018 VP.n2167 a_400_38200# 0.06fF
C9019 VP.n2168 a_400_38200# 0.06fF
C9020 VP.n2169 a_400_38200# 0.06fF
C9021 VP.n2170 a_400_38200# 0.06fF
C9022 VP.n2171 a_400_38200# 0.03fF
C9023 VP.n2172 a_400_38200# 0.05fF
C9024 VP.n2173 a_400_38200# 0.07fF
C9025 VP.n2174 a_400_38200# 0.19fF
C9026 VP.n2175 a_400_38200# 0.59fF
C9027 VP.n2176 a_400_38200# 0.34fF
C9028 VP.n2177 a_400_38200# 0.04fF
C9029 VP.n2178 a_400_38200# 0.02fF
C9030 VP.n2179 a_400_38200# 0.06fF
C9031 VP.n2180 a_400_38200# 0.30fF
C9032 VP.n2181 a_400_38200# 1.93fF
C9033 VP.n2182 a_400_38200# 0.12fF
C9034 VP.t1285 a_400_38200# 0.02fF
C9035 VP.n2183 a_400_38200# 0.14fF
C9036 VP.t567 a_400_38200# 0.02fF
C9037 VP.n2185 a_400_38200# 0.24fF
C9038 VP.n2186 a_400_38200# 0.35fF
C9039 VP.n2187 a_400_38200# 0.60fF
C9040 VP.n2188 a_400_38200# 0.72fF
C9041 VP.n2189 a_400_38200# 1.24fF
C9042 VP.n2190 a_400_38200# 0.54fF
C9043 VP.n2191 a_400_38200# 0.22fF
C9044 VP.n2192 a_400_38200# 1.73fF
C9045 VP.t54 a_400_38200# 0.02fF
C9046 VP.n2193 a_400_38200# 0.12fF
C9047 VP.n2194 a_400_38200# 0.14fF
C9048 VP.t1141 a_400_38200# 0.02fF
C9049 VP.n2196 a_400_38200# 0.24fF
C9050 VP.n2197 a_400_38200# 0.91fF
C9051 VP.n2198 a_400_38200# 0.05fF
C9052 VP.n2199 a_400_38200# 0.10fF
C9053 VP.n2200 a_400_38200# 0.06fF
C9054 VP.n2201 a_400_38200# 0.06fF
C9055 VP.n2202 a_400_38200# 0.28fF
C9056 VP.n2203 a_400_38200# 0.03fF
C9057 VP.n2204 a_400_38200# 0.15fF
C9058 VP.n2205 a_400_38200# 0.08fF
C9059 VP.n2206 a_400_38200# 0.14fF
C9060 VP.n2207 a_400_38200# 0.03fF
C9061 VP.n2208 a_400_38200# 0.06fF
C9062 VP.n2209 a_400_38200# 0.06fF
C9063 VP.n2210 a_400_38200# 0.06fF
C9064 VP.n2211 a_400_38200# 0.06fF
C9065 VP.n2212 a_400_38200# 0.03fF
C9066 VP.n2213 a_400_38200# 0.05fF
C9067 VP.n2214 a_400_38200# 0.07fF
C9068 VP.n2215 a_400_38200# 0.19fF
C9069 VP.n2216 a_400_38200# 0.59fF
C9070 VP.n2217 a_400_38200# 0.34fF
C9071 VP.n2218 a_400_38200# 0.04fF
C9072 VP.n2219 a_400_38200# 0.02fF
C9073 VP.n2220 a_400_38200# 0.06fF
C9074 VP.n2221 a_400_38200# 0.30fF
C9075 VP.n2222 a_400_38200# 1.93fF
C9076 VP.n2223 a_400_38200# 0.12fF
C9077 VP.t841 a_400_38200# 0.02fF
C9078 VP.n2224 a_400_38200# 0.14fF
C9079 VP.t99 a_400_38200# 0.02fF
C9080 VP.n2226 a_400_38200# 0.24fF
C9081 VP.n2227 a_400_38200# 0.35fF
C9082 VP.n2228 a_400_38200# 0.60fF
C9083 VP.n2229 a_400_38200# 0.71fF
C9084 VP.n2230 a_400_38200# 1.24fF
C9085 VP.n2231 a_400_38200# 0.54fF
C9086 VP.n2232 a_400_38200# 0.21fF
C9087 VP.n2233 a_400_38200# 1.73fF
C9088 VP.t940 a_400_38200# 0.02fF
C9089 VP.n2234 a_400_38200# 0.12fF
C9090 VP.n2235 a_400_38200# 0.14fF
C9091 VP.t692 a_400_38200# 0.02fF
C9092 VP.n2237 a_400_38200# 0.24fF
C9093 VP.n2238 a_400_38200# 0.91fF
C9094 VP.n2239 a_400_38200# 0.05fF
C9095 VP.n2240 a_400_38200# 0.04fF
C9096 VP.n2241 a_400_38200# 0.10fF
C9097 VP.n2242 a_400_38200# 0.59fF
C9098 VP.n2243 a_400_38200# 1.71fF
C9099 VP.n2244 a_400_38200# 0.12fF
C9100 VP.t1104 a_400_38200# 0.02fF
C9101 VP.n2245 a_400_38200# 0.14fF
C9102 VP.t395 a_400_38200# 0.02fF
C9103 VP.n2247 a_400_38200# 0.24fF
C9104 VP.n2248 a_400_38200# 0.35fF
C9105 VP.n2249 a_400_38200# 0.60fF
C9106 VP.n2250 a_400_38200# 0.05fF
C9107 VP.n2251 a_400_38200# 0.71fF
C9108 VP.n2252 a_400_38200# 1.49fF
C9109 VP.n2253 a_400_38200# 0.06fF
C9110 VP.n2254 a_400_38200# 0.19fF
C9111 VP.n2255 a_400_38200# 0.05fF
C9112 VP.n2256 a_400_38200# 0.16fF
C9113 VP.n2257 a_400_38200# 0.10fF
C9114 VP.n2258 a_400_38200# 0.09fF
C9115 VP.n2259 a_400_38200# 0.09fF
C9116 VP.n2260 a_400_38200# 0.14fF
C9117 VP.n2262 a_400_38200# 2.51fF
C9118 VP.n2263 a_400_38200# 1.88fF
C9119 VP.t449 a_400_38200# 0.02fF
C9120 VP.n2264 a_400_38200# 0.12fF
C9121 VP.n2265 a_400_38200# 0.14fF
C9122 VP.t972 a_400_38200# 0.02fF
C9123 VP.n2267 a_400_38200# 0.24fF
C9124 VP.n2268 a_400_38200# 0.91fF
C9125 VP.n2269 a_400_38200# 0.05fF
C9126 VP.t53 a_400_38200# 35.17fF
C9127 VP.t408 a_400_38200# 0.02fF
C9128 VP.n2270 a_400_38200# 1.21fF
C9129 VP.n2271 a_400_38200# 0.25fF
C9130 VP.n2272 a_400_38200# 26.29fF
C9131 VP.n2273 a_400_38200# 26.29fF
C9132 VP.n2274 a_400_38200# 0.76fF
C9133 VP.n2275 a_400_38200# 0.27fF
C9134 VP.n2276 a_400_38200# 0.59fF
C9135 VP.n2277 a_400_38200# 0.10fF
C9136 VP.n2278 a_400_38200# 3.02fF
C9137 VP.t98 a_400_38200# 15.72fF
C9138 VP.n2279 a_400_38200# 1.15fF
C9139 VP.n2281 a_400_38200# 13.70fF
C9140 VP.n2283 a_400_38200# 1.99fF
C9141 VP.n2284 a_400_38200# 4.39fF
C9142 VP.n2285 a_400_38200# 0.03fF
C9143 VP.n2286 a_400_38200# 0.05fF
C9144 VP.n2287 a_400_38200# 0.07fF
C9145 VP.n2288 a_400_38200# 0.03fF
C9146 VP.n2289 a_400_38200# 0.06fF
C9147 VP.n2290 a_400_38200# 0.06fF
C9148 VP.n2291 a_400_38200# 0.06fF
C9149 VP.n2292 a_400_38200# 0.07fF
C9150 VP.n2293 a_400_38200# 0.57fF
C9151 VP.n2294 a_400_38200# 1.88fF
C9152 VP.n2295 a_400_38200# 0.92fF
C9153 VP.n2296 a_400_38200# 2.63fF
C9154 VP.n2297 a_400_38200# 0.10fF
C9155 VP.n2298 a_400_38200# 0.28fF
C9156 VP.n2299 a_400_38200# 0.15fF
C9157 VP.n2300 a_400_38200# 0.08fF
C9158 VP.n2301 a_400_38200# 0.14fF
C9159 VP.n2302 a_400_38200# 0.06fF
C9160 VP.n2303 a_400_38200# 0.06fF
C9161 VP.n2304 a_400_38200# 0.03fF
C9162 VP.n2305 a_400_38200# 0.05fF
C9163 VP.n2306 a_400_38200# 0.07fF
C9164 VP.n2307 a_400_38200# 0.19fF
C9165 VP.n2308 a_400_38200# 0.59fF
C9166 VP.n2309 a_400_38200# 0.34fF
C9167 VP.n2310 a_400_38200# 0.04fF
C9168 VP.n2311 a_400_38200# 0.02fF
C9169 VP.n2312 a_400_38200# 0.06fF
C9170 VP.n2313 a_400_38200# 0.30fF
C9171 VP.n2314 a_400_38200# 0.12fF
C9172 VP.t1288 a_400_38200# 0.02fF
C9173 VP.n2315 a_400_38200# 0.14fF
C9174 VP.n2317 a_400_38200# 0.02fF
C9175 VP.n2318 a_400_38200# 0.32fF
C9176 VP.n2319 a_400_38200# 0.08fF
C9177 VP.n2320 a_400_38200# 0.09fF
C9178 VP.n2321 a_400_38200# 0.05fF
C9179 VP.n2322 a_400_38200# 0.04fF
C9180 VP.n2323 a_400_38200# 0.05fF
C9181 VP.n2324 a_400_38200# 0.04fF
C9182 VP.n2325 a_400_38200# 0.12fF
C9183 VP.n2326 a_400_38200# 0.09fF
C9184 VP.n2327 a_400_38200# 0.14fF
C9185 VP.n2328 a_400_38200# 0.56fF
C9186 VP.n2329 a_400_38200# 0.19fF
C9187 VP.n2330 a_400_38200# 1.93fF
C9188 VP.n2331 a_400_38200# 0.12fF
C9189 VP.t1018 a_400_38200# 0.02fF
C9190 VP.n2332 a_400_38200# 0.14fF
C9191 VP.t310 a_400_38200# 0.02fF
C9192 VP.n2334 a_400_38200# 0.24fF
C9193 VP.n2335 a_400_38200# 0.35fF
C9194 VP.n2336 a_400_38200# 0.60fF
C9195 VP.n2337 a_400_38200# 2.72fF
C9196 VP.n2338 a_400_38200# 2.19fF
C9197 VP.t1183 a_400_38200# 0.02fF
C9198 VP.n2339 a_400_38200# 0.24fF
C9199 VP.n2340 a_400_38200# 0.91fF
C9200 VP.n2341 a_400_38200# 0.05fF
C9201 VP.t115 a_400_38200# 0.02fF
C9202 VP.n2342 a_400_38200# 0.12fF
C9203 VP.n2343 a_400_38200# 0.14fF
C9204 VP.n2345 a_400_38200# 0.10fF
C9205 VP.n2346 a_400_38200# 0.28fF
C9206 VP.n2347 a_400_38200# 0.15fF
C9207 VP.n2348 a_400_38200# 0.08fF
C9208 VP.n2349 a_400_38200# 0.14fF
C9209 VP.n2350 a_400_38200# 0.06fF
C9210 VP.n2351 a_400_38200# 0.06fF
C9211 VP.n2352 a_400_38200# 0.03fF
C9212 VP.n2353 a_400_38200# 0.05fF
C9213 VP.n2354 a_400_38200# 0.07fF
C9214 VP.n2355 a_400_38200# 0.19fF
C9215 VP.n2356 a_400_38200# 0.59fF
C9216 VP.n2357 a_400_38200# 0.34fF
C9217 VP.n2358 a_400_38200# 0.04fF
C9218 VP.n2359 a_400_38200# 0.02fF
C9219 VP.n2360 a_400_38200# 0.06fF
C9220 VP.n2361 a_400_38200# 0.30fF
C9221 VP.n2362 a_400_38200# 1.93fF
C9222 VP.n2363 a_400_38200# 0.12fF
C9223 VP.t216 a_400_38200# 0.02fF
C9224 VP.n2364 a_400_38200# 0.14fF
C9225 VP.t806 a_400_38200# 0.02fF
C9226 VP.n2366 a_400_38200# 0.24fF
C9227 VP.n2367 a_400_38200# 0.35fF
C9228 VP.n2368 a_400_38200# 0.60fF
C9229 VP.n2369 a_400_38200# 2.39fF
C9230 VP.n2370 a_400_38200# 1.79fF
C9231 VP.t373 a_400_38200# 0.02fF
C9232 VP.n2371 a_400_38200# 0.24fF
C9233 VP.n2372 a_400_38200# 0.91fF
C9234 VP.n2373 a_400_38200# 0.05fF
C9235 VP.t562 a_400_38200# 0.02fF
C9236 VP.n2374 a_400_38200# 0.12fF
C9237 VP.n2375 a_400_38200# 0.14fF
C9238 VP.n2377 a_400_38200# 0.10fF
C9239 VP.n2378 a_400_38200# 0.28fF
C9240 VP.n2379 a_400_38200# 0.15fF
C9241 VP.n2380 a_400_38200# 0.08fF
C9242 VP.n2381 a_400_38200# 0.14fF
C9243 VP.n2382 a_400_38200# 0.06fF
C9244 VP.n2383 a_400_38200# 0.06fF
C9245 VP.n2384 a_400_38200# 0.03fF
C9246 VP.n2385 a_400_38200# 0.05fF
C9247 VP.n2386 a_400_38200# 0.07fF
C9248 VP.n2387 a_400_38200# 0.19fF
C9249 VP.n2388 a_400_38200# 0.59fF
C9250 VP.n2389 a_400_38200# 0.34fF
C9251 VP.n2390 a_400_38200# 0.04fF
C9252 VP.n2391 a_400_38200# 0.02fF
C9253 VP.n2392 a_400_38200# 0.06fF
C9254 VP.n2393 a_400_38200# 0.30fF
C9255 VP.n2394 a_400_38200# 1.93fF
C9256 VP.n2395 a_400_38200# 0.12fF
C9257 VP.t663 a_400_38200# 0.02fF
C9258 VP.n2396 a_400_38200# 0.14fF
C9259 VP.t1251 a_400_38200# 0.02fF
C9260 VP.n2398 a_400_38200# 0.24fF
C9261 VP.n2399 a_400_38200# 0.35fF
C9262 VP.n2400 a_400_38200# 0.60fF
C9263 VP.n2401 a_400_38200# 2.47fF
C9264 VP.n2402 a_400_38200# 2.20fF
C9265 VP.t825 a_400_38200# 0.02fF
C9266 VP.n2403 a_400_38200# 0.24fF
C9267 VP.n2404 a_400_38200# 0.91fF
C9268 VP.n2405 a_400_38200# 0.05fF
C9269 VP.t1005 a_400_38200# 0.02fF
C9270 VP.n2406 a_400_38200# 0.12fF
C9271 VP.n2407 a_400_38200# 0.14fF
C9272 VP.n2409 a_400_38200# 0.10fF
C9273 VP.n2410 a_400_38200# 0.28fF
C9274 VP.n2411 a_400_38200# 0.15fF
C9275 VP.n2412 a_400_38200# 0.08fF
C9276 VP.n2413 a_400_38200# 0.14fF
C9277 VP.n2414 a_400_38200# 0.06fF
C9278 VP.n2415 a_400_38200# 0.06fF
C9279 VP.n2416 a_400_38200# 0.03fF
C9280 VP.n2417 a_400_38200# 0.05fF
C9281 VP.n2418 a_400_38200# 0.07fF
C9282 VP.n2419 a_400_38200# 0.19fF
C9283 VP.n2420 a_400_38200# 0.59fF
C9284 VP.n2421 a_400_38200# 0.34fF
C9285 VP.n2422 a_400_38200# 0.04fF
C9286 VP.n2423 a_400_38200# 0.02fF
C9287 VP.n2424 a_400_38200# 0.06fF
C9288 VP.n2425 a_400_38200# 0.30fF
C9289 VP.n2426 a_400_38200# 1.93fF
C9290 VP.n2427 a_400_38200# 0.12fF
C9291 VP.t1106 a_400_38200# 0.02fF
C9292 VP.n2428 a_400_38200# 0.14fF
C9293 VP.t396 a_400_38200# 0.02fF
C9294 VP.n2430 a_400_38200# 0.24fF
C9295 VP.n2431 a_400_38200# 0.35fF
C9296 VP.n2432 a_400_38200# 0.60fF
C9297 VP.n2433 a_400_38200# 2.47fF
C9298 VP.n2434 a_400_38200# 2.20fF
C9299 VP.t1271 a_400_38200# 0.02fF
C9300 VP.n2435 a_400_38200# 0.24fF
C9301 VP.n2436 a_400_38200# 0.91fF
C9302 VP.n2437 a_400_38200# 0.05fF
C9303 VP.t146 a_400_38200# 0.02fF
C9304 VP.n2438 a_400_38200# 0.12fF
C9305 VP.n2439 a_400_38200# 0.14fF
C9306 VP.n2441 a_400_38200# 0.10fF
C9307 VP.n2442 a_400_38200# 0.28fF
C9308 VP.n2443 a_400_38200# 0.15fF
C9309 VP.n2444 a_400_38200# 0.08fF
C9310 VP.n2445 a_400_38200# 0.14fF
C9311 VP.n2446 a_400_38200# 0.06fF
C9312 VP.n2447 a_400_38200# 0.06fF
C9313 VP.n2448 a_400_38200# 0.03fF
C9314 VP.n2449 a_400_38200# 0.05fF
C9315 VP.n2450 a_400_38200# 0.07fF
C9316 VP.n2451 a_400_38200# 0.19fF
C9317 VP.n2452 a_400_38200# 0.59fF
C9318 VP.n2453 a_400_38200# 0.34fF
C9319 VP.n2454 a_400_38200# 0.04fF
C9320 VP.n2455 a_400_38200# 0.02fF
C9321 VP.n2456 a_400_38200# 0.06fF
C9322 VP.n2457 a_400_38200# 0.30fF
C9323 VP.n2458 a_400_38200# 1.93fF
C9324 VP.n2459 a_400_38200# 0.12fF
C9325 VP.t252 a_400_38200# 0.02fF
C9326 VP.n2460 a_400_38200# 0.14fF
C9327 VP.t846 a_400_38200# 0.02fF
C9328 VP.n2462 a_400_38200# 0.24fF
C9329 VP.n2463 a_400_38200# 0.35fF
C9330 VP.n2464 a_400_38200# 0.60fF
C9331 VP.n2465 a_400_38200# 2.47fF
C9332 VP.n2466 a_400_38200# 2.20fF
C9333 VP.t416 a_400_38200# 0.02fF
C9334 VP.n2467 a_400_38200# 0.24fF
C9335 VP.n2468 a_400_38200# 0.91fF
C9336 VP.n2469 a_400_38200# 0.05fF
C9337 VP.t611 a_400_38200# 0.02fF
C9338 VP.n2470 a_400_38200# 0.12fF
C9339 VP.n2471 a_400_38200# 0.14fF
C9340 VP.n2473 a_400_38200# 0.10fF
C9341 VP.n2474 a_400_38200# 0.28fF
C9342 VP.n2475 a_400_38200# 0.15fF
C9343 VP.n2476 a_400_38200# 0.08fF
C9344 VP.n2477 a_400_38200# 0.14fF
C9345 VP.n2478 a_400_38200# 0.06fF
C9346 VP.n2479 a_400_38200# 0.06fF
C9347 VP.n2480 a_400_38200# 0.03fF
C9348 VP.n2481 a_400_38200# 0.05fF
C9349 VP.n2482 a_400_38200# 0.07fF
C9350 VP.n2483 a_400_38200# 0.19fF
C9351 VP.n2484 a_400_38200# 0.59fF
C9352 VP.n2485 a_400_38200# 0.34fF
C9353 VP.n2486 a_400_38200# 0.04fF
C9354 VP.n2487 a_400_38200# 0.02fF
C9355 VP.n2488 a_400_38200# 0.06fF
C9356 VP.n2489 a_400_38200# 0.30fF
C9357 VP.n2490 a_400_38200# 1.93fF
C9358 VP.n2491 a_400_38200# 0.12fF
C9359 VP.t697 a_400_38200# 0.02fF
C9360 VP.n2492 a_400_38200# 0.14fF
C9361 VP.t1232 a_400_38200# 0.02fF
C9362 VP.n2494 a_400_38200# 0.24fF
C9363 VP.n2495 a_400_38200# 0.35fF
C9364 VP.n2496 a_400_38200# 0.60fF
C9365 VP.n2497 a_400_38200# 0.07fF
C9366 VP.n2498 a_400_38200# 0.72fF
C9367 VP.n2499 a_400_38200# 0.09fF
C9368 VP.n2500 a_400_38200# 0.16fF
C9369 VP.n2501 a_400_38200# 0.98fF
C9370 VP.n2502 a_400_38200# 0.15fF
C9371 VP.n2504 a_400_38200# 1.72fF
C9372 VP.t803 a_400_38200# 0.02fF
C9373 VP.n2505 a_400_38200# 0.24fF
C9374 VP.n2506 a_400_38200# 0.91fF
C9375 VP.n2507 a_400_38200# 0.05fF
C9376 VP.t1058 a_400_38200# 0.02fF
C9377 VP.n2508 a_400_38200# 0.12fF
C9378 VP.n2509 a_400_38200# 0.14fF
C9379 VP.n2511 a_400_38200# 0.10fF
C9380 VP.n2512 a_400_38200# 0.28fF
C9381 VP.n2513 a_400_38200# 0.15fF
C9382 VP.n2514 a_400_38200# 0.08fF
C9383 VP.n2515 a_400_38200# 0.14fF
C9384 VP.n2516 a_400_38200# 0.06fF
C9385 VP.n2517 a_400_38200# 0.06fF
C9386 VP.n2518 a_400_38200# 0.03fF
C9387 VP.n2519 a_400_38200# 0.05fF
C9388 VP.n2520 a_400_38200# 0.07fF
C9389 VP.n2521 a_400_38200# 0.19fF
C9390 VP.n2522 a_400_38200# 0.59fF
C9391 VP.n2523 a_400_38200# 0.34fF
C9392 VP.n2524 a_400_38200# 0.04fF
C9393 VP.n2525 a_400_38200# 0.02fF
C9394 VP.n2526 a_400_38200# 0.06fF
C9395 VP.n2527 a_400_38200# 0.30fF
C9396 VP.n2528 a_400_38200# 1.93fF
C9397 VP.n2529 a_400_38200# 0.12fF
C9398 VP.t392 a_400_38200# 0.02fF
C9399 VP.n2530 a_400_38200# 0.14fF
C9400 VP.t977 a_400_38200# 0.02fF
C9401 VP.n2532 a_400_38200# 0.24fF
C9402 VP.n2533 a_400_38200# 0.35fF
C9403 VP.n2534 a_400_38200# 0.60fF
C9404 VP.n2535 a_400_38200# 0.07fF
C9405 VP.n2536 a_400_38200# 0.72fF
C9406 VP.n2537 a_400_38200# 0.09fF
C9407 VP.n2538 a_400_38200# 0.16fF
C9408 VP.n2539 a_400_38200# 0.98fF
C9409 VP.n2540 a_400_38200# 0.15fF
C9410 VP.n2542 a_400_38200# 1.72fF
C9411 VP.t550 a_400_38200# 0.02fF
C9412 VP.n2543 a_400_38200# 0.24fF
C9413 VP.n2544 a_400_38200# 0.91fF
C9414 VP.n2545 a_400_38200# 0.05fF
C9415 VP.t811 a_400_38200# 0.02fF
C9416 VP.n2546 a_400_38200# 0.12fF
C9417 VP.n2547 a_400_38200# 0.14fF
C9418 VP.n2549 a_400_38200# 0.10fF
C9419 VP.n2550 a_400_38200# 0.28fF
C9420 VP.n2551 a_400_38200# 0.15fF
C9421 VP.n2552 a_400_38200# 0.08fF
C9422 VP.n2553 a_400_38200# 0.14fF
C9423 VP.n2554 a_400_38200# 0.06fF
C9424 VP.n2555 a_400_38200# 0.06fF
C9425 VP.n2556 a_400_38200# 0.03fF
C9426 VP.n2557 a_400_38200# 0.05fF
C9427 VP.n2558 a_400_38200# 0.07fF
C9428 VP.n2559 a_400_38200# 0.19fF
C9429 VP.n2560 a_400_38200# 0.59fF
C9430 VP.n2561 a_400_38200# 0.34fF
C9431 VP.n2562 a_400_38200# 0.04fF
C9432 VP.n2563 a_400_38200# 0.02fF
C9433 VP.n2564 a_400_38200# 0.06fF
C9434 VP.n2565 a_400_38200# 0.30fF
C9435 VP.n2566 a_400_38200# 1.93fF
C9436 VP.n2567 a_400_38200# 0.12fF
C9437 VP.t844 a_400_38200# 0.02fF
C9438 VP.n2568 a_400_38200# 0.14fF
C9439 VP.t101 a_400_38200# 0.02fF
C9440 VP.n2570 a_400_38200# 0.24fF
C9441 VP.n2571 a_400_38200# 0.35fF
C9442 VP.n2572 a_400_38200# 0.60fF
C9443 VP.n2573 a_400_38200# 0.07fF
C9444 VP.n2574 a_400_38200# 0.72fF
C9445 VP.n2575 a_400_38200# 0.09fF
C9446 VP.n2576 a_400_38200# 0.16fF
C9447 VP.n2577 a_400_38200# 0.98fF
C9448 VP.n2578 a_400_38200# 0.15fF
C9449 VP.n2580 a_400_38200# 1.72fF
C9450 VP.t994 a_400_38200# 0.02fF
C9451 VP.n2581 a_400_38200# 0.24fF
C9452 VP.n2582 a_400_38200# 0.91fF
C9453 VP.n2583 a_400_38200# 0.05fF
C9454 VP.t1255 a_400_38200# 0.02fF
C9455 VP.n2584 a_400_38200# 0.12fF
C9456 VP.n2585 a_400_38200# 0.14fF
C9457 VP.n2587 a_400_38200# 15.28fF
C9458 VP.t103 a_400_38200# 0.02fF
C9459 VP.n2588 a_400_38200# 0.95fF
C9460 VP.n2589 a_400_38200# 0.70fF
C9461 VP.t558 a_400_38200# 0.02fF
C9462 VP.n2590 a_400_38200# 1.21fF
C9463 VP.n2591 a_400_38200# 0.31fF
C9464 VP.n2592 a_400_38200# 0.04fF
C9465 VP.n2593 a_400_38200# 0.88fF
C9466 VP.n2594 a_400_38200# 0.48fF
C9467 VP.n2595 a_400_38200# 0.88fF
C9468 VP.n2596 a_400_38200# 0.60fF
C9469 VP.n2597 a_400_38200# 2.33fF
C9470 VP.n2598 a_400_38200# 0.59fF
C9471 VP.n2599 a_400_38200# 0.02fF
C9472 VP.n2600 a_400_38200# 0.96fF
C9473 VP.t60 a_400_38200# 15.72fF
C9474 VP.n2601 a_400_38200# 15.42fF
C9475 VP.n2603 a_400_38200# 0.38fF
C9476 VP.n2604 a_400_38200# 0.23fF
C9477 VP.n2605 a_400_38200# 3.28fF
C9478 VP.n2606 a_400_38200# 1.42fF
C9479 VP.n2607 a_400_38200# 0.16fF
C9480 VP.n2608 a_400_38200# 2.20fF
C9481 VP.n2609 a_400_38200# 3.70fF
C9482 VP.n2610 a_400_38200# 0.25fF
C9483 VP.n2611 a_400_38200# 0.06fF
C9484 VP.n2612 a_400_38200# 0.09fF
C9485 VP.n2613 a_400_38200# 0.09fF
C9486 VP.n2614 a_400_38200# 0.43fF
C9487 VP.n2615 a_400_38200# 0.69fF
C9488 VP.n2616 a_400_38200# 0.14fF
C9489 VP.n2617 a_400_38200# 0.07fF
C9490 VP.n2618 a_400_38200# 0.72fF
C9491 VP.n2619 a_400_38200# 1.81fF
C9492 VP.n2620 a_400_38200# 0.12fF
C9493 VP.t166 a_400_38200# 0.02fF
C9494 VP.n2621 a_400_38200# 0.14fF
C9495 VP.t764 a_400_38200# 0.02fF
C9496 VP.n2623 a_400_38200# 0.24fF
C9497 VP.n2624 a_400_38200# 0.35fF
C9498 VP.n2625 a_400_38200# 0.60fF
C9499 VP.n2626 a_400_38200# 2.30fF
C9500 VP.t582 a_400_38200# 0.02fF
C9501 VP.n2627 a_400_38200# 0.12fF
C9502 VP.n2628 a_400_38200# 0.14fF
C9503 VP.t337 a_400_38200# 0.02fF
C9504 VP.n2630 a_400_38200# 0.24fF
C9505 VP.n2631 a_400_38200# 0.91fF
C9506 VP.n2632 a_400_38200# 0.05fF
C9507 VP.n2633 a_400_38200# 0.10fF
C9508 VP.n2634 a_400_38200# 0.10fF
C9509 VP.n2635 a_400_38200# 0.18fF
C9510 VP.n2636 a_400_38200# 0.09fF
C9511 VP.n2637 a_400_38200# 0.04fF
C9512 VP.n2638 a_400_38200# 0.26fF
C9513 VP.n2639 a_400_38200# 1.17fF
C9514 VP.n2640 a_400_38200# 0.06fF
C9515 VP.n2641 a_400_38200# 0.44fF
C9516 VP.n2642 a_400_38200# 0.13fF
C9517 VP.n2643 a_400_38200# 0.02fF
C9518 VP.n2644 a_400_38200# 1.81fF
C9519 VP.n2645 a_400_38200# 0.12fF
C9520 VP.t626 a_400_38200# 0.02fF
C9521 VP.n2646 a_400_38200# 0.14fF
C9522 VP.t1211 a_400_38200# 0.02fF
C9523 VP.n2648 a_400_38200# 0.24fF
C9524 VP.n2649 a_400_38200# 0.35fF
C9525 VP.n2650 a_400_38200# 0.60fF
C9526 VP.n2651 a_400_38200# 2.28fF
C9527 VP.t1030 a_400_38200# 0.02fF
C9528 VP.n2652 a_400_38200# 0.12fF
C9529 VP.n2653 a_400_38200# 0.14fF
C9530 VP.t785 a_400_38200# 0.02fF
C9531 VP.n2655 a_400_38200# 0.24fF
C9532 VP.n2656 a_400_38200# 0.91fF
C9533 VP.n2657 a_400_38200# 0.05fF
C9534 VP.n2658 a_400_38200# 1.93fF
C9535 VP.t357 a_400_38200# 0.02fF
C9536 VP.n2659 a_400_38200# 0.24fF
C9537 VP.n2660 a_400_38200# 0.35fF
C9538 VP.n2661 a_400_38200# 0.60fF
C9539 VP.n2662 a_400_38200# 0.12fF
C9540 VP.t1071 a_400_38200# 0.02fF
C9541 VP.n2663 a_400_38200# 0.14fF
C9542 VP.n2665 a_400_38200# 0.04fF
C9543 VP.n2666 a_400_38200# 0.02fF
C9544 VP.n2667 a_400_38200# 0.06fF
C9545 VP.n2668 a_400_38200# 0.30fF
C9546 VP.n2669 a_400_38200# 0.10fF
C9547 VP.n2670 a_400_38200# 0.28fF
C9548 VP.n2671 a_400_38200# 0.15fF
C9549 VP.n2672 a_400_38200# 0.08fF
C9550 VP.n2673 a_400_38200# 0.14fF
C9551 VP.n2674 a_400_38200# 0.06fF
C9552 VP.n2675 a_400_38200# 0.06fF
C9553 VP.n2676 a_400_38200# 0.03fF
C9554 VP.n2677 a_400_38200# 0.05fF
C9555 VP.n2678 a_400_38200# 0.07fF
C9556 VP.n2679 a_400_38200# 0.19fF
C9557 VP.n2680 a_400_38200# 0.59fF
C9558 VP.n2681 a_400_38200# 0.34fF
C9559 VP.n2682 a_400_38200# 2.18fF
C9560 VP.t92 a_400_38200# 0.02fF
C9561 VP.n2683 a_400_38200# 0.12fF
C9562 VP.n2684 a_400_38200# 0.14fF
C9563 VP.t1229 a_400_38200# 0.02fF
C9564 VP.n2686 a_400_38200# 0.24fF
C9565 VP.n2687 a_400_38200# 0.91fF
C9566 VP.n2688 a_400_38200# 0.05fF
C9567 VP.t385 a_400_38200# 0.02fF
C9568 VP.n2689 a_400_38200# 0.01fF
C9569 VP.n2690 a_400_38200# 0.26fF
C9570 VP.t91 a_400_38200# 35.17fF
C9571 VP.t398 a_400_38200# 0.02fF
C9572 VP.n2691 a_400_38200# 0.12fF
C9573 VP.n2692 a_400_38200# 0.14fF
C9574 VP.t124 a_400_38200# 0.02fF
C9575 VP.n2694 a_400_38200# 0.24fF
C9576 VP.n2695 a_400_38200# 0.91fF
C9577 VP.n2696 a_400_38200# 0.05fF
C9578 VP.t570 a_400_38200# 0.02fF
C9579 VP.n2697 a_400_38200# 0.24fF
C9580 VP.n2698 a_400_38200# 0.35fF
C9581 VP.n2699 a_400_38200# 0.60fF
C9582 VP.n2700 a_400_38200# 0.04fF
C9583 VP.n2701 a_400_38200# 0.08fF
C9584 VP.n2702 a_400_38200# 0.72fF
C9585 VP.n2703 a_400_38200# 0.09fF
C9586 VP.n2704 a_400_38200# 0.00fF
C9587 VP.n2705 a_400_38200# 0.98fF
C9588 VP.n2706 a_400_38200# 0.19fF
C9589 VP.n2708 a_400_38200# 1.72fF
C9590 VP.n2709 a_400_38200# 1.96fF
C9591 VP.n2710 a_400_38200# 1.04fF
C9592 VP.n2711 a_400_38200# 0.05fF
C9593 VP.n2712 a_400_38200# 0.03fF
C9594 VP.n2713 a_400_38200# 0.06fF
C9595 VP.n2714 a_400_38200# 0.06fF
C9596 VP.n2715 a_400_38200# 0.06fF
C9597 VP.n2716 a_400_38200# 0.07fF
C9598 VP.n2717 a_400_38200# 0.03fF
C9599 VP.n2718 a_400_38200# 0.05fF
C9600 VP.n2719 a_400_38200# 0.07fF
C9601 VP.n2720 a_400_38200# 0.19fF
C9602 VP.n2721 a_400_38200# 0.60fF
C9603 VP.n2722 a_400_38200# 0.76fF
C9604 VP.n2723 a_400_38200# 0.40fF
C9605 VP.n2724 a_400_38200# 0.03fF
C9606 VP.n2725 a_400_38200# 0.01fF
C9607 VP.t1274 a_400_38200# 0.02fF
C9608 VP.n2726 a_400_38200# 0.25fF
C9609 VP.t1128 a_400_38200# 0.02fF
C9610 VP.n2727 a_400_38200# 0.95fF
C9611 VP.n2728 a_400_38200# 0.70fF
C9612 VP.n2729 a_400_38200# 1.93fF
C9613 VP.n2730 a_400_38200# 2.96fF
C9614 VP.n2731 a_400_38200# 2.27fF
C9615 VP.t263 a_400_38200# 0.02fF
C9616 VP.n2732 a_400_38200# 0.24fF
C9617 VP.n2733 a_400_38200# 0.35fF
C9618 VP.n2734 a_400_38200# 0.60fF
C9619 VP.n2735 a_400_38200# 0.12fF
C9620 VP.t983 a_400_38200# 0.02fF
C9621 VP.n2736 a_400_38200# 0.14fF
C9622 VP.n2738 a_400_38200# 0.04fF
C9623 VP.n2739 a_400_38200# 0.02fF
C9624 VP.n2740 a_400_38200# 0.06fF
C9625 VP.n2741 a_400_38200# 0.30fF
C9626 VP.n2742 a_400_38200# 0.10fF
C9627 VP.n2743 a_400_38200# 0.28fF
C9628 VP.n2744 a_400_38200# 0.06fF
C9629 VP.n2745 a_400_38200# 0.06fF
C9630 VP.n2746 a_400_38200# 0.03fF
C9631 VP.n2747 a_400_38200# 0.15fF
C9632 VP.n2748 a_400_38200# 0.08fF
C9633 VP.n2749 a_400_38200# 0.14fF
C9634 VP.n2750 a_400_38200# 0.03fF
C9635 VP.n2751 a_400_38200# 0.06fF
C9636 VP.n2752 a_400_38200# 0.06fF
C9637 VP.n2753 a_400_38200# 0.06fF
C9638 VP.n2754 a_400_38200# 0.06fF
C9639 VP.n2755 a_400_38200# 0.03fF
C9640 VP.n2756 a_400_38200# 0.05fF
C9641 VP.n2757 a_400_38200# 0.07fF
C9642 VP.n2758 a_400_38200# 0.19fF
C9643 VP.n2759 a_400_38200# 0.59fF
C9644 VP.n2760 a_400_38200# 0.34fF
C9645 VP.n2761 a_400_38200# 1.88fF
C9646 VP.t850 a_400_38200# 0.02fF
C9647 VP.n2762 a_400_38200# 0.24fF
C9648 VP.n2763 a_400_38200# 0.91fF
C9649 VP.n2764 a_400_38200# 0.05fF
C9650 VP.t1085 a_400_38200# 0.02fF
C9651 VP.n2765 a_400_38200# 0.12fF
C9652 VP.n2766 a_400_38200# 0.14fF
C9653 VP.n2768 a_400_38200# 0.19fF
C9654 VP.n2769 a_400_38200# 0.10fF
C9655 VP.n2770 a_400_38200# 0.10fF
C9656 VP.n2771 a_400_38200# 0.18fF
C9657 VP.n2772 a_400_38200# 0.09fF
C9658 VP.n2773 a_400_38200# 0.04fF
C9659 VP.n2774 a_400_38200# 0.19fF
C9660 VP.n2775 a_400_38200# 0.26fF
C9661 VP.n2776 a_400_38200# 1.17fF
C9662 VP.n2777 a_400_38200# 0.06fF
C9663 VP.n2778 a_400_38200# 0.44fF
C9664 VP.n2779 a_400_38200# 0.13fF
C9665 VP.n2780 a_400_38200# 0.02fF
C9666 VP.n2781 a_400_38200# 1.81fF
C9667 VP.n2782 a_400_38200# 0.12fF
C9668 VP.t608 a_400_38200# 0.02fF
C9669 VP.n2783 a_400_38200# 0.14fF
C9670 VP.t1120 a_400_38200# 0.02fF
C9671 VP.n2785 a_400_38200# 0.24fF
C9672 VP.n2786 a_400_38200# 0.35fF
C9673 VP.n2787 a_400_38200# 0.60fF
C9674 VP.n2788 a_400_38200# 3.18fF
C9675 VP.n2789 a_400_38200# 2.06fF
C9676 VP.n2790 a_400_38200# 1.98fF
C9677 VP.t400 a_400_38200# 0.02fF
C9678 VP.n2791 a_400_38200# 0.24fF
C9679 VP.n2792 a_400_38200# 0.91fF
C9680 VP.n2793 a_400_38200# 0.05fF
C9681 VP.t642 a_400_38200# 0.02fF
C9682 VP.n2794 a_400_38200# 0.12fF
C9683 VP.n2795 a_400_38200# 0.14fF
C9684 VP.n2797 a_400_38200# 0.16fF
C9685 VP.n2798 a_400_38200# 0.19fF
C9686 VP.n2799 a_400_38200# 0.09fF
C9687 VP.n2800 a_400_38200# 0.04fF
C9688 VP.n2801 a_400_38200# 0.14fF
C9689 VP.n2802 a_400_38200# 0.64fF
C9690 VP.n2803 a_400_38200# 1.32fF
C9691 VP.n2804 a_400_38200# 1.81fF
C9692 VP.n2805 a_400_38200# 0.12fF
C9693 VP.t142 a_400_38200# 0.02fF
C9694 VP.n2806 a_400_38200# 0.14fF
C9695 VP.t740 a_400_38200# 0.02fF
C9696 VP.n2808 a_400_38200# 0.24fF
C9697 VP.n2809 a_400_38200# 0.35fF
C9698 VP.n2810 a_400_38200# 0.60fF
C9699 VP.n2811 a_400_38200# 2.97fF
C9700 VP.n2812 a_400_38200# 2.27fF
C9701 VP.n2813 a_400_38200# 2.00fF
C9702 VP.t1319 a_400_38200# 0.02fF
C9703 VP.n2814 a_400_38200# 0.24fF
C9704 VP.n2815 a_400_38200# 0.91fF
C9705 VP.n2816 a_400_38200# 0.05fF
C9706 VP.t192 a_400_38200# 0.02fF
C9707 VP.n2817 a_400_38200# 0.12fF
C9708 VP.n2818 a_400_38200# 0.14fF
C9709 VP.n2820 a_400_38200# 0.24fF
C9710 VP.t1114 a_400_38200# 0.02fF
C9711 VP.n2821 a_400_38200# 0.36fF
C9712 VP.n2822 a_400_38200# 0.36fF
C9713 VP.n2823 a_400_38200# 0.67fF
C9714 VP.n2824 a_400_38200# 0.11fF
C9715 VP.n2825 a_400_38200# 1.52fF
C9716 VP.n2826 a_400_38200# 0.05fF
C9717 VP.n2827 a_400_38200# 0.06fF
C9718 VP.n2828 a_400_38200# 0.22fF
C9719 VP.n2829 a_400_38200# 0.14fF
C9720 VP.n2830 a_400_38200# 0.28fF
C9721 VP.n2831 a_400_38200# 0.15fF
C9722 VP.n2832 a_400_38200# 0.39fF
C9723 VP.n2833 a_400_38200# 1.27fF
C9724 VP.n2834 a_400_38200# 2.05fF
C9725 VP.n2835 a_400_38200# 2.75fF
C9726 VP.n2836 a_400_38200# 0.75fF
C9727 VP.n2837 a_400_38200# 0.24fF
C9728 VP.t541 a_400_38200# 0.02fF
C9729 VP.n2838 a_400_38200# 0.35fF
C9730 VP.n2839 a_400_38200# 0.63fF
C9731 VP.n2840 a_400_38200# 0.40fF
C9732 VP.n2841 a_400_38200# 0.40fF
C9733 VP.n2842 a_400_38200# 0.12fF
C9734 VP.t1259 a_400_38200# 0.02fF
C9735 VP.n2843 a_400_38200# 0.14fF
C9736 VP.t596 a_400_38200# 0.02fF
C9737 VP.n2845 a_400_38200# 0.12fF
C9738 VP.n2846 a_400_38200# 0.14fF
C9739 VP.n2848 a_400_38200# 15.28fF
C9740 VP.n2849 a_400_38200# 0.10fF
C9741 VP.n2850 a_400_38200# 0.28fF
C9742 VP.n2851 a_400_38200# 0.06fF
C9743 VP.n2852 a_400_38200# 0.06fF
C9744 VP.n2853 a_400_38200# 0.03fF
C9745 VP.n2854 a_400_38200# 0.15fF
C9746 VP.n2855 a_400_38200# 0.08fF
C9747 VP.n2856 a_400_38200# 0.14fF
C9748 VP.n2857 a_400_38200# 0.03fF
C9749 VP.n2858 a_400_38200# 0.06fF
C9750 VP.n2859 a_400_38200# 0.06fF
C9751 VP.n2860 a_400_38200# 0.06fF
C9752 VP.n2861 a_400_38200# 0.06fF
C9753 VP.n2862 a_400_38200# 0.03fF
C9754 VP.n2863 a_400_38200# 0.05fF
C9755 VP.n2864 a_400_38200# 0.07fF
C9756 VP.n2865 a_400_38200# 0.19fF
C9757 VP.n2866 a_400_38200# 0.59fF
C9758 VP.n2867 a_400_38200# 0.34fF
C9759 VP.n2868 a_400_38200# 0.04fF
C9760 VP.n2869 a_400_38200# 0.02fF
C9761 VP.n2870 a_400_38200# 0.06fF
C9762 VP.n2871 a_400_38200# 0.30fF
C9763 VP.n2872 a_400_38200# 1.93fF
C9764 VP.n2873 a_400_38200# 0.12fF
C9765 VP.t829 a_400_38200# 0.02fF
C9766 VP.n2874 a_400_38200# 0.14fF
C9767 VP.t84 a_400_38200# 0.02fF
C9768 VP.n2876 a_400_38200# 0.24fF
C9769 VP.n2877 a_400_38200# 0.35fF
C9770 VP.n2878 a_400_38200# 0.60fF
C9771 VP.n2879 a_400_38200# 0.07fF
C9772 VP.n2880 a_400_38200# 0.72fF
C9773 VP.n2881 a_400_38200# 0.20fF
C9774 VP.n2882 a_400_38200# 0.19fF
C9775 VP.n2883 a_400_38200# 0.10fF
C9776 VP.n2884 a_400_38200# 0.11fF
C9777 VP.n2885 a_400_38200# 0.09fF
C9778 VP.n2886 a_400_38200# 0.16fF
C9779 VP.n2887 a_400_38200# 0.10fF
C9780 VP.n2888 a_400_38200# 0.11fF
C9781 VP.n2889 a_400_38200# 0.19fF
C9782 VP.n2890 a_400_38200# 0.20fF
C9783 VP.n2891 a_400_38200# 0.98fF
C9784 VP.n2892 a_400_38200# 0.15fF
C9785 VP.n2894 a_400_38200# 1.72fF
C9786 VP.t858 a_400_38200# 0.02fF
C9787 VP.n2895 a_400_38200# 0.12fF
C9788 VP.n2896 a_400_38200# 0.14fF
C9789 VP.t681 a_400_38200# 0.02fF
C9790 VP.n2898 a_400_38200# 0.24fF
C9791 VP.n2899 a_400_38200# 0.91fF
C9792 VP.n2900 a_400_38200# 0.05fF
C9793 VP.n2901 a_400_38200# 0.10fF
C9794 VP.n2902 a_400_38200# 0.28fF
C9795 VP.n2903 a_400_38200# 0.06fF
C9796 VP.n2904 a_400_38200# 0.06fF
C9797 VP.n2905 a_400_38200# 0.03fF
C9798 VP.n2906 a_400_38200# 0.15fF
C9799 VP.n2907 a_400_38200# 0.08fF
C9800 VP.n2908 a_400_38200# 0.14fF
C9801 VP.n2909 a_400_38200# 0.03fF
C9802 VP.n2910 a_400_38200# 0.06fF
C9803 VP.n2911 a_400_38200# 0.06fF
C9804 VP.n2912 a_400_38200# 0.06fF
C9805 VP.n2913 a_400_38200# 0.06fF
C9806 VP.n2914 a_400_38200# 0.03fF
C9807 VP.n2915 a_400_38200# 0.05fF
C9808 VP.n2916 a_400_38200# 0.07fF
C9809 VP.n2917 a_400_38200# 0.19fF
C9810 VP.n2918 a_400_38200# 0.59fF
C9811 VP.n2919 a_400_38200# 0.34fF
C9812 VP.n2920 a_400_38200# 0.04fF
C9813 VP.n2921 a_400_38200# 0.02fF
C9814 VP.n2922 a_400_38200# 0.06fF
C9815 VP.n2923 a_400_38200# 0.30fF
C9816 VP.n2924 a_400_38200# 1.93fF
C9817 VP.n2925 a_400_38200# 0.12fF
C9818 VP.t377 a_400_38200# 0.02fF
C9819 VP.n2926 a_400_38200# 0.14fF
C9820 VP.t963 a_400_38200# 0.02fF
C9821 VP.n2928 a_400_38200# 0.24fF
C9822 VP.n2929 a_400_38200# 0.35fF
C9823 VP.n2930 a_400_38200# 0.60fF
C9824 VP.n2931 a_400_38200# 0.07fF
C9825 VP.n2932 a_400_38200# 0.72fF
C9826 VP.n2933 a_400_38200# 0.20fF
C9827 VP.n2934 a_400_38200# 0.19fF
C9828 VP.n2935 a_400_38200# 0.10fF
C9829 VP.n2936 a_400_38200# 0.11fF
C9830 VP.n2937 a_400_38200# 0.09fF
C9831 VP.n2938 a_400_38200# 0.16fF
C9832 VP.n2939 a_400_38200# 0.10fF
C9833 VP.n2940 a_400_38200# 0.11fF
C9834 VP.n2941 a_400_38200# 0.19fF
C9835 VP.n2942 a_400_38200# 0.20fF
C9836 VP.n2943 a_400_38200# 0.98fF
C9837 VP.n2944 a_400_38200# 0.15fF
C9838 VP.n2946 a_400_38200# 1.72fF
C9839 VP.t411 a_400_38200# 0.02fF
C9840 VP.n2947 a_400_38200# 0.12fF
C9841 VP.n2948 a_400_38200# 0.14fF
C9842 VP.t238 a_400_38200# 0.02fF
C9843 VP.n2950 a_400_38200# 0.24fF
C9844 VP.n2951 a_400_38200# 0.91fF
C9845 VP.n2952 a_400_38200# 0.05fF
C9846 VP.n2953 a_400_38200# 0.10fF
C9847 VP.n2954 a_400_38200# 0.28fF
C9848 VP.n2955 a_400_38200# 0.06fF
C9849 VP.n2956 a_400_38200# 0.06fF
C9850 VP.n2957 a_400_38200# 0.03fF
C9851 VP.n2958 a_400_38200# 0.15fF
C9852 VP.n2959 a_400_38200# 0.08fF
C9853 VP.n2960 a_400_38200# 0.14fF
C9854 VP.n2961 a_400_38200# 0.03fF
C9855 VP.n2962 a_400_38200# 0.06fF
C9856 VP.n2963 a_400_38200# 0.06fF
C9857 VP.n2964 a_400_38200# 0.06fF
C9858 VP.n2965 a_400_38200# 0.06fF
C9859 VP.n2966 a_400_38200# 0.03fF
C9860 VP.n2967 a_400_38200# 0.05fF
C9861 VP.n2968 a_400_38200# 0.07fF
C9862 VP.n2969 a_400_38200# 0.19fF
C9863 VP.n2970 a_400_38200# 0.59fF
C9864 VP.n2971 a_400_38200# 0.34fF
C9865 VP.n2972 a_400_38200# 0.04fF
C9866 VP.n2973 a_400_38200# 0.02fF
C9867 VP.n2974 a_400_38200# 0.06fF
C9868 VP.n2975 a_400_38200# 0.30fF
C9869 VP.n2976 a_400_38200# 1.93fF
C9870 VP.n2977 a_400_38200# 0.12fF
C9871 VP.t630 a_400_38200# 0.02fF
C9872 VP.n2978 a_400_38200# 0.14fF
C9873 VP.t1215 a_400_38200# 0.02fF
C9874 VP.n2980 a_400_38200# 0.24fF
C9875 VP.n2981 a_400_38200# 0.35fF
C9876 VP.n2982 a_400_38200# 0.60fF
C9877 VP.n2983 a_400_38200# 0.07fF
C9878 VP.n2984 a_400_38200# 0.72fF
C9879 VP.n2985 a_400_38200# 0.20fF
C9880 VP.n2986 a_400_38200# 0.19fF
C9881 VP.n2987 a_400_38200# 0.10fF
C9882 VP.n2988 a_400_38200# 0.11fF
C9883 VP.n2989 a_400_38200# 0.09fF
C9884 VP.n2990 a_400_38200# 0.16fF
C9885 VP.n2991 a_400_38200# 0.10fF
C9886 VP.n2992 a_400_38200# 0.11fF
C9887 VP.n2993 a_400_38200# 0.19fF
C9888 VP.n2994 a_400_38200# 0.20fF
C9889 VP.n2995 a_400_38200# 0.98fF
C9890 VP.n2996 a_400_38200# 0.15fF
C9891 VP.n2998 a_400_38200# 1.72fF
C9892 VP.t1267 a_400_38200# 0.02fF
C9893 VP.n2999 a_400_38200# 0.12fF
C9894 VP.n3000 a_400_38200# 0.14fF
C9895 VP.t492 a_400_38200# 0.02fF
C9896 VP.n3002 a_400_38200# 0.24fF
C9897 VP.n3003 a_400_38200# 0.91fF
C9898 VP.n3004 a_400_38200# 0.05fF
C9899 VP.n3005 a_400_38200# 0.10fF
C9900 VP.n3006 a_400_38200# 0.28fF
C9901 VP.n3007 a_400_38200# 0.06fF
C9902 VP.n3008 a_400_38200# 0.06fF
C9903 VP.n3009 a_400_38200# 0.03fF
C9904 VP.n3010 a_400_38200# 0.15fF
C9905 VP.n3011 a_400_38200# 0.08fF
C9906 VP.n3012 a_400_38200# 0.14fF
C9907 VP.n3013 a_400_38200# 0.03fF
C9908 VP.n3014 a_400_38200# 0.06fF
C9909 VP.n3015 a_400_38200# 0.06fF
C9910 VP.n3016 a_400_38200# 0.06fF
C9911 VP.n3017 a_400_38200# 0.06fF
C9912 VP.n3018 a_400_38200# 0.03fF
C9913 VP.n3019 a_400_38200# 0.05fF
C9914 VP.n3020 a_400_38200# 0.07fF
C9915 VP.n3021 a_400_38200# 0.19fF
C9916 VP.n3022 a_400_38200# 0.59fF
C9917 VP.n3023 a_400_38200# 0.34fF
C9918 VP.n3024 a_400_38200# 0.04fF
C9919 VP.n3025 a_400_38200# 0.02fF
C9920 VP.n3026 a_400_38200# 0.06fF
C9921 VP.n3027 a_400_38200# 0.30fF
C9922 VP.n3028 a_400_38200# 1.93fF
C9923 VP.n3029 a_400_38200# 0.12fF
C9924 VP.t174 a_400_38200# 0.02fF
C9925 VP.n3030 a_400_38200# 0.14fF
C9926 VP.t768 a_400_38200# 0.02fF
C9927 VP.n3032 a_400_38200# 0.24fF
C9928 VP.n3033 a_400_38200# 0.35fF
C9929 VP.n3034 a_400_38200# 0.60fF
C9930 VP.n3035 a_400_38200# 0.72fF
C9931 VP.n3036 a_400_38200# 1.24fF
C9932 VP.n3037 a_400_38200# 0.54fF
C9933 VP.n3038 a_400_38200# 0.22fF
C9934 VP.n3039 a_400_38200# 1.73fF
C9935 VP.t268 a_400_38200# 0.02fF
C9936 VP.n3040 a_400_38200# 0.12fF
C9937 VP.n3041 a_400_38200# 0.14fF
C9938 VP.t1342 a_400_38200# 0.02fF
C9939 VP.n3043 a_400_38200# 0.24fF
C9940 VP.n3044 a_400_38200# 0.91fF
C9941 VP.n3045 a_400_38200# 0.05fF
C9942 VP.n3046 a_400_38200# 0.10fF
C9943 VP.n3047 a_400_38200# 0.28fF
C9944 VP.n3048 a_400_38200# 0.06fF
C9945 VP.n3049 a_400_38200# 0.06fF
C9946 VP.n3050 a_400_38200# 0.03fF
C9947 VP.n3051 a_400_38200# 0.15fF
C9948 VP.n3052 a_400_38200# 0.08fF
C9949 VP.n3053 a_400_38200# 0.14fF
C9950 VP.n3054 a_400_38200# 0.03fF
C9951 VP.n3055 a_400_38200# 0.06fF
C9952 VP.n3056 a_400_38200# 0.06fF
C9953 VP.n3057 a_400_38200# 0.06fF
C9954 VP.n3058 a_400_38200# 0.06fF
C9955 VP.n3059 a_400_38200# 0.03fF
C9956 VP.n3060 a_400_38200# 0.05fF
C9957 VP.n3061 a_400_38200# 0.07fF
C9958 VP.n3062 a_400_38200# 0.19fF
C9959 VP.n3063 a_400_38200# 0.59fF
C9960 VP.n3064 a_400_38200# 0.34fF
C9961 VP.n3065 a_400_38200# 0.04fF
C9962 VP.n3066 a_400_38200# 0.02fF
C9963 VP.n3067 a_400_38200# 0.06fF
C9964 VP.n3068 a_400_38200# 0.30fF
C9965 VP.n3069 a_400_38200# 1.93fF
C9966 VP.n3070 a_400_38200# 0.12fF
C9967 VP.t1024 a_400_38200# 0.02fF
C9968 VP.n3071 a_400_38200# 0.14fF
C9969 VP.t315 a_400_38200# 0.02fF
C9970 VP.n3073 a_400_38200# 0.24fF
C9971 VP.n3074 a_400_38200# 0.35fF
C9972 VP.n3075 a_400_38200# 0.60fF
C9973 VP.n3076 a_400_38200# 0.72fF
C9974 VP.n3077 a_400_38200# 1.24fF
C9975 VP.n3078 a_400_38200# 0.54fF
C9976 VP.n3079 a_400_38200# 0.22fF
C9977 VP.n3080 a_400_38200# 1.73fF
C9978 VP.t1124 a_400_38200# 0.02fF
C9979 VP.n3081 a_400_38200# 0.12fF
C9980 VP.n3082 a_400_38200# 0.14fF
C9981 VP.t893 a_400_38200# 0.02fF
C9982 VP.n3084 a_400_38200# 0.24fF
C9983 VP.n3085 a_400_38200# 0.91fF
C9984 VP.n3086 a_400_38200# 0.05fF
C9985 VP.n3087 a_400_38200# 0.10fF
C9986 VP.n3088 a_400_38200# 0.28fF
C9987 VP.n3089 a_400_38200# 0.06fF
C9988 VP.n3090 a_400_38200# 0.06fF
C9989 VP.n3091 a_400_38200# 0.03fF
C9990 VP.n3092 a_400_38200# 0.15fF
C9991 VP.n3093 a_400_38200# 0.08fF
C9992 VP.n3094 a_400_38200# 0.14fF
C9993 VP.n3095 a_400_38200# 0.03fF
C9994 VP.n3096 a_400_38200# 0.06fF
C9995 VP.n3097 a_400_38200# 0.06fF
C9996 VP.n3098 a_400_38200# 0.06fF
C9997 VP.n3099 a_400_38200# 0.06fF
C9998 VP.n3100 a_400_38200# 0.03fF
C9999 VP.n3101 a_400_38200# 0.05fF
C10000 VP.n3102 a_400_38200# 0.07fF
C10001 VP.n3103 a_400_38200# 0.19fF
C10002 VP.n3104 a_400_38200# 0.59fF
C10003 VP.n3105 a_400_38200# 0.34fF
C10004 VP.n3106 a_400_38200# 0.04fF
C10005 VP.n3107 a_400_38200# 0.02fF
C10006 VP.n3108 a_400_38200# 0.06fF
C10007 VP.n3109 a_400_38200# 0.30fF
C10008 VP.n3110 a_400_38200# 1.93fF
C10009 VP.n3111 a_400_38200# 0.12fF
C10010 VP.t576 a_400_38200# 0.02fF
C10011 VP.n3112 a_400_38200# 0.14fF
C10012 VP.t1158 a_400_38200# 0.02fF
C10013 VP.n3114 a_400_38200# 0.24fF
C10014 VP.n3115 a_400_38200# 0.35fF
C10015 VP.n3116 a_400_38200# 0.60fF
C10016 VP.n3117 a_400_38200# 0.72fF
C10017 VP.n3118 a_400_38200# 1.24fF
C10018 VP.n3119 a_400_38200# 0.54fF
C10019 VP.n3120 a_400_38200# 0.22fF
C10020 VP.n3121 a_400_38200# 1.73fF
C10021 VP.t677 a_400_38200# 0.02fF
C10022 VP.n3122 a_400_38200# 0.12fF
C10023 VP.n3123 a_400_38200# 0.14fF
C10024 VP.t442 a_400_38200# 0.02fF
C10025 VP.n3125 a_400_38200# 0.24fF
C10026 VP.n3126 a_400_38200# 0.91fF
C10027 VP.n3127 a_400_38200# 0.05fF
C10028 VP.n3128 a_400_38200# 0.10fF
C10029 VP.n3129 a_400_38200# 0.28fF
C10030 VP.n3130 a_400_38200# 0.06fF
C10031 VP.n3131 a_400_38200# 0.06fF
C10032 VP.n3132 a_400_38200# 0.03fF
C10033 VP.n3133 a_400_38200# 0.15fF
C10034 VP.n3134 a_400_38200# 0.08fF
C10035 VP.n3135 a_400_38200# 0.14fF
C10036 VP.n3136 a_400_38200# 0.03fF
C10037 VP.n3137 a_400_38200# 0.06fF
C10038 VP.n3138 a_400_38200# 0.06fF
C10039 VP.n3139 a_400_38200# 0.06fF
C10040 VP.n3140 a_400_38200# 0.06fF
C10041 VP.n3141 a_400_38200# 0.03fF
C10042 VP.n3142 a_400_38200# 0.05fF
C10043 VP.n3143 a_400_38200# 0.07fF
C10044 VP.n3144 a_400_38200# 0.19fF
C10045 VP.n3145 a_400_38200# 0.59fF
C10046 VP.n3146 a_400_38200# 0.34fF
C10047 VP.n3147 a_400_38200# 0.04fF
C10048 VP.n3148 a_400_38200# 0.02fF
C10049 VP.n3149 a_400_38200# 0.06fF
C10050 VP.n3150 a_400_38200# 0.30fF
C10051 VP.n3151 a_400_38200# 1.93fF
C10052 VP.n3152 a_400_38200# 0.12fF
C10053 VP.t109 a_400_38200# 0.02fF
C10054 VP.n3153 a_400_38200# 0.14fF
C10055 VP.t708 a_400_38200# 0.02fF
C10056 VP.n3155 a_400_38200# 0.24fF
C10057 VP.n3156 a_400_38200# 0.35fF
C10058 VP.n3157 a_400_38200# 0.60fF
C10059 VP.n3158 a_400_38200# 0.71fF
C10060 VP.n3159 a_400_38200# 1.39fF
C10061 VP.n3160 a_400_38200# 0.54fF
C10062 VP.n3161 a_400_38200# 0.21fF
C10063 VP.n3162 a_400_38200# 1.73fF
C10064 VP.t230 a_400_38200# 0.02fF
C10065 VP.n3163 a_400_38200# 0.12fF
C10066 VP.n3164 a_400_38200# 0.14fF
C10067 VP.t1296 a_400_38200# 0.02fF
C10068 VP.n3166 a_400_38200# 0.24fF
C10069 VP.n3167 a_400_38200# 0.91fF
C10070 VP.n3168 a_400_38200# 0.05fF
C10071 VP.n3169 a_400_38200# 0.06fF
C10072 VP.n3170 a_400_38200# 0.06fF
C10073 VP.n3171 a_400_38200# 0.03fF
C10074 VP.n3172 a_400_38200# 0.10fF
C10075 VP.n3173 a_400_38200# 0.17fF
C10076 VP.n3174 a_400_38200# 0.10fF
C10077 VP.n3175 a_400_38200# 0.13fF
C10078 VP.n3176 a_400_38200# 0.02fF
C10079 VP.n3177 a_400_38200# 0.04fF
C10080 VP.n3178 a_400_38200# 0.06fF
C10081 VP.n3179 a_400_38200# 0.05fF
C10082 VP.n3180 a_400_38200# 0.03fF
C10083 VP.n3181 a_400_38200# 0.04fF
C10084 VP.n3182 a_400_38200# 0.20fF
C10085 VP.n3183 a_400_38200# 0.17fF
C10086 VP.n3184 a_400_38200# 0.04fF
C10087 VP.n3185 a_400_38200# 0.02fF
C10088 VP.n3186 a_400_38200# 0.03fF
C10089 VP.n3187 a_400_38200# 0.03fF
C10090 VP.n3188 a_400_38200# 0.14fF
C10091 VP.n3189 a_400_38200# 0.02fF
C10092 VP.n3190 a_400_38200# 0.07fF
C10093 VP.n3191 a_400_38200# 0.13fF
C10094 VP.n3192 a_400_38200# 0.55fF
C10095 VP.n3193 a_400_38200# 0.10fF
C10096 VP.n3194 a_400_38200# 1.93fF
C10097 VP.n3195 a_400_38200# 0.12fF
C10098 VP.t1003 a_400_38200# 0.02fF
C10099 VP.n3196 a_400_38200# 0.14fF
C10100 VP.t288 a_400_38200# 0.02fF
C10101 VP.n3198 a_400_38200# 0.24fF
C10102 VP.n3199 a_400_38200# 0.35fF
C10103 VP.n3200 a_400_38200# 0.60fF
C10104 VP.n3201 a_400_38200# 0.18fF
C10105 VP.n3202 a_400_38200# 0.45fF
C10106 VP.n3203 a_400_38200# 0.06fF
C10107 VP.n3204 a_400_38200# 0.01fF
C10108 VP.n3205 a_400_38200# 0.01fF
C10109 VP.n3206 a_400_38200# 0.04fF
C10110 VP.n3207 a_400_38200# 0.02fF
C10111 VP.n3208 a_400_38200# 0.07fF
C10112 VP.n3209 a_400_38200# 0.04fF
C10113 VP.n3210 a_400_38200# 0.14fF
C10114 VP.n3211 a_400_38200# 0.53fF
C10115 VP.n3212 a_400_38200# 1.62fF
C10116 VP.n3213 a_400_38200# 1.95fF
C10117 VP.t1047 a_400_38200# 0.02fF
C10118 VP.n3214 a_400_38200# 0.12fF
C10119 VP.n3215 a_400_38200# 0.14fF
C10120 VP.t869 a_400_38200# 0.02fF
C10121 VP.n3217 a_400_38200# 0.24fF
C10122 VP.n3218 a_400_38200# 0.91fF
C10123 VP.n3219 a_400_38200# 0.05fF
C10124 VP.t108 a_400_38200# 35.17fF
C10125 VP.t556 a_400_38200# 0.02fF
C10126 VP.n3220 a_400_38200# 1.21fF
C10127 VP.n3221 a_400_38200# 0.25fF
C10128 VP.n3222 a_400_38200# 26.29fF
C10129 VP.n3223 a_400_38200# 26.29fF
C10130 VP.n3224 a_400_38200# 0.76fF
C10131 VP.n3225 a_400_38200# 0.27fF
C10132 VP.n3226 a_400_38200# 0.59fF
C10133 VP.n3227 a_400_38200# 0.10fF
C10134 VP.n3228 a_400_38200# 3.02fF
C10135 VP.t83 a_400_38200# 15.72fF
C10136 VP.n3229 a_400_38200# 1.15fF
C10137 VP.n3231 a_400_38200# 13.70fF
C10138 VP.n3233 a_400_38200# 1.99fF
C10139 VP.n3234 a_400_38200# 4.39fF
C10140 VP.n3235 a_400_38200# 0.03fF
C10141 VP.n3236 a_400_38200# 0.05fF
C10142 VP.n3237 a_400_38200# 0.07fF
C10143 VP.n3238 a_400_38200# 0.03fF
C10144 VP.n3239 a_400_38200# 0.06fF
C10145 VP.n3240 a_400_38200# 0.06fF
C10146 VP.n3241 a_400_38200# 0.06fF
C10147 VP.n3242 a_400_38200# 0.07fF
C10148 VP.n3243 a_400_38200# 0.57fF
C10149 VP.n3244 a_400_38200# 1.88fF
C10150 VP.n3245 a_400_38200# 0.92fF
C10151 VP.n3246 a_400_38200# 2.63fF
C10152 VP.n3247 a_400_38200# 0.10fF
C10153 VP.n3248 a_400_38200# 0.28fF
C10154 VP.n3249 a_400_38200# 0.15fF
C10155 VP.n3250 a_400_38200# 0.08fF
C10156 VP.n3251 a_400_38200# 0.14fF
C10157 VP.n3252 a_400_38200# 0.06fF
C10158 VP.n3253 a_400_38200# 0.06fF
C10159 VP.n3254 a_400_38200# 0.03fF
C10160 VP.n3255 a_400_38200# 0.05fF
C10161 VP.n3256 a_400_38200# 0.07fF
C10162 VP.n3257 a_400_38200# 0.19fF
C10163 VP.n3258 a_400_38200# 0.59fF
C10164 VP.n3259 a_400_38200# 0.34fF
C10165 VP.n3260 a_400_38200# 0.04fF
C10166 VP.n3261 a_400_38200# 0.02fF
C10167 VP.n3262 a_400_38200# 0.06fF
C10168 VP.n3263 a_400_38200# 0.30fF
C10169 VP.n3264 a_400_38200# 0.12fF
C10170 VP.t113 a_400_38200# 0.02fF
C10171 VP.n3265 a_400_38200# 0.14fF
C10172 VP.n3267 a_400_38200# 1.93fF
C10173 VP.t949 a_400_38200# 0.02fF
C10174 VP.n3268 a_400_38200# 0.24fF
C10175 VP.n3269 a_400_38200# 0.35fF
C10176 VP.n3270 a_400_38200# 0.60fF
C10177 VP.n3271 a_400_38200# 0.12fF
C10178 VP.t366 a_400_38200# 0.02fF
C10179 VP.n3272 a_400_38200# 0.14fF
C10180 VP.n3274 a_400_38200# 0.04fF
C10181 VP.n3275 a_400_38200# 0.02fF
C10182 VP.n3276 a_400_38200# 0.06fF
C10183 VP.n3277 a_400_38200# 0.30fF
C10184 VP.n3278 a_400_38200# 0.10fF
C10185 VP.n3279 a_400_38200# 0.28fF
C10186 VP.n3280 a_400_38200# 0.15fF
C10187 VP.n3281 a_400_38200# 0.08fF
C10188 VP.n3282 a_400_38200# 0.14fF
C10189 VP.n3283 a_400_38200# 0.06fF
C10190 VP.n3284 a_400_38200# 0.06fF
C10191 VP.n3285 a_400_38200# 0.03fF
C10192 VP.n3286 a_400_38200# 0.05fF
C10193 VP.n3287 a_400_38200# 0.07fF
C10194 VP.n3288 a_400_38200# 0.19fF
C10195 VP.n3289 a_400_38200# 0.59fF
C10196 VP.n3290 a_400_38200# 0.34fF
C10197 VP.n3291 a_400_38200# 2.18fF
C10198 VP.t518 a_400_38200# 0.02fF
C10199 VP.n3292 a_400_38200# 0.24fF
C10200 VP.n3293 a_400_38200# 0.91fF
C10201 VP.n3294 a_400_38200# 0.05fF
C10202 VP.t701 a_400_38200# 0.02fF
C10203 VP.n3295 a_400_38200# 0.12fF
C10204 VP.n3296 a_400_38200# 0.14fF
C10205 VP.n3298 a_400_38200# 0.10fF
C10206 VP.n3299 a_400_38200# 0.10fF
C10207 VP.n3300 a_400_38200# 0.18fF
C10208 VP.n3301 a_400_38200# 0.09fF
C10209 VP.n3302 a_400_38200# 0.04fF
C10210 VP.n3303 a_400_38200# 0.26fF
C10211 VP.n3304 a_400_38200# 1.17fF
C10212 VP.n3305 a_400_38200# 0.06fF
C10213 VP.n3306 a_400_38200# 0.44fF
C10214 VP.n3307 a_400_38200# 0.13fF
C10215 VP.n3308 a_400_38200# 0.02fF
C10216 VP.n3309 a_400_38200# 1.81fF
C10217 VP.n3310 a_400_38200# 0.12fF
C10218 VP.t1221 a_400_38200# 0.02fF
C10219 VP.n3311 a_400_38200# 0.14fF
C10220 VP.t503 a_400_38200# 0.02fF
C10221 VP.n3313 a_400_38200# 0.24fF
C10222 VP.n3314 a_400_38200# 0.35fF
C10223 VP.n3315 a_400_38200# 0.60fF
C10224 VP.n3316 a_400_38200# 2.28fF
C10225 VP.t38 a_400_38200# 0.02fF
C10226 VP.n3317 a_400_38200# 0.24fF
C10227 VP.n3318 a_400_38200# 0.91fF
C10228 VP.n3319 a_400_38200# 0.05fF
C10229 VP.t258 a_400_38200# 0.02fF
C10230 VP.n3320 a_400_38200# 0.12fF
C10231 VP.n3321 a_400_38200# 0.14fF
C10232 VP.n3323 a_400_38200# 0.06fF
C10233 VP.n3324 a_400_38200# 0.09fF
C10234 VP.n3325 a_400_38200# 0.09fF
C10235 VP.n3326 a_400_38200# 1.45fF
C10236 VP.n3327 a_400_38200# 0.14fF
C10237 VP.n3328 a_400_38200# 0.07fF
C10238 VP.n3329 a_400_38200# 0.72fF
C10239 VP.n3330 a_400_38200# 1.81fF
C10240 VP.n3331 a_400_38200# 0.12fF
C10241 VP.t774 a_400_38200# 0.02fF
C10242 VP.n3332 a_400_38200# 0.14fF
C10243 VP.t13 a_400_38200# 0.02fF
C10244 VP.n3334 a_400_38200# 0.24fF
C10245 VP.n3335 a_400_38200# 0.35fF
C10246 VP.n3336 a_400_38200# 0.60fF
C10247 VP.n3337 a_400_38200# 2.30fF
C10248 VP.t929 a_400_38200# 0.02fF
C10249 VP.n3338 a_400_38200# 0.24fF
C10250 VP.n3339 a_400_38200# 0.91fF
C10251 VP.n3340 a_400_38200# 0.05fF
C10252 VP.t1179 a_400_38200# 0.02fF
C10253 VP.n3341 a_400_38200# 0.12fF
C10254 VP.n3342 a_400_38200# 0.14fF
C10255 VP.n3344 a_400_38200# 0.06fF
C10256 VP.n3345 a_400_38200# 0.25fF
C10257 VP.n3346 a_400_38200# 0.45fF
C10258 VP.n3347 a_400_38200# 0.03fF
C10259 VP.n3348 a_400_38200# 0.05fF
C10260 VP.n3349 a_400_38200# 0.07fF
C10261 VP.n3350 a_400_38200# 0.06fF
C10262 VP.n3351 a_400_38200# 0.06fF
C10263 VP.n3352 a_400_38200# 0.19fF
C10264 VP.n3353 a_400_38200# 0.59fF
C10265 VP.n3354 a_400_38200# 0.34fF
C10266 VP.n3355 a_400_38200# 0.05fF
C10267 VP.n3356 a_400_38200# 0.30fF
C10268 VP.n3357 a_400_38200# 1.93fF
C10269 VP.n3358 a_400_38200# 0.12fF
C10270 VP.t323 a_400_38200# 0.02fF
C10271 VP.n3359 a_400_38200# 0.14fF
C10272 VP.t914 a_400_38200# 0.02fF
C10273 VP.n3361 a_400_38200# 0.24fF
C10274 VP.n3362 a_400_38200# 0.35fF
C10275 VP.n3363 a_400_38200# 0.60fF
C10276 VP.n3364 a_400_38200# 2.04fF
C10277 VP.t484 a_400_38200# 0.02fF
C10278 VP.n3365 a_400_38200# 0.24fF
C10279 VP.n3366 a_400_38200# 0.91fF
C10280 VP.n3367 a_400_38200# 0.05fF
C10281 VP.t727 a_400_38200# 0.02fF
C10282 VP.n3368 a_400_38200# 0.12fF
C10283 VP.n3369 a_400_38200# 0.14fF
C10284 VP.n3371 a_400_38200# 0.24fF
C10285 VP.t1332 a_400_38200# 0.02fF
C10286 VP.n3372 a_400_38200# 0.36fF
C10287 VP.n3373 a_400_38200# 0.36fF
C10288 VP.n3374 a_400_38200# 0.67fF
C10289 VP.n3375 a_400_38200# 0.06fF
C10290 VP.n3376 a_400_38200# 0.11fF
C10291 VP.n3377 a_400_38200# 0.03fF
C10292 VP.n3378 a_400_38200# 0.09fF
C10293 VP.n3379 a_400_38200# 0.05fF
C10294 VP.n3380 a_400_38200# 0.11fF
C10295 VP.n3381 a_400_38200# 0.09fF
C10296 VP.n3382 a_400_38200# 0.09fF
C10297 VP.n3383 a_400_38200# 0.02fF
C10298 VP.n3384 a_400_38200# 0.46fF
C10299 VP.n3385 a_400_38200# 1.81fF
C10300 VP.n3386 a_400_38200# 1.19fF
C10301 VP.n3387 a_400_38200# 0.24fF
C10302 VP.t463 a_400_38200# 0.02fF
C10303 VP.n3388 a_400_38200# 0.35fF
C10304 VP.n3389 a_400_38200# 0.63fF
C10305 VP.n3390 a_400_38200# 0.40fF
C10306 VP.n3391 a_400_38200# 0.40fF
C10307 VP.n3392 a_400_38200# 0.12fF
C10308 VP.t1167 a_400_38200# 0.02fF
C10309 VP.n3393 a_400_38200# 0.14fF
C10310 VP.t277 a_400_38200# 0.02fF
C10311 VP.n3395 a_400_38200# 0.12fF
C10312 VP.n3396 a_400_38200# 0.14fF
C10313 VP.n3398 a_400_38200# 0.88fF
C10314 VP.n3399 a_400_38200# 0.48fF
C10315 VP.n3400 a_400_38200# 0.88fF
C10316 VP.n3401 a_400_38200# 0.60fF
C10317 VP.n3402 a_400_38200# 2.33fF
C10318 VP.n3403 a_400_38200# 0.59fF
C10319 VP.n3404 a_400_38200# 0.02fF
C10320 VP.n3405 a_400_38200# 0.96fF
C10321 VP.t12 a_400_38200# 15.72fF
C10322 VP.n3406 a_400_38200# 15.42fF
C10323 VP.n3408 a_400_38200# 0.38fF
C10324 VP.n3409 a_400_38200# 0.23fF
C10325 VP.n3410 a_400_38200# 3.42fF
C10326 VP.n3411 a_400_38200# 0.21fF
C10327 VP.n3412 a_400_38200# 1.08fF
C10328 VP.n3413 a_400_38200# 0.03fF
C10329 VP.n3414 a_400_38200# 0.09fF
C10330 VP.n3415 a_400_38200# 0.43fF
C10331 VP.n3416 a_400_38200# 0.37fF
C10332 VP.t698 a_400_38200# 0.02fF
C10333 VP.n3417 a_400_38200# 0.64fF
C10334 VP.n3418 a_400_38200# 0.60fF
C10335 VP.n3419 a_400_38200# 2.32fF
C10336 VP.n3420 a_400_38200# 4.93fF
C10337 VP.t269 a_400_38200# 0.02fF
C10338 VP.n3421 a_400_38200# 1.19fF
C10339 VP.n3422 a_400_38200# 0.05fF
C10340 VP.t530 a_400_38200# 0.02fF
C10341 VP.n3423 a_400_38200# 0.01fF
C10342 VP.n3424 a_400_38200# 0.26fF
C10343 VP.n3426 a_400_38200# 15.28fF
C10344 VP.n3427 a_400_38200# 0.10fF
C10345 VP.n3428 a_400_38200# 0.28fF
C10346 VP.n3429 a_400_38200# 0.15fF
C10347 VP.n3430 a_400_38200# 0.08fF
C10348 VP.n3431 a_400_38200# 0.14fF
C10349 VP.n3432 a_400_38200# 0.06fF
C10350 VP.n3433 a_400_38200# 0.06fF
C10351 VP.n3434 a_400_38200# 0.03fF
C10352 VP.n3435 a_400_38200# 0.05fF
C10353 VP.n3436 a_400_38200# 0.07fF
C10354 VP.n3437 a_400_38200# 0.19fF
C10355 VP.n3438 a_400_38200# 0.59fF
C10356 VP.n3439 a_400_38200# 0.34fF
C10357 VP.n3440 a_400_38200# 0.04fF
C10358 VP.n3441 a_400_38200# 0.02fF
C10359 VP.n3442 a_400_38200# 0.06fF
C10360 VP.n3443 a_400_38200# 0.30fF
C10361 VP.n3444 a_400_38200# 1.93fF
C10362 VP.n3445 a_400_38200# 0.12fF
C10363 VP.t986 a_400_38200# 0.02fF
C10364 VP.n3446 a_400_38200# 0.14fF
C10365 VP.t267 a_400_38200# 0.02fF
C10366 VP.n3448 a_400_38200# 0.24fF
C10367 VP.n3449 a_400_38200# 0.35fF
C10368 VP.n3450 a_400_38200# 0.60fF
C10369 VP.n3451 a_400_38200# 0.07fF
C10370 VP.n3452 a_400_38200# 0.72fF
C10371 VP.n3453 a_400_38200# 0.09fF
C10372 VP.n3454 a_400_38200# 0.16fF
C10373 VP.n3455 a_400_38200# 0.98fF
C10374 VP.n3456 a_400_38200# 0.15fF
C10375 VP.n3458 a_400_38200# 1.72fF
C10376 VP.t73 a_400_38200# 0.02fF
C10377 VP.n3459 a_400_38200# 0.12fF
C10378 VP.n3460 a_400_38200# 0.14fF
C10379 VP.t1139 a_400_38200# 0.02fF
C10380 VP.n3462 a_400_38200# 0.24fF
C10381 VP.n3463 a_400_38200# 0.91fF
C10382 VP.n3464 a_400_38200# 0.05fF
C10383 VP.n3465 a_400_38200# 0.10fF
C10384 VP.n3466 a_400_38200# 0.28fF
C10385 VP.n3467 a_400_38200# 0.15fF
C10386 VP.n3468 a_400_38200# 0.08fF
C10387 VP.n3469 a_400_38200# 0.14fF
C10388 VP.n3470 a_400_38200# 0.06fF
C10389 VP.n3471 a_400_38200# 0.06fF
C10390 VP.n3472 a_400_38200# 0.03fF
C10391 VP.n3473 a_400_38200# 0.05fF
C10392 VP.n3474 a_400_38200# 0.07fF
C10393 VP.n3475 a_400_38200# 0.19fF
C10394 VP.n3476 a_400_38200# 0.59fF
C10395 VP.n3477 a_400_38200# 0.34fF
C10396 VP.n3478 a_400_38200# 0.04fF
C10397 VP.n3479 a_400_38200# 0.02fF
C10398 VP.n3480 a_400_38200# 0.06fF
C10399 VP.n3481 a_400_38200# 0.30fF
C10400 VP.n3482 a_400_38200# 1.93fF
C10401 VP.n3483 a_400_38200# 0.12fF
C10402 VP.t538 a_400_38200# 0.02fF
C10403 VP.n3484 a_400_38200# 0.14fF
C10404 VP.t1122 a_400_38200# 0.02fF
C10405 VP.n3486 a_400_38200# 0.24fF
C10406 VP.n3487 a_400_38200# 0.35fF
C10407 VP.n3488 a_400_38200# 0.60fF
C10408 VP.n3489 a_400_38200# 0.07fF
C10409 VP.n3490 a_400_38200# 0.72fF
C10410 VP.n3491 a_400_38200# 0.09fF
C10411 VP.n3492 a_400_38200# 0.16fF
C10412 VP.n3493 a_400_38200# 0.98fF
C10413 VP.n3494 a_400_38200# 0.15fF
C10414 VP.n3496 a_400_38200# 1.72fF
C10415 VP.t955 a_400_38200# 0.02fF
C10416 VP.n3497 a_400_38200# 0.12fF
C10417 VP.n3498 a_400_38200# 0.14fF
C10418 VP.t690 a_400_38200# 0.02fF
C10419 VP.n3500 a_400_38200# 0.24fF
C10420 VP.n3501 a_400_38200# 0.91fF
C10421 VP.n3502 a_400_38200# 0.05fF
C10422 VP.n3503 a_400_38200# 0.10fF
C10423 VP.n3504 a_400_38200# 0.28fF
C10424 VP.n3505 a_400_38200# 0.15fF
C10425 VP.n3506 a_400_38200# 0.08fF
C10426 VP.n3507 a_400_38200# 0.14fF
C10427 VP.n3508 a_400_38200# 0.06fF
C10428 VP.n3509 a_400_38200# 0.06fF
C10429 VP.n3510 a_400_38200# 0.03fF
C10430 VP.n3511 a_400_38200# 0.05fF
C10431 VP.n3512 a_400_38200# 0.07fF
C10432 VP.n3513 a_400_38200# 0.19fF
C10433 VP.n3514 a_400_38200# 0.59fF
C10434 VP.n3515 a_400_38200# 0.34fF
C10435 VP.n3516 a_400_38200# 0.04fF
C10436 VP.n3517 a_400_38200# 0.02fF
C10437 VP.n3518 a_400_38200# 0.06fF
C10438 VP.n3519 a_400_38200# 0.30fF
C10439 VP.n3520 a_400_38200# 1.93fF
C10440 VP.n3521 a_400_38200# 0.12fF
C10441 VP.t854 a_400_38200# 0.02fF
C10442 VP.n3522 a_400_38200# 0.14fF
C10443 VP.t41 a_400_38200# 0.02fF
C10444 VP.n3524 a_400_38200# 0.24fF
C10445 VP.n3525 a_400_38200# 0.35fF
C10446 VP.n3526 a_400_38200# 0.60fF
C10447 VP.n3527 a_400_38200# 2.47fF
C10448 VP.n3528 a_400_38200# 2.20fF
C10449 VP.t1204 a_400_38200# 0.02fF
C10450 VP.n3529 a_400_38200# 0.12fF
C10451 VP.n3530 a_400_38200# 0.14fF
C10452 VP.t946 a_400_38200# 0.02fF
C10453 VP.n3532 a_400_38200# 0.24fF
C10454 VP.n3533 a_400_38200# 0.91fF
C10455 VP.n3534 a_400_38200# 0.05fF
C10456 VP.n3535 a_400_38200# 0.10fF
C10457 VP.n3536 a_400_38200# 0.28fF
C10458 VP.n3537 a_400_38200# 0.15fF
C10459 VP.n3538 a_400_38200# 0.08fF
C10460 VP.n3539 a_400_38200# 0.14fF
C10461 VP.n3540 a_400_38200# 0.06fF
C10462 VP.n3541 a_400_38200# 0.06fF
C10463 VP.n3542 a_400_38200# 0.03fF
C10464 VP.n3543 a_400_38200# 0.05fF
C10465 VP.n3544 a_400_38200# 0.07fF
C10466 VP.n3545 a_400_38200# 0.19fF
C10467 VP.n3546 a_400_38200# 0.59fF
C10468 VP.n3547 a_400_38200# 0.34fF
C10469 VP.n3548 a_400_38200# 0.04fF
C10470 VP.n3549 a_400_38200# 0.02fF
C10471 VP.n3550 a_400_38200# 0.06fF
C10472 VP.n3551 a_400_38200# 0.30fF
C10473 VP.n3552 a_400_38200# 1.93fF
C10474 VP.n3553 a_400_38200# 0.12fF
C10475 VP.t404 a_400_38200# 0.02fF
C10476 VP.n3554 a_400_38200# 0.14fF
C10477 VP.t989 a_400_38200# 0.02fF
C10478 VP.n3556 a_400_38200# 0.24fF
C10479 VP.n3557 a_400_38200# 0.35fF
C10480 VP.n3558 a_400_38200# 0.60fF
C10481 VP.n3559 a_400_38200# 2.47fF
C10482 VP.n3560 a_400_38200# 2.20fF
C10483 VP.t756 a_400_38200# 0.02fF
C10484 VP.n3561 a_400_38200# 0.12fF
C10485 VP.n3562 a_400_38200# 0.14fF
C10486 VP.t561 a_400_38200# 0.02fF
C10487 VP.n3564 a_400_38200# 0.24fF
C10488 VP.n3565 a_400_38200# 0.91fF
C10489 VP.n3566 a_400_38200# 0.05fF
C10490 VP.n3567 a_400_38200# 0.10fF
C10491 VP.n3568 a_400_38200# 0.28fF
C10492 VP.n3569 a_400_38200# 0.15fF
C10493 VP.n3570 a_400_38200# 0.08fF
C10494 VP.n3571 a_400_38200# 0.14fF
C10495 VP.n3572 a_400_38200# 0.06fF
C10496 VP.n3573 a_400_38200# 0.06fF
C10497 VP.n3574 a_400_38200# 0.03fF
C10498 VP.n3575 a_400_38200# 0.05fF
C10499 VP.n3576 a_400_38200# 0.07fF
C10500 VP.n3577 a_400_38200# 0.19fF
C10501 VP.n3578 a_400_38200# 0.59fF
C10502 VP.n3579 a_400_38200# 0.34fF
C10503 VP.n3580 a_400_38200# 0.04fF
C10504 VP.n3581 a_400_38200# 0.02fF
C10505 VP.n3582 a_400_38200# 0.06fF
C10506 VP.n3583 a_400_38200# 0.30fF
C10507 VP.n3584 a_400_38200# 1.93fF
C10508 VP.n3585 a_400_38200# 0.12fF
C10509 VP.t1260 a_400_38200# 0.02fF
C10510 VP.n3586 a_400_38200# 0.14fF
C10511 VP.t543 a_400_38200# 0.02fF
C10512 VP.n3588 a_400_38200# 0.24fF
C10513 VP.n3589 a_400_38200# 0.35fF
C10514 VP.n3590 a_400_38200# 0.60fF
C10515 VP.n3591 a_400_38200# 2.47fF
C10516 VP.n3592 a_400_38200# 2.20fF
C10517 VP.t302 a_400_38200# 0.02fF
C10518 VP.n3593 a_400_38200# 0.12fF
C10519 VP.n3594 a_400_38200# 0.14fF
C10520 VP.t90 a_400_38200# 0.02fF
C10521 VP.n3596 a_400_38200# 0.24fF
C10522 VP.n3597 a_400_38200# 0.91fF
C10523 VP.n3598 a_400_38200# 0.05fF
C10524 VP.n3599 a_400_38200# 0.10fF
C10525 VP.n3600 a_400_38200# 0.28fF
C10526 VP.n3601 a_400_38200# 0.15fF
C10527 VP.n3602 a_400_38200# 0.08fF
C10528 VP.n3603 a_400_38200# 0.14fF
C10529 VP.n3604 a_400_38200# 0.06fF
C10530 VP.n3605 a_400_38200# 0.06fF
C10531 VP.n3606 a_400_38200# 0.03fF
C10532 VP.n3607 a_400_38200# 0.05fF
C10533 VP.n3608 a_400_38200# 0.07fF
C10534 VP.n3609 a_400_38200# 0.19fF
C10535 VP.n3610 a_400_38200# 0.59fF
C10536 VP.n3611 a_400_38200# 0.34fF
C10537 VP.n3612 a_400_38200# 0.04fF
C10538 VP.n3613 a_400_38200# 0.02fF
C10539 VP.n3614 a_400_38200# 0.06fF
C10540 VP.n3615 a_400_38200# 0.30fF
C10541 VP.n3616 a_400_38200# 1.93fF
C10542 VP.n3617 a_400_38200# 0.12fF
C10543 VP.t815 a_400_38200# 0.02fF
C10544 VP.n3618 a_400_38200# 0.14fF
C10545 VP.t65 a_400_38200# 0.02fF
C10546 VP.n3620 a_400_38200# 0.24fF
C10547 VP.n3621 a_400_38200# 0.35fF
C10548 VP.n3622 a_400_38200# 0.60fF
C10549 VP.n3623 a_400_38200# 2.39fF
C10550 VP.n3624 a_400_38200# 1.79fF
C10551 VP.t1150 a_400_38200# 0.02fF
C10552 VP.n3625 a_400_38200# 0.12fF
C10553 VP.n3626 a_400_38200# 0.14fF
C10554 VP.t966 a_400_38200# 0.02fF
C10555 VP.n3628 a_400_38200# 0.24fF
C10556 VP.n3629 a_400_38200# 0.91fF
C10557 VP.n3630 a_400_38200# 0.05fF
C10558 VP.t72 a_400_38200# 34.79fF
C10559 VP.t547 a_400_38200# 0.02fF
C10560 VP.n3631 a_400_38200# 0.12fF
C10561 VP.n3632 a_400_38200# 0.14fF
C10562 VP.t284 a_400_38200# 0.02fF
C10563 VP.n3634 a_400_38200# 0.24fF
C10564 VP.n3635 a_400_38200# 0.91fF
C10565 VP.n3636 a_400_38200# 0.05fF
C10566 VP.t713 a_400_38200# 0.02fF
C10567 VP.n3637 a_400_38200# 0.24fF
C10568 VP.n3638 a_400_38200# 0.35fF
C10569 VP.n3639 a_400_38200# 0.60fF
C10570 VP.n3640 a_400_38200# 0.04fF
C10571 VP.n3641 a_400_38200# 0.08fF
C10572 VP.n3642 a_400_38200# 0.72fF
C10573 VP.n3643 a_400_38200# 0.09fF
C10574 VP.n3644 a_400_38200# 0.00fF
C10575 VP.n3645 a_400_38200# 0.98fF
C10576 VP.n3646 a_400_38200# 0.19fF
C10577 VP.n3648 a_400_38200# 1.72fF
C10578 VP.n3649 a_400_38200# 1.96fF
C10579 VP.n3650 a_400_38200# 1.04fF
C10580 VP.n3651 a_400_38200# 0.05fF
C10581 VP.n3652 a_400_38200# 0.03fF
C10582 VP.n3653 a_400_38200# 0.06fF
C10583 VP.n3654 a_400_38200# 0.06fF
C10584 VP.n3655 a_400_38200# 0.06fF
C10585 VP.n3656 a_400_38200# 0.07fF
C10586 VP.n3657 a_400_38200# 0.03fF
C10587 VP.n3658 a_400_38200# 0.05fF
C10588 VP.n3659 a_400_38200# 0.07fF
C10589 VP.n3660 a_400_38200# 0.19fF
C10590 VP.n3661 a_400_38200# 0.60fF
C10591 VP.n3662 a_400_38200# 0.76fF
C10592 VP.n3663 a_400_38200# 0.40fF
C10593 VP.n3664 a_400_38200# 0.03fF
C10594 VP.n3665 a_400_38200# 0.01fF
C10595 VP.t95 a_400_38200# 0.02fF
C10596 VP.n3666 a_400_38200# 0.25fF
C10597 VP.t1021 a_400_38200# 0.02fF
C10598 VP.n3667 a_400_38200# 0.95fF
C10599 VP.n3668 a_400_38200# 0.70fF
C10600 VP.n3669 a_400_38200# 1.93fF
C10601 VP.n3670 a_400_38200# 2.97fF
C10602 VP.n3671 a_400_38200# 2.27fF
C10603 VP.t864 a_400_38200# 0.02fF
C10604 VP.n3672 a_400_38200# 0.24fF
C10605 VP.n3673 a_400_38200# 0.35fF
C10606 VP.n3674 a_400_38200# 0.60fF
C10607 VP.n3675 a_400_38200# 0.12fF
C10608 VP.t272 a_400_38200# 0.02fF
C10609 VP.n3676 a_400_38200# 0.14fF
C10610 VP.n3678 a_400_38200# 0.04fF
C10611 VP.n3679 a_400_38200# 0.02fF
C10612 VP.n3680 a_400_38200# 0.06fF
C10613 VP.n3681 a_400_38200# 0.30fF
C10614 VP.n3682 a_400_38200# 0.10fF
C10615 VP.n3683 a_400_38200# 0.06fF
C10616 VP.n3684 a_400_38200# 0.06fF
C10617 VP.n3685 a_400_38200# 0.28fF
C10618 VP.n3686 a_400_38200# 0.03fF
C10619 VP.n3687 a_400_38200# 0.15fF
C10620 VP.n3688 a_400_38200# 0.08fF
C10621 VP.n3689 a_400_38200# 0.14fF
C10622 VP.n3690 a_400_38200# 0.03fF
C10623 VP.n3691 a_400_38200# 0.06fF
C10624 VP.n3692 a_400_38200# 0.06fF
C10625 VP.n3693 a_400_38200# 0.06fF
C10626 VP.n3694 a_400_38200# 0.06fF
C10627 VP.n3695 a_400_38200# 0.03fF
C10628 VP.n3696 a_400_38200# 0.05fF
C10629 VP.n3697 a_400_38200# 0.07fF
C10630 VP.n3698 a_400_38200# 0.19fF
C10631 VP.n3699 a_400_38200# 0.59fF
C10632 VP.n3700 a_400_38200# 0.34fF
C10633 VP.n3701 a_400_38200# 1.88fF
C10634 VP.t1193 a_400_38200# 0.02fF
C10635 VP.n3702 a_400_38200# 0.24fF
C10636 VP.n3703 a_400_38200# 0.91fF
C10637 VP.n3704 a_400_38200# 0.05fF
C10638 VP.t381 a_400_38200# 0.02fF
C10639 VP.n3705 a_400_38200# 0.12fF
C10640 VP.n3706 a_400_38200# 0.14fF
C10641 VP.n3708 a_400_38200# 0.19fF
C10642 VP.n3709 a_400_38200# 0.10fF
C10643 VP.n3710 a_400_38200# 0.10fF
C10644 VP.n3711 a_400_38200# 0.18fF
C10645 VP.n3712 a_400_38200# 0.09fF
C10646 VP.n3713 a_400_38200# 0.04fF
C10647 VP.n3714 a_400_38200# 0.19fF
C10648 VP.n3715 a_400_38200# 0.26fF
C10649 VP.n3716 a_400_38200# 1.17fF
C10650 VP.n3717 a_400_38200# 0.06fF
C10651 VP.n3718 a_400_38200# 0.44fF
C10652 VP.n3719 a_400_38200# 0.13fF
C10653 VP.n3720 a_400_38200# 0.02fF
C10654 VP.n3721 a_400_38200# 1.81fF
C10655 VP.n3722 a_400_38200# 0.12fF
C10656 VP.t1126 a_400_38200# 0.02fF
C10657 VP.n3723 a_400_38200# 0.14fF
C10658 VP.t420 a_400_38200# 0.02fF
C10659 VP.n3725 a_400_38200# 0.24fF
C10660 VP.n3726 a_400_38200# 0.35fF
C10661 VP.n3727 a_400_38200# 0.60fF
C10662 VP.n3728 a_400_38200# 3.18fF
C10663 VP.n3729 a_400_38200# 2.06fF
C10664 VP.n3730 a_400_38200# 1.98fF
C10665 VP.t738 a_400_38200# 0.02fF
C10666 VP.n3731 a_400_38200# 0.24fF
C10667 VP.n3732 a_400_38200# 0.91fF
C10668 VP.n3733 a_400_38200# 0.05fF
C10669 VP.t1237 a_400_38200# 0.02fF
C10670 VP.n3734 a_400_38200# 0.12fF
C10671 VP.n3735 a_400_38200# 0.14fF
C10672 VP.n3737 a_400_38200# 0.16fF
C10673 VP.n3738 a_400_38200# 0.19fF
C10674 VP.n3739 a_400_38200# 0.09fF
C10675 VP.n3740 a_400_38200# 0.04fF
C10676 VP.n3741 a_400_38200# 0.14fF
C10677 VP.n3742 a_400_38200# 0.64fF
C10678 VP.n3743 a_400_38200# 1.32fF
C10679 VP.n3744 a_400_38200# 1.81fF
C10680 VP.n3745 a_400_38200# 0.12fF
C10681 VP.t754 a_400_38200# 0.02fF
C10682 VP.n3746 a_400_38200# 0.14fF
C10683 VP.t1275 a_400_38200# 0.02fF
C10684 VP.n3748 a_400_38200# 0.24fF
C10685 VP.n3749 a_400_38200# 0.35fF
C10686 VP.n3750 a_400_38200# 0.60fF
C10687 VP.n3751 a_400_38200# 2.97fF
C10688 VP.n3752 a_400_38200# 2.27fF
C10689 VP.n3753 a_400_38200# 2.00fF
C10690 VP.t286 a_400_38200# 0.02fF
C10691 VP.n3754 a_400_38200# 0.24fF
C10692 VP.n3755 a_400_38200# 0.91fF
C10693 VP.n3756 a_400_38200# 0.05fF
C10694 VP.t793 a_400_38200# 0.02fF
C10695 VP.n3757 a_400_38200# 0.12fF
C10696 VP.n3758 a_400_38200# 0.14fF
C10697 VP.n3760 a_400_38200# 0.24fF
C10698 VP.t770 a_400_38200# 0.02fF
C10699 VP.n3761 a_400_38200# 0.36fF
C10700 VP.n3762 a_400_38200# 0.36fF
C10701 VP.n3763 a_400_38200# 0.67fF
C10702 VP.n3764 a_400_38200# 0.19fF
C10703 VP.n3765 a_400_38200# 0.03fF
C10704 VP.n3766 a_400_38200# 0.24fF
C10705 VP.n3767 a_400_38200# 0.99fF
C10706 VP.n3768 a_400_38200# 0.12fF
C10707 VP.n3769 a_400_38200# 0.19fF
C10708 VP.n3770 a_400_38200# 0.09fF
C10709 VP.n3771 a_400_38200# 0.18fF
C10710 VP.n3772 a_400_38200# 0.09fF
C10711 VP.n3773 a_400_38200# 0.08fF
C10712 VP.n3774 a_400_38200# 0.39fF
C10713 VP.n3775 a_400_38200# 0.24fF
C10714 VP.n3776 a_400_38200# 0.13fF
C10715 VP.n3777 a_400_38200# 0.02fF
C10716 VP.n3778 a_400_38200# 1.81fF
C10717 VP.n3779 a_400_38200# 2.96fF
C10718 VP.n3780 a_400_38200# 2.27fF
C10719 VP.n3781 a_400_38200# 0.74fF
C10720 VP.n3782 a_400_38200# 0.24fF
C10721 VP.t440 a_400_38200# 0.02fF
C10722 VP.n3783 a_400_38200# 0.35fF
C10723 VP.n3784 a_400_38200# 0.63fF
C10724 VP.n3785 a_400_38200# 0.40fF
C10725 VP.n3786 a_400_38200# 0.40fF
C10726 VP.n3787 a_400_38200# 0.12fF
C10727 VP.t1147 a_400_38200# 0.02fF
C10728 VP.n3788 a_400_38200# 0.14fF
C10729 VP.t1194 a_400_38200# 0.02fF
C10730 VP.n3790 a_400_38200# 0.12fF
C10731 VP.n3791 a_400_38200# 0.14fF
C10732 VP.n3793 a_400_38200# 15.28fF
C10733 VP.n3794 a_400_38200# 0.10fF
C10734 VP.n3795 a_400_38200# 0.06fF
C10735 VP.n3796 a_400_38200# 0.06fF
C10736 VP.n3797 a_400_38200# 0.28fF
C10737 VP.n3798 a_400_38200# 0.03fF
C10738 VP.n3799 a_400_38200# 0.15fF
C10739 VP.n3800 a_400_38200# 0.08fF
C10740 VP.n3801 a_400_38200# 0.14fF
C10741 VP.n3802 a_400_38200# 0.03fF
C10742 VP.n3803 a_400_38200# 0.06fF
C10743 VP.n3804 a_400_38200# 0.06fF
C10744 VP.n3805 a_400_38200# 0.06fF
C10745 VP.n3806 a_400_38200# 0.06fF
C10746 VP.n3807 a_400_38200# 0.03fF
C10747 VP.n3808 a_400_38200# 0.05fF
C10748 VP.n3809 a_400_38200# 0.07fF
C10749 VP.n3810 a_400_38200# 0.19fF
C10750 VP.n3811 a_400_38200# 0.59fF
C10751 VP.n3812 a_400_38200# 0.34fF
C10752 VP.n3813 a_400_38200# 0.04fF
C10753 VP.n3814 a_400_38200# 0.02fF
C10754 VP.n3815 a_400_38200# 0.06fF
C10755 VP.n3816 a_400_38200# 0.30fF
C10756 VP.n3817 a_400_38200# 1.93fF
C10757 VP.n3818 a_400_38200# 0.12fF
C10758 VP.t970 a_400_38200# 0.02fF
C10759 VP.n3819 a_400_38200# 0.14fF
C10760 VP.t251 a_400_38200# 0.02fF
C10761 VP.n3821 a_400_38200# 0.24fF
C10762 VP.n3822 a_400_38200# 0.35fF
C10763 VP.n3823 a_400_38200# 0.60fF
C10764 VP.n3824 a_400_38200# 0.07fF
C10765 VP.n3825 a_400_38200# 0.72fF
C10766 VP.n3826 a_400_38200# 0.20fF
C10767 VP.n3827 a_400_38200# 0.19fF
C10768 VP.n3828 a_400_38200# 0.10fF
C10769 VP.n3829 a_400_38200# 0.11fF
C10770 VP.n3830 a_400_38200# 0.09fF
C10771 VP.n3831 a_400_38200# 0.16fF
C10772 VP.n3832 a_400_38200# 0.10fF
C10773 VP.n3833 a_400_38200# 0.11fF
C10774 VP.n3834 a_400_38200# 0.19fF
C10775 VP.n3835 a_400_38200# 0.20fF
C10776 VP.n3836 a_400_38200# 0.98fF
C10777 VP.n3837 a_400_38200# 0.15fF
C10778 VP.n3839 a_400_38200# 1.72fF
C10779 VP.t1001 a_400_38200# 0.02fF
C10780 VP.n3840 a_400_38200# 0.12fF
C10781 VP.n3841 a_400_38200# 0.14fF
C10782 VP.t574 a_400_38200# 0.02fF
C10783 VP.n3843 a_400_38200# 0.24fF
C10784 VP.n3844 a_400_38200# 0.91fF
C10785 VP.n3845 a_400_38200# 0.05fF
C10786 VP.n3846 a_400_38200# 0.10fF
C10787 VP.n3847 a_400_38200# 0.28fF
C10788 VP.n3848 a_400_38200# 0.06fF
C10789 VP.n3849 a_400_38200# 0.06fF
C10790 VP.n3850 a_400_38200# 0.03fF
C10791 VP.n3851 a_400_38200# 0.15fF
C10792 VP.n3852 a_400_38200# 0.08fF
C10793 VP.n3853 a_400_38200# 0.14fF
C10794 VP.n3854 a_400_38200# 0.03fF
C10795 VP.n3855 a_400_38200# 0.06fF
C10796 VP.n3856 a_400_38200# 0.06fF
C10797 VP.n3857 a_400_38200# 0.06fF
C10798 VP.n3858 a_400_38200# 0.06fF
C10799 VP.n3859 a_400_38200# 0.03fF
C10800 VP.n3860 a_400_38200# 0.05fF
C10801 VP.n3861 a_400_38200# 0.07fF
C10802 VP.n3862 a_400_38200# 0.19fF
C10803 VP.n3863 a_400_38200# 0.59fF
C10804 VP.n3864 a_400_38200# 0.34fF
C10805 VP.n3865 a_400_38200# 0.04fF
C10806 VP.n3866 a_400_38200# 0.02fF
C10807 VP.n3867 a_400_38200# 0.06fF
C10808 VP.n3868 a_400_38200# 0.30fF
C10809 VP.n3869 a_400_38200# 1.93fF
C10810 VP.n3870 a_400_38200# 0.12fF
C10811 VP.t522 a_400_38200# 0.02fF
C10812 VP.n3871 a_400_38200# 0.14fF
C10813 VP.t1105 a_400_38200# 0.02fF
C10814 VP.n3873 a_400_38200# 0.24fF
C10815 VP.n3874 a_400_38200# 0.35fF
C10816 VP.n3875 a_400_38200# 0.60fF
C10817 VP.n3876 a_400_38200# 0.07fF
C10818 VP.n3877 a_400_38200# 0.72fF
C10819 VP.n3878 a_400_38200# 0.20fF
C10820 VP.n3879 a_400_38200# 0.19fF
C10821 VP.n3880 a_400_38200# 0.10fF
C10822 VP.n3881 a_400_38200# 0.11fF
C10823 VP.n3882 a_400_38200# 0.09fF
C10824 VP.n3883 a_400_38200# 0.16fF
C10825 VP.n3884 a_400_38200# 0.10fF
C10826 VP.n3885 a_400_38200# 0.11fF
C10827 VP.n3886 a_400_38200# 0.19fF
C10828 VP.n3887 a_400_38200# 0.20fF
C10829 VP.n3888 a_400_38200# 0.98fF
C10830 VP.n3889 a_400_38200# 0.15fF
C10831 VP.n3891 a_400_38200# 1.72fF
C10832 VP.t557 a_400_38200# 0.02fF
C10833 VP.n3892 a_400_38200# 0.12fF
C10834 VP.n3893 a_400_38200# 0.14fF
C10835 VP.t106 a_400_38200# 0.02fF
C10836 VP.n3895 a_400_38200# 0.24fF
C10837 VP.n3896 a_400_38200# 0.91fF
C10838 VP.n3897 a_400_38200# 0.05fF
C10839 VP.n3898 a_400_38200# 0.10fF
C10840 VP.n3899 a_400_38200# 0.06fF
C10841 VP.n3900 a_400_38200# 0.06fF
C10842 VP.n3901 a_400_38200# 0.28fF
C10843 VP.n3902 a_400_38200# 0.03fF
C10844 VP.n3903 a_400_38200# 0.15fF
C10845 VP.n3904 a_400_38200# 0.08fF
C10846 VP.n3905 a_400_38200# 0.14fF
C10847 VP.n3906 a_400_38200# 0.03fF
C10848 VP.n3907 a_400_38200# 0.06fF
C10849 VP.n3908 a_400_38200# 0.06fF
C10850 VP.n3909 a_400_38200# 0.06fF
C10851 VP.n3910 a_400_38200# 0.06fF
C10852 VP.n3911 a_400_38200# 0.03fF
C10853 VP.n3912 a_400_38200# 0.05fF
C10854 VP.n3913 a_400_38200# 0.07fF
C10855 VP.n3914 a_400_38200# 0.19fF
C10856 VP.n3915 a_400_38200# 0.59fF
C10857 VP.n3916 a_400_38200# 0.34fF
C10858 VP.n3917 a_400_38200# 0.04fF
C10859 VP.n3918 a_400_38200# 0.02fF
C10860 VP.n3919 a_400_38200# 0.06fF
C10861 VP.n3920 a_400_38200# 0.30fF
C10862 VP.n3921 a_400_38200# 1.93fF
C10863 VP.n3922 a_400_38200# 0.12fF
C10864 VP.t777 a_400_38200# 0.02fF
C10865 VP.n3923 a_400_38200# 0.14fF
C10866 VP.t21 a_400_38200# 0.02fF
C10867 VP.n3925 a_400_38200# 0.24fF
C10868 VP.n3926 a_400_38200# 0.35fF
C10869 VP.n3927 a_400_38200# 0.60fF
C10870 VP.n3928 a_400_38200# 0.72fF
C10871 VP.n3929 a_400_38200# 1.24fF
C10872 VP.n3930 a_400_38200# 0.54fF
C10873 VP.n3931 a_400_38200# 0.22fF
C10874 VP.n3932 a_400_38200# 1.73fF
C10875 VP.t86 a_400_38200# 0.02fF
C10876 VP.n3933 a_400_38200# 0.12fF
C10877 VP.n3934 a_400_38200# 0.14fF
C10878 VP.t380 a_400_38200# 0.02fF
C10879 VP.n3936 a_400_38200# 0.24fF
C10880 VP.n3937 a_400_38200# 0.91fF
C10881 VP.n3938 a_400_38200# 0.05fF
C10882 VP.n3939 a_400_38200# 0.10fF
C10883 VP.n3940 a_400_38200# 0.06fF
C10884 VP.n3941 a_400_38200# 0.06fF
C10885 VP.n3942 a_400_38200# 0.28fF
C10886 VP.n3943 a_400_38200# 0.03fF
C10887 VP.n3944 a_400_38200# 0.15fF
C10888 VP.n3945 a_400_38200# 0.08fF
C10889 VP.n3946 a_400_38200# 0.14fF
C10890 VP.n3947 a_400_38200# 0.03fF
C10891 VP.n3948 a_400_38200# 0.06fF
C10892 VP.n3949 a_400_38200# 0.06fF
C10893 VP.n3950 a_400_38200# 0.06fF
C10894 VP.n3951 a_400_38200# 0.06fF
C10895 VP.n3952 a_400_38200# 0.03fF
C10896 VP.n3953 a_400_38200# 0.05fF
C10897 VP.n3954 a_400_38200# 0.07fF
C10898 VP.n3955 a_400_38200# 0.19fF
C10899 VP.n3956 a_400_38200# 0.59fF
C10900 VP.n3957 a_400_38200# 0.34fF
C10901 VP.n3958 a_400_38200# 0.04fF
C10902 VP.n3959 a_400_38200# 0.02fF
C10903 VP.n3960 a_400_38200# 0.06fF
C10904 VP.n3961 a_400_38200# 0.30fF
C10905 VP.n3962 a_400_38200# 1.93fF
C10906 VP.n3963 a_400_38200# 0.12fF
C10907 VP.t328 a_400_38200# 0.02fF
C10908 VP.n3964 a_400_38200# 0.14fF
C10909 VP.t918 a_400_38200# 0.02fF
C10910 VP.n3966 a_400_38200# 0.24fF
C10911 VP.n3967 a_400_38200# 0.35fF
C10912 VP.n3968 a_400_38200# 0.60fF
C10913 VP.n3969 a_400_38200# 0.72fF
C10914 VP.n3970 a_400_38200# 1.24fF
C10915 VP.n3971 a_400_38200# 0.54fF
C10916 VP.n3972 a_400_38200# 0.22fF
C10917 VP.n3973 a_400_38200# 1.73fF
C10918 VP.t422 a_400_38200# 0.02fF
C10919 VP.n3974 a_400_38200# 0.12fF
C10920 VP.n3975 a_400_38200# 0.14fF
C10921 VP.t1235 a_400_38200# 0.02fF
C10922 VP.n3977 a_400_38200# 0.24fF
C10923 VP.n3978 a_400_38200# 0.91fF
C10924 VP.n3979 a_400_38200# 0.05fF
C10925 VP.n3980 a_400_38200# 0.10fF
C10926 VP.n3981 a_400_38200# 0.28fF
C10927 VP.n3982 a_400_38200# 0.06fF
C10928 VP.n3983 a_400_38200# 0.06fF
C10929 VP.n3984 a_400_38200# 0.03fF
C10930 VP.n3985 a_400_38200# 0.15fF
C10931 VP.n3986 a_400_38200# 0.08fF
C10932 VP.n3987 a_400_38200# 0.14fF
C10933 VP.n3988 a_400_38200# 0.03fF
C10934 VP.n3989 a_400_38200# 0.06fF
C10935 VP.n3990 a_400_38200# 0.06fF
C10936 VP.n3991 a_400_38200# 0.06fF
C10937 VP.n3992 a_400_38200# 0.06fF
C10938 VP.n3993 a_400_38200# 0.03fF
C10939 VP.n3994 a_400_38200# 0.05fF
C10940 VP.n3995 a_400_38200# 0.07fF
C10941 VP.n3996 a_400_38200# 0.19fF
C10942 VP.n3997 a_400_38200# 0.59fF
C10943 VP.n3998 a_400_38200# 0.34fF
C10944 VP.n3999 a_400_38200# 0.04fF
C10945 VP.n4000 a_400_38200# 0.02fF
C10946 VP.n4001 a_400_38200# 0.06fF
C10947 VP.n4002 a_400_38200# 0.30fF
C10948 VP.n4003 a_400_38200# 1.93fF
C10949 VP.n4004 a_400_38200# 0.12fF
C10950 VP.t1172 a_400_38200# 0.02fF
C10951 VP.n4005 a_400_38200# 0.14fF
C10952 VP.t467 a_400_38200# 0.02fF
C10953 VP.n4007 a_400_38200# 0.24fF
C10954 VP.n4008 a_400_38200# 0.35fF
C10955 VP.n4009 a_400_38200# 0.60fF
C10956 VP.n4010 a_400_38200# 0.72fF
C10957 VP.n4011 a_400_38200# 1.24fF
C10958 VP.n4012 a_400_38200# 0.54fF
C10959 VP.n4013 a_400_38200# 0.22fF
C10960 VP.n4014 a_400_38200# 1.73fF
C10961 VP.t1277 a_400_38200# 0.02fF
C10962 VP.n4015 a_400_38200# 0.12fF
C10963 VP.n4016 a_400_38200# 0.14fF
C10964 VP.t790 a_400_38200# 0.02fF
C10965 VP.n4018 a_400_38200# 0.24fF
C10966 VP.n4019 a_400_38200# 0.91fF
C10967 VP.n4020 a_400_38200# 0.05fF
C10968 VP.n4021 a_400_38200# 0.10fF
C10969 VP.n4022 a_400_38200# 0.28fF
C10970 VP.n4023 a_400_38200# 0.06fF
C10971 VP.n4024 a_400_38200# 0.06fF
C10972 VP.n4025 a_400_38200# 0.03fF
C10973 VP.n4026 a_400_38200# 0.15fF
C10974 VP.n4027 a_400_38200# 0.08fF
C10975 VP.n4028 a_400_38200# 0.14fF
C10976 VP.n4029 a_400_38200# 0.03fF
C10977 VP.n4030 a_400_38200# 0.06fF
C10978 VP.n4031 a_400_38200# 0.06fF
C10979 VP.n4032 a_400_38200# 0.06fF
C10980 VP.n4033 a_400_38200# 0.06fF
C10981 VP.n4034 a_400_38200# 0.03fF
C10982 VP.n4035 a_400_38200# 0.05fF
C10983 VP.n4036 a_400_38200# 0.07fF
C10984 VP.n4037 a_400_38200# 0.19fF
C10985 VP.n4038 a_400_38200# 0.59fF
C10986 VP.n4039 a_400_38200# 0.34fF
C10987 VP.n4040 a_400_38200# 0.04fF
C10988 VP.n4041 a_400_38200# 0.02fF
C10989 VP.n4042 a_400_38200# 0.06fF
C10990 VP.n4043 a_400_38200# 0.30fF
C10991 VP.n4044 a_400_38200# 1.93fF
C10992 VP.n4045 a_400_38200# 0.12fF
C10993 VP.t718 a_400_38200# 0.02fF
C10994 VP.n4046 a_400_38200# 0.14fF
C10995 VP.t1314 a_400_38200# 0.02fF
C10996 VP.n4048 a_400_38200# 0.24fF
C10997 VP.n4049 a_400_38200# 0.35fF
C10998 VP.n4050 a_400_38200# 0.60fF
C10999 VP.n4051 a_400_38200# 0.71fF
C11000 VP.n4052 a_400_38200# 1.39fF
C11001 VP.n4053 a_400_38200# 0.54fF
C11002 VP.n4054 a_400_38200# 0.21fF
C11003 VP.n4055 a_400_38200# 1.73fF
C11004 VP.t832 a_400_38200# 0.02fF
C11005 VP.n4056 a_400_38200# 0.12fF
C11006 VP.n4057 a_400_38200# 0.14fF
C11007 VP.t344 a_400_38200# 0.02fF
C11008 VP.n4059 a_400_38200# 0.24fF
C11009 VP.n4060 a_400_38200# 0.91fF
C11010 VP.n4061 a_400_38200# 0.05fF
C11011 VP.n4062 a_400_38200# 0.06fF
C11012 VP.n4063 a_400_38200# 0.06fF
C11013 VP.n4064 a_400_38200# 0.03fF
C11014 VP.n4065 a_400_38200# 0.10fF
C11015 VP.n4066 a_400_38200# 0.17fF
C11016 VP.n4067 a_400_38200# 0.10fF
C11017 VP.n4068 a_400_38200# 0.13fF
C11018 VP.n4069 a_400_38200# 0.02fF
C11019 VP.n4070 a_400_38200# 0.04fF
C11020 VP.n4071 a_400_38200# 0.06fF
C11021 VP.n4072 a_400_38200# 0.09fF
C11022 VP.n4073 a_400_38200# 0.10fF
C11023 VP.n4074 a_400_38200# 0.05fF
C11024 VP.n4075 a_400_38200# 0.19fF
C11025 VP.n4076 a_400_38200# 0.16fF
C11026 VP.n4077 a_400_38200# 0.04fF
C11027 VP.n4078 a_400_38200# 0.05fF
C11028 VP.n4079 a_400_38200# 0.04fF
C11029 VP.n4080 a_400_38200# 0.12fF
C11030 VP.n4081 a_400_38200# 0.09fF
C11031 VP.n4082 a_400_38200# 0.14fF
C11032 VP.n4083 a_400_38200# 0.56fF
C11033 VP.n4084 a_400_38200# 0.10fF
C11034 VP.n4085 a_400_38200# 1.93fF
C11035 VP.n4086 a_400_38200# 0.12fF
C11036 VP.t299 a_400_38200# 0.02fF
C11037 VP.n4087 a_400_38200# 0.14fF
C11038 VP.t890 a_400_38200# 0.02fF
C11039 VP.n4089 a_400_38200# 0.24fF
C11040 VP.n4090 a_400_38200# 0.35fF
C11041 VP.n4091 a_400_38200# 0.60fF
C11042 VP.n4092 a_400_38200# 2.23fF
C11043 VP.n4093 a_400_38200# 0.18fF
C11044 VP.n4094 a_400_38200# 0.45fF
C11045 VP.n4095 a_400_38200# 0.06fF
C11046 VP.n4096 a_400_38200# 0.01fF
C11047 VP.n4097 a_400_38200# 0.01fF
C11048 VP.n4098 a_400_38200# 0.04fF
C11049 VP.n4099 a_400_38200# 0.02fF
C11050 VP.n4100 a_400_38200# 0.07fF
C11051 VP.n4101 a_400_38200# 0.04fF
C11052 VP.n4102 a_400_38200# 0.14fF
C11053 VP.n4103 a_400_38200# 0.45fF
C11054 VP.n4104 a_400_38200# 1.46fF
C11055 VP.n4105 a_400_38200# 1.78fF
C11056 VP.t346 a_400_38200# 0.02fF
C11057 VP.n4106 a_400_38200# 0.12fF
C11058 VP.n4107 a_400_38200# 0.14fF
C11059 VP.t1216 a_400_38200# 0.02fF
C11060 VP.n4109 a_400_38200# 0.24fF
C11061 VP.n4110 a_400_38200# 0.91fF
C11062 VP.n4111 a_400_38200# 0.05fF
C11063 VP.n4112 a_400_38200# 1.92fF
C11064 VP.n4113 a_400_38200# 2.51fF
C11065 VP.t684 a_400_38200# 0.02fF
C11066 VP.n4114 a_400_38200# 0.24fF
C11067 VP.n4115 a_400_38200# 0.35fF
C11068 VP.n4116 a_400_38200# 0.60fF
C11069 VP.n4117 a_400_38200# 0.12fF
C11070 VP.t77 a_400_38200# 0.02fF
C11071 VP.n4118 a_400_38200# 0.14fF
C11072 VP.n4120 a_400_38200# 0.06fF
C11073 VP.n4121 a_400_38200# 0.30fF
C11074 VP.n4122 a_400_38200# 0.20fF
C11075 VP.n4123 a_400_38200# 0.09fF
C11076 VP.n4124 a_400_38200# 0.26fF
C11077 VP.n4125 a_400_38200# 0.22fF
C11078 VP.n4126 a_400_38200# 0.19fF
C11079 VP.n4127 a_400_38200# 0.05fF
C11080 VP.n4128 a_400_38200# 0.13fF
C11081 VP.n4129 a_400_38200# 0.09fF
C11082 VP.n4130 a_400_38200# 0.09fF
C11083 VP.n4131 a_400_38200# 0.07fF
C11084 VP.n4132 a_400_38200# 0.71fF
C11085 VP.n4133 a_400_38200# 0.24fF
C11086 VP.n4134 a_400_38200# 1.88fF
C11087 VP.t741 a_400_38200# 0.02fF
C11088 VP.n4135 a_400_38200# 0.12fF
C11089 VP.n4136 a_400_38200# 0.14fF
C11090 VP.t1006 a_400_38200# 0.02fF
C11091 VP.n4138 a_400_38200# 0.24fF
C11092 VP.n4139 a_400_38200# 0.91fF
C11093 VP.n4140 a_400_38200# 0.05fF
C11094 VP.t76 a_400_38200# 35.17fF
C11095 VP.t696 a_400_38200# 0.02fF
C11096 VP.n4141 a_400_38200# 1.21fF
C11097 VP.n4142 a_400_38200# 0.25fF
C11098 VP.n4143 a_400_38200# 26.29fF
C11099 VP.n4144 a_400_38200# 26.29fF
C11100 VP.n4145 a_400_38200# 0.76fF
C11101 VP.n4146 a_400_38200# 0.27fF
C11102 VP.n4147 a_400_38200# 0.59fF
C11103 VP.n4148 a_400_38200# 0.10fF
C11104 VP.n4149 a_400_38200# 3.02fF
C11105 VP.t20 a_400_38200# 15.72fF
C11106 VP.n4150 a_400_38200# 1.15fF
C11107 VP.n4152 a_400_38200# 13.70fF
C11108 VP.n4154 a_400_38200# 1.99fF
C11109 VP.n4155 a_400_38200# 4.39fF
C11110 VP.n4156 a_400_38200# 0.03fF
C11111 VP.n4157 a_400_38200# 0.05fF
C11112 VP.n4158 a_400_38200# 0.07fF
C11113 VP.n4159 a_400_38200# 0.03fF
C11114 VP.n4160 a_400_38200# 0.06fF
C11115 VP.n4161 a_400_38200# 0.06fF
C11116 VP.n4162 a_400_38200# 0.06fF
C11117 VP.n4163 a_400_38200# 0.07fF
C11118 VP.n4164 a_400_38200# 0.57fF
C11119 VP.n4165 a_400_38200# 1.88fF
C11120 VP.n4166 a_400_38200# 0.92fF
C11121 VP.n4167 a_400_38200# 2.63fF
C11122 VP.n4168 a_400_38200# 0.10fF
C11123 VP.n4169 a_400_38200# 0.28fF
C11124 VP.n4170 a_400_38200# 0.15fF
C11125 VP.n4171 a_400_38200# 0.08fF
C11126 VP.n4172 a_400_38200# 0.14fF
C11127 VP.n4173 a_400_38200# 0.06fF
C11128 VP.n4174 a_400_38200# 0.06fF
C11129 VP.n4175 a_400_38200# 0.03fF
C11130 VP.n4176 a_400_38200# 0.05fF
C11131 VP.n4177 a_400_38200# 0.07fF
C11132 VP.n4178 a_400_38200# 0.19fF
C11133 VP.n4179 a_400_38200# 0.59fF
C11134 VP.n4180 a_400_38200# 0.34fF
C11135 VP.n4181 a_400_38200# 0.04fF
C11136 VP.n4182 a_400_38200# 0.02fF
C11137 VP.n4183 a_400_38200# 0.06fF
C11138 VP.n4184 a_400_38200# 0.30fF
C11139 VP.n4185 a_400_38200# 0.12fF
C11140 VP.t1328 a_400_38200# 0.02fF
C11141 VP.n4186 a_400_38200# 0.14fF
C11142 VP.n4188 a_400_38200# 1.93fF
C11143 VP.t1289 a_400_38200# 0.02fF
C11144 VP.n4189 a_400_38200# 0.24fF
C11145 VP.n4190 a_400_38200# 0.35fF
C11146 VP.n4191 a_400_38200# 0.60fF
C11147 VP.n4192 a_400_38200# 0.12fF
C11148 VP.t693 a_400_38200# 0.02fF
C11149 VP.n4193 a_400_38200# 0.14fF
C11150 VP.n4195 a_400_38200# 0.04fF
C11151 VP.n4196 a_400_38200# 0.02fF
C11152 VP.n4197 a_400_38200# 0.06fF
C11153 VP.n4198 a_400_38200# 0.30fF
C11154 VP.n4199 a_400_38200# 0.10fF
C11155 VP.n4200 a_400_38200# 0.28fF
C11156 VP.n4201 a_400_38200# 0.15fF
C11157 VP.n4202 a_400_38200# 0.08fF
C11158 VP.n4203 a_400_38200# 0.14fF
C11159 VP.n4204 a_400_38200# 0.06fF
C11160 VP.n4205 a_400_38200# 0.06fF
C11161 VP.n4206 a_400_38200# 0.03fF
C11162 VP.n4207 a_400_38200# 0.05fF
C11163 VP.n4208 a_400_38200# 0.07fF
C11164 VP.n4209 a_400_38200# 0.19fF
C11165 VP.n4210 a_400_38200# 0.59fF
C11166 VP.n4211 a_400_38200# 0.34fF
C11167 VP.n4212 a_400_38200# 2.18fF
C11168 VP.t859 a_400_38200# 0.02fF
C11169 VP.n4213 a_400_38200# 0.24fF
C11170 VP.n4214 a_400_38200# 0.91fF
C11171 VP.n4215 a_400_38200# 0.05fF
C11172 VP.t1055 a_400_38200# 0.02fF
C11173 VP.n4216 a_400_38200# 0.12fF
C11174 VP.n4217 a_400_38200# 0.14fF
C11175 VP.n4219 a_400_38200# 0.10fF
C11176 VP.n4220 a_400_38200# 0.10fF
C11177 VP.n4221 a_400_38200# 0.18fF
C11178 VP.n4222 a_400_38200# 0.09fF
C11179 VP.n4223 a_400_38200# 0.04fF
C11180 VP.n4224 a_400_38200# 0.26fF
C11181 VP.n4225 a_400_38200# 1.17fF
C11182 VP.n4226 a_400_38200# 0.06fF
C11183 VP.n4227 a_400_38200# 0.44fF
C11184 VP.n4228 a_400_38200# 0.13fF
C11185 VP.n4229 a_400_38200# 0.02fF
C11186 VP.n4230 a_400_38200# 1.81fF
C11187 VP.n4231 a_400_38200# 0.12fF
C11188 VP.t250 a_400_38200# 0.02fF
C11189 VP.n4232 a_400_38200# 0.14fF
C11190 VP.t845 a_400_38200# 0.02fF
C11191 VP.n4234 a_400_38200# 0.24fF
C11192 VP.n4235 a_400_38200# 0.35fF
C11193 VP.n4236 a_400_38200# 0.60fF
C11194 VP.n4237 a_400_38200# 2.28fF
C11195 VP.t413 a_400_38200# 0.02fF
C11196 VP.n4238 a_400_38200# 0.24fF
C11197 VP.n4239 a_400_38200# 0.91fF
C11198 VP.n4240 a_400_38200# 0.05fF
C11199 VP.t607 a_400_38200# 0.02fF
C11200 VP.n4241 a_400_38200# 0.12fF
C11201 VP.n4242 a_400_38200# 0.14fF
C11202 VP.n4244 a_400_38200# 0.06fF
C11203 VP.n4245 a_400_38200# 0.09fF
C11204 VP.n4246 a_400_38200# 0.09fF
C11205 VP.n4247 a_400_38200# 1.45fF
C11206 VP.n4248 a_400_38200# 0.14fF
C11207 VP.n4249 a_400_38200# 0.07fF
C11208 VP.n4250 a_400_38200# 0.72fF
C11209 VP.n4251 a_400_38200# 1.81fF
C11210 VP.n4252 a_400_38200# 0.12fF
C11211 VP.t1103 a_400_38200# 0.02fF
C11212 VP.n4253 a_400_38200# 0.14fF
C11213 VP.t394 a_400_38200# 0.02fF
C11214 VP.n4255 a_400_38200# 0.24fF
C11215 VP.n4256 a_400_38200# 0.35fF
C11216 VP.n4257 a_400_38200# 0.60fF
C11217 VP.n4258 a_400_38200# 2.30fF
C11218 VP.t1268 a_400_38200# 0.02fF
C11219 VP.n4259 a_400_38200# 0.24fF
C11220 VP.n4260 a_400_38200# 0.91fF
C11221 VP.n4261 a_400_38200# 0.05fF
C11222 VP.t141 a_400_38200# 0.02fF
C11223 VP.n4262 a_400_38200# 0.12fF
C11224 VP.n4263 a_400_38200# 0.14fF
C11225 VP.n4265 a_400_38200# 0.06fF
C11226 VP.n4266 a_400_38200# 0.25fF
C11227 VP.n4267 a_400_38200# 0.45fF
C11228 VP.n4268 a_400_38200# 0.03fF
C11229 VP.n4269 a_400_38200# 0.05fF
C11230 VP.n4270 a_400_38200# 0.07fF
C11231 VP.n4271 a_400_38200# 0.06fF
C11232 VP.n4272 a_400_38200# 0.06fF
C11233 VP.n4273 a_400_38200# 0.19fF
C11234 VP.n4274 a_400_38200# 0.59fF
C11235 VP.n4275 a_400_38200# 0.34fF
C11236 VP.n4276 a_400_38200# 0.05fF
C11237 VP.n4277 a_400_38200# 0.30fF
C11238 VP.n4278 a_400_38200# 1.93fF
C11239 VP.n4279 a_400_38200# 0.12fF
C11240 VP.t661 a_400_38200# 0.02fF
C11241 VP.n4280 a_400_38200# 0.14fF
C11242 VP.t1250 a_400_38200# 0.02fF
C11243 VP.n4282 a_400_38200# 0.24fF
C11244 VP.n4283 a_400_38200# 0.35fF
C11245 VP.n4284 a_400_38200# 0.60fF
C11246 VP.n4285 a_400_38200# 2.04fF
C11247 VP.t823 a_400_38200# 0.02fF
C11248 VP.n4286 a_400_38200# 0.24fF
C11249 VP.n4287 a_400_38200# 0.91fF
C11250 VP.n4288 a_400_38200# 0.05fF
C11251 VP.t1075 a_400_38200# 0.02fF
C11252 VP.n4289 a_400_38200# 0.12fF
C11253 VP.n4290 a_400_38200# 0.14fF
C11254 VP.n4292 a_400_38200# 0.24fF
C11255 VP.t372 a_400_38200# 0.02fF
C11256 VP.n4293 a_400_38200# 0.36fF
C11257 VP.n4294 a_400_38200# 0.36fF
C11258 VP.n4295 a_400_38200# 0.67fF
C11259 VP.n4296 a_400_38200# 0.06fF
C11260 VP.n4297 a_400_38200# 0.09fF
C11261 VP.n4298 a_400_38200# 0.09fF
C11262 VP.n4299 a_400_38200# 0.43fF
C11263 VP.n4300 a_400_38200# 0.69fF
C11264 VP.n4301 a_400_38200# 0.14fF
C11265 VP.n4302 a_400_38200# 0.07fF
C11266 VP.n4303 a_400_38200# 0.72fF
C11267 VP.n4304 a_400_38200# 1.81fF
C11268 VP.n4305 a_400_38200# 1.06fF
C11269 VP.n4306 a_400_38200# 0.24fF
C11270 VP.t805 a_400_38200# 0.02fF
C11271 VP.n4307 a_400_38200# 0.35fF
C11272 VP.n4308 a_400_38200# 0.63fF
C11273 VP.n4309 a_400_38200# 0.40fF
C11274 VP.n4310 a_400_38200# 0.40fF
C11275 VP.n4311 a_400_38200# 0.12fF
C11276 VP.t213 a_400_38200# 0.02fF
C11277 VP.n4312 a_400_38200# 0.14fF
C11278 VP.t632 a_400_38200# 0.02fF
C11279 VP.n4314 a_400_38200# 0.12fF
C11280 VP.n4315 a_400_38200# 0.14fF
C11281 VP.n4317 a_400_38200# 0.31fF
C11282 VP.n4318 a_400_38200# 0.04fF
C11283 VP.n4319 a_400_38200# 0.88fF
C11284 VP.n4320 a_400_38200# 0.48fF
C11285 VP.n4321 a_400_38200# 0.88fF
C11286 VP.n4322 a_400_38200# 0.60fF
C11287 VP.n4323 a_400_38200# 2.33fF
C11288 VP.n4324 a_400_38200# 0.59fF
C11289 VP.n4325 a_400_38200# 0.02fF
C11290 VP.n4326 a_400_38200# 0.96fF
C11291 VP.t105 a_400_38200# 15.72fF
C11292 VP.n4327 a_400_38200# 15.42fF
C11293 VP.n4329 a_400_38200# 0.38fF
C11294 VP.n4330 a_400_38200# 0.23fF
C11295 VP.n4331 a_400_38200# 3.28fF
C11296 VP.n4332 a_400_38200# 1.41fF
C11297 VP.n4333 a_400_38200# 0.30fF
C11298 VP.t602 a_400_38200# 0.02fF
C11299 VP.n4334 a_400_38200# 0.64fF
C11300 VP.n4335 a_400_38200# 0.60fF
C11301 VP.n4336 a_400_38200# 1.88fF
C11302 VP.n4337 a_400_38200# 4.64fF
C11303 VP.t164 a_400_38200# 0.02fF
C11304 VP.n4338 a_400_38200# 1.19fF
C11305 VP.n4339 a_400_38200# 0.05fF
C11306 VP.t423 a_400_38200# 0.02fF
C11307 VP.n4340 a_400_38200# 0.01fF
C11308 VP.n4341 a_400_38200# 0.26fF
C11309 VP.n4343 a_400_38200# 15.28fF
C11310 VP.n4344 a_400_38200# 0.10fF
C11311 VP.n4345 a_400_38200# 0.28fF
C11312 VP.n4346 a_400_38200# 0.15fF
C11313 VP.n4347 a_400_38200# 0.08fF
C11314 VP.n4348 a_400_38200# 0.14fF
C11315 VP.n4349 a_400_38200# 0.06fF
C11316 VP.n4350 a_400_38200# 0.06fF
C11317 VP.n4351 a_400_38200# 0.03fF
C11318 VP.n4352 a_400_38200# 0.05fF
C11319 VP.n4353 a_400_38200# 0.07fF
C11320 VP.n4354 a_400_38200# 0.19fF
C11321 VP.n4355 a_400_38200# 0.59fF
C11322 VP.n4356 a_400_38200# 0.34fF
C11323 VP.n4357 a_400_38200# 0.04fF
C11324 VP.n4358 a_400_38200# 0.02fF
C11325 VP.n4359 a_400_38200# 0.06fF
C11326 VP.n4360 a_400_38200# 0.30fF
C11327 VP.n4361 a_400_38200# 1.93fF
C11328 VP.n4362 a_400_38200# 0.12fF
C11329 VP.t877 a_400_38200# 0.02fF
C11330 VP.n4363 a_400_38200# 0.14fF
C11331 VP.t158 a_400_38200# 0.02fF
C11332 VP.n4365 a_400_38200# 0.24fF
C11333 VP.n4366 a_400_38200# 0.35fF
C11334 VP.n4367 a_400_38200# 0.60fF
C11335 VP.n4368 a_400_38200# 0.07fF
C11336 VP.n4369 a_400_38200# 0.72fF
C11337 VP.n4370 a_400_38200# 0.09fF
C11338 VP.n4371 a_400_38200# 0.16fF
C11339 VP.n4372 a_400_38200# 0.98fF
C11340 VP.n4373 a_400_38200# 0.15fF
C11341 VP.n4375 a_400_38200# 1.72fF
C11342 VP.t1293 a_400_38200# 0.02fF
C11343 VP.n4376 a_400_38200# 0.12fF
C11344 VP.n4377 a_400_38200# 0.14fF
C11345 VP.t1038 a_400_38200# 0.02fF
C11346 VP.n4379 a_400_38200# 0.24fF
C11347 VP.n4380 a_400_38200# 0.91fF
C11348 VP.n4381 a_400_38200# 0.05fF
C11349 VP.n4382 a_400_38200# 0.10fF
C11350 VP.n4383 a_400_38200# 0.28fF
C11351 VP.n4384 a_400_38200# 0.15fF
C11352 VP.n4385 a_400_38200# 0.08fF
C11353 VP.n4386 a_400_38200# 0.14fF
C11354 VP.n4387 a_400_38200# 0.06fF
C11355 VP.n4388 a_400_38200# 0.06fF
C11356 VP.n4389 a_400_38200# 0.03fF
C11357 VP.n4390 a_400_38200# 0.05fF
C11358 VP.n4391 a_400_38200# 0.07fF
C11359 VP.n4392 a_400_38200# 0.19fF
C11360 VP.n4393 a_400_38200# 0.59fF
C11361 VP.n4394 a_400_38200# 0.34fF
C11362 VP.n4395 a_400_38200# 0.04fF
C11363 VP.n4396 a_400_38200# 0.02fF
C11364 VP.n4397 a_400_38200# 0.06fF
C11365 VP.n4398 a_400_38200# 0.30fF
C11366 VP.n4399 a_400_38200# 1.93fF
C11367 VP.n4400 a_400_38200# 0.12fF
C11368 VP.t429 a_400_38200# 0.02fF
C11369 VP.n4401 a_400_38200# 0.14fF
C11370 VP.t1011 a_400_38200# 0.02fF
C11371 VP.n4403 a_400_38200# 0.24fF
C11372 VP.n4404 a_400_38200# 0.35fF
C11373 VP.n4405 a_400_38200# 0.60fF
C11374 VP.n4406 a_400_38200# 2.47fF
C11375 VP.n4407 a_400_38200# 2.20fF
C11376 VP.t848 a_400_38200# 0.02fF
C11377 VP.n4408 a_400_38200# 0.12fF
C11378 VP.n4409 a_400_38200# 0.14fF
C11379 VP.t588 a_400_38200# 0.02fF
C11380 VP.n4411 a_400_38200# 0.24fF
C11381 VP.n4412 a_400_38200# 0.91fF
C11382 VP.n4413 a_400_38200# 0.05fF
C11383 VP.n4414 a_400_38200# 0.10fF
C11384 VP.n4415 a_400_38200# 0.28fF
C11385 VP.n4416 a_400_38200# 0.15fF
C11386 VP.n4417 a_400_38200# 0.08fF
C11387 VP.n4418 a_400_38200# 0.14fF
C11388 VP.n4419 a_400_38200# 0.06fF
C11389 VP.n4420 a_400_38200# 0.06fF
C11390 VP.n4421 a_400_38200# 0.03fF
C11391 VP.n4422 a_400_38200# 0.05fF
C11392 VP.n4423 a_400_38200# 0.07fF
C11393 VP.n4424 a_400_38200# 0.19fF
C11394 VP.n4425 a_400_38200# 0.59fF
C11395 VP.n4426 a_400_38200# 0.34fF
C11396 VP.n4427 a_400_38200# 0.04fF
C11397 VP.n4428 a_400_38200# 0.02fF
C11398 VP.n4429 a_400_38200# 0.06fF
C11399 VP.n4430 a_400_38200# 0.30fF
C11400 VP.n4431 a_400_38200# 1.93fF
C11401 VP.n4432 a_400_38200# 0.12fF
C11402 VP.t746 a_400_38200# 0.02fF
C11403 VP.n4433 a_400_38200# 0.14fF
C11404 VP.t1269 a_400_38200# 0.02fF
C11405 VP.n4435 a_400_38200# 0.24fF
C11406 VP.n4436 a_400_38200# 0.35fF
C11407 VP.n4437 a_400_38200# 0.60fF
C11408 VP.n4438 a_400_38200# 2.47fF
C11409 VP.n4439 a_400_38200# 2.20fF
C11410 VP.t1093 a_400_38200# 0.02fF
C11411 VP.n4440 a_400_38200# 0.12fF
C11412 VP.n4441 a_400_38200# 0.14fF
C11413 VP.t840 a_400_38200# 0.02fF
C11414 VP.n4443 a_400_38200# 0.24fF
C11415 VP.n4444 a_400_38200# 0.91fF
C11416 VP.n4445 a_400_38200# 0.05fF
C11417 VP.n4446 a_400_38200# 0.10fF
C11418 VP.n4447 a_400_38200# 0.28fF
C11419 VP.n4448 a_400_38200# 0.15fF
C11420 VP.n4449 a_400_38200# 0.08fF
C11421 VP.n4450 a_400_38200# 0.14fF
C11422 VP.n4451 a_400_38200# 0.06fF
C11423 VP.n4452 a_400_38200# 0.06fF
C11424 VP.n4453 a_400_38200# 0.03fF
C11425 VP.n4454 a_400_38200# 0.05fF
C11426 VP.n4455 a_400_38200# 0.07fF
C11427 VP.n4456 a_400_38200# 0.19fF
C11428 VP.n4457 a_400_38200# 0.59fF
C11429 VP.n4458 a_400_38200# 0.34fF
C11430 VP.n4459 a_400_38200# 0.04fF
C11431 VP.n4460 a_400_38200# 0.02fF
C11432 VP.n4461 a_400_38200# 0.06fF
C11433 VP.n4462 a_400_38200# 0.30fF
C11434 VP.n4463 a_400_38200# 1.93fF
C11435 VP.n4464 a_400_38200# 0.12fF
C11436 VP.t292 a_400_38200# 0.02fF
C11437 VP.n4465 a_400_38200# 0.14fF
C11438 VP.t883 a_400_38200# 0.02fF
C11439 VP.n4467 a_400_38200# 0.24fF
C11440 VP.n4468 a_400_38200# 0.35fF
C11441 VP.n4469 a_400_38200# 0.60fF
C11442 VP.n4470 a_400_38200# 2.47fF
C11443 VP.n4471 a_400_38200# 2.20fF
C11444 VP.t650 a_400_38200# 0.02fF
C11445 VP.n4472 a_400_38200# 0.12fF
C11446 VP.n4473 a_400_38200# 0.14fF
C11447 VP.t456 a_400_38200# 0.02fF
C11448 VP.n4475 a_400_38200# 0.24fF
C11449 VP.n4476 a_400_38200# 0.91fF
C11450 VP.n4477 a_400_38200# 0.05fF
C11451 VP.n4478 a_400_38200# 0.10fF
C11452 VP.n4479 a_400_38200# 0.28fF
C11453 VP.n4480 a_400_38200# 0.15fF
C11454 VP.n4481 a_400_38200# 0.08fF
C11455 VP.n4482 a_400_38200# 0.14fF
C11456 VP.n4483 a_400_38200# 0.06fF
C11457 VP.n4484 a_400_38200# 0.06fF
C11458 VP.n4485 a_400_38200# 0.03fF
C11459 VP.n4486 a_400_38200# 0.05fF
C11460 VP.n4487 a_400_38200# 0.07fF
C11461 VP.n4488 a_400_38200# 0.19fF
C11462 VP.n4489 a_400_38200# 0.59fF
C11463 VP.n4490 a_400_38200# 0.34fF
C11464 VP.n4491 a_400_38200# 0.04fF
C11465 VP.n4492 a_400_38200# 0.02fF
C11466 VP.n4493 a_400_38200# 0.06fF
C11467 VP.n4494 a_400_38200# 0.30fF
C11468 VP.n4495 a_400_38200# 1.93fF
C11469 VP.n4496 a_400_38200# 0.12fF
C11470 VP.t1143 a_400_38200# 0.02fF
C11471 VP.n4497 a_400_38200# 0.14fF
C11472 VP.t433 a_400_38200# 0.02fF
C11473 VP.n4499 a_400_38200# 0.24fF
C11474 VP.n4500 a_400_38200# 0.35fF
C11475 VP.n4501 a_400_38200# 0.60fF
C11476 VP.n4502 a_400_38200# 2.39fF
C11477 VP.n4503 a_400_38200# 1.79fF
C11478 VP.t203 a_400_38200# 0.02fF
C11479 VP.n4504 a_400_38200# 0.12fF
C11480 VP.n4505 a_400_38200# 0.14fF
C11481 VP.t1306 a_400_38200# 0.02fF
C11482 VP.n4507 a_400_38200# 0.24fF
C11483 VP.n4508 a_400_38200# 0.91fF
C11484 VP.n4509 a_400_38200# 0.05fF
C11485 VP.n4510 a_400_38200# 1.93fF
C11486 VP.t354 a_400_38200# 0.02fF
C11487 VP.n4511 a_400_38200# 0.24fF
C11488 VP.n4512 a_400_38200# 0.35fF
C11489 VP.n4513 a_400_38200# 0.60fF
C11490 VP.n4514 a_400_38200# 0.12fF
C11491 VP.t1068 a_400_38200# 0.02fF
C11492 VP.n4515 a_400_38200# 0.14fF
C11493 VP.n4517 a_400_38200# 0.02fF
C11494 VP.n4518 a_400_38200# 0.32fF
C11495 VP.n4519 a_400_38200# 0.04fF
C11496 VP.n4520 a_400_38200# 0.05fF
C11497 VP.n4521 a_400_38200# 0.04fF
C11498 VP.n4522 a_400_38200# 0.12fF
C11499 VP.n4523 a_400_38200# 0.09fF
C11500 VP.n4524 a_400_38200# 0.14fF
C11501 VP.n4525 a_400_38200# 0.08fF
C11502 VP.n4526 a_400_38200# 0.09fF
C11503 VP.n4527 a_400_38200# 0.07fF
C11504 VP.n4528 a_400_38200# 0.56fF
C11505 VP.n4529 a_400_38200# 0.20fF
C11506 VP.n4530 a_400_38200# 2.19fF
C11507 VP.t176 a_400_38200# 0.02fF
C11508 VP.n4531 a_400_38200# 0.12fF
C11509 VP.n4532 a_400_38200# 0.14fF
C11510 VP.t1227 a_400_38200# 0.02fF
C11511 VP.n4534 a_400_38200# 0.24fF
C11512 VP.n4535 a_400_38200# 0.91fF
C11513 VP.n4536 a_400_38200# 0.05fF
C11514 VP.t140 a_400_38200# 34.79fF
C11515 VP.t438 a_400_38200# 0.02fF
C11516 VP.n4537 a_400_38200# 0.12fF
C11517 VP.n4538 a_400_38200# 0.14fF
C11518 VP.t188 a_400_38200# 0.02fF
C11519 VP.n4540 a_400_38200# 0.24fF
C11520 VP.n4541 a_400_38200# 0.91fF
C11521 VP.n4542 a_400_38200# 0.05fF
C11522 VP.t621 a_400_38200# 0.02fF
C11523 VP.n4543 a_400_38200# 0.24fF
C11524 VP.n4544 a_400_38200# 0.35fF
C11525 VP.n4545 a_400_38200# 0.60fF
C11526 VP.n4546 a_400_38200# 0.04fF
C11527 VP.n4547 a_400_38200# 0.08fF
C11528 VP.n4548 a_400_38200# 0.72fF
C11529 VP.n4549 a_400_38200# 0.09fF
C11530 VP.n4550 a_400_38200# 0.00fF
C11531 VP.n4551 a_400_38200# 0.98fF
C11532 VP.n4552 a_400_38200# 0.19fF
C11533 VP.n4554 a_400_38200# 1.72fF
C11534 VP.n4555 a_400_38200# 1.96fF
C11535 VP.n4556 a_400_38200# 1.04fF
C11536 VP.n4557 a_400_38200# 0.05fF
C11537 VP.n4558 a_400_38200# 0.03fF
C11538 VP.n4559 a_400_38200# 0.06fF
C11539 VP.n4560 a_400_38200# 0.06fF
C11540 VP.n4561 a_400_38200# 0.06fF
C11541 VP.n4562 a_400_38200# 0.07fF
C11542 VP.n4563 a_400_38200# 0.03fF
C11543 VP.n4564 a_400_38200# 0.05fF
C11544 VP.n4565 a_400_38200# 0.07fF
C11545 VP.n4566 a_400_38200# 0.19fF
C11546 VP.n4567 a_400_38200# 0.60fF
C11547 VP.n4568 a_400_38200# 0.76fF
C11548 VP.n4569 a_400_38200# 0.40fF
C11549 VP.n4570 a_400_38200# 0.03fF
C11550 VP.n4571 a_400_38200# 0.01fF
C11551 VP.t1311 a_400_38200# 0.02fF
C11552 VP.n4572 a_400_38200# 0.25fF
C11553 VP.t1169 a_400_38200# 0.02fF
C11554 VP.n4573 a_400_38200# 0.95fF
C11555 VP.n4574 a_400_38200# 0.70fF
C11556 VP.n4575 a_400_38200# 1.93fF
C11557 VP.n4576 a_400_38200# 2.97fF
C11558 VP.n4577 a_400_38200# 2.27fF
C11559 VP.t1212 a_400_38200# 0.02fF
C11560 VP.n4578 a_400_38200# 0.24fF
C11561 VP.n4579 a_400_38200# 0.35fF
C11562 VP.n4580 a_400_38200# 0.60fF
C11563 VP.t711 a_400_38200# 0.02fF
C11564 VP.n4581 a_400_38200# 0.12fF
C11565 VP.n4582 a_400_38200# 0.14fF
C11566 VP.n4584 a_400_38200# 0.12fF
C11567 VP.t627 a_400_38200# 0.02fF
C11568 VP.n4585 a_400_38200# 0.14fF
C11569 VP.n4587 a_400_38200# 0.04fF
C11570 VP.n4588 a_400_38200# 0.02fF
C11571 VP.n4589 a_400_38200# 0.06fF
C11572 VP.n4590 a_400_38200# 0.30fF
C11573 VP.n4591 a_400_38200# 0.10fF
C11574 VP.n4592 a_400_38200# 0.28fF
C11575 VP.n4593 a_400_38200# 0.06fF
C11576 VP.n4594 a_400_38200# 0.06fF
C11577 VP.n4595 a_400_38200# 0.03fF
C11578 VP.n4596 a_400_38200# 0.15fF
C11579 VP.n4597 a_400_38200# 0.08fF
C11580 VP.n4598 a_400_38200# 0.14fF
C11581 VP.n4599 a_400_38200# 0.03fF
C11582 VP.n4600 a_400_38200# 0.06fF
C11583 VP.n4601 a_400_38200# 0.06fF
C11584 VP.n4602 a_400_38200# 0.06fF
C11585 VP.n4603 a_400_38200# 0.06fF
C11586 VP.n4604 a_400_38200# 0.03fF
C11587 VP.n4605 a_400_38200# 0.05fF
C11588 VP.n4606 a_400_38200# 0.07fF
C11589 VP.n4607 a_400_38200# 0.19fF
C11590 VP.n4608 a_400_38200# 0.59fF
C11591 VP.n4609 a_400_38200# 0.34fF
C11592 VP.n4610 a_400_38200# 1.88fF
C11593 VP.t490 a_400_38200# 0.02fF
C11594 VP.n4611 a_400_38200# 0.24fF
C11595 VP.n4612 a_400_38200# 0.91fF
C11596 VP.n4613 a_400_38200# 0.05fF
C11597 VP.n4614 a_400_38200# 0.19fF
C11598 VP.n4615 a_400_38200# 0.10fF
C11599 VP.n4616 a_400_38200# 0.10fF
C11600 VP.n4617 a_400_38200# 0.18fF
C11601 VP.n4618 a_400_38200# 0.09fF
C11602 VP.n4619 a_400_38200# 0.04fF
C11603 VP.n4620 a_400_38200# 0.19fF
C11604 VP.n4621 a_400_38200# 0.26fF
C11605 VP.n4622 a_400_38200# 1.17fF
C11606 VP.n4623 a_400_38200# 0.06fF
C11607 VP.n4624 a_400_38200# 0.44fF
C11608 VP.n4625 a_400_38200# 0.13fF
C11609 VP.n4626 a_400_38200# 0.02fF
C11610 VP.n4627 a_400_38200# 1.81fF
C11611 VP.n4628 a_400_38200# 0.12fF
C11612 VP.t170 a_400_38200# 0.02fF
C11613 VP.n4629 a_400_38200# 0.14fF
C11614 VP.t765 a_400_38200# 0.02fF
C11615 VP.n4631 a_400_38200# 0.24fF
C11616 VP.n4632 a_400_38200# 0.35fF
C11617 VP.n4633 a_400_38200# 0.60fF
C11618 VP.n4634 a_400_38200# 3.18fF
C11619 VP.n4635 a_400_38200# 2.06fF
C11620 VP.n4636 a_400_38200# 1.98fF
C11621 VP.t1340 a_400_38200# 0.02fF
C11622 VP.n4637 a_400_38200# 0.24fF
C11623 VP.n4638 a_400_38200# 0.91fF
C11624 VP.n4639 a_400_38200# 0.05fF
C11625 VP.t265 a_400_38200# 0.02fF
C11626 VP.n4640 a_400_38200# 0.12fF
C11627 VP.n4641 a_400_38200# 0.14fF
C11628 VP.n4643 a_400_38200# 0.16fF
C11629 VP.n4644 a_400_38200# 0.19fF
C11630 VP.n4645 a_400_38200# 0.09fF
C11631 VP.n4646 a_400_38200# 0.04fF
C11632 VP.n4647 a_400_38200# 0.14fF
C11633 VP.n4648 a_400_38200# 0.64fF
C11634 VP.n4649 a_400_38200# 1.32fF
C11635 VP.n4650 a_400_38200# 1.81fF
C11636 VP.n4651 a_400_38200# 0.12fF
C11637 VP.t1019 a_400_38200# 0.02fF
C11638 VP.n4652 a_400_38200# 0.14fF
C11639 VP.t311 a_400_38200# 0.02fF
C11640 VP.n4654 a_400_38200# 0.24fF
C11641 VP.n4655 a_400_38200# 0.35fF
C11642 VP.n4656 a_400_38200# 0.60fF
C11643 VP.n4657 a_400_38200# 2.97fF
C11644 VP.n4658 a_400_38200# 2.27fF
C11645 VP.n4659 a_400_38200# 2.00fF
C11646 VP.t889 a_400_38200# 0.02fF
C11647 VP.n4660 a_400_38200# 0.24fF
C11648 VP.n4661 a_400_38200# 0.91fF
C11649 VP.n4662 a_400_38200# 0.05fF
C11650 VP.t1121 a_400_38200# 0.02fF
C11651 VP.n4663 a_400_38200# 0.12fF
C11652 VP.n4664 a_400_38200# 0.14fF
C11653 VP.n4666 a_400_38200# 0.24fF
C11654 VP.t23 a_400_38200# 0.02fF
C11655 VP.n4667 a_400_38200# 0.36fF
C11656 VP.n4668 a_400_38200# 0.36fF
C11657 VP.n4669 a_400_38200# 0.67fF
C11658 VP.n4670 a_400_38200# 0.16fF
C11659 VP.n4671 a_400_38200# 0.19fF
C11660 VP.n4672 a_400_38200# 0.09fF
C11661 VP.n4673 a_400_38200# 0.04fF
C11662 VP.n4674 a_400_38200# 0.14fF
C11663 VP.n4675 a_400_38200# 0.64fF
C11664 VP.n4676 a_400_38200# 1.32fF
C11665 VP.n4677 a_400_38200# 1.81fF
C11666 VP.n4678 a_400_38200# 2.97fF
C11667 VP.n4679 a_400_38200# 2.27fF
C11668 VP.n4680 a_400_38200# 0.75fF
C11669 VP.n4681 a_400_38200# 0.24fF
C11670 VP.t789 a_400_38200# 0.02fF
C11671 VP.n4682 a_400_38200# 0.35fF
C11672 VP.n4683 a_400_38200# 0.63fF
C11673 VP.n4684 a_400_38200# 0.40fF
C11674 VP.n4685 a_400_38200# 0.40fF
C11675 VP.n4686 a_400_38200# 0.12fF
C11676 VP.t199 a_400_38200# 0.02fF
C11677 VP.n4687 a_400_38200# 0.14fF
C11678 VP.t229 a_400_38200# 0.02fF
C11679 VP.n4689 a_400_38200# 0.12fF
C11680 VP.n4690 a_400_38200# 0.14fF
C11681 VP.n4692 a_400_38200# 0.09fF
C11682 VP.n4693 a_400_38200# 0.03fF
C11683 VP.n4694 a_400_38200# 0.04fF
C11684 VP.n4695 a_400_38200# 0.37fF
C11685 VP.n4696 a_400_38200# 0.11fF
C11686 VP.n4697 a_400_38200# 0.05fF
C11687 VP.n4698 a_400_38200# 0.08fF
C11688 VP.n4699 a_400_38200# 0.10fF
C11689 VP.n4700 a_400_38200# 0.06fF
C11690 VP.n4701 a_400_38200# 0.08fF
C11691 VP.n4702 a_400_38200# 0.19fF
C11692 VP.n4703 a_400_38200# 0.06fF
C11693 VP.n4704 a_400_38200# 0.15fF
C11694 VP.n4705 a_400_38200# 0.14fF
C11695 VP.n4706 a_400_38200# 0.13fF
C11696 VP.n4707 a_400_38200# 0.12fF
C11697 VP.n4708 a_400_38200# 0.05fF
C11698 VP.n4709 a_400_38200# 0.17fF
C11699 VP.n4710 a_400_38200# 0.26fF
C11700 VP.n4711 a_400_38200# 0.37fF
C11701 VP.n4712 a_400_38200# 0.27fF
C11702 VP.n4713 a_400_38200# 2.05fF
C11703 VP.n4714 a_400_38200# 0.12fF
C11704 VP.t1294 a_400_38200# 0.02fF
C11705 VP.n4715 a_400_38200# 0.14fF
C11706 VP.t579 a_400_38200# 0.02fF
C11707 VP.n4717 a_400_38200# 0.24fF
C11708 VP.n4718 a_400_38200# 0.35fF
C11709 VP.n4719 a_400_38200# 0.60fF
C11710 VP.n4720 a_400_38200# 2.87fF
C11711 VP.n4721 a_400_38200# 2.00fF
C11712 VP.t1151 a_400_38200# 0.02fF
C11713 VP.n4722 a_400_38200# 0.24fF
C11714 VP.n4723 a_400_38200# 0.91fF
C11715 VP.n4724 a_400_38200# 0.05fF
C11716 VP.t640 a_400_38200# 0.02fF
C11717 VP.n4725 a_400_38200# 0.12fF
C11718 VP.n4726 a_400_38200# 0.14fF
C11719 VP.n4728 a_400_38200# 15.28fF
C11720 VP.n4729 a_400_38200# 0.10fF
C11721 VP.n4730 a_400_38200# 0.28fF
C11722 VP.n4731 a_400_38200# 0.06fF
C11723 VP.n4732 a_400_38200# 0.06fF
C11724 VP.n4733 a_400_38200# 0.03fF
C11725 VP.n4734 a_400_38200# 0.15fF
C11726 VP.n4735 a_400_38200# 0.08fF
C11727 VP.n4736 a_400_38200# 0.14fF
C11728 VP.n4737 a_400_38200# 0.03fF
C11729 VP.n4738 a_400_38200# 0.06fF
C11730 VP.n4739 a_400_38200# 0.06fF
C11731 VP.n4740 a_400_38200# 0.06fF
C11732 VP.n4741 a_400_38200# 0.06fF
C11733 VP.n4742 a_400_38200# 0.03fF
C11734 VP.n4743 a_400_38200# 0.05fF
C11735 VP.n4744 a_400_38200# 0.07fF
C11736 VP.n4745 a_400_38200# 0.19fF
C11737 VP.n4746 a_400_38200# 0.59fF
C11738 VP.n4747 a_400_38200# 0.34fF
C11739 VP.n4748 a_400_38200# 0.04fF
C11740 VP.n4749 a_400_38200# 0.02fF
C11741 VP.n4750 a_400_38200# 0.06fF
C11742 VP.n4751 a_400_38200# 0.30fF
C11743 VP.n4752 a_400_38200# 1.93fF
C11744 VP.n4753 a_400_38200# 0.12fF
C11745 VP.t863 a_400_38200# 0.02fF
C11746 VP.n4754 a_400_38200# 0.14fF
C11747 VP.t132 a_400_38200# 0.02fF
C11748 VP.n4756 a_400_38200# 0.24fF
C11749 VP.n4757 a_400_38200# 0.35fF
C11750 VP.n4758 a_400_38200# 0.60fF
C11751 VP.n4759 a_400_38200# 0.07fF
C11752 VP.n4760 a_400_38200# 0.72fF
C11753 VP.n4761 a_400_38200# 0.20fF
C11754 VP.n4762 a_400_38200# 0.19fF
C11755 VP.n4763 a_400_38200# 0.10fF
C11756 VP.n4764 a_400_38200# 0.11fF
C11757 VP.n4765 a_400_38200# 0.09fF
C11758 VP.n4766 a_400_38200# 0.16fF
C11759 VP.n4767 a_400_38200# 0.10fF
C11760 VP.n4768 a_400_38200# 0.11fF
C11761 VP.n4769 a_400_38200# 0.19fF
C11762 VP.n4770 a_400_38200# 0.20fF
C11763 VP.n4771 a_400_38200# 0.98fF
C11764 VP.n4772 a_400_38200# 0.15fF
C11765 VP.n4774 a_400_38200# 1.72fF
C11766 VP.t904 a_400_38200# 0.02fF
C11767 VP.n4775 a_400_38200# 0.12fF
C11768 VP.n4776 a_400_38200# 0.14fF
C11769 VP.t717 a_400_38200# 0.02fF
C11770 VP.n4778 a_400_38200# 0.24fF
C11771 VP.n4779 a_400_38200# 0.91fF
C11772 VP.n4780 a_400_38200# 0.05fF
C11773 VP.n4781 a_400_38200# 0.10fF
C11774 VP.n4782 a_400_38200# 0.06fF
C11775 VP.n4783 a_400_38200# 0.06fF
C11776 VP.n4784 a_400_38200# 0.28fF
C11777 VP.n4785 a_400_38200# 0.03fF
C11778 VP.n4786 a_400_38200# 0.15fF
C11779 VP.n4787 a_400_38200# 0.08fF
C11780 VP.n4788 a_400_38200# 0.14fF
C11781 VP.n4789 a_400_38200# 0.03fF
C11782 VP.n4790 a_400_38200# 0.06fF
C11783 VP.n4791 a_400_38200# 0.06fF
C11784 VP.n4792 a_400_38200# 0.06fF
C11785 VP.n4793 a_400_38200# 0.06fF
C11786 VP.n4794 a_400_38200# 0.03fF
C11787 VP.n4795 a_400_38200# 0.05fF
C11788 VP.n4796 a_400_38200# 0.07fF
C11789 VP.n4797 a_400_38200# 0.19fF
C11790 VP.n4798 a_400_38200# 0.59fF
C11791 VP.n4799 a_400_38200# 0.34fF
C11792 VP.n4800 a_400_38200# 0.04fF
C11793 VP.n4801 a_400_38200# 0.02fF
C11794 VP.n4802 a_400_38200# 0.06fF
C11795 VP.n4803 a_400_38200# 0.30fF
C11796 VP.n4804 a_400_38200# 1.93fF
C11797 VP.n4805 a_400_38200# 0.12fF
C11798 VP.t417 a_400_38200# 0.02fF
C11799 VP.n4806 a_400_38200# 0.14fF
C11800 VP.t998 a_400_38200# 0.02fF
C11801 VP.n4808 a_400_38200# 0.24fF
C11802 VP.n4809 a_400_38200# 0.35fF
C11803 VP.n4810 a_400_38200# 0.60fF
C11804 VP.n4811 a_400_38200# 0.72fF
C11805 VP.n4812 a_400_38200# 1.24fF
C11806 VP.n4813 a_400_38200# 0.54fF
C11807 VP.n4814 a_400_38200# 0.22fF
C11808 VP.n4815 a_400_38200# 1.73fF
C11809 VP.t452 a_400_38200# 0.02fF
C11810 VP.n4816 a_400_38200# 0.12fF
C11811 VP.n4817 a_400_38200# 0.14fF
C11812 VP.t271 a_400_38200# 0.02fF
C11813 VP.n4819 a_400_38200# 0.24fF
C11814 VP.n4820 a_400_38200# 0.91fF
C11815 VP.n4821 a_400_38200# 0.05fF
C11816 VP.n4822 a_400_38200# 0.10fF
C11817 VP.n4823 a_400_38200# 0.06fF
C11818 VP.n4824 a_400_38200# 0.06fF
C11819 VP.n4825 a_400_38200# 0.28fF
C11820 VP.n4826 a_400_38200# 0.03fF
C11821 VP.n4827 a_400_38200# 0.15fF
C11822 VP.n4828 a_400_38200# 0.08fF
C11823 VP.n4829 a_400_38200# 0.14fF
C11824 VP.n4830 a_400_38200# 0.03fF
C11825 VP.n4831 a_400_38200# 0.06fF
C11826 VP.n4832 a_400_38200# 0.06fF
C11827 VP.n4833 a_400_38200# 0.06fF
C11828 VP.n4834 a_400_38200# 0.06fF
C11829 VP.n4835 a_400_38200# 0.03fF
C11830 VP.n4836 a_400_38200# 0.05fF
C11831 VP.n4837 a_400_38200# 0.07fF
C11832 VP.n4838 a_400_38200# 0.19fF
C11833 VP.n4839 a_400_38200# 0.59fF
C11834 VP.n4840 a_400_38200# 0.34fF
C11835 VP.n4841 a_400_38200# 0.04fF
C11836 VP.n4842 a_400_38200# 0.02fF
C11837 VP.n4843 a_400_38200# 0.06fF
C11838 VP.n4844 a_400_38200# 0.30fF
C11839 VP.n4845 a_400_38200# 1.93fF
C11840 VP.n4846 a_400_38200# 0.12fF
C11841 VP.t665 a_400_38200# 0.02fF
C11842 VP.n4847 a_400_38200# 0.14fF
C11843 VP.t1252 a_400_38200# 0.02fF
C11844 VP.n4849 a_400_38200# 0.24fF
C11845 VP.n4850 a_400_38200# 0.35fF
C11846 VP.n4851 a_400_38200# 0.60fF
C11847 VP.n4852 a_400_38200# 0.72fF
C11848 VP.n4853 a_400_38200# 1.24fF
C11849 VP.n4854 a_400_38200# 0.54fF
C11850 VP.n4855 a_400_38200# 0.22fF
C11851 VP.n4856 a_400_38200# 1.73fF
C11852 VP.t1302 a_400_38200# 0.02fF
C11853 VP.n4857 a_400_38200# 0.12fF
C11854 VP.n4858 a_400_38200# 0.14fF
C11855 VP.t526 a_400_38200# 0.02fF
C11856 VP.n4860 a_400_38200# 0.24fF
C11857 VP.n4861 a_400_38200# 0.91fF
C11858 VP.n4862 a_400_38200# 0.05fF
C11859 VP.n4863 a_400_38200# 0.10fF
C11860 VP.n4864 a_400_38200# 0.28fF
C11861 VP.n4865 a_400_38200# 0.06fF
C11862 VP.n4866 a_400_38200# 0.06fF
C11863 VP.n4867 a_400_38200# 0.03fF
C11864 VP.n4868 a_400_38200# 0.15fF
C11865 VP.n4869 a_400_38200# 0.08fF
C11866 VP.n4870 a_400_38200# 0.14fF
C11867 VP.n4871 a_400_38200# 0.03fF
C11868 VP.n4872 a_400_38200# 0.06fF
C11869 VP.n4873 a_400_38200# 0.06fF
C11870 VP.n4874 a_400_38200# 0.06fF
C11871 VP.n4875 a_400_38200# 0.06fF
C11872 VP.n4876 a_400_38200# 0.03fF
C11873 VP.n4877 a_400_38200# 0.05fF
C11874 VP.n4878 a_400_38200# 0.07fF
C11875 VP.n4879 a_400_38200# 0.19fF
C11876 VP.n4880 a_400_38200# 0.59fF
C11877 VP.n4881 a_400_38200# 0.34fF
C11878 VP.n4882 a_400_38200# 0.04fF
C11879 VP.n4883 a_400_38200# 0.02fF
C11880 VP.n4884 a_400_38200# 0.06fF
C11881 VP.n4885 a_400_38200# 0.30fF
C11882 VP.n4886 a_400_38200# 1.93fF
C11883 VP.n4887 a_400_38200# 0.12fF
C11884 VP.t218 a_400_38200# 0.02fF
C11885 VP.n4888 a_400_38200# 0.14fF
C11886 VP.t807 a_400_38200# 0.02fF
C11887 VP.n4890 a_400_38200# 0.24fF
C11888 VP.n4891 a_400_38200# 0.35fF
C11889 VP.n4892 a_400_38200# 0.60fF
C11890 VP.n4893 a_400_38200# 0.72fF
C11891 VP.n4894 a_400_38200# 1.24fF
C11892 VP.n4895 a_400_38200# 0.54fF
C11893 VP.n4896 a_400_38200# 0.22fF
C11894 VP.n4897 a_400_38200# 1.73fF
C11895 VP.t317 a_400_38200# 0.02fF
C11896 VP.n4898 a_400_38200# 0.12fF
C11897 VP.n4899 a_400_38200# 0.14fF
C11898 VP.t47 a_400_38200# 0.02fF
C11899 VP.n4901 a_400_38200# 0.24fF
C11900 VP.n4902 a_400_38200# 0.91fF
C11901 VP.n4903 a_400_38200# 0.05fF
C11902 VP.n4904 a_400_38200# 0.10fF
C11903 VP.n4905 a_400_38200# 0.06fF
C11904 VP.n4906 a_400_38200# 0.06fF
C11905 VP.n4907 a_400_38200# 0.28fF
C11906 VP.n4908 a_400_38200# 0.03fF
C11907 VP.n4909 a_400_38200# 0.15fF
C11908 VP.n4910 a_400_38200# 0.08fF
C11909 VP.n4911 a_400_38200# 0.14fF
C11910 VP.n4912 a_400_38200# 0.03fF
C11911 VP.n4913 a_400_38200# 0.06fF
C11912 VP.n4914 a_400_38200# 0.06fF
C11913 VP.n4915 a_400_38200# 0.06fF
C11914 VP.n4916 a_400_38200# 0.06fF
C11915 VP.n4917 a_400_38200# 0.03fF
C11916 VP.n4918 a_400_38200# 0.05fF
C11917 VP.n4919 a_400_38200# 0.07fF
C11918 VP.n4920 a_400_38200# 0.19fF
C11919 VP.n4921 a_400_38200# 0.59fF
C11920 VP.n4922 a_400_38200# 0.34fF
C11921 VP.n4923 a_400_38200# 0.04fF
C11922 VP.n4924 a_400_38200# 0.02fF
C11923 VP.n4925 a_400_38200# 0.06fF
C11924 VP.n4926 a_400_38200# 0.30fF
C11925 VP.n4927 a_400_38200# 1.93fF
C11926 VP.n4928 a_400_38200# 0.12fF
C11927 VP.t1072 a_400_38200# 0.02fF
C11928 VP.n4929 a_400_38200# 0.14fF
C11929 VP.t358 a_400_38200# 0.02fF
C11930 VP.n4931 a_400_38200# 0.24fF
C11931 VP.n4932 a_400_38200# 0.35fF
C11932 VP.n4933 a_400_38200# 0.60fF
C11933 VP.n4934 a_400_38200# 0.71fF
C11934 VP.n4935 a_400_38200# 1.39fF
C11935 VP.n4936 a_400_38200# 0.54fF
C11936 VP.n4937 a_400_38200# 0.21fF
C11937 VP.n4938 a_400_38200# 1.73fF
C11938 VP.t1160 a_400_38200# 0.02fF
C11939 VP.n4939 a_400_38200# 0.12fF
C11940 VP.n4940 a_400_38200# 0.14fF
C11941 VP.t936 a_400_38200# 0.02fF
C11942 VP.n4942 a_400_38200# 0.24fF
C11943 VP.n4943 a_400_38200# 0.91fF
C11944 VP.n4944 a_400_38200# 0.05fF
C11945 VP.n4945 a_400_38200# 0.06fF
C11946 VP.n4946 a_400_38200# 0.06fF
C11947 VP.n4947 a_400_38200# 0.03fF
C11948 VP.n4948 a_400_38200# 0.10fF
C11949 VP.n4949 a_400_38200# 0.17fF
C11950 VP.n4950 a_400_38200# 0.10fF
C11951 VP.n4951 a_400_38200# 0.13fF
C11952 VP.n4952 a_400_38200# 0.02fF
C11953 VP.n4953 a_400_38200# 0.04fF
C11954 VP.n4954 a_400_38200# 0.06fF
C11955 VP.n4955 a_400_38200# 0.09fF
C11956 VP.n4956 a_400_38200# 0.10fF
C11957 VP.n4957 a_400_38200# 0.05fF
C11958 VP.n4958 a_400_38200# 0.19fF
C11959 VP.n4959 a_400_38200# 0.16fF
C11960 VP.n4960 a_400_38200# 0.04fF
C11961 VP.n4961 a_400_38200# 0.05fF
C11962 VP.n4962 a_400_38200# 0.04fF
C11963 VP.n4963 a_400_38200# 0.12fF
C11964 VP.n4964 a_400_38200# 0.09fF
C11965 VP.n4965 a_400_38200# 0.14fF
C11966 VP.n4966 a_400_38200# 0.56fF
C11967 VP.n4967 a_400_38200# 0.10fF
C11968 VP.n4968 a_400_38200# 1.93fF
C11969 VP.n4969 a_400_38200# 0.12fF
C11970 VP.t647 a_400_38200# 0.02fF
C11971 VP.n4970 a_400_38200# 0.14fF
C11972 VP.t1156 a_400_38200# 0.02fF
C11973 VP.n4972 a_400_38200# 0.24fF
C11974 VP.n4973 a_400_38200# 0.35fF
C11975 VP.n4974 a_400_38200# 0.60fF
C11976 VP.n4975 a_400_38200# 2.23fF
C11977 VP.n4976 a_400_38200# 0.18fF
C11978 VP.n4977 a_400_38200# 0.45fF
C11979 VP.n4978 a_400_38200# 0.06fF
C11980 VP.n4979 a_400_38200# 0.01fF
C11981 VP.n4980 a_400_38200# 0.01fF
C11982 VP.n4981 a_400_38200# 0.04fF
C11983 VP.n4982 a_400_38200# 0.02fF
C11984 VP.n4983 a_400_38200# 0.07fF
C11985 VP.n4984 a_400_38200# 0.04fF
C11986 VP.n4985 a_400_38200# 0.14fF
C11987 VP.n4986 a_400_38200# 0.45fF
C11988 VP.n4987 a_400_38200# 1.46fF
C11989 VP.n4988 a_400_38200# 1.78fF
C11990 VP.t675 a_400_38200# 0.02fF
C11991 VP.n4989 a_400_38200# 0.12fF
C11992 VP.n4990 a_400_38200# 0.14fF
C11993 VP.t439 a_400_38200# 0.02fF
C11994 VP.n4992 a_400_38200# 0.24fF
C11995 VP.n4993 a_400_38200# 0.91fF
C11996 VP.n4994 a_400_38200# 0.05fF
C11997 VP.n4995 a_400_38200# 1.93fF
C11998 VP.n4996 a_400_38200# 2.72fF
C11999 VP.n4997 a_400_38200# 0.18fF
C12000 VP.n4998 a_400_38200# 0.45fF
C12001 VP.n4999 a_400_38200# 0.06fF
C12002 VP.n5000 a_400_38200# 0.01fF
C12003 VP.n5001 a_400_38200# 0.01fF
C12004 VP.n5002 a_400_38200# 0.04fF
C12005 VP.n5003 a_400_38200# 0.02fF
C12006 VP.n5004 a_400_38200# 0.07fF
C12007 VP.n5005 a_400_38200# 0.04fF
C12008 VP.n5006 a_400_38200# 0.14fF
C12009 VP.n5007 a_400_38200# 0.53fF
C12010 VP.n5008 a_400_38200# 1.62fF
C12011 VP.t343 a_400_38200# 0.02fF
C12012 VP.n5009 a_400_38200# 0.24fF
C12013 VP.n5010 a_400_38200# 0.35fF
C12014 VP.n5011 a_400_38200# 0.60fF
C12015 VP.n5012 a_400_38200# 0.12fF
C12016 VP.t1052 a_400_38200# 0.02fF
C12017 VP.n5013 a_400_38200# 0.14fF
C12018 VP.n5015 a_400_38200# 0.10fF
C12019 VP.n5016 a_400_38200# 0.17fF
C12020 VP.n5017 a_400_38200# 0.06fF
C12021 VP.n5018 a_400_38200# 0.06fF
C12022 VP.n5019 a_400_38200# 0.03fF
C12023 VP.n5020 a_400_38200# 0.10fF
C12024 VP.n5021 a_400_38200# 0.13fF
C12025 VP.n5022 a_400_38200# 0.14fF
C12026 VP.n5023 a_400_38200# 0.04fF
C12027 VP.n5024 a_400_38200# 0.02fF
C12028 VP.n5025 a_400_38200# 0.03fF
C12029 VP.n5026 a_400_38200# 0.03fF
C12030 VP.n5027 a_400_38200# 0.05fF
C12031 VP.n5028 a_400_38200# 0.03fF
C12032 VP.n5029 a_400_38200# 0.04fF
C12033 VP.n5030 a_400_38200# 0.20fF
C12034 VP.n5031 a_400_38200# 0.14fF
C12035 VP.n5032 a_400_38200# 0.02fF
C12036 VP.n5033 a_400_38200# 0.07fF
C12037 VP.n5034 a_400_38200# 0.13fF
C12038 VP.n5035 a_400_38200# 0.04fF
C12039 VP.n5036 a_400_38200# 0.02fF
C12040 VP.n5037 a_400_38200# 0.06fF
C12041 VP.n5038 a_400_38200# 0.55fF
C12042 VP.n5039 a_400_38200# 0.10fF
C12043 VP.n5040 a_400_38200# 1.95fF
C12044 VP.t1083 a_400_38200# 0.02fF
C12045 VP.n5041 a_400_38200# 0.12fF
C12046 VP.n5042 a_400_38200# 0.14fF
C12047 VP.t920 a_400_38200# 0.02fF
C12048 VP.n5044 a_400_38200# 0.24fF
C12049 VP.n5045 a_400_38200# 0.91fF
C12050 VP.n5046 a_400_38200# 0.05fF
C12051 VP.t169 a_400_38200# 35.17fF
C12052 VP.t599 a_400_38200# 0.02fF
C12053 VP.n5047 a_400_38200# 1.21fF
C12054 VP.n5048 a_400_38200# 0.25fF
C12055 VP.n5049 a_400_38200# 26.29fF
C12056 VP.n5050 a_400_38200# 26.29fF
C12057 VP.n5051 a_400_38200# 0.76fF
C12058 VP.n5052 a_400_38200# 0.27fF
C12059 VP.n5053 a_400_38200# 0.59fF
C12060 VP.n5054 a_400_38200# 0.10fF
C12061 VP.n5055 a_400_38200# 3.02fF
C12062 VP.t131 a_400_38200# 15.72fF
C12063 VP.n5056 a_400_38200# 1.15fF
C12064 VP.n5058 a_400_38200# 13.70fF
C12065 VP.n5060 a_400_38200# 1.99fF
C12066 VP.n5061 a_400_38200# 4.39fF
C12067 VP.n5062 a_400_38200# 0.03fF
C12068 VP.n5063 a_400_38200# 0.05fF
C12069 VP.n5064 a_400_38200# 0.07fF
C12070 VP.n5065 a_400_38200# 0.03fF
C12071 VP.n5066 a_400_38200# 0.06fF
C12072 VP.n5067 a_400_38200# 0.06fF
C12073 VP.n5068 a_400_38200# 0.06fF
C12074 VP.n5069 a_400_38200# 0.07fF
C12075 VP.n5070 a_400_38200# 0.57fF
C12076 VP.n5071 a_400_38200# 1.88fF
C12077 VP.n5072 a_400_38200# 0.92fF
C12078 VP.n5073 a_400_38200# 2.63fF
C12079 VP.n5074 a_400_38200# 0.10fF
C12080 VP.n5075 a_400_38200# 0.28fF
C12081 VP.n5076 a_400_38200# 0.15fF
C12082 VP.n5077 a_400_38200# 0.08fF
C12083 VP.n5078 a_400_38200# 0.14fF
C12084 VP.n5079 a_400_38200# 0.06fF
C12085 VP.n5080 a_400_38200# 0.06fF
C12086 VP.n5081 a_400_38200# 0.03fF
C12087 VP.n5082 a_400_38200# 0.05fF
C12088 VP.n5083 a_400_38200# 0.07fF
C12089 VP.n5084 a_400_38200# 0.19fF
C12090 VP.n5085 a_400_38200# 0.59fF
C12091 VP.n5086 a_400_38200# 0.34fF
C12092 VP.n5087 a_400_38200# 0.04fF
C12093 VP.n5088 a_400_38200# 0.02fF
C12094 VP.n5089 a_400_38200# 0.06fF
C12095 VP.n5090 a_400_38200# 0.30fF
C12096 VP.n5091 a_400_38200# 0.12fF
C12097 VP.t173 a_400_38200# 0.02fF
C12098 VP.n5092 a_400_38200# 0.14fF
C12099 VP.n5094 a_400_38200# 1.93fF
C12100 VP.t580 a_400_38200# 0.02fF
C12101 VP.n5095 a_400_38200# 0.24fF
C12102 VP.n5096 a_400_38200# 0.35fF
C12103 VP.n5097 a_400_38200# 0.60fF
C12104 VP.n5098 a_400_38200# 0.12fF
C12105 VP.t1297 a_400_38200# 0.02fF
C12106 VP.n5099 a_400_38200# 0.14fF
C12107 VP.n5101 a_400_38200# 0.04fF
C12108 VP.n5102 a_400_38200# 0.02fF
C12109 VP.n5103 a_400_38200# 0.06fF
C12110 VP.n5104 a_400_38200# 0.30fF
C12111 VP.n5105 a_400_38200# 0.10fF
C12112 VP.n5106 a_400_38200# 0.28fF
C12113 VP.n5107 a_400_38200# 0.15fF
C12114 VP.n5108 a_400_38200# 0.08fF
C12115 VP.n5109 a_400_38200# 0.14fF
C12116 VP.n5110 a_400_38200# 0.06fF
C12117 VP.n5111 a_400_38200# 0.06fF
C12118 VP.n5112 a_400_38200# 0.03fF
C12119 VP.n5113 a_400_38200# 0.05fF
C12120 VP.n5114 a_400_38200# 0.07fF
C12121 VP.n5115 a_400_38200# 0.19fF
C12122 VP.n5116 a_400_38200# 0.59fF
C12123 VP.n5117 a_400_38200# 0.34fF
C12124 VP.n5118 a_400_38200# 2.18fF
C12125 VP.t139 a_400_38200# 0.02fF
C12126 VP.n5119 a_400_38200# 0.24fF
C12127 VP.n5120 a_400_38200# 0.91fF
C12128 VP.n5121 a_400_38200# 0.05fF
C12129 VP.t351 a_400_38200# 0.02fF
C12130 VP.n5122 a_400_38200# 0.12fF
C12131 VP.n5123 a_400_38200# 0.14fF
C12132 VP.n5125 a_400_38200# 0.10fF
C12133 VP.n5126 a_400_38200# 0.10fF
C12134 VP.n5127 a_400_38200# 0.18fF
C12135 VP.n5128 a_400_38200# 0.09fF
C12136 VP.n5129 a_400_38200# 0.04fF
C12137 VP.n5130 a_400_38200# 0.26fF
C12138 VP.n5131 a_400_38200# 1.17fF
C12139 VP.n5132 a_400_38200# 0.06fF
C12140 VP.n5133 a_400_38200# 0.44fF
C12141 VP.n5134 a_400_38200# 0.13fF
C12142 VP.n5135 a_400_38200# 0.02fF
C12143 VP.n5136 a_400_38200# 1.81fF
C12144 VP.n5137 a_400_38200# 0.12fF
C12145 VP.t852 a_400_38200# 0.02fF
C12146 VP.n5138 a_400_38200# 0.14fF
C12147 VP.t114 a_400_38200# 0.02fF
C12148 VP.n5140 a_400_38200# 0.24fF
C12149 VP.n5141 a_400_38200# 0.35fF
C12150 VP.n5142 a_400_38200# 0.60fF
C12151 VP.n5143 a_400_38200# 2.28fF
C12152 VP.t1002 a_400_38200# 0.02fF
C12153 VP.n5144 a_400_38200# 0.24fF
C12154 VP.n5145 a_400_38200# 0.91fF
C12155 VP.n5146 a_400_38200# 0.05fF
C12156 VP.t1202 a_400_38200# 0.02fF
C12157 VP.n5147 a_400_38200# 0.12fF
C12158 VP.n5148 a_400_38200# 0.14fF
C12159 VP.n5150 a_400_38200# 0.06fF
C12160 VP.n5151 a_400_38200# 0.09fF
C12161 VP.n5152 a_400_38200# 0.09fF
C12162 VP.n5153 a_400_38200# 1.45fF
C12163 VP.n5154 a_400_38200# 0.14fF
C12164 VP.n5155 a_400_38200# 0.07fF
C12165 VP.n5156 a_400_38200# 0.72fF
C12166 VP.n5157 a_400_38200# 1.81fF
C12167 VP.n5158 a_400_38200# 0.12fF
C12168 VP.t403 a_400_38200# 0.02fF
C12169 VP.n5159 a_400_38200# 0.14fF
C12170 VP.t987 a_400_38200# 0.02fF
C12171 VP.n5161 a_400_38200# 0.24fF
C12172 VP.n5162 a_400_38200# 0.35fF
C12173 VP.n5163 a_400_38200# 0.60fF
C12174 VP.n5164 a_400_38200# 2.30fF
C12175 VP.t559 a_400_38200# 0.02fF
C12176 VP.n5165 a_400_38200# 0.24fF
C12177 VP.n5166 a_400_38200# 0.91fF
C12178 VP.n5167 a_400_38200# 0.05fF
C12179 VP.t752 a_400_38200# 0.02fF
C12180 VP.n5168 a_400_38200# 0.12fF
C12181 VP.n5169 a_400_38200# 0.14fF
C12182 VP.n5171 a_400_38200# 0.06fF
C12183 VP.n5172 a_400_38200# 0.25fF
C12184 VP.n5173 a_400_38200# 0.45fF
C12185 VP.n5174 a_400_38200# 0.03fF
C12186 VP.n5175 a_400_38200# 0.05fF
C12187 VP.n5176 a_400_38200# 0.07fF
C12188 VP.n5177 a_400_38200# 0.06fF
C12189 VP.n5178 a_400_38200# 0.06fF
C12190 VP.n5179 a_400_38200# 0.19fF
C12191 VP.n5180 a_400_38200# 0.59fF
C12192 VP.n5181 a_400_38200# 0.34fF
C12193 VP.n5182 a_400_38200# 0.05fF
C12194 VP.n5183 a_400_38200# 0.30fF
C12195 VP.n5184 a_400_38200# 1.93fF
C12196 VP.n5185 a_400_38200# 0.12fF
C12197 VP.t1257 a_400_38200# 0.02fF
C12198 VP.n5186 a_400_38200# 0.14fF
C12199 VP.t540 a_400_38200# 0.02fF
C12200 VP.n5188 a_400_38200# 0.24fF
C12201 VP.n5189 a_400_38200# 0.35fF
C12202 VP.n5190 a_400_38200# 0.60fF
C12203 VP.n5191 a_400_38200# 2.04fF
C12204 VP.t87 a_400_38200# 0.02fF
C12205 VP.n5192 a_400_38200# 0.24fF
C12206 VP.n5193 a_400_38200# 0.91fF
C12207 VP.n5194 a_400_38200# 0.05fF
C12208 VP.t297 a_400_38200# 0.02fF
C12209 VP.n5195 a_400_38200# 0.12fF
C12210 VP.n5196 a_400_38200# 0.14fF
C12211 VP.n5198 a_400_38200# 0.24fF
C12212 VP.t965 a_400_38200# 0.02fF
C12213 VP.n5199 a_400_38200# 0.36fF
C12214 VP.n5200 a_400_38200# 0.36fF
C12215 VP.n5201 a_400_38200# 0.67fF
C12216 VP.n5202 a_400_38200# 0.06fF
C12217 VP.n5203 a_400_38200# 0.09fF
C12218 VP.n5204 a_400_38200# 0.09fF
C12219 VP.n5205 a_400_38200# 1.45fF
C12220 VP.n5206 a_400_38200# 0.14fF
C12221 VP.n5207 a_400_38200# 0.07fF
C12222 VP.n5208 a_400_38200# 0.72fF
C12223 VP.n5209 a_400_38200# 1.81fF
C12224 VP.n5210 a_400_38200# 1.06fF
C12225 VP.n5211 a_400_38200# 0.24fF
C12226 VP.t64 a_400_38200# 0.02fF
C12227 VP.n5212 a_400_38200# 0.35fF
C12228 VP.n5213 a_400_38200# 0.63fF
C12229 VP.n5214 a_400_38200# 0.40fF
C12230 VP.n5215 a_400_38200# 0.40fF
C12231 VP.n5216 a_400_38200# 0.12fF
C12232 VP.t813 a_400_38200# 0.02fF
C12233 VP.n5217 a_400_38200# 0.14fF
C12234 VP.t1224 a_400_38200# 0.02fF
C12235 VP.n5219 a_400_38200# 0.12fF
C12236 VP.n5220 a_400_38200# 0.14fF
C12237 VP.n5222 a_400_38200# 1.93fF
C12238 VP.t947 a_400_38200# 0.02fF
C12239 VP.n5223 a_400_38200# 0.24fF
C12240 VP.n5224 a_400_38200# 0.35fF
C12241 VP.n5225 a_400_38200# 0.60fF
C12242 VP.n5226 a_400_38200# 0.12fF
C12243 VP.t362 a_400_38200# 0.02fF
C12244 VP.n5227 a_400_38200# 0.14fF
C12245 VP.n5229 a_400_38200# 0.07fF
C12246 VP.n5230 a_400_38200# 0.30fF
C12247 VP.n5231 a_400_38200# 0.06fF
C12248 VP.n5232 a_400_38200# 0.25fF
C12249 VP.n5233 a_400_38200# 0.45fF
C12250 VP.n5234 a_400_38200# 0.06fF
C12251 VP.n5235 a_400_38200# 0.06fF
C12252 VP.n5236 a_400_38200# 0.03fF
C12253 VP.n5237 a_400_38200# 0.05fF
C12254 VP.n5238 a_400_38200# 0.07fF
C12255 VP.n5239 a_400_38200# 0.19fF
C12256 VP.n5240 a_400_38200# 0.59fF
C12257 VP.n5241 a_400_38200# 0.34fF
C12258 VP.n5242 a_400_38200# 2.04fF
C12259 VP.t517 a_400_38200# 0.02fF
C12260 VP.n5243 a_400_38200# 0.24fF
C12261 VP.n5244 a_400_38200# 0.91fF
C12262 VP.n5245 a_400_38200# 0.05fF
C12263 VP.t779 a_400_38200# 0.02fF
C12264 VP.n5246 a_400_38200# 0.12fF
C12265 VP.n5247 a_400_38200# 0.14fF
C12266 VP.n5249 a_400_38200# 1.81fF
C12267 VP.t501 a_400_38200# 0.02fF
C12268 VP.n5250 a_400_38200# 0.24fF
C12269 VP.n5251 a_400_38200# 0.35fF
C12270 VP.n5252 a_400_38200# 0.60fF
C12271 VP.n5253 a_400_38200# 0.12fF
C12272 VP.t1218 a_400_38200# 0.02fF
C12273 VP.n5254 a_400_38200# 0.14fF
C12274 VP.n5256 a_400_38200# 0.03fF
C12275 VP.n5257 a_400_38200# 0.09fF
C12276 VP.n5258 a_400_38200# 0.09fF
C12277 VP.n5259 a_400_38200# 0.05fF
C12278 VP.n5260 a_400_38200# 0.11fF
C12279 VP.n5261 a_400_38200# 0.09fF
C12280 VP.n5262 a_400_38200# 0.02fF
C12281 VP.n5263 a_400_38200# 0.03fF
C12282 VP.n5264 a_400_38200# 0.11fF
C12283 VP.n5265 a_400_38200# 1.39fF
C12284 VP.n5266 a_400_38200# 0.06fF
C12285 VP.n5267 a_400_38200# 0.37fF
C12286 VP.n5268 a_400_38200# 2.30fF
C12287 VP.t36 a_400_38200# 0.02fF
C12288 VP.n5269 a_400_38200# 0.24fF
C12289 VP.n5270 a_400_38200# 0.91fF
C12290 VP.n5271 a_400_38200# 0.05fF
C12291 VP.t330 a_400_38200# 0.02fF
C12292 VP.n5272 a_400_38200# 0.12fF
C12293 VP.n5273 a_400_38200# 0.14fF
C12294 VP.n5275 a_400_38200# 0.88fF
C12295 VP.n5276 a_400_38200# 0.48fF
C12296 VP.n5277 a_400_38200# 0.88fF
C12297 VP.n5278 a_400_38200# 0.60fF
C12298 VP.n5279 a_400_38200# 2.33fF
C12299 VP.n5280 a_400_38200# 0.59fF
C12300 VP.n5281 a_400_38200# 0.02fF
C12301 VP.n5282 a_400_38200# 0.96fF
C12302 VP.t22 a_400_38200# 15.72fF
C12303 VP.n5283 a_400_38200# 15.42fF
C12304 VP.n5285 a_400_38200# 0.38fF
C12305 VP.n5286 a_400_38200# 0.23fF
C12306 VP.n5287 a_400_38200# 3.42fF
C12307 VP.n5288 a_400_38200# 0.21fF
C12308 VP.n5289 a_400_38200# 1.08fF
C12309 VP.n5290 a_400_38200# 0.03fF
C12310 VP.n5291 a_400_38200# 0.09fF
C12311 VP.n5292 a_400_38200# 0.43fF
C12312 VP.n5293 a_400_38200# 0.37fF
C12313 VP.t748 a_400_38200# 0.02fF
C12314 VP.n5294 a_400_38200# 0.64fF
C12315 VP.n5295 a_400_38200# 0.60fF
C12316 VP.n5296 a_400_38200# 2.32fF
C12317 VP.n5297 a_400_38200# 4.93fF
C12318 VP.t320 a_400_38200# 0.02fF
C12319 VP.n5298 a_400_38200# 1.19fF
C12320 VP.n5299 a_400_38200# 0.05fF
C12321 VP.t568 a_400_38200# 0.02fF
C12322 VP.n5300 a_400_38200# 0.01fF
C12323 VP.n5301 a_400_38200# 0.26fF
C12324 VP.n5303 a_400_38200# 15.28fF
C12325 VP.n5304 a_400_38200# 0.10fF
C12326 VP.n5305 a_400_38200# 0.28fF
C12327 VP.n5306 a_400_38200# 0.15fF
C12328 VP.n5307 a_400_38200# 0.08fF
C12329 VP.n5308 a_400_38200# 0.14fF
C12330 VP.n5309 a_400_38200# 0.06fF
C12331 VP.n5310 a_400_38200# 0.06fF
C12332 VP.n5311 a_400_38200# 0.03fF
C12333 VP.n5312 a_400_38200# 0.05fF
C12334 VP.n5313 a_400_38200# 0.07fF
C12335 VP.n5314 a_400_38200# 0.19fF
C12336 VP.n5315 a_400_38200# 0.59fF
C12337 VP.n5316 a_400_38200# 0.34fF
C12338 VP.n5317 a_400_38200# 0.04fF
C12339 VP.n5318 a_400_38200# 0.02fF
C12340 VP.n5319 a_400_38200# 0.06fF
C12341 VP.n5320 a_400_38200# 0.30fF
C12342 VP.n5321 a_400_38200# 1.93fF
C12343 VP.n5322 a_400_38200# 0.12fF
C12344 VP.t1023 a_400_38200# 0.02fF
C12345 VP.n5323 a_400_38200# 0.14fF
C12346 VP.t313 a_400_38200# 0.02fF
C12347 VP.n5325 a_400_38200# 0.24fF
C12348 VP.n5326 a_400_38200# 0.35fF
C12349 VP.n5327 a_400_38200# 0.60fF
C12350 VP.n5328 a_400_38200# 2.47fF
C12351 VP.n5329 a_400_38200# 2.20fF
C12352 VP.t120 a_400_38200# 0.02fF
C12353 VP.n5330 a_400_38200# 0.12fF
C12354 VP.n5331 a_400_38200# 0.14fF
C12355 VP.t1185 a_400_38200# 0.02fF
C12356 VP.n5333 a_400_38200# 0.24fF
C12357 VP.n5334 a_400_38200# 0.91fF
C12358 VP.n5335 a_400_38200# 0.05fF
C12359 VP.n5336 a_400_38200# 0.10fF
C12360 VP.n5337 a_400_38200# 0.28fF
C12361 VP.n5338 a_400_38200# 0.15fF
C12362 VP.n5339 a_400_38200# 0.08fF
C12363 VP.n5340 a_400_38200# 0.14fF
C12364 VP.n5341 a_400_38200# 0.06fF
C12365 VP.n5342 a_400_38200# 0.06fF
C12366 VP.n5343 a_400_38200# 0.03fF
C12367 VP.n5344 a_400_38200# 0.05fF
C12368 VP.n5345 a_400_38200# 0.07fF
C12369 VP.n5346 a_400_38200# 0.19fF
C12370 VP.n5347 a_400_38200# 0.59fF
C12371 VP.n5348 a_400_38200# 0.34fF
C12372 VP.n5349 a_400_38200# 0.04fF
C12373 VP.n5350 a_400_38200# 0.02fF
C12374 VP.n5351 a_400_38200# 0.06fF
C12375 VP.n5352 a_400_38200# 0.30fF
C12376 VP.n5353 a_400_38200# 1.93fF
C12377 VP.n5354 a_400_38200# 0.12fF
C12378 VP.t575 a_400_38200# 0.02fF
C12379 VP.n5355 a_400_38200# 0.14fF
C12380 VP.t1157 a_400_38200# 0.02fF
C12381 VP.n5357 a_400_38200# 0.24fF
C12382 VP.n5358 a_400_38200# 0.35fF
C12383 VP.n5359 a_400_38200# 0.60fF
C12384 VP.n5360 a_400_38200# 2.47fF
C12385 VP.n5361 a_400_38200# 2.20fF
C12386 VP.t991 a_400_38200# 0.02fF
C12387 VP.n5362 a_400_38200# 0.12fF
C12388 VP.n5363 a_400_38200# 0.14fF
C12389 VP.t732 a_400_38200# 0.02fF
C12390 VP.n5365 a_400_38200# 0.24fF
C12391 VP.n5366 a_400_38200# 0.91fF
C12392 VP.n5367 a_400_38200# 0.05fF
C12393 VP.n5368 a_400_38200# 0.10fF
C12394 VP.n5369 a_400_38200# 0.28fF
C12395 VP.n5370 a_400_38200# 0.15fF
C12396 VP.n5371 a_400_38200# 0.08fF
C12397 VP.n5372 a_400_38200# 0.14fF
C12398 VP.n5373 a_400_38200# 0.06fF
C12399 VP.n5374 a_400_38200# 0.06fF
C12400 VP.n5375 a_400_38200# 0.03fF
C12401 VP.n5376 a_400_38200# 0.05fF
C12402 VP.n5377 a_400_38200# 0.07fF
C12403 VP.n5378 a_400_38200# 0.19fF
C12404 VP.n5379 a_400_38200# 0.59fF
C12405 VP.n5380 a_400_38200# 0.34fF
C12406 VP.n5381 a_400_38200# 0.04fF
C12407 VP.n5382 a_400_38200# 0.02fF
C12408 VP.n5383 a_400_38200# 0.06fF
C12409 VP.n5384 a_400_38200# 0.30fF
C12410 VP.n5385 a_400_38200# 1.93fF
C12411 VP.n5386 a_400_38200# 0.12fF
C12412 VP.t895 a_400_38200# 0.02fF
C12413 VP.n5387 a_400_38200# 0.14fF
C12414 VP.t88 a_400_38200# 0.02fF
C12415 VP.n5389 a_400_38200# 0.24fF
C12416 VP.n5390 a_400_38200# 0.35fF
C12417 VP.n5391 a_400_38200# 0.60fF
C12418 VP.n5392 a_400_38200# 2.47fF
C12419 VP.n5393 a_400_38200# 2.20fF
C12420 VP.t1244 a_400_38200# 0.02fF
C12421 VP.n5394 a_400_38200# 0.12fF
C12422 VP.n5395 a_400_38200# 0.14fF
C12423 VP.t981 a_400_38200# 0.02fF
C12424 VP.n5397 a_400_38200# 0.24fF
C12425 VP.n5398 a_400_38200# 0.91fF
C12426 VP.n5399 a_400_38200# 0.05fF
C12427 VP.n5400 a_400_38200# 0.10fF
C12428 VP.n5401 a_400_38200# 0.28fF
C12429 VP.n5402 a_400_38200# 0.15fF
C12430 VP.n5403 a_400_38200# 0.08fF
C12431 VP.n5404 a_400_38200# 0.14fF
C12432 VP.n5405 a_400_38200# 0.06fF
C12433 VP.n5406 a_400_38200# 0.06fF
C12434 VP.n5407 a_400_38200# 0.03fF
C12435 VP.n5408 a_400_38200# 0.05fF
C12436 VP.n5409 a_400_38200# 0.07fF
C12437 VP.n5410 a_400_38200# 0.19fF
C12438 VP.n5411 a_400_38200# 0.59fF
C12439 VP.n5412 a_400_38200# 0.34fF
C12440 VP.n5413 a_400_38200# 0.04fF
C12441 VP.n5414 a_400_38200# 0.02fF
C12442 VP.n5415 a_400_38200# 0.06fF
C12443 VP.n5416 a_400_38200# 0.30fF
C12444 VP.n5417 a_400_38200# 1.93fF
C12445 VP.n5418 a_400_38200# 0.12fF
C12446 VP.t443 a_400_38200# 0.02fF
C12447 VP.n5419 a_400_38200# 0.14fF
C12448 VP.t1028 a_400_38200# 0.02fF
C12449 VP.n5421 a_400_38200# 0.24fF
C12450 VP.n5422 a_400_38200# 0.35fF
C12451 VP.n5423 a_400_38200# 0.60fF
C12452 VP.n5424 a_400_38200# 2.39fF
C12453 VP.n5425 a_400_38200# 1.79fF
C12454 VP.t798 a_400_38200# 0.02fF
C12455 VP.n5426 a_400_38200# 0.12fF
C12456 VP.n5427 a_400_38200# 0.14fF
C12457 VP.t606 a_400_38200# 0.02fF
C12458 VP.n5429 a_400_38200# 0.24fF
C12459 VP.n5430 a_400_38200# 0.91fF
C12460 VP.n5431 a_400_38200# 0.05fF
C12461 VP.t119 a_400_38200# 34.79fF
C12462 VP.t586 a_400_38200# 0.02fF
C12463 VP.n5432 a_400_38200# 0.12fF
C12464 VP.n5433 a_400_38200# 0.14fF
C12465 VP.t339 a_400_38200# 0.02fF
C12466 VP.n5435 a_400_38200# 0.24fF
C12467 VP.n5436 a_400_38200# 0.91fF
C12468 VP.n5437 a_400_38200# 0.05fF
C12469 VP.t766 a_400_38200# 0.02fF
C12470 VP.n5438 a_400_38200# 0.24fF
C12471 VP.n5439 a_400_38200# 0.35fF
C12472 VP.n5440 a_400_38200# 0.60fF
C12473 VP.n5441 a_400_38200# 0.04fF
C12474 VP.n5442 a_400_38200# 0.08fF
C12475 VP.n5443 a_400_38200# 0.72fF
C12476 VP.n5444 a_400_38200# 0.09fF
C12477 VP.n5445 a_400_38200# 0.00fF
C12478 VP.n5446 a_400_38200# 0.98fF
C12479 VP.n5447 a_400_38200# 0.19fF
C12480 VP.n5449 a_400_38200# 1.72fF
C12481 VP.n5450 a_400_38200# 1.96fF
C12482 VP.n5451 a_400_38200# 1.04fF
C12483 VP.n5452 a_400_38200# 0.05fF
C12484 VP.n5453 a_400_38200# 0.03fF
C12485 VP.n5454 a_400_38200# 0.06fF
C12486 VP.n5455 a_400_38200# 0.06fF
C12487 VP.n5456 a_400_38200# 0.06fF
C12488 VP.n5457 a_400_38200# 0.07fF
C12489 VP.n5458 a_400_38200# 0.03fF
C12490 VP.n5459 a_400_38200# 0.05fF
C12491 VP.n5460 a_400_38200# 0.07fF
C12492 VP.n5461 a_400_38200# 0.19fF
C12493 VP.n5462 a_400_38200# 0.60fF
C12494 VP.n5463 a_400_38200# 0.76fF
C12495 VP.n5464 a_400_38200# 0.40fF
C12496 VP.n5465 a_400_38200# 0.03fF
C12497 VP.n5466 a_400_38200# 0.01fF
C12498 VP.t303 a_400_38200# 0.02fF
C12499 VP.n5467 a_400_38200# 0.25fF
C12500 VP.t1323 a_400_38200# 0.02fF
C12501 VP.n5468 a_400_38200# 0.95fF
C12502 VP.n5469 a_400_38200# 0.70fF
C12503 VP.n5470 a_400_38200# 1.93fF
C12504 VP.n5471 a_400_38200# 2.97fF
C12505 VP.n5472 a_400_38200# 2.27fF
C12506 VP.t504 a_400_38200# 0.02fF
C12507 VP.n5473 a_400_38200# 0.24fF
C12508 VP.n5474 a_400_38200# 0.35fF
C12509 VP.n5475 a_400_38200# 0.60fF
C12510 VP.n5476 a_400_38200# 0.12fF
C12511 VP.t27 a_400_38200# 0.02fF
C12512 VP.n5477 a_400_38200# 0.14fF
C12513 VP.n5479 a_400_38200# 0.04fF
C12514 VP.n5480 a_400_38200# 0.02fF
C12515 VP.n5481 a_400_38200# 0.06fF
C12516 VP.n5482 a_400_38200# 0.30fF
C12517 VP.n5483 a_400_38200# 0.10fF
C12518 VP.n5484 a_400_38200# 0.28fF
C12519 VP.n5485 a_400_38200# 0.06fF
C12520 VP.n5486 a_400_38200# 0.06fF
C12521 VP.n5487 a_400_38200# 0.03fF
C12522 VP.n5488 a_400_38200# 0.15fF
C12523 VP.n5489 a_400_38200# 0.08fF
C12524 VP.n5490 a_400_38200# 0.14fF
C12525 VP.n5491 a_400_38200# 0.03fF
C12526 VP.n5492 a_400_38200# 0.06fF
C12527 VP.n5493 a_400_38200# 0.06fF
C12528 VP.n5494 a_400_38200# 0.06fF
C12529 VP.n5495 a_400_38200# 0.06fF
C12530 VP.n5496 a_400_38200# 0.03fF
C12531 VP.n5497 a_400_38200# 0.05fF
C12532 VP.n5498 a_400_38200# 0.07fF
C12533 VP.n5499 a_400_38200# 0.19fF
C12534 VP.n5500 a_400_38200# 0.59fF
C12535 VP.n5501 a_400_38200# 0.34fF
C12536 VP.n5502 a_400_38200# 1.88fF
C12537 VP.t1080 a_400_38200# 0.02fF
C12538 VP.n5503 a_400_38200# 0.24fF
C12539 VP.n5504 a_400_38200# 0.91fF
C12540 VP.n5505 a_400_38200# 0.05fF
C12541 VP.t151 a_400_38200# 0.02fF
C12542 VP.n5506 a_400_38200# 0.12fF
C12543 VP.n5507 a_400_38200# 0.14fF
C12544 VP.n5509 a_400_38200# 0.19fF
C12545 VP.n5510 a_400_38200# 0.10fF
C12546 VP.n5511 a_400_38200# 0.10fF
C12547 VP.n5512 a_400_38200# 0.18fF
C12548 VP.n5513 a_400_38200# 0.09fF
C12549 VP.n5514 a_400_38200# 0.04fF
C12550 VP.n5515 a_400_38200# 0.19fF
C12551 VP.n5516 a_400_38200# 0.26fF
C12552 VP.n5517 a_400_38200# 1.17fF
C12553 VP.n5518 a_400_38200# 0.06fF
C12554 VP.n5519 a_400_38200# 0.44fF
C12555 VP.n5520 a_400_38200# 0.13fF
C12556 VP.n5521 a_400_38200# 0.02fF
C12557 VP.n5522 a_400_38200# 1.81fF
C12558 VP.n5523 a_400_38200# 0.12fF
C12559 VP.t923 a_400_38200# 0.02fF
C12560 VP.n5524 a_400_38200# 0.14fF
C12561 VP.t15 a_400_38200# 0.02fF
C12562 VP.n5526 a_400_38200# 0.24fF
C12563 VP.n5527 a_400_38200# 0.35fF
C12564 VP.n5528 a_400_38200# 0.60fF
C12565 VP.n5529 a_400_38200# 3.18fF
C12566 VP.n5530 a_400_38200# 2.06fF
C12567 VP.n5531 a_400_38200# 1.98fF
C12568 VP.t638 a_400_38200# 0.02fF
C12569 VP.n5532 a_400_38200# 0.24fF
C12570 VP.n5533 a_400_38200# 0.91fF
C12571 VP.n5534 a_400_38200# 0.05fF
C12572 VP.t1009 a_400_38200# 0.02fF
C12573 VP.n5535 a_400_38200# 0.12fF
C12574 VP.n5536 a_400_38200# 0.14fF
C12575 VP.n5538 a_400_38200# 0.16fF
C12576 VP.n5539 a_400_38200# 0.19fF
C12577 VP.n5540 a_400_38200# 0.09fF
C12578 VP.n5541 a_400_38200# 0.04fF
C12579 VP.n5542 a_400_38200# 0.14fF
C12580 VP.n5543 a_400_38200# 0.64fF
C12581 VP.n5544 a_400_38200# 1.32fF
C12582 VP.n5545 a_400_38200# 1.81fF
C12583 VP.n5546 a_400_38200# 0.12fF
C12584 VP.t473 a_400_38200# 0.02fF
C12585 VP.n5547 a_400_38200# 0.14fF
C12586 VP.t915 a_400_38200# 0.02fF
C12587 VP.n5549 a_400_38200# 0.24fF
C12588 VP.n5550 a_400_38200# 0.35fF
C12589 VP.n5551 a_400_38200# 0.60fF
C12590 VP.n5552 a_400_38200# 2.97fF
C12591 VP.n5553 a_400_38200# 2.27fF
C12592 VP.n5554 a_400_38200# 2.00fF
C12593 VP.t187 a_400_38200# 0.02fF
C12594 VP.n5555 a_400_38200# 0.24fF
C12595 VP.n5556 a_400_38200# 0.91fF
C12596 VP.n5557 a_400_38200# 0.05fF
C12597 VP.t565 a_400_38200# 0.02fF
C12598 VP.n5558 a_400_38200# 0.12fF
C12599 VP.n5559 a_400_38200# 0.14fF
C12600 VP.n5561 a_400_38200# 0.24fF
C12601 VP.t587 a_400_38200# 0.02fF
C12602 VP.n5562 a_400_38200# 0.36fF
C12603 VP.n5563 a_400_38200# 0.36fF
C12604 VP.n5564 a_400_38200# 0.67fF
C12605 VP.n5565 a_400_38200# 0.16fF
C12606 VP.n5566 a_400_38200# 0.19fF
C12607 VP.n5567 a_400_38200# 0.09fF
C12608 VP.n5568 a_400_38200# 0.04fF
C12609 VP.n5569 a_400_38200# 0.14fF
C12610 VP.n5570 a_400_38200# 0.64fF
C12611 VP.n5571 a_400_38200# 1.32fF
C12612 VP.n5572 a_400_38200# 1.81fF
C12613 VP.n5573 a_400_38200# 2.97fF
C12614 VP.n5574 a_400_38200# 2.27fF
C12615 VP.n5575 a_400_38200# 0.75fF
C12616 VP.n5576 a_400_38200# 0.24fF
C12617 VP.t1312 a_400_38200# 0.02fF
C12618 VP.n5577 a_400_38200# 0.35fF
C12619 VP.n5578 a_400_38200# 0.63fF
C12620 VP.n5579 a_400_38200# 0.40fF
C12621 VP.n5580 a_400_38200# 0.40fF
C12622 VP.n5581 a_400_38200# 0.12fF
C12623 VP.t939 a_400_38200# 0.02fF
C12624 VP.n5582 a_400_38200# 0.14fF
C12625 VP.t974 a_400_38200# 0.02fF
C12626 VP.n5584 a_400_38200# 0.12fF
C12627 VP.n5585 a_400_38200# 0.14fF
C12628 VP.n5587 a_400_38200# 0.03fF
C12629 VP.n5588 a_400_38200# 0.19fF
C12630 VP.n5589 a_400_38200# 0.24fF
C12631 VP.n5590 a_400_38200# 0.98fF
C12632 VP.n5591 a_400_38200# 0.12fF
C12633 VP.n5592 a_400_38200# 0.19fF
C12634 VP.n5593 a_400_38200# 0.09fF
C12635 VP.n5594 a_400_38200# 0.18fF
C12636 VP.n5595 a_400_38200# 0.09fF
C12637 VP.n5596 a_400_38200# 0.08fF
C12638 VP.n5597 a_400_38200# 0.39fF
C12639 VP.n5598 a_400_38200# 0.24fF
C12640 VP.n5599 a_400_38200# 0.13fF
C12641 VP.n5600 a_400_38200# 0.02fF
C12642 VP.n5601 a_400_38200# 1.81fF
C12643 VP.n5602 a_400_38200# 0.12fF
C12644 VP.t1345 a_400_38200# 0.02fF
C12645 VP.n5603 a_400_38200# 0.14fF
C12646 VP.t488 a_400_38200# 0.02fF
C12647 VP.n5605 a_400_38200# 0.24fF
C12648 VP.n5606 a_400_38200# 0.35fF
C12649 VP.n5607 a_400_38200# 0.60fF
C12650 VP.n5608 a_400_38200# 3.17fF
C12651 VP.n5609 a_400_38200# 2.27fF
C12652 VP.n5610 a_400_38200# 1.98fF
C12653 VP.t1064 a_400_38200# 0.02fF
C12654 VP.n5611 a_400_38200# 0.24fF
C12655 VP.n5612 a_400_38200# 0.91fF
C12656 VP.n5613 a_400_38200# 0.05fF
C12657 VP.t44 a_400_38200# 0.02fF
C12658 VP.n5614 a_400_38200# 0.12fF
C12659 VP.n5615 a_400_38200# 0.14fF
C12660 VP.n5617 a_400_38200# 15.28fF
C12661 VP.n5618 a_400_38200# 0.10fF
C12662 VP.n5619 a_400_38200# 0.28fF
C12663 VP.n5620 a_400_38200# 0.06fF
C12664 VP.n5621 a_400_38200# 0.06fF
C12665 VP.n5622 a_400_38200# 0.03fF
C12666 VP.n5623 a_400_38200# 0.15fF
C12667 VP.n5624 a_400_38200# 0.08fF
C12668 VP.n5625 a_400_38200# 0.14fF
C12669 VP.n5626 a_400_38200# 0.03fF
C12670 VP.n5627 a_400_38200# 0.06fF
C12671 VP.n5628 a_400_38200# 0.06fF
C12672 VP.n5629 a_400_38200# 0.06fF
C12673 VP.n5630 a_400_38200# 0.06fF
C12674 VP.n5631 a_400_38200# 0.03fF
C12675 VP.n5632 a_400_38200# 0.05fF
C12676 VP.n5633 a_400_38200# 0.07fF
C12677 VP.n5634 a_400_38200# 0.19fF
C12678 VP.n5635 a_400_38200# 0.59fF
C12679 VP.n5636 a_400_38200# 0.34fF
C12680 VP.n5637 a_400_38200# 0.04fF
C12681 VP.n5638 a_400_38200# 0.02fF
C12682 VP.n5639 a_400_38200# 0.06fF
C12683 VP.n5640 a_400_38200# 0.30fF
C12684 VP.n5641 a_400_38200# 1.93fF
C12685 VP.n5642 a_400_38200# 0.12fF
C12686 VP.t1149 a_400_38200# 0.02fF
C12687 VP.n5643 a_400_38200# 0.14fF
C12688 VP.t291 a_400_38200# 0.02fF
C12689 VP.n5645 a_400_38200# 0.24fF
C12690 VP.n5646 a_400_38200# 0.35fF
C12691 VP.n5647 a_400_38200# 0.60fF
C12692 VP.n5648 a_400_38200# 0.56fF
C12693 VP.n5649 a_400_38200# 1.24fF
C12694 VP.n5650 a_400_38200# 0.54fF
C12695 VP.n5651 a_400_38200# 0.22fF
C12696 VP.n5652 a_400_38200# 1.73fF
C12697 VP.t1198 a_400_38200# 0.02fF
C12698 VP.n5653 a_400_38200# 0.12fF
C12699 VP.n5654 a_400_38200# 0.14fF
C12700 VP.t872 a_400_38200# 0.02fF
C12701 VP.n5656 a_400_38200# 0.24fF
C12702 VP.n5657 a_400_38200# 0.91fF
C12703 VP.n5658 a_400_38200# 0.05fF
C12704 VP.n5659 a_400_38200# 0.10fF
C12705 VP.n5660 a_400_38200# 0.06fF
C12706 VP.n5661 a_400_38200# 0.06fF
C12707 VP.n5662 a_400_38200# 0.28fF
C12708 VP.n5663 a_400_38200# 0.03fF
C12709 VP.n5664 a_400_38200# 0.15fF
C12710 VP.n5665 a_400_38200# 0.08fF
C12711 VP.n5666 a_400_38200# 0.14fF
C12712 VP.n5667 a_400_38200# 0.03fF
C12713 VP.n5668 a_400_38200# 0.06fF
C12714 VP.n5669 a_400_38200# 0.06fF
C12715 VP.n5670 a_400_38200# 0.06fF
C12716 VP.n5671 a_400_38200# 0.06fF
C12717 VP.n5672 a_400_38200# 0.03fF
C12718 VP.n5673 a_400_38200# 0.05fF
C12719 VP.n5674 a_400_38200# 0.07fF
C12720 VP.n5675 a_400_38200# 0.19fF
C12721 VP.n5676 a_400_38200# 0.59fF
C12722 VP.n5677 a_400_38200# 0.34fF
C12723 VP.n5678 a_400_38200# 0.04fF
C12724 VP.n5679 a_400_38200# 0.02fF
C12725 VP.n5680 a_400_38200# 0.06fF
C12726 VP.n5681 a_400_38200# 0.30fF
C12727 VP.n5682 a_400_38200# 1.93fF
C12728 VP.n5683 a_400_38200# 0.12fF
C12729 VP.t702 a_400_38200# 0.02fF
C12730 VP.n5684 a_400_38200# 0.14fF
C12731 VP.t1142 a_400_38200# 0.02fF
C12732 VP.n5686 a_400_38200# 0.24fF
C12733 VP.n5687 a_400_38200# 0.35fF
C12734 VP.n5688 a_400_38200# 0.60fF
C12735 VP.n5689 a_400_38200# 0.72fF
C12736 VP.n5690 a_400_38200# 1.24fF
C12737 VP.n5691 a_400_38200# 0.54fF
C12738 VP.n5692 a_400_38200# 0.22fF
C12739 VP.n5693 a_400_38200# 1.73fF
C12740 VP.t747 a_400_38200# 0.02fF
C12741 VP.n5694 a_400_38200# 0.12fF
C12742 VP.n5695 a_400_38200# 0.14fF
C12743 VP.t426 a_400_38200# 0.02fF
C12744 VP.n5697 a_400_38200# 0.24fF
C12745 VP.n5698 a_400_38200# 0.91fF
C12746 VP.n5699 a_400_38200# 0.05fF
C12747 VP.n5700 a_400_38200# 0.10fF
C12748 VP.n5701 a_400_38200# 0.28fF
C12749 VP.n5702 a_400_38200# 0.06fF
C12750 VP.n5703 a_400_38200# 0.06fF
C12751 VP.n5704 a_400_38200# 0.03fF
C12752 VP.n5705 a_400_38200# 0.15fF
C12753 VP.n5706 a_400_38200# 0.08fF
C12754 VP.n5707 a_400_38200# 0.14fF
C12755 VP.n5708 a_400_38200# 0.03fF
C12756 VP.n5709 a_400_38200# 0.06fF
C12757 VP.n5710 a_400_38200# 0.06fF
C12758 VP.n5711 a_400_38200# 0.06fF
C12759 VP.n5712 a_400_38200# 0.06fF
C12760 VP.n5713 a_400_38200# 0.03fF
C12761 VP.n5714 a_400_38200# 0.05fF
C12762 VP.n5715 a_400_38200# 0.07fF
C12763 VP.n5716 a_400_38200# 0.19fF
C12764 VP.n5717 a_400_38200# 0.59fF
C12765 VP.n5718 a_400_38200# 0.34fF
C12766 VP.n5719 a_400_38200# 0.04fF
C12767 VP.n5720 a_400_38200# 0.02fF
C12768 VP.n5721 a_400_38200# 0.06fF
C12769 VP.n5722 a_400_38200# 0.30fF
C12770 VP.n5723 a_400_38200# 1.93fF
C12771 VP.n5724 a_400_38200# 0.12fF
C12772 VP.t958 a_400_38200# 0.02fF
C12773 VP.n5725 a_400_38200# 0.14fF
C12774 VP.t66 a_400_38200# 0.02fF
C12775 VP.n5727 a_400_38200# 0.24fF
C12776 VP.n5728 a_400_38200# 0.35fF
C12777 VP.n5729 a_400_38200# 0.60fF
C12778 VP.n5730 a_400_38200# 0.72fF
C12779 VP.n5731 a_400_38200# 1.24fF
C12780 VP.n5732 a_400_38200# 0.54fF
C12781 VP.n5733 a_400_38200# 0.22fF
C12782 VP.n5734 a_400_38200# 1.73fF
C12783 VP.t293 a_400_38200# 0.02fF
C12784 VP.n5735 a_400_38200# 0.12fF
C12785 VP.n5736 a_400_38200# 0.14fF
C12786 VP.t672 a_400_38200# 0.02fF
C12787 VP.n5738 a_400_38200# 0.24fF
C12788 VP.n5739 a_400_38200# 0.91fF
C12789 VP.n5740 a_400_38200# 0.05fF
C12790 VP.n5741 a_400_38200# 0.10fF
C12791 VP.n5742 a_400_38200# 0.06fF
C12792 VP.n5743 a_400_38200# 0.06fF
C12793 VP.n5744 a_400_38200# 0.28fF
C12794 VP.n5745 a_400_38200# 0.03fF
C12795 VP.n5746 a_400_38200# 0.15fF
C12796 VP.n5747 a_400_38200# 0.08fF
C12797 VP.n5748 a_400_38200# 0.14fF
C12798 VP.n5749 a_400_38200# 0.03fF
C12799 VP.n5750 a_400_38200# 0.06fF
C12800 VP.n5751 a_400_38200# 0.06fF
C12801 VP.n5752 a_400_38200# 0.06fF
C12802 VP.n5753 a_400_38200# 0.06fF
C12803 VP.n5754 a_400_38200# 0.03fF
C12804 VP.n5755 a_400_38200# 0.05fF
C12805 VP.n5756 a_400_38200# 0.07fF
C12806 VP.n5757 a_400_38200# 0.19fF
C12807 VP.n5758 a_400_38200# 0.59fF
C12808 VP.n5759 a_400_38200# 0.34fF
C12809 VP.n5760 a_400_38200# 0.04fF
C12810 VP.n5761 a_400_38200# 0.02fF
C12811 VP.n5762 a_400_38200# 0.06fF
C12812 VP.n5763 a_400_38200# 0.30fF
C12813 VP.n5764 a_400_38200# 1.93fF
C12814 VP.n5765 a_400_38200# 0.12fF
C12815 VP.t510 a_400_38200# 0.02fF
C12816 VP.n5766 a_400_38200# 0.14fF
C12817 VP.t950 a_400_38200# 0.02fF
C12818 VP.n5768 a_400_38200# 0.24fF
C12819 VP.n5769 a_400_38200# 0.35fF
C12820 VP.n5770 a_400_38200# 0.60fF
C12821 VP.n5771 a_400_38200# 0.71fF
C12822 VP.n5772 a_400_38200# 1.39fF
C12823 VP.n5773 a_400_38200# 0.54fF
C12824 VP.n5774 a_400_38200# 0.21fF
C12825 VP.n5775 a_400_38200# 1.73fF
C12826 VP.t615 a_400_38200# 0.02fF
C12827 VP.n5776 a_400_38200# 0.12fF
C12828 VP.n5777 a_400_38200# 0.14fF
C12829 VP.t225 a_400_38200# 0.02fF
C12830 VP.n5779 a_400_38200# 0.24fF
C12831 VP.n5780 a_400_38200# 0.91fF
C12832 VP.n5781 a_400_38200# 0.05fF
C12833 VP.n5782 a_400_38200# 0.06fF
C12834 VP.n5783 a_400_38200# 0.06fF
C12835 VP.n5784 a_400_38200# 0.03fF
C12836 VP.n5785 a_400_38200# 0.10fF
C12837 VP.n5786 a_400_38200# 0.17fF
C12838 VP.n5787 a_400_38200# 0.10fF
C12839 VP.n5788 a_400_38200# 0.13fF
C12840 VP.n5789 a_400_38200# 0.02fF
C12841 VP.n5790 a_400_38200# 0.04fF
C12842 VP.n5791 a_400_38200# 0.06fF
C12843 VP.n5792 a_400_38200# 0.09fF
C12844 VP.n5793 a_400_38200# 0.10fF
C12845 VP.n5794 a_400_38200# 0.05fF
C12846 VP.n5795 a_400_38200# 0.19fF
C12847 VP.n5796 a_400_38200# 0.16fF
C12848 VP.n5797 a_400_38200# 0.04fF
C12849 VP.n5798 a_400_38200# 0.05fF
C12850 VP.n5799 a_400_38200# 0.04fF
C12851 VP.n5800 a_400_38200# 0.12fF
C12852 VP.n5801 a_400_38200# 0.09fF
C12853 VP.n5802 a_400_38200# 0.14fF
C12854 VP.n5803 a_400_38200# 0.56fF
C12855 VP.n5804 a_400_38200# 0.10fF
C12856 VP.n5805 a_400_38200# 1.93fF
C12857 VP.n5806 a_400_38200# 0.12fF
C12858 VP.t1321 a_400_38200# 0.02fF
C12859 VP.n5807 a_400_38200# 0.14fF
C12860 VP.t464 a_400_38200# 0.02fF
C12861 VP.n5809 a_400_38200# 0.24fF
C12862 VP.n5810 a_400_38200# 0.35fF
C12863 VP.n5811 a_400_38200# 0.60fF
C12864 VP.n5812 a_400_38200# 2.23fF
C12865 VP.n5813 a_400_38200# 0.18fF
C12866 VP.n5814 a_400_38200# 0.45fF
C12867 VP.n5815 a_400_38200# 0.06fF
C12868 VP.n5816 a_400_38200# 0.01fF
C12869 VP.n5817 a_400_38200# 0.01fF
C12870 VP.n5818 a_400_38200# 0.04fF
C12871 VP.n5819 a_400_38200# 0.02fF
C12872 VP.n5820 a_400_38200# 0.07fF
C12873 VP.n5821 a_400_38200# 0.04fF
C12874 VP.n5822 a_400_38200# 0.14fF
C12875 VP.n5823 a_400_38200# 0.45fF
C12876 VP.n5824 a_400_38200# 1.46fF
C12877 VP.n5825 a_400_38200# 1.78fF
C12878 VP.t97 a_400_38200# 0.02fF
C12879 VP.n5826 a_400_38200# 0.12fF
C12880 VP.n5827 a_400_38200# 0.14fF
C12881 VP.t1036 a_400_38200# 0.02fF
C12882 VP.n5829 a_400_38200# 0.24fF
C12883 VP.n5830 a_400_38200# 0.91fF
C12884 VP.n5831 a_400_38200# 0.05fF
C12885 VP.n5832 a_400_38200# 1.93fF
C12886 VP.n5833 a_400_38200# 2.23fF
C12887 VP.n5834 a_400_38200# 0.18fF
C12888 VP.n5835 a_400_38200# 0.45fF
C12889 VP.n5836 a_400_38200# 0.06fF
C12890 VP.n5837 a_400_38200# 0.01fF
C12891 VP.n5838 a_400_38200# 0.01fF
C12892 VP.n5839 a_400_38200# 0.04fF
C12893 VP.n5840 a_400_38200# 0.02fF
C12894 VP.n5841 a_400_38200# 0.07fF
C12895 VP.n5842 a_400_38200# 0.04fF
C12896 VP.n5843 a_400_38200# 0.14fF
C12897 VP.n5844 a_400_38200# 0.45fF
C12898 VP.n5845 a_400_38200# 1.46fF
C12899 VP.t934 a_400_38200# 0.02fF
C12900 VP.n5846 a_400_38200# 0.24fF
C12901 VP.n5847 a_400_38200# 0.35fF
C12902 VP.n5848 a_400_38200# 0.60fF
C12903 VP.n5849 a_400_38200# 0.12fF
C12904 VP.t494 a_400_38200# 0.02fF
C12905 VP.n5850 a_400_38200# 0.14fF
C12906 VP.n5852 a_400_38200# 0.10fF
C12907 VP.n5853 a_400_38200# 0.17fF
C12908 VP.n5854 a_400_38200# 0.06fF
C12909 VP.n5855 a_400_38200# 0.06fF
C12910 VP.n5856 a_400_38200# 0.03fF
C12911 VP.n5857 a_400_38200# 0.10fF
C12912 VP.n5858 a_400_38200# 0.13fF
C12913 VP.n5859 a_400_38200# 0.13fF
C12914 VP.n5860 a_400_38200# 0.04fF
C12915 VP.n5861 a_400_38200# 0.05fF
C12916 VP.n5862 a_400_38200# 0.04fF
C12917 VP.n5863 a_400_38200# 0.09fF
C12918 VP.n5864 a_400_38200# 0.09fF
C12919 VP.n5865 a_400_38200# 0.05fF
C12920 VP.n5866 a_400_38200# 0.19fF
C12921 VP.n5867 a_400_38200# 0.12fF
C12922 VP.n5868 a_400_38200# 0.09fF
C12923 VP.n5869 a_400_38200# 0.14fF
C12924 VP.n5870 a_400_38200# 0.04fF
C12925 VP.n5871 a_400_38200# 0.02fF
C12926 VP.n5872 a_400_38200# 0.06fF
C12927 VP.n5873 a_400_38200# 0.56fF
C12928 VP.n5874 a_400_38200# 0.10fF
C12929 VP.n5875 a_400_38200# 1.78fF
C12930 VP.t525 a_400_38200# 0.02fF
C12931 VP.n5876 a_400_38200# 0.12fF
C12932 VP.n5877 a_400_38200# 0.14fF
C12933 VP.t209 a_400_38200# 0.02fF
C12934 VP.n5879 a_400_38200# 0.24fF
C12935 VP.n5880 a_400_38200# 0.91fF
C12936 VP.n5881 a_400_38200# 0.05fF
C12937 VP.n5882 a_400_38200# 1.92fF
C12938 VP.n5883 a_400_38200# 2.51fF
C12939 VP.t722 a_400_38200# 0.02fF
C12940 VP.n5884 a_400_38200# 0.24fF
C12941 VP.n5885 a_400_38200# 0.35fF
C12942 VP.n5886 a_400_38200# 0.60fF
C12943 VP.n5887 a_400_38200# 0.12fF
C12944 VP.t280 a_400_38200# 0.02fF
C12945 VP.n5888 a_400_38200# 0.14fF
C12946 VP.n5890 a_400_38200# 0.06fF
C12947 VP.n5891 a_400_38200# 0.30fF
C12948 VP.n5892 a_400_38200# 0.20fF
C12949 VP.n5893 a_400_38200# 0.09fF
C12950 VP.n5894 a_400_38200# 0.26fF
C12951 VP.n5895 a_400_38200# 0.22fF
C12952 VP.n5896 a_400_38200# 0.19fF
C12953 VP.n5897 a_400_38200# 0.05fF
C12954 VP.n5898 a_400_38200# 0.13fF
C12955 VP.n5899 a_400_38200# 0.09fF
C12956 VP.n5900 a_400_38200# 0.09fF
C12957 VP.n5901 a_400_38200# 0.07fF
C12958 VP.n5902 a_400_38200# 0.71fF
C12959 VP.n5903 a_400_38200# 0.24fF
C12960 VP.n5904 a_400_38200# 1.88fF
C12961 VP.t933 a_400_38200# 0.02fF
C12962 VP.n5905 a_400_38200# 0.12fF
C12963 VP.n5906 a_400_38200# 0.14fF
C12964 VP.t1305 a_400_38200# 0.02fF
C12965 VP.n5908 a_400_38200# 0.24fF
C12966 VP.n5909 a_400_38200# 0.91fF
C12967 VP.n5910 a_400_38200# 0.05fF
C12968 VP.t26 a_400_38200# 35.17fF
C12969 VP.t744 a_400_38200# 0.02fF
C12970 VP.n5911 a_400_38200# 1.21fF
C12971 VP.n5912 a_400_38200# 0.25fF
C12972 VP.n5913 a_400_38200# 26.29fF
C12973 VP.n5914 a_400_38200# 26.29fF
C12974 VP.n5915 a_400_38200# 0.76fF
C12975 VP.n5916 a_400_38200# 0.27fF
C12976 VP.n5917 a_400_38200# 0.59fF
C12977 VP.n5918 a_400_38200# 0.10fF
C12978 VP.n5919 a_400_38200# 3.02fF
C12979 VP.t14 a_400_38200# 15.72fF
C12980 VP.n5920 a_400_38200# 1.15fF
C12981 VP.n5922 a_400_38200# 13.70fF
C12982 VP.n5924 a_400_38200# 1.99fF
C12983 VP.n5925 a_400_38200# 4.39fF
C12984 VP.n5926 a_400_38200# 0.03fF
C12985 VP.n5927 a_400_38200# 0.05fF
C12986 VP.n5928 a_400_38200# 0.07fF
C12987 VP.n5929 a_400_38200# 0.03fF
C12988 VP.n5930 a_400_38200# 0.06fF
C12989 VP.n5931 a_400_38200# 0.06fF
C12990 VP.n5932 a_400_38200# 0.06fF
C12991 VP.n5933 a_400_38200# 0.07fF
C12992 VP.n5934 a_400_38200# 0.57fF
C12993 VP.n5935 a_400_38200# 1.88fF
C12994 VP.n5936 a_400_38200# 0.92fF
C12995 VP.n5937 a_400_38200# 2.63fF
C12996 VP.n5938 a_400_38200# 0.10fF
C12997 VP.n5939 a_400_38200# 0.28fF
C12998 VP.n5940 a_400_38200# 0.15fF
C12999 VP.n5941 a_400_38200# 0.08fF
C13000 VP.n5942 a_400_38200# 0.14fF
C13001 VP.n5943 a_400_38200# 0.06fF
C13002 VP.n5944 a_400_38200# 0.06fF
C13003 VP.n5945 a_400_38200# 0.03fF
C13004 VP.n5946 a_400_38200# 0.05fF
C13005 VP.n5947 a_400_38200# 0.07fF
C13006 VP.n5948 a_400_38200# 0.19fF
C13007 VP.n5949 a_400_38200# 0.59fF
C13008 VP.n5950 a_400_38200# 0.34fF
C13009 VP.n5951 a_400_38200# 0.04fF
C13010 VP.n5952 a_400_38200# 0.02fF
C13011 VP.n5953 a_400_38200# 0.06fF
C13012 VP.n5954 a_400_38200# 0.30fF
C13013 VP.n5955 a_400_38200# 0.12fF
C13014 VP.t327 a_400_38200# 0.02fF
C13015 VP.n5956 a_400_38200# 0.14fF
C13016 VP.n5958 a_400_38200# 1.93fF
C13017 VP.t1177 a_400_38200# 0.02fF
C13018 VP.n5959 a_400_38200# 0.24fF
C13019 VP.n5960 a_400_38200# 0.35fF
C13020 VP.n5961 a_400_38200# 0.60fF
C13021 VP.n5962 a_400_38200# 0.12fF
C13022 VP.t592 a_400_38200# 0.02fF
C13023 VP.n5963 a_400_38200# 0.14fF
C13024 VP.n5965 a_400_38200# 0.04fF
C13025 VP.n5966 a_400_38200# 0.02fF
C13026 VP.n5967 a_400_38200# 0.06fF
C13027 VP.n5968 a_400_38200# 0.30fF
C13028 VP.n5969 a_400_38200# 0.10fF
C13029 VP.n5970 a_400_38200# 0.28fF
C13030 VP.n5971 a_400_38200# 0.15fF
C13031 VP.n5972 a_400_38200# 0.08fF
C13032 VP.n5973 a_400_38200# 0.14fF
C13033 VP.n5974 a_400_38200# 0.06fF
C13034 VP.n5975 a_400_38200# 0.06fF
C13035 VP.n5976 a_400_38200# 0.03fF
C13036 VP.n5977 a_400_38200# 0.05fF
C13037 VP.n5978 a_400_38200# 0.07fF
C13038 VP.n5979 a_400_38200# 0.19fF
C13039 VP.n5980 a_400_38200# 0.59fF
C13040 VP.n5981 a_400_38200# 0.34fF
C13041 VP.n5982 a_400_38200# 2.18fF
C13042 VP.t901 a_400_38200# 0.02fF
C13043 VP.n5983 a_400_38200# 0.24fF
C13044 VP.n5984 a_400_38200# 0.91fF
C13045 VP.n5985 a_400_38200# 0.05fF
C13046 VP.t942 a_400_38200# 0.02fF
C13047 VP.n5986 a_400_38200# 0.12fF
C13048 VP.n5987 a_400_38200# 0.14fF
C13049 VP.n5989 a_400_38200# 0.10fF
C13050 VP.n5990 a_400_38200# 0.10fF
C13051 VP.n5991 a_400_38200# 0.18fF
C13052 VP.n5992 a_400_38200# 0.09fF
C13053 VP.n5993 a_400_38200# 0.04fF
C13054 VP.n5994 a_400_38200# 0.26fF
C13055 VP.n5995 a_400_38200# 1.17fF
C13056 VP.n5996 a_400_38200# 0.06fF
C13057 VP.n5997 a_400_38200# 0.44fF
C13058 VP.n5998 a_400_38200# 0.13fF
C13059 VP.n5999 a_400_38200# 0.02fF
C13060 VP.n6000 a_400_38200# 1.81fF
C13061 VP.n6001 a_400_38200# 0.12fF
C13062 VP.t125 a_400_38200# 0.02fF
C13063 VP.n6002 a_400_38200# 0.14fF
C13064 VP.t725 a_400_38200# 0.02fF
C13065 VP.n6004 a_400_38200# 0.24fF
C13066 VP.n6005 a_400_38200# 0.35fF
C13067 VP.n6006 a_400_38200# 0.60fF
C13068 VP.n6007 a_400_38200# 2.28fF
C13069 VP.t448 a_400_38200# 0.02fF
C13070 VP.n6008 a_400_38200# 0.24fF
C13071 VP.n6009 a_400_38200# 0.91fF
C13072 VP.n6010 a_400_38200# 0.05fF
C13073 VP.t497 a_400_38200# 0.02fF
C13074 VP.n6011 a_400_38200# 0.12fF
C13075 VP.n6012 a_400_38200# 0.14fF
C13076 VP.n6014 a_400_38200# 0.06fF
C13077 VP.n6015 a_400_38200# 0.09fF
C13078 VP.n6016 a_400_38200# 0.09fF
C13079 VP.n6017 a_400_38200# 1.45fF
C13080 VP.n6018 a_400_38200# 0.14fF
C13081 VP.n6019 a_400_38200# 0.07fF
C13082 VP.n6020 a_400_38200# 0.72fF
C13083 VP.n6021 a_400_38200# 1.81fF
C13084 VP.n6022 a_400_38200# 0.12fF
C13085 VP.t995 a_400_38200# 0.02fF
C13086 VP.n6023 a_400_38200# 0.14fF
C13087 VP.t276 a_400_38200# 0.02fF
C13088 VP.n6025 a_400_38200# 0.24fF
C13089 VP.n6026 a_400_38200# 0.35fF
C13090 VP.n6027 a_400_38200# 0.60fF
C13091 VP.n6028 a_400_38200# 2.30fF
C13092 VP.t1301 a_400_38200# 0.02fF
C13093 VP.n6029 a_400_38200# 0.24fF
C13094 VP.n6030 a_400_38200# 0.91fF
C13095 VP.n6031 a_400_38200# 0.05fF
C13096 VP.t1348 a_400_38200# 0.02fF
C13097 VP.n6032 a_400_38200# 0.12fF
C13098 VP.n6033 a_400_38200# 0.14fF
C13099 VP.n6035 a_400_38200# 0.06fF
C13100 VP.n6036 a_400_38200# 0.25fF
C13101 VP.n6037 a_400_38200# 0.45fF
C13102 VP.n6038 a_400_38200# 0.03fF
C13103 VP.n6039 a_400_38200# 0.05fF
C13104 VP.n6040 a_400_38200# 0.07fF
C13105 VP.n6041 a_400_38200# 0.06fF
C13106 VP.n6042 a_400_38200# 0.06fF
C13107 VP.n6043 a_400_38200# 0.19fF
C13108 VP.n6044 a_400_38200# 0.59fF
C13109 VP.n6045 a_400_38200# 0.34fF
C13110 VP.n6046 a_400_38200# 0.05fF
C13111 VP.n6047 a_400_38200# 0.30fF
C13112 VP.n6048 a_400_38200# 1.93fF
C13113 VP.n6049 a_400_38200# 0.12fF
C13114 VP.t549 a_400_38200# 0.02fF
C13115 VP.n6050 a_400_38200# 0.14fF
C13116 VP.t1131 a_400_38200# 0.02fF
C13117 VP.n6052 a_400_38200# 0.24fF
C13118 VP.n6053 a_400_38200# 0.35fF
C13119 VP.n6054 a_400_38200# 0.60fF
C13120 VP.n6055 a_400_38200# 2.23fF
C13121 VP.n6056 a_400_38200# 2.04fF
C13122 VP.t855 a_400_38200# 0.02fF
C13123 VP.n6057 a_400_38200# 0.24fF
C13124 VP.n6058 a_400_38200# 0.91fF
C13125 VP.n6059 a_400_38200# 0.05fF
C13126 VP.t902 a_400_38200# 0.02fF
C13127 VP.n6060 a_400_38200# 0.12fF
C13128 VP.n6061 a_400_38200# 0.14fF
C13129 VP.n6063 a_400_38200# 0.24fF
C13130 VP.t406 a_400_38200# 0.02fF
C13131 VP.n6064 a_400_38200# 0.36fF
C13132 VP.n6065 a_400_38200# 0.36fF
C13133 VP.n6066 a_400_38200# 0.67fF
C13134 VP.n6067 a_400_38200# 0.06fF
C13135 VP.n6068 a_400_38200# 0.09fF
C13136 VP.n6069 a_400_38200# 0.09fF
C13137 VP.n6070 a_400_38200# 1.45fF
C13138 VP.n6071 a_400_38200# 0.14fF
C13139 VP.n6072 a_400_38200# 0.07fF
C13140 VP.n6073 a_400_38200# 0.72fF
C13141 VP.n6074 a_400_38200# 1.81fF
C13142 VP.n6075 a_400_38200# 1.06fF
C13143 VP.n6076 a_400_38200# 0.24fF
C13144 VP.t683 a_400_38200# 0.02fF
C13145 VP.n6077 a_400_38200# 0.35fF
C13146 VP.n6078 a_400_38200# 0.63fF
C13147 VP.n6079 a_400_38200# 0.40fF
C13148 VP.n6080 a_400_38200# 0.40fF
C13149 VP.n6081 a_400_38200# 0.12fF
C13150 VP.t75 a_400_38200# 0.02fF
C13151 VP.n6082 a_400_38200# 0.14fF
C13152 VP.t450 a_400_38200# 0.02fF
C13153 VP.n6084 a_400_38200# 0.12fF
C13154 VP.n6085 a_400_38200# 0.14fF
C13155 VP.n6087 a_400_38200# 1.93fF
C13156 VP.n6088 a_400_38200# 2.23fF
C13157 VP.t239 a_400_38200# 0.02fF
C13158 VP.n6089 a_400_38200# 0.24fF
C13159 VP.n6090 a_400_38200# 0.35fF
C13160 VP.n6091 a_400_38200# 0.60fF
C13161 VP.n6092 a_400_38200# 0.12fF
C13162 VP.t957 a_400_38200# 0.02fF
C13163 VP.n6093 a_400_38200# 0.14fF
C13164 VP.n6095 a_400_38200# 0.07fF
C13165 VP.n6096 a_400_38200# 0.30fF
C13166 VP.n6097 a_400_38200# 0.06fF
C13167 VP.n6098 a_400_38200# 0.25fF
C13168 VP.n6099 a_400_38200# 0.45fF
C13169 VP.n6100 a_400_38200# 0.06fF
C13170 VP.n6101 a_400_38200# 0.06fF
C13171 VP.n6102 a_400_38200# 0.03fF
C13172 VP.n6103 a_400_38200# 0.05fF
C13173 VP.n6104 a_400_38200# 0.07fF
C13174 VP.n6105 a_400_38200# 0.19fF
C13175 VP.n6106 a_400_38200# 0.59fF
C13176 VP.n6107 a_400_38200# 0.34fF
C13177 VP.n6108 a_400_38200# 2.04fF
C13178 VP.t1262 a_400_38200# 0.02fF
C13179 VP.n6109 a_400_38200# 0.24fF
C13180 VP.n6110 a_400_38200# 0.91fF
C13181 VP.n6111 a_400_38200# 0.05fF
C13182 VP.t33 a_400_38200# 0.02fF
C13183 VP.n6112 a_400_38200# 0.12fF
C13184 VP.n6113 a_400_38200# 0.14fF
C13185 VP.n6115 a_400_38200# 0.06fF
C13186 VP.n6116 a_400_38200# 0.09fF
C13187 VP.n6117 a_400_38200# 0.09fF
C13188 VP.n6118 a_400_38200# 0.43fF
C13189 VP.n6119 a_400_38200# 0.69fF
C13190 VP.n6120 a_400_38200# 0.14fF
C13191 VP.n6121 a_400_38200# 0.07fF
C13192 VP.n6122 a_400_38200# 0.72fF
C13193 VP.n6123 a_400_38200# 1.81fF
C13194 VP.n6124 a_400_38200# 0.12fF
C13195 VP.t509 a_400_38200# 0.02fF
C13196 VP.n6125 a_400_38200# 0.14fF
C13197 VP.t1094 a_400_38200# 0.02fF
C13198 VP.n6127 a_400_38200# 0.24fF
C13199 VP.n6128 a_400_38200# 0.35fF
C13200 VP.n6129 a_400_38200# 0.60fF
C13201 VP.n6130 a_400_38200# 2.30fF
C13202 VP.t817 a_400_38200# 0.02fF
C13203 VP.n6131 a_400_38200# 0.24fF
C13204 VP.n6132 a_400_38200# 0.91fF
C13205 VP.n6133 a_400_38200# 0.05fF
C13206 VP.t925 a_400_38200# 0.02fF
C13207 VP.n6134 a_400_38200# 0.12fF
C13208 VP.n6135 a_400_38200# 0.14fF
C13209 VP.n6137 a_400_38200# 0.31fF
C13210 VP.n6138 a_400_38200# 0.04fF
C13211 VP.n6139 a_400_38200# 0.88fF
C13212 VP.n6140 a_400_38200# 0.48fF
C13213 VP.n6141 a_400_38200# 0.88fF
C13214 VP.n6142 a_400_38200# 0.60fF
C13215 VP.n6143 a_400_38200# 2.33fF
C13216 VP.n6144 a_400_38200# 0.59fF
C13217 VP.n6145 a_400_38200# 0.02fF
C13218 VP.n6146 a_400_38200# 0.96fF
C13219 VP.t186 a_400_38200# 15.72fF
C13220 VP.n6147 a_400_38200# 15.42fF
C13221 VP.n6149 a_400_38200# 0.38fF
C13222 VP.n6150 a_400_38200# 0.23fF
C13223 VP.n6151 a_400_38200# 3.28fF
C13224 VP.n6152 a_400_38200# 1.41fF
C13225 VP.n6153 a_400_38200# 0.30fF
C13226 VP.t897 a_400_38200# 0.02fF
C13227 VP.n6154 a_400_38200# 0.64fF
C13228 VP.n6155 a_400_38200# 0.60fF
C13229 VP.n6156 a_400_38200# 1.88fF
C13230 VP.n6157 a_400_38200# 4.64fF
C13231 VP.t618 a_400_38200# 0.02fF
C13232 VP.n6158 a_400_38200# 1.19fF
C13233 VP.n6159 a_400_38200# 0.05fF
C13234 VP.t709 a_400_38200# 0.02fF
C13235 VP.n6160 a_400_38200# 0.01fF
C13236 VP.n6161 a_400_38200# 0.26fF
C13237 VP.n6163 a_400_38200# 15.28fF
C13238 VP.n6164 a_400_38200# 0.10fF
C13239 VP.n6165 a_400_38200# 0.28fF
C13240 VP.n6166 a_400_38200# 0.15fF
C13241 VP.n6167 a_400_38200# 0.08fF
C13242 VP.n6168 a_400_38200# 0.14fF
C13243 VP.n6169 a_400_38200# 0.06fF
C13244 VP.n6170 a_400_38200# 0.06fF
C13245 VP.n6171 a_400_38200# 0.03fF
C13246 VP.n6172 a_400_38200# 0.05fF
C13247 VP.n6173 a_400_38200# 0.07fF
C13248 VP.n6174 a_400_38200# 0.19fF
C13249 VP.n6175 a_400_38200# 0.59fF
C13250 VP.n6176 a_400_38200# 0.34fF
C13251 VP.n6177 a_400_38200# 0.04fF
C13252 VP.n6178 a_400_38200# 0.02fF
C13253 VP.n6179 a_400_38200# 0.06fF
C13254 VP.n6180 a_400_38200# 0.30fF
C13255 VP.n6181 a_400_38200# 1.93fF
C13256 VP.n6182 a_400_38200# 0.12fF
C13257 VP.t1171 a_400_38200# 0.02fF
C13258 VP.n6183 a_400_38200# 0.14fF
C13259 VP.t466 a_400_38200# 0.02fF
C13260 VP.n6185 a_400_38200# 0.24fF
C13261 VP.n6186 a_400_38200# 0.35fF
C13262 VP.n6187 a_400_38200# 0.60fF
C13263 VP.n6188 a_400_38200# 2.47fF
C13264 VP.n6189 a_400_38200# 2.20fF
C13265 VP.t279 a_400_38200# 0.02fF
C13266 VP.n6190 a_400_38200# 0.12fF
C13267 VP.n6191 a_400_38200# 0.14fF
C13268 VP.t178 a_400_38200# 0.02fF
C13269 VP.n6193 a_400_38200# 0.24fF
C13270 VP.n6194 a_400_38200# 0.91fF
C13271 VP.n6195 a_400_38200# 0.05fF
C13272 VP.n6196 a_400_38200# 0.10fF
C13273 VP.n6197 a_400_38200# 0.28fF
C13274 VP.n6198 a_400_38200# 0.15fF
C13275 VP.n6199 a_400_38200# 0.08fF
C13276 VP.n6200 a_400_38200# 0.14fF
C13277 VP.n6201 a_400_38200# 0.06fF
C13278 VP.n6202 a_400_38200# 0.06fF
C13279 VP.n6203 a_400_38200# 0.03fF
C13280 VP.n6204 a_400_38200# 0.05fF
C13281 VP.n6205 a_400_38200# 0.07fF
C13282 VP.n6206 a_400_38200# 0.19fF
C13283 VP.n6207 a_400_38200# 0.59fF
C13284 VP.n6208 a_400_38200# 0.34fF
C13285 VP.n6209 a_400_38200# 0.04fF
C13286 VP.n6210 a_400_38200# 0.02fF
C13287 VP.n6211 a_400_38200# 0.06fF
C13288 VP.n6212 a_400_38200# 0.30fF
C13289 VP.n6213 a_400_38200# 1.93fF
C13290 VP.n6214 a_400_38200# 0.12fF
C13291 VP.t719 a_400_38200# 0.02fF
C13292 VP.n6215 a_400_38200# 0.14fF
C13293 VP.t1313 a_400_38200# 0.02fF
C13294 VP.n6217 a_400_38200# 0.24fF
C13295 VP.n6218 a_400_38200# 0.35fF
C13296 VP.n6219 a_400_38200# 0.60fF
C13297 VP.n6220 a_400_38200# 2.47fF
C13298 VP.n6221 a_400_38200# 2.20fF
C13299 VP.t1133 a_400_38200# 0.02fF
C13300 VP.n6222 a_400_38200# 0.12fF
C13301 VP.n6223 a_400_38200# 0.14fF
C13302 VP.t1029 a_400_38200# 0.02fF
C13303 VP.n6225 a_400_38200# 0.24fF
C13304 VP.n6226 a_400_38200# 0.91fF
C13305 VP.n6227 a_400_38200# 0.05fF
C13306 VP.n6228 a_400_38200# 0.10fF
C13307 VP.n6229 a_400_38200# 0.28fF
C13308 VP.n6230 a_400_38200# 0.15fF
C13309 VP.n6231 a_400_38200# 0.08fF
C13310 VP.n6232 a_400_38200# 0.14fF
C13311 VP.n6233 a_400_38200# 0.06fF
C13312 VP.n6234 a_400_38200# 0.06fF
C13313 VP.n6235 a_400_38200# 0.03fF
C13314 VP.n6236 a_400_38200# 0.05fF
C13315 VP.n6237 a_400_38200# 0.07fF
C13316 VP.n6238 a_400_38200# 0.19fF
C13317 VP.n6239 a_400_38200# 0.59fF
C13318 VP.n6240 a_400_38200# 0.34fF
C13319 VP.n6241 a_400_38200# 0.04fF
C13320 VP.n6242 a_400_38200# 0.02fF
C13321 VP.n6243 a_400_38200# 0.06fF
C13322 VP.n6244 a_400_38200# 0.30fF
C13323 VP.n6245 a_400_38200# 1.93fF
C13324 VP.n6246 a_400_38200# 0.12fF
C13325 VP.t1041 a_400_38200# 0.02fF
C13326 VP.n6247 a_400_38200# 0.14fF
C13327 VP.t255 a_400_38200# 0.02fF
C13328 VP.n6249 a_400_38200# 0.24fF
C13329 VP.n6250 a_400_38200# 0.35fF
C13330 VP.n6251 a_400_38200# 0.60fF
C13331 VP.n6252 a_400_38200# 2.39fF
C13332 VP.n6253 a_400_38200# 1.79fF
C13333 VP.t55 a_400_38200# 0.02fF
C13334 VP.n6254 a_400_38200# 0.12fF
C13335 VP.n6255 a_400_38200# 0.14fF
C13336 VP.t1280 a_400_38200# 0.02fF
C13337 VP.n6257 a_400_38200# 0.24fF
C13338 VP.n6258 a_400_38200# 0.91fF
C13339 VP.n6259 a_400_38200# 0.05fF
C13340 VP.n6260 a_400_38200# 1.93fF
C13341 VP.n6261 a_400_38200# 2.72fF
C13342 VP.t651 a_400_38200# 0.02fF
C13343 VP.n6262 a_400_38200# 0.24fF
C13344 VP.n6263 a_400_38200# 0.35fF
C13345 VP.n6264 a_400_38200# 0.60fF
C13346 VP.n6265 a_400_38200# 0.12fF
C13347 VP.t25 a_400_38200# 0.02fF
C13348 VP.n6266 a_400_38200# 0.14fF
C13349 VP.n6268 a_400_38200# 0.02fF
C13350 VP.n6269 a_400_38200# 0.32fF
C13351 VP.n6270 a_400_38200# 0.04fF
C13352 VP.n6271 a_400_38200# 0.05fF
C13353 VP.n6272 a_400_38200# 0.04fF
C13354 VP.n6273 a_400_38200# 0.12fF
C13355 VP.n6274 a_400_38200# 0.09fF
C13356 VP.n6275 a_400_38200# 0.14fF
C13357 VP.n6276 a_400_38200# 0.08fF
C13358 VP.n6277 a_400_38200# 0.09fF
C13359 VP.n6278 a_400_38200# 0.07fF
C13360 VP.n6279 a_400_38200# 0.56fF
C13361 VP.n6280 a_400_38200# 0.20fF
C13362 VP.n6281 a_400_38200# 2.19fF
C13363 VP.t477 a_400_38200# 0.02fF
C13364 VP.n6282 a_400_38200# 0.12fF
C13365 VP.n6283 a_400_38200# 0.14fF
C13366 VP.t367 a_400_38200# 0.02fF
C13367 VP.n6285 a_400_38200# 0.24fF
C13368 VP.n6286 a_400_38200# 0.91fF
C13369 VP.n6287 a_400_38200# 0.05fF
C13370 VP.t24 a_400_38200# 34.79fF
C13371 VP.t730 a_400_38200# 0.02fF
C13372 VP.n6288 a_400_38200# 0.12fF
C13373 VP.n6289 a_400_38200# 0.14fF
C13374 VP.t634 a_400_38200# 0.02fF
C13375 VP.n6291 a_400_38200# 0.24fF
C13376 VP.n6292 a_400_38200# 0.91fF
C13377 VP.n6293 a_400_38200# 0.05fF
C13378 VP.t916 a_400_38200# 0.02fF
C13379 VP.n6294 a_400_38200# 0.24fF
C13380 VP.n6295 a_400_38200# 0.35fF
C13381 VP.n6296 a_400_38200# 0.60fF
C13382 VP.n6297 a_400_38200# 0.04fF
C13383 VP.n6298 a_400_38200# 0.08fF
C13384 VP.n6299 a_400_38200# 0.72fF
C13385 VP.n6300 a_400_38200# 0.09fF
C13386 VP.n6301 a_400_38200# 0.00fF
C13387 VP.n6302 a_400_38200# 1.22fF
C13388 VP.n6303 a_400_38200# 0.19fF
C13389 VP.n6305 a_400_38200# 1.72fF
C13390 VP.n6306 a_400_38200# 1.96fF
C13391 VP.n6307 a_400_38200# 1.04fF
C13392 VP.n6308 a_400_38200# 0.05fF
C13393 VP.n6309 a_400_38200# 0.03fF
C13394 VP.n6310 a_400_38200# 0.06fF
C13395 VP.n6311 a_400_38200# 0.06fF
C13396 VP.n6312 a_400_38200# 0.06fF
C13397 VP.n6313 a_400_38200# 0.07fF
C13398 VP.n6314 a_400_38200# 0.03fF
C13399 VP.n6315 a_400_38200# 0.05fF
C13400 VP.n6316 a_400_38200# 0.07fF
C13401 VP.n6317 a_400_38200# 0.19fF
C13402 VP.n6318 a_400_38200# 0.60fF
C13403 VP.n6319 a_400_38200# 0.76fF
C13404 VP.n6320 a_400_38200# 0.40fF
C13405 VP.n6321 a_400_38200# 0.03fF
C13406 VP.n6322 a_400_38200# 0.01fF
C13407 VP.t454 a_400_38200# 0.02fF
C13408 VP.n6323 a_400_38200# 0.25fF
C13409 VP.t162 a_400_38200# 0.02fF
C13410 VP.n6324 a_400_38200# 0.95fF
C13411 VP.n6325 a_400_38200# 0.70fF
C13412 VP.n6326 a_400_38200# 1.93fF
C13413 VP.n6327 a_400_38200# 2.97fF
C13414 VP.n6328 a_400_38200# 2.27fF
C13415 VP.t1246 a_400_38200# 0.02fF
C13416 VP.n6329 a_400_38200# 0.24fF
C13417 VP.n6330 a_400_38200# 0.35fF
C13418 VP.n6331 a_400_38200# 0.60fF
C13419 VP.n6332 a_400_38200# 0.12fF
C13420 VP.t658 a_400_38200# 0.02fF
C13421 VP.n6333 a_400_38200# 0.14fF
C13422 VP.n6335 a_400_38200# 0.04fF
C13423 VP.n6336 a_400_38200# 0.02fF
C13424 VP.n6337 a_400_38200# 0.06fF
C13425 VP.n6338 a_400_38200# 0.30fF
C13426 VP.n6339 a_400_38200# 0.10fF
C13427 VP.n6340 a_400_38200# 0.28fF
C13428 VP.n6341 a_400_38200# 0.06fF
C13429 VP.n6342 a_400_38200# 0.06fF
C13430 VP.n6343 a_400_38200# 0.03fF
C13431 VP.n6344 a_400_38200# 0.15fF
C13432 VP.n6345 a_400_38200# 0.08fF
C13433 VP.n6346 a_400_38200# 0.14fF
C13434 VP.n6347 a_400_38200# 0.03fF
C13435 VP.n6348 a_400_38200# 0.06fF
C13436 VP.n6349 a_400_38200# 0.06fF
C13437 VP.n6350 a_400_38200# 0.06fF
C13438 VP.n6351 a_400_38200# 0.06fF
C13439 VP.n6352 a_400_38200# 0.03fF
C13440 VP.n6353 a_400_38200# 0.05fF
C13441 VP.n6354 a_400_38200# 0.07fF
C13442 VP.n6355 a_400_38200# 0.19fF
C13443 VP.n6356 a_400_38200# 0.59fF
C13444 VP.n6357 a_400_38200# 0.34fF
C13445 VP.n6358 a_400_38200# 1.88fF
C13446 VP.t375 a_400_38200# 0.02fF
C13447 VP.n6359 a_400_38200# 0.24fF
C13448 VP.n6360 a_400_38200# 0.91fF
C13449 VP.n6361 a_400_38200# 0.05fF
C13450 VP.t760 a_400_38200# 0.02fF
C13451 VP.n6362 a_400_38200# 0.12fF
C13452 VP.n6363 a_400_38200# 0.14fF
C13453 VP.n6365 a_400_38200# 0.19fF
C13454 VP.n6366 a_400_38200# 0.10fF
C13455 VP.n6367 a_400_38200# 0.10fF
C13456 VP.n6368 a_400_38200# 0.18fF
C13457 VP.n6369 a_400_38200# 0.09fF
C13458 VP.n6370 a_400_38200# 0.04fF
C13459 VP.n6371 a_400_38200# 0.19fF
C13460 VP.n6372 a_400_38200# 0.26fF
C13461 VP.n6373 a_400_38200# 1.17fF
C13462 VP.n6374 a_400_38200# 0.06fF
C13463 VP.n6375 a_400_38200# 0.44fF
C13464 VP.n6376 a_400_38200# 0.13fF
C13465 VP.n6377 a_400_38200# 0.02fF
C13466 VP.n6378 a_400_38200# 1.81fF
C13467 VP.n6379 a_400_38200# 0.12fF
C13468 VP.t212 a_400_38200# 0.02fF
C13469 VP.n6380 a_400_38200# 0.14fF
C13470 VP.t801 a_400_38200# 0.02fF
C13471 VP.n6382 a_400_38200# 0.24fF
C13472 VP.n6383 a_400_38200# 0.35fF
C13473 VP.n6384 a_400_38200# 0.60fF
C13474 VP.n6385 a_400_38200# 3.18fF
C13475 VP.n6386 a_400_38200# 2.06fF
C13476 VP.n6387 a_400_38200# 1.98fF
C13477 VP.t1231 a_400_38200# 0.02fF
C13478 VP.n6388 a_400_38200# 0.24fF
C13479 VP.n6389 a_400_38200# 0.91fF
C13480 VP.n6390 a_400_38200# 0.05fF
C13481 VP.t307 a_400_38200# 0.02fF
C13482 VP.n6391 a_400_38200# 0.12fF
C13483 VP.n6392 a_400_38200# 0.14fF
C13484 VP.n6394 a_400_38200# 0.16fF
C13485 VP.n6395 a_400_38200# 0.19fF
C13486 VP.n6396 a_400_38200# 0.09fF
C13487 VP.n6397 a_400_38200# 0.04fF
C13488 VP.n6398 a_400_38200# 0.14fF
C13489 VP.n6399 a_400_38200# 0.64fF
C13490 VP.n6400 a_400_38200# 1.32fF
C13491 VP.n6401 a_400_38200# 1.81fF
C13492 VP.n6402 a_400_38200# 0.12fF
C13493 VP.t1067 a_400_38200# 0.02fF
C13494 VP.n6403 a_400_38200# 0.14fF
C13495 VP.t353 a_400_38200# 0.02fF
C13496 VP.n6405 a_400_38200# 0.24fF
C13497 VP.n6406 a_400_38200# 0.35fF
C13498 VP.n6407 a_400_38200# 0.60fF
C13499 VP.n6408 a_400_38200# 2.97fF
C13500 VP.n6409 a_400_38200# 2.27fF
C13501 VP.n6410 a_400_38200# 2.00fF
C13502 VP.t786 a_400_38200# 0.02fF
C13503 VP.n6411 a_400_38200# 0.24fF
C13504 VP.n6412 a_400_38200# 0.91fF
C13505 VP.n6413 a_400_38200# 0.05fF
C13506 VP.t1154 a_400_38200# 0.02fF
C13507 VP.n6414 a_400_38200# 0.12fF
C13508 VP.n6415 a_400_38200# 0.14fF
C13509 VP.n6417 a_400_38200# 0.24fF
C13510 VP.t1184 a_400_38200# 0.02fF
C13511 VP.n6418 a_400_38200# 0.36fF
C13512 VP.n6419 a_400_38200# 0.36fF
C13513 VP.n6420 a_400_38200# 0.67fF
C13514 VP.n6421 a_400_38200# 0.16fF
C13515 VP.n6422 a_400_38200# 0.19fF
C13516 VP.n6423 a_400_38200# 0.09fF
C13517 VP.n6424 a_400_38200# 0.04fF
C13518 VP.n6425 a_400_38200# 0.14fF
C13519 VP.n6426 a_400_38200# 0.64fF
C13520 VP.n6427 a_400_38200# 1.32fF
C13521 VP.n6428 a_400_38200# 1.81fF
C13522 VP.n6429 a_400_38200# 2.97fF
C13523 VP.n6430 a_400_38200# 2.27fF
C13524 VP.n6431 a_400_38200# 0.75fF
C13525 VP.n6432 a_400_38200# 0.24fF
C13526 VP.t757 a_400_38200# 0.02fF
C13527 VP.n6433 a_400_38200# 0.35fF
C13528 VP.n6434 a_400_38200# 0.63fF
C13529 VP.n6435 a_400_38200# 0.40fF
C13530 VP.n6436 a_400_38200# 0.40fF
C13531 VP.n6437 a_400_38200# 0.12fF
C13532 VP.t160 a_400_38200# 0.02fF
C13533 VP.n6438 a_400_38200# 0.14fF
C13534 VP.t261 a_400_38200# 0.02fF
C13535 VP.n6440 a_400_38200# 0.12fF
C13536 VP.n6441 a_400_38200# 0.14fF
C13537 VP.n6443 a_400_38200# 0.16fF
C13538 VP.n6444 a_400_38200# 0.19fF
C13539 VP.n6445 a_400_38200# 0.09fF
C13540 VP.n6446 a_400_38200# 0.04fF
C13541 VP.n6447 a_400_38200# 0.14fF
C13542 VP.n6448 a_400_38200# 0.64fF
C13543 VP.n6449 a_400_38200# 1.32fF
C13544 VP.n6450 a_400_38200# 1.81fF
C13545 VP.n6451 a_400_38200# 0.12fF
C13546 VP.t641 a_400_38200# 0.02fF
C13547 VP.n6452 a_400_38200# 0.14fF
C13548 VP.t1228 a_400_38200# 0.02fF
C13549 VP.n6454 a_400_38200# 0.24fF
C13550 VP.n6455 a_400_38200# 0.35fF
C13551 VP.n6456 a_400_38200# 0.60fF
C13552 VP.n6457 a_400_38200# 2.97fF
C13553 VP.n6458 a_400_38200# 2.27fF
C13554 VP.n6459 a_400_38200# 2.00fF
C13555 VP.t356 a_400_38200# 0.02fF
C13556 VP.n6460 a_400_38200# 0.24fF
C13557 VP.n6461 a_400_38200# 0.91fF
C13558 VP.n6462 a_400_38200# 0.05fF
C13559 VP.t670 a_400_38200# 0.02fF
C13560 VP.n6463 a_400_38200# 0.12fF
C13561 VP.n6464 a_400_38200# 0.14fF
C13562 VP.n6466 a_400_38200# 0.09fF
C13563 VP.n6467 a_400_38200# 0.03fF
C13564 VP.n6468 a_400_38200# 0.04fF
C13565 VP.n6469 a_400_38200# 0.37fF
C13566 VP.n6470 a_400_38200# 0.11fF
C13567 VP.n6471 a_400_38200# 0.05fF
C13568 VP.n6472 a_400_38200# 0.08fF
C13569 VP.n6473 a_400_38200# 0.10fF
C13570 VP.n6474 a_400_38200# 0.06fF
C13571 VP.n6475 a_400_38200# 0.08fF
C13572 VP.n6476 a_400_38200# 0.19fF
C13573 VP.n6477 a_400_38200# 0.06fF
C13574 VP.n6478 a_400_38200# 0.15fF
C13575 VP.n6479 a_400_38200# 0.14fF
C13576 VP.n6480 a_400_38200# 0.13fF
C13577 VP.n6481 a_400_38200# 0.12fF
C13578 VP.n6482 a_400_38200# 0.05fF
C13579 VP.n6483 a_400_38200# 0.17fF
C13580 VP.n6484 a_400_38200# 0.26fF
C13581 VP.n6485 a_400_38200# 0.37fF
C13582 VP.n6486 a_400_38200# 0.27fF
C13583 VP.n6487 a_400_38200# 2.05fF
C13584 VP.n6488 a_400_38200# 0.12fF
C13585 VP.t434 a_400_38200# 0.02fF
C13586 VP.n6489 a_400_38200# 0.14fF
C13587 VP.t1015 a_400_38200# 0.02fF
C13588 VP.n6491 a_400_38200# 0.24fF
C13589 VP.n6492 a_400_38200# 0.35fF
C13590 VP.n6493 a_400_38200# 0.60fF
C13591 VP.n6494 a_400_38200# 2.87fF
C13592 VP.n6495 a_400_38200# 2.00fF
C13593 VP.t137 a_400_38200# 0.02fF
C13594 VP.n6496 a_400_38200# 0.24fF
C13595 VP.n6497 a_400_38200# 0.91fF
C13596 VP.n6498 a_400_38200# 0.05fF
C13597 VP.t1078 a_400_38200# 0.02fF
C13598 VP.n6499 a_400_38200# 0.12fF
C13599 VP.n6500 a_400_38200# 0.14fF
C13600 VP.n6502 a_400_38200# 15.28fF
C13601 VP.n6503 a_400_38200# 0.10fF
C13602 VP.n6504 a_400_38200# 0.28fF
C13603 VP.n6505 a_400_38200# 0.06fF
C13604 VP.n6506 a_400_38200# 0.06fF
C13605 VP.n6507 a_400_38200# 0.03fF
C13606 VP.n6508 a_400_38200# 0.15fF
C13607 VP.n6509 a_400_38200# 0.08fF
C13608 VP.n6510 a_400_38200# 0.14fF
C13609 VP.n6511 a_400_38200# 0.03fF
C13610 VP.n6512 a_400_38200# 0.06fF
C13611 VP.n6513 a_400_38200# 0.06fF
C13612 VP.n6514 a_400_38200# 0.06fF
C13613 VP.n6515 a_400_38200# 0.06fF
C13614 VP.n6516 a_400_38200# 0.03fF
C13615 VP.n6517 a_400_38200# 0.05fF
C13616 VP.n6518 a_400_38200# 0.07fF
C13617 VP.n6519 a_400_38200# 0.19fF
C13618 VP.n6520 a_400_38200# 0.59fF
C13619 VP.n6521 a_400_38200# 0.34fF
C13620 VP.n6522 a_400_38200# 0.04fF
C13621 VP.n6523 a_400_38200# 0.02fF
C13622 VP.n6524 a_400_38200# 0.06fF
C13623 VP.n6525 a_400_38200# 0.30fF
C13624 VP.n6526 a_400_38200# 1.93fF
C13625 VP.n6527 a_400_38200# 0.12fF
C13626 VP.t1304 a_400_38200# 0.02fF
C13627 VP.n6528 a_400_38200# 0.14fF
C13628 VP.t590 a_400_38200# 0.02fF
C13629 VP.n6530 a_400_38200# 0.24fF
C13630 VP.n6531 a_400_38200# 0.35fF
C13631 VP.n6532 a_400_38200# 0.60fF
C13632 VP.n6533 a_400_38200# 0.56fF
C13633 VP.n6534 a_400_38200# 1.24fF
C13634 VP.n6535 a_400_38200# 0.54fF
C13635 VP.n6536 a_400_38200# 0.22fF
C13636 VP.n6537 a_400_38200# 1.73fF
C13637 VP.t1344 a_400_38200# 0.02fF
C13638 VP.n6538 a_400_38200# 0.12fF
C13639 VP.n6539 a_400_38200# 0.14fF
C13640 VP.t1013 a_400_38200# 0.02fF
C13641 VP.n6541 a_400_38200# 0.24fF
C13642 VP.n6542 a_400_38200# 0.91fF
C13643 VP.n6543 a_400_38200# 0.05fF
C13644 VP.n6544 a_400_38200# 0.10fF
C13645 VP.n6545 a_400_38200# 0.28fF
C13646 VP.n6546 a_400_38200# 0.06fF
C13647 VP.n6547 a_400_38200# 0.06fF
C13648 VP.n6548 a_400_38200# 0.03fF
C13649 VP.n6549 a_400_38200# 0.15fF
C13650 VP.n6550 a_400_38200# 0.08fF
C13651 VP.n6551 a_400_38200# 0.14fF
C13652 VP.n6552 a_400_38200# 0.03fF
C13653 VP.n6553 a_400_38200# 0.06fF
C13654 VP.n6554 a_400_38200# 0.06fF
C13655 VP.n6555 a_400_38200# 0.06fF
C13656 VP.n6556 a_400_38200# 0.06fF
C13657 VP.n6557 a_400_38200# 0.03fF
C13658 VP.n6558 a_400_38200# 0.05fF
C13659 VP.n6559 a_400_38200# 0.07fF
C13660 VP.n6560 a_400_38200# 0.19fF
C13661 VP.n6561 a_400_38200# 0.59fF
C13662 VP.n6562 a_400_38200# 0.34fF
C13663 VP.n6563 a_400_38200# 0.04fF
C13664 VP.n6564 a_400_38200# 0.02fF
C13665 VP.n6565 a_400_38200# 0.06fF
C13666 VP.n6566 a_400_38200# 0.30fF
C13667 VP.n6567 a_400_38200# 1.93fF
C13668 VP.n6568 a_400_38200# 0.12fF
C13669 VP.t857 a_400_38200# 0.02fF
C13670 VP.n6569 a_400_38200# 0.14fF
C13671 VP.t123 a_400_38200# 0.02fF
C13672 VP.n6571 a_400_38200# 0.24fF
C13673 VP.n6572 a_400_38200# 0.35fF
C13674 VP.n6573 a_400_38200# 0.60fF
C13675 VP.n6574 a_400_38200# 0.72fF
C13676 VP.n6575 a_400_38200# 1.24fF
C13677 VP.n6576 a_400_38200# 0.54fF
C13678 VP.n6577 a_400_38200# 0.22fF
C13679 VP.n6578 a_400_38200# 1.73fF
C13680 VP.t896 a_400_38200# 0.02fF
C13681 VP.n6579 a_400_38200# 0.12fF
C13682 VP.n6580 a_400_38200# 0.14fF
C13683 VP.t569 a_400_38200# 0.02fF
C13684 VP.n6582 a_400_38200# 0.24fF
C13685 VP.n6583 a_400_38200# 0.91fF
C13686 VP.n6584 a_400_38200# 0.05fF
C13687 VP.n6585 a_400_38200# 0.10fF
C13688 VP.n6586 a_400_38200# 0.28fF
C13689 VP.n6587 a_400_38200# 0.06fF
C13690 VP.n6588 a_400_38200# 0.06fF
C13691 VP.n6589 a_400_38200# 0.03fF
C13692 VP.n6590 a_400_38200# 0.15fF
C13693 VP.n6591 a_400_38200# 0.08fF
C13694 VP.n6592 a_400_38200# 0.14fF
C13695 VP.n6593 a_400_38200# 0.03fF
C13696 VP.n6594 a_400_38200# 0.06fF
C13697 VP.n6595 a_400_38200# 0.06fF
C13698 VP.n6596 a_400_38200# 0.06fF
C13699 VP.n6597 a_400_38200# 0.06fF
C13700 VP.n6598 a_400_38200# 0.03fF
C13701 VP.n6599 a_400_38200# 0.05fF
C13702 VP.n6600 a_400_38200# 0.07fF
C13703 VP.n6601 a_400_38200# 0.19fF
C13704 VP.n6602 a_400_38200# 0.59fF
C13705 VP.n6603 a_400_38200# 0.34fF
C13706 VP.n6604 a_400_38200# 0.04fF
C13707 VP.n6605 a_400_38200# 0.02fF
C13708 VP.n6606 a_400_38200# 0.06fF
C13709 VP.n6607 a_400_38200# 0.30fF
C13710 VP.n6608 a_400_38200# 1.93fF
C13711 VP.n6609 a_400_38200# 0.12fF
C13712 VP.t1100 a_400_38200# 0.02fF
C13713 VP.n6610 a_400_38200# 0.14fF
C13714 VP.t389 a_400_38200# 0.02fF
C13715 VP.n6612 a_400_38200# 0.24fF
C13716 VP.n6613 a_400_38200# 0.35fF
C13717 VP.n6614 a_400_38200# 0.60fF
C13718 VP.n6615 a_400_38200# 0.71fF
C13719 VP.n6616 a_400_38200# 1.39fF
C13720 VP.n6617 a_400_38200# 0.54fF
C13721 VP.n6618 a_400_38200# 0.21fF
C13722 VP.n6619 a_400_38200# 1.73fF
C13723 VP.t444 a_400_38200# 0.02fF
C13724 VP.n6620 a_400_38200# 0.12fF
C13725 VP.n6621 a_400_38200# 0.14fF
C13726 VP.t826 a_400_38200# 0.02fF
C13727 VP.n6623 a_400_38200# 0.24fF
C13728 VP.n6624 a_400_38200# 0.91fF
C13729 VP.n6625 a_400_38200# 0.05fF
C13730 VP.n6626 a_400_38200# 0.06fF
C13731 VP.n6627 a_400_38200# 0.06fF
C13732 VP.n6628 a_400_38200# 0.03fF
C13733 VP.n6629 a_400_38200# 0.10fF
C13734 VP.n6630 a_400_38200# 0.17fF
C13735 VP.n6631 a_400_38200# 0.10fF
C13736 VP.n6632 a_400_38200# 0.13fF
C13737 VP.n6633 a_400_38200# 0.02fF
C13738 VP.n6634 a_400_38200# 0.04fF
C13739 VP.n6635 a_400_38200# 0.06fF
C13740 VP.n6636 a_400_38200# 0.09fF
C13741 VP.n6637 a_400_38200# 0.10fF
C13742 VP.n6638 a_400_38200# 0.05fF
C13743 VP.n6639 a_400_38200# 0.19fF
C13744 VP.n6640 a_400_38200# 0.16fF
C13745 VP.n6641 a_400_38200# 0.04fF
C13746 VP.n6642 a_400_38200# 0.05fF
C13747 VP.n6643 a_400_38200# 0.04fF
C13748 VP.n6644 a_400_38200# 0.12fF
C13749 VP.n6645 a_400_38200# 0.09fF
C13750 VP.n6646 a_400_38200# 0.14fF
C13751 VP.n6647 a_400_38200# 0.56fF
C13752 VP.n6648 a_400_38200# 0.10fF
C13753 VP.n6649 a_400_38200# 1.93fF
C13754 VP.n6650 a_400_38200# 0.12fF
C13755 VP.t622 a_400_38200# 0.02fF
C13756 VP.n6651 a_400_38200# 0.14fF
C13757 VP.t1206 a_400_38200# 0.02fF
C13758 VP.n6653 a_400_38200# 0.24fF
C13759 VP.n6654 a_400_38200# 0.35fF
C13760 VP.n6655 a_400_38200# 0.60fF
C13761 VP.n6656 a_400_38200# 0.18fF
C13762 VP.n6657 a_400_38200# 0.45fF
C13763 VP.n6658 a_400_38200# 0.06fF
C13764 VP.n6659 a_400_38200# 0.01fF
C13765 VP.n6660 a_400_38200# 0.01fF
C13766 VP.n6661 a_400_38200# 0.04fF
C13767 VP.n6662 a_400_38200# 0.02fF
C13768 VP.n6663 a_400_38200# 0.07fF
C13769 VP.n6664 a_400_38200# 0.04fF
C13770 VP.n6665 a_400_38200# 0.14fF
C13771 VP.n6666 a_400_38200# 0.45fF
C13772 VP.n6667 a_400_38200# 1.46fF
C13773 VP.n6668 a_400_38200# 1.78fF
C13774 VP.t705 a_400_38200# 0.02fF
C13775 VP.n6669 a_400_38200# 0.12fF
C13776 VP.n6670 a_400_38200# 0.14fF
C13777 VP.t338 a_400_38200# 0.02fF
C13778 VP.n6672 a_400_38200# 0.24fF
C13779 VP.n6673 a_400_38200# 0.91fF
C13780 VP.n6674 a_400_38200# 0.05fF
C13781 VP.n6675 a_400_38200# 1.93fF
C13782 VP.n6676 a_400_38200# 0.18fF
C13783 VP.n6677 a_400_38200# 0.45fF
C13784 VP.n6678 a_400_38200# 0.06fF
C13785 VP.n6679 a_400_38200# 0.01fF
C13786 VP.n6680 a_400_38200# 0.01fF
C13787 VP.n6681 a_400_38200# 0.04fF
C13788 VP.n6682 a_400_38200# 0.02fF
C13789 VP.n6683 a_400_38200# 0.07fF
C13790 VP.n6684 a_400_38200# 0.04fF
C13791 VP.n6685 a_400_38200# 0.14fF
C13792 VP.n6686 a_400_38200# 0.45fF
C13793 VP.n6687 a_400_38200# 1.46fF
C13794 VP.t304 a_400_38200# 0.02fF
C13795 VP.n6688 a_400_38200# 0.24fF
C13796 VP.n6689 a_400_38200# 0.35fF
C13797 VP.n6690 a_400_38200# 0.60fF
C13798 VP.n6691 a_400_38200# 0.12fF
C13799 VP.t1084 a_400_38200# 0.02fF
C13800 VP.n6692 a_400_38200# 0.14fF
C13801 VP.n6694 a_400_38200# 0.10fF
C13802 VP.n6695 a_400_38200# 0.17fF
C13803 VP.n6696 a_400_38200# 0.06fF
C13804 VP.n6697 a_400_38200# 0.06fF
C13805 VP.n6698 a_400_38200# 0.03fF
C13806 VP.n6699 a_400_38200# 0.10fF
C13807 VP.n6700 a_400_38200# 0.13fF
C13808 VP.n6701 a_400_38200# 0.13fF
C13809 VP.n6702 a_400_38200# 0.04fF
C13810 VP.n6703 a_400_38200# 0.05fF
C13811 VP.n6704 a_400_38200# 0.04fF
C13812 VP.n6705 a_400_38200# 0.09fF
C13813 VP.n6706 a_400_38200# 0.09fF
C13814 VP.n6707 a_400_38200# 0.05fF
C13815 VP.n6708 a_400_38200# 0.19fF
C13816 VP.n6709 a_400_38200# 0.12fF
C13817 VP.n6710 a_400_38200# 0.09fF
C13818 VP.n6711 a_400_38200# 0.14fF
C13819 VP.n6712 a_400_38200# 0.04fF
C13820 VP.n6713 a_400_38200# 0.02fF
C13821 VP.n6714 a_400_38200# 0.06fF
C13822 VP.n6715 a_400_38200# 0.56fF
C13823 VP.n6716 a_400_38200# 0.10fF
C13824 VP.n6717 a_400_38200# 1.78fF
C13825 VP.t1116 a_400_38200# 0.02fF
C13826 VP.n6718 a_400_38200# 0.12fF
C13827 VP.n6719 a_400_38200# 0.14fF
C13828 VP.t731 a_400_38200# 0.02fF
C13829 VP.n6721 a_400_38200# 0.24fF
C13830 VP.n6722 a_400_38200# 0.91fF
C13831 VP.n6723 a_400_38200# 0.05fF
C13832 VP.n6724 a_400_38200# 1.93fF
C13833 VP.n6725 a_400_38200# 0.18fF
C13834 VP.n6726 a_400_38200# 0.45fF
C13835 VP.n6727 a_400_38200# 0.06fF
C13836 VP.n6728 a_400_38200# 0.01fF
C13837 VP.n6729 a_400_38200# 0.01fF
C13838 VP.n6730 a_400_38200# 0.04fF
C13839 VP.n6731 a_400_38200# 0.02fF
C13840 VP.n6732 a_400_38200# 0.07fF
C13841 VP.n6733 a_400_38200# 0.04fF
C13842 VP.n6734 a_400_38200# 0.14fF
C13843 VP.n6735 a_400_38200# 0.53fF
C13844 VP.n6736 a_400_38200# 1.62fF
C13845 VP.t783 a_400_38200# 0.02fF
C13846 VP.n6737 a_400_38200# 0.24fF
C13847 VP.n6738 a_400_38200# 0.35fF
C13848 VP.n6739 a_400_38200# 0.60fF
C13849 VP.n6740 a_400_38200# 0.12fF
C13850 VP.t191 a_400_38200# 0.02fF
C13851 VP.n6741 a_400_38200# 0.14fF
C13852 VP.n6743 a_400_38200# 0.10fF
C13853 VP.n6744 a_400_38200# 0.17fF
C13854 VP.n6745 a_400_38200# 0.06fF
C13855 VP.n6746 a_400_38200# 0.06fF
C13856 VP.n6747 a_400_38200# 0.03fF
C13857 VP.n6748 a_400_38200# 0.10fF
C13858 VP.n6749 a_400_38200# 0.13fF
C13859 VP.n6750 a_400_38200# 0.14fF
C13860 VP.n6751 a_400_38200# 0.04fF
C13861 VP.n6752 a_400_38200# 0.02fF
C13862 VP.n6753 a_400_38200# 0.03fF
C13863 VP.n6754 a_400_38200# 0.03fF
C13864 VP.n6755 a_400_38200# 0.05fF
C13865 VP.n6756 a_400_38200# 0.03fF
C13866 VP.n6757 a_400_38200# 0.04fF
C13867 VP.n6758 a_400_38200# 0.20fF
C13868 VP.n6759 a_400_38200# 0.14fF
C13869 VP.n6760 a_400_38200# 0.02fF
C13870 VP.n6761 a_400_38200# 0.07fF
C13871 VP.n6762 a_400_38200# 0.13fF
C13872 VP.n6763 a_400_38200# 0.04fF
C13873 VP.n6764 a_400_38200# 0.02fF
C13874 VP.n6765 a_400_38200# 0.06fF
C13875 VP.n6766 a_400_38200# 0.55fF
C13876 VP.n6767 a_400_38200# 0.10fF
C13877 VP.n6768 a_400_38200# 1.95fF
C13878 VP.t223 a_400_38200# 0.02fF
C13879 VP.n6769 a_400_38200# 0.12fF
C13880 VP.n6770 a_400_38200# 0.14fF
C13881 VP.t1210 a_400_38200# 0.02fF
C13882 VP.n6772 a_400_38200# 0.24fF
C13883 VP.n6773 a_400_38200# 0.91fF
C13884 VP.n6774 a_400_38200# 0.05fF
C13885 VP.t159 a_400_38200# 35.17fF
C13886 VP.t1040 a_400_38200# 0.02fF
C13887 VP.n6775 a_400_38200# 1.21fF
C13888 VP.n6776 a_400_38200# 0.25fF
C13889 VP.n6777 a_400_38200# 26.29fF
C13890 VP.n6778 a_400_38200# 26.29fF
C13891 VP.n6779 a_400_38200# 0.76fF
C13892 VP.n6780 a_400_38200# 0.27fF
C13893 VP.n6781 a_400_38200# 0.59fF
C13894 VP.n6782 a_400_38200# 0.10fF
C13895 VP.n6783 a_400_38200# 3.02fF
C13896 VP.t122 a_400_38200# 15.72fF
C13897 VP.n6784 a_400_38200# 1.15fF
C13898 VP.n6786 a_400_38200# 13.70fF
C13899 VP.n6788 a_400_38200# 1.99fF
C13900 VP.n6789 a_400_38200# 4.39fF
C13901 VP.n6790 a_400_38200# 0.03fF
C13902 VP.n6791 a_400_38200# 0.05fF
C13903 VP.n6792 a_400_38200# 0.07fF
C13904 VP.n6793 a_400_38200# 0.03fF
C13905 VP.n6794 a_400_38200# 0.06fF
C13906 VP.n6795 a_400_38200# 0.06fF
C13907 VP.n6796 a_400_38200# 0.06fF
C13908 VP.n6797 a_400_38200# 0.07fF
C13909 VP.n6798 a_400_38200# 0.57fF
C13910 VP.n6799 a_400_38200# 1.88fF
C13911 VP.n6800 a_400_38200# 0.92fF
C13912 VP.n6801 a_400_38200# 2.63fF
C13913 VP.n6802 a_400_38200# 0.10fF
C13914 VP.n6803 a_400_38200# 0.28fF
C13915 VP.n6804 a_400_38200# 0.15fF
C13916 VP.n6805 a_400_38200# 0.08fF
C13917 VP.n6806 a_400_38200# 0.14fF
C13918 VP.n6807 a_400_38200# 0.06fF
C13919 VP.n6808 a_400_38200# 0.06fF
C13920 VP.n6809 a_400_38200# 0.03fF
C13921 VP.n6810 a_400_38200# 0.05fF
C13922 VP.n6811 a_400_38200# 0.07fF
C13923 VP.n6812 a_400_38200# 0.19fF
C13924 VP.n6813 a_400_38200# 0.59fF
C13925 VP.n6814 a_400_38200# 0.34fF
C13926 VP.n6815 a_400_38200# 0.04fF
C13927 VP.n6816 a_400_38200# 0.02fF
C13928 VP.n6817 a_400_38200# 0.06fF
C13929 VP.n6818 a_400_38200# 0.30fF
C13930 VP.n6819 a_400_38200# 0.12fF
C13931 VP.t476 a_400_38200# 0.02fF
C13932 VP.n6820 a_400_38200# 0.14fF
C13933 VP.n6822 a_400_38200# 1.93fF
C13934 VP.t407 a_400_38200# 0.02fF
C13935 VP.n6823 a_400_38200# 0.24fF
C13936 VP.n6824 a_400_38200# 0.35fF
C13937 VP.n6825 a_400_38200# 0.60fF
C13938 VP.n6826 a_400_38200# 0.12fF
C13939 VP.t1190 a_400_38200# 0.02fF
C13940 VP.n6827 a_400_38200# 0.14fF
C13941 VP.n6829 a_400_38200# 0.04fF
C13942 VP.n6830 a_400_38200# 0.02fF
C13943 VP.n6831 a_400_38200# 0.06fF
C13944 VP.n6832 a_400_38200# 0.30fF
C13945 VP.n6833 a_400_38200# 0.10fF
C13946 VP.n6834 a_400_38200# 0.28fF
C13947 VP.n6835 a_400_38200# 0.15fF
C13948 VP.n6836 a_400_38200# 0.08fF
C13949 VP.n6837 a_400_38200# 0.14fF
C13950 VP.n6838 a_400_38200# 0.06fF
C13951 VP.n6839 a_400_38200# 0.06fF
C13952 VP.n6840 a_400_38200# 0.03fF
C13953 VP.n6841 a_400_38200# 0.05fF
C13954 VP.n6842 a_400_38200# 0.07fF
C13955 VP.n6843 a_400_38200# 0.19fF
C13956 VP.n6844 a_400_38200# 0.59fF
C13957 VP.n6845 a_400_38200# 0.34fF
C13958 VP.n6846 a_400_38200# 2.18fF
C13959 VP.t100 a_400_38200# 0.02fF
C13960 VP.n6847 a_400_38200# 0.24fF
C13961 VP.n6848 a_400_38200# 0.91fF
C13962 VP.n6849 a_400_38200# 0.05fF
C13963 VP.t232 a_400_38200# 0.02fF
C13964 VP.n6850 a_400_38200# 0.12fF
C13965 VP.n6851 a_400_38200# 0.14fF
C13966 VP.n6853 a_400_38200# 0.10fF
C13967 VP.n6854 a_400_38200# 0.10fF
C13968 VP.n6855 a_400_38200# 0.18fF
C13969 VP.n6856 a_400_38200# 0.09fF
C13970 VP.n6857 a_400_38200# 0.04fF
C13971 VP.n6858 a_400_38200# 0.26fF
C13972 VP.n6859 a_400_38200# 1.17fF
C13973 VP.n6860 a_400_38200# 0.06fF
C13974 VP.n6861 a_400_38200# 0.44fF
C13975 VP.n6862 a_400_38200# 0.13fF
C13976 VP.n6863 a_400_38200# 0.02fF
C13977 VP.n6864 a_400_38200# 1.81fF
C13978 VP.n6865 a_400_38200# 0.12fF
C13979 VP.t736 a_400_38200# 0.02fF
C13980 VP.n6866 a_400_38200# 0.14fF
C13981 VP.t1326 a_400_38200# 0.02fF
C13982 VP.n6868 a_400_38200# 0.24fF
C13983 VP.n6869 a_400_38200# 0.35fF
C13984 VP.n6870 a_400_38200# 0.60fF
C13985 VP.n6871 a_400_38200# 2.28fF
C13986 VP.t1046 a_400_38200# 0.02fF
C13987 VP.n6872 a_400_38200# 0.24fF
C13988 VP.n6873 a_400_38200# 0.91fF
C13989 VP.n6874 a_400_38200# 0.05fF
C13990 VP.t1087 a_400_38200# 0.02fF
C13991 VP.n6875 a_400_38200# 0.12fF
C13992 VP.n6876 a_400_38200# 0.14fF
C13993 VP.n6878 a_400_38200# 0.06fF
C13994 VP.n6879 a_400_38200# 0.09fF
C13995 VP.n6880 a_400_38200# 0.09fF
C13996 VP.n6881 a_400_38200# 1.45fF
C13997 VP.n6882 a_400_38200# 0.14fF
C13998 VP.n6883 a_400_38200# 0.07fF
C13999 VP.n6884 a_400_38200# 0.72fF
C14000 VP.n6885 a_400_38200# 1.81fF
C14001 VP.n6886 a_400_38200# 0.12fF
C14002 VP.t285 a_400_38200# 0.02fF
C14003 VP.n6887 a_400_38200# 0.14fF
C14004 VP.t875 a_400_38200# 0.02fF
C14005 VP.n6889 a_400_38200# 0.24fF
C14006 VP.n6890 a_400_38200# 0.35fF
C14007 VP.n6891 a_400_38200# 0.60fF
C14008 VP.n6892 a_400_38200# 2.30fF
C14009 VP.t597 a_400_38200# 0.02fF
C14010 VP.n6893 a_400_38200# 0.24fF
C14011 VP.n6894 a_400_38200# 0.91fF
C14012 VP.n6895 a_400_38200# 0.05fF
C14013 VP.t644 a_400_38200# 0.02fF
C14014 VP.n6896 a_400_38200# 0.12fF
C14015 VP.n6897 a_400_38200# 0.14fF
C14016 VP.n6899 a_400_38200# 0.06fF
C14017 VP.n6900 a_400_38200# 0.25fF
C14018 VP.n6901 a_400_38200# 0.45fF
C14019 VP.n6902 a_400_38200# 0.03fF
C14020 VP.n6903 a_400_38200# 0.05fF
C14021 VP.n6904 a_400_38200# 0.07fF
C14022 VP.n6905 a_400_38200# 0.06fF
C14023 VP.n6906 a_400_38200# 0.06fF
C14024 VP.n6907 a_400_38200# 0.19fF
C14025 VP.n6908 a_400_38200# 0.59fF
C14026 VP.n6909 a_400_38200# 0.34fF
C14027 VP.n6910 a_400_38200# 0.05fF
C14028 VP.n6911 a_400_38200# 0.30fF
C14029 VP.n6912 a_400_38200# 1.93fF
C14030 VP.n6913 a_400_38200# 0.12fF
C14031 VP.t1137 a_400_38200# 0.02fF
C14032 VP.n6914 a_400_38200# 0.14fF
C14033 VP.t428 a_400_38200# 0.02fF
C14034 VP.n6916 a_400_38200# 0.24fF
C14035 VP.n6917 a_400_38200# 0.35fF
C14036 VP.n6918 a_400_38200# 0.60fF
C14037 VP.n6919 a_400_38200# 2.23fF
C14038 VP.n6920 a_400_38200# 2.04fF
C14039 VP.t129 a_400_38200# 0.02fF
C14040 VP.n6921 a_400_38200# 0.24fF
C14041 VP.n6922 a_400_38200# 0.91fF
C14042 VP.n6923 a_400_38200# 0.05fF
C14043 VP.t196 a_400_38200# 0.02fF
C14044 VP.n6924 a_400_38200# 0.12fF
C14045 VP.n6925 a_400_38200# 0.14fF
C14046 VP.n6927 a_400_38200# 0.24fF
C14047 VP.t996 a_400_38200# 0.02fF
C14048 VP.n6928 a_400_38200# 0.36fF
C14049 VP.n6929 a_400_38200# 0.36fF
C14050 VP.n6930 a_400_38200# 0.67fF
C14051 VP.n6931 a_400_38200# 0.06fF
C14052 VP.n6932 a_400_38200# 0.09fF
C14053 VP.n6933 a_400_38200# 0.09fF
C14054 VP.n6934 a_400_38200# 1.45fF
C14055 VP.n6935 a_400_38200# 0.14fF
C14056 VP.n6936 a_400_38200# 0.07fF
C14057 VP.n6937 a_400_38200# 0.72fF
C14058 VP.n6938 a_400_38200# 1.81fF
C14059 VP.n6939 a_400_38200# 1.06fF
C14060 VP.n6940 a_400_38200# 0.24fF
C14061 VP.t1284 a_400_38200# 0.02fF
C14062 VP.n6941 a_400_38200# 0.35fF
C14063 VP.n6942 a_400_38200# 0.63fF
C14064 VP.n6943 a_400_38200# 0.40fF
C14065 VP.n6944 a_400_38200# 0.40fF
C14066 VP.n6945 a_400_38200# 0.12fF
C14067 VP.t689 a_400_38200# 0.02fF
C14068 VP.n6946 a_400_38200# 0.14fF
C14069 VP.t1049 a_400_38200# 0.02fF
C14070 VP.n6948 a_400_38200# 0.12fF
C14071 VP.n6949 a_400_38200# 0.14fF
C14072 VP.n6951 a_400_38200# 1.93fF
C14073 VP.n6952 a_400_38200# 2.23fF
C14074 VP.t839 a_400_38200# 0.02fF
C14075 VP.n6953 a_400_38200# 0.24fF
C14076 VP.n6954 a_400_38200# 0.35fF
C14077 VP.n6955 a_400_38200# 0.60fF
C14078 VP.n6956 a_400_38200# 0.12fF
C14079 VP.t245 a_400_38200# 0.02fF
C14080 VP.n6957 a_400_38200# 0.14fF
C14081 VP.n6959 a_400_38200# 0.07fF
C14082 VP.n6960 a_400_38200# 0.30fF
C14083 VP.n6961 a_400_38200# 0.06fF
C14084 VP.n6962 a_400_38200# 0.25fF
C14085 VP.n6963 a_400_38200# 0.45fF
C14086 VP.n6964 a_400_38200# 0.06fF
C14087 VP.n6965 a_400_38200# 0.06fF
C14088 VP.n6966 a_400_38200# 0.03fF
C14089 VP.n6967 a_400_38200# 0.05fF
C14090 VP.n6968 a_400_38200# 0.07fF
C14091 VP.n6969 a_400_38200# 0.19fF
C14092 VP.n6970 a_400_38200# 0.59fF
C14093 VP.n6971 a_400_38200# 0.34fF
C14094 VP.n6972 a_400_38200# 2.04fF
C14095 VP.t551 a_400_38200# 0.02fF
C14096 VP.n6973 a_400_38200# 0.24fF
C14097 VP.n6974 a_400_38200# 0.91fF
C14098 VP.n6975 a_400_38200# 0.05fF
C14099 VP.t600 a_400_38200# 0.02fF
C14100 VP.n6976 a_400_38200# 0.12fF
C14101 VP.n6977 a_400_38200# 0.14fF
C14102 VP.n6979 a_400_38200# 0.06fF
C14103 VP.n6980 a_400_38200# 0.09fF
C14104 VP.n6981 a_400_38200# 0.09fF
C14105 VP.n6982 a_400_38200# 1.45fF
C14106 VP.n6983 a_400_38200# 0.14fF
C14107 VP.n6984 a_400_38200# 0.07fF
C14108 VP.n6985 a_400_38200# 0.72fF
C14109 VP.n6986 a_400_38200# 1.81fF
C14110 VP.n6987 a_400_38200# 0.12fF
C14111 VP.t1099 a_400_38200# 0.02fF
C14112 VP.n6988 a_400_38200# 0.14fF
C14113 VP.t388 a_400_38200# 0.02fF
C14114 VP.n6990 a_400_38200# 0.24fF
C14115 VP.n6991 a_400_38200# 0.35fF
C14116 VP.n6992 a_400_38200# 0.60fF
C14117 VP.n6993 a_400_38200# 2.30fF
C14118 VP.t79 a_400_38200# 0.02fF
C14119 VP.n6994 a_400_38200# 0.24fF
C14120 VP.n6995 a_400_38200# 0.91fF
C14121 VP.n6996 a_400_38200# 0.05fF
C14122 VP.t215 a_400_38200# 0.02fF
C14123 VP.n6997 a_400_38200# 0.12fF
C14124 VP.n6998 a_400_38200# 0.14fF
C14125 VP.n7000 a_400_38200# 1.93fF
C14126 VP.n7001 a_400_38200# 2.23fF
C14127 VP.t1245 a_400_38200# 0.02fF
C14128 VP.n7002 a_400_38200# 0.24fF
C14129 VP.n7003 a_400_38200# 0.35fF
C14130 VP.n7004 a_400_38200# 0.60fF
C14131 VP.n7005 a_400_38200# 0.12fF
C14132 VP.t657 a_400_38200# 0.02fF
C14133 VP.n7006 a_400_38200# 0.14fF
C14134 VP.n7008 a_400_38200# 0.07fF
C14135 VP.n7009 a_400_38200# 0.30fF
C14136 VP.n7010 a_400_38200# 0.06fF
C14137 VP.n7011 a_400_38200# 0.25fF
C14138 VP.n7012 a_400_38200# 0.45fF
C14139 VP.n7013 a_400_38200# 0.06fF
C14140 VP.n7014 a_400_38200# 0.06fF
C14141 VP.n7015 a_400_38200# 0.03fF
C14142 VP.n7016 a_400_38200# 0.05fF
C14143 VP.n7017 a_400_38200# 0.07fF
C14144 VP.n7018 a_400_38200# 0.19fF
C14145 VP.n7019 a_400_38200# 0.59fF
C14146 VP.n7020 a_400_38200# 0.34fF
C14147 VP.n7021 a_400_38200# 2.04fF
C14148 VP.t960 a_400_38200# 0.02fF
C14149 VP.n7022 a_400_38200# 0.24fF
C14150 VP.n7023 a_400_38200# 0.91fF
C14151 VP.n7024 a_400_38200# 0.05fF
C14152 VP.t1069 a_400_38200# 0.02fF
C14153 VP.n7025 a_400_38200# 0.12fF
C14154 VP.n7026 a_400_38200# 0.14fF
C14155 VP.n7028 a_400_38200# 1.81fF
C14156 VP.t799 a_400_38200# 0.02fF
C14157 VP.n7029 a_400_38200# 0.24fF
C14158 VP.n7030 a_400_38200# 0.35fF
C14159 VP.n7031 a_400_38200# 0.60fF
C14160 VP.n7032 a_400_38200# 0.12fF
C14161 VP.t211 a_400_38200# 0.02fF
C14162 VP.n7033 a_400_38200# 0.14fF
C14163 VP.n7035 a_400_38200# 0.03fF
C14164 VP.n7036 a_400_38200# 0.09fF
C14165 VP.n7037 a_400_38200# 0.09fF
C14166 VP.n7038 a_400_38200# 0.05fF
C14167 VP.n7039 a_400_38200# 0.11fF
C14168 VP.n7040 a_400_38200# 0.09fF
C14169 VP.n7041 a_400_38200# 0.02fF
C14170 VP.n7042 a_400_38200# 0.03fF
C14171 VP.n7043 a_400_38200# 0.11fF
C14172 VP.n7044 a_400_38200# 1.39fF
C14173 VP.n7045 a_400_38200# 0.06fF
C14174 VP.n7046 a_400_38200# 0.37fF
C14175 VP.n7047 a_400_38200# 2.30fF
C14176 VP.t513 a_400_38200# 0.02fF
C14177 VP.n7048 a_400_38200# 0.24fF
C14178 VP.n7049 a_400_38200# 0.91fF
C14179 VP.n7050 a_400_38200# 0.05fF
C14180 VP.t625 a_400_38200# 0.02fF
C14181 VP.n7051 a_400_38200# 0.12fF
C14182 VP.n7052 a_400_38200# 0.14fF
C14183 VP.n7054 a_400_38200# 0.88fF
C14184 VP.n7055 a_400_38200# 0.48fF
C14185 VP.n7056 a_400_38200# 0.88fF
C14186 VP.n7057 a_400_38200# 0.60fF
C14187 VP.n7058 a_400_38200# 2.33fF
C14188 VP.n7059 a_400_38200# 0.59fF
C14189 VP.n7060 a_400_38200# 0.02fF
C14190 VP.n7061 a_400_38200# 0.96fF
C14191 VP.t136 a_400_38200# 15.72fF
C14192 VP.n7062 a_400_38200# 15.42fF
C14193 VP.n7064 a_400_38200# 0.38fF
C14194 VP.n7065 a_400_38200# 0.23fF
C14195 VP.n7066 a_400_38200# 3.42fF
C14196 VP.n7067 a_400_38200# 0.21fF
C14197 VP.n7068 a_400_38200# 1.08fF
C14198 VP.n7069 a_400_38200# 0.03fF
C14199 VP.n7070 a_400_38200# 0.09fF
C14200 VP.n7071 a_400_38200# 0.43fF
C14201 VP.n7072 a_400_38200# 0.37fF
C14202 VP.t1043 a_400_38200# 0.02fF
C14203 VP.n7073 a_400_38200# 0.64fF
C14204 VP.n7074 a_400_38200# 0.60fF
C14205 VP.n7075 a_400_38200# 2.32fF
C14206 VP.n7076 a_400_38200# 4.93fF
C14207 VP.t763 a_400_38200# 0.02fF
C14208 VP.n7077 a_400_38200# 1.19fF
C14209 VP.n7078 a_400_38200# 0.05fF
C14210 VP.t865 a_400_38200# 0.02fF
C14211 VP.n7079 a_400_38200# 0.01fF
C14212 VP.n7080 a_400_38200# 0.26fF
C14213 VP.n7082 a_400_38200# 15.28fF
C14214 VP.n7083 a_400_38200# 0.10fF
C14215 VP.n7084 a_400_38200# 0.28fF
C14216 VP.n7085 a_400_38200# 0.15fF
C14217 VP.n7086 a_400_38200# 0.08fF
C14218 VP.n7087 a_400_38200# 0.14fF
C14219 VP.n7088 a_400_38200# 0.06fF
C14220 VP.n7089 a_400_38200# 0.06fF
C14221 VP.n7090 a_400_38200# 0.03fF
C14222 VP.n7091 a_400_38200# 0.05fF
C14223 VP.n7092 a_400_38200# 0.07fF
C14224 VP.n7093 a_400_38200# 0.19fF
C14225 VP.n7094 a_400_38200# 0.59fF
C14226 VP.n7095 a_400_38200# 0.34fF
C14227 VP.n7096 a_400_38200# 0.04fF
C14228 VP.n7097 a_400_38200# 0.02fF
C14229 VP.n7098 a_400_38200# 0.06fF
C14230 VP.n7099 a_400_38200# 0.30fF
C14231 VP.n7100 a_400_38200# 1.93fF
C14232 VP.n7101 a_400_38200# 0.12fF
C14233 VP.t1324 a_400_38200# 0.02fF
C14234 VP.n7102 a_400_38200# 0.14fF
C14235 VP.t613 a_400_38200# 0.02fF
C14236 VP.n7104 a_400_38200# 0.24fF
C14237 VP.n7105 a_400_38200# 0.35fF
C14238 VP.n7106 a_400_38200# 0.60fF
C14239 VP.n7107 a_400_38200# 2.47fF
C14240 VP.n7108 a_400_38200# 2.20fF
C14241 VP.t432 a_400_38200# 0.02fF
C14242 VP.n7109 a_400_38200# 0.12fF
C14243 VP.n7110 a_400_38200# 0.14fF
C14244 VP.t333 a_400_38200# 0.02fF
C14245 VP.n7112 a_400_38200# 0.24fF
C14246 VP.n7113 a_400_38200# 0.91fF
C14247 VP.n7114 a_400_38200# 0.05fF
C14248 VP.n7115 a_400_38200# 0.10fF
C14249 VP.n7116 a_400_38200# 0.28fF
C14250 VP.n7117 a_400_38200# 0.15fF
C14251 VP.n7118 a_400_38200# 0.08fF
C14252 VP.n7119 a_400_38200# 0.14fF
C14253 VP.n7120 a_400_38200# 0.06fF
C14254 VP.n7121 a_400_38200# 0.06fF
C14255 VP.n7122 a_400_38200# 0.03fF
C14256 VP.n7123 a_400_38200# 0.05fF
C14257 VP.n7124 a_400_38200# 0.07fF
C14258 VP.n7125 a_400_38200# 0.19fF
C14259 VP.n7126 a_400_38200# 0.59fF
C14260 VP.n7127 a_400_38200# 0.34fF
C14261 VP.n7128 a_400_38200# 0.04fF
C14262 VP.n7129 a_400_38200# 0.02fF
C14263 VP.n7130 a_400_38200# 0.06fF
C14264 VP.n7131 a_400_38200# 0.30fF
C14265 VP.n7132 a_400_38200# 1.93fF
C14266 VP.n7133 a_400_38200# 0.12fF
C14267 VP.t873 a_400_38200# 0.02fF
C14268 VP.n7134 a_400_38200# 0.14fF
C14269 VP.t150 a_400_38200# 0.02fF
C14270 VP.n7136 a_400_38200# 0.24fF
C14271 VP.n7137 a_400_38200# 0.35fF
C14272 VP.n7138 a_400_38200# 0.60fF
C14273 VP.n7139 a_400_38200# 2.39fF
C14274 VP.n7140 a_400_38200# 1.79fF
C14275 VP.t1287 a_400_38200# 0.02fF
C14276 VP.n7141 a_400_38200# 0.12fF
C14277 VP.n7142 a_400_38200# 0.14fF
C14278 VP.t1178 a_400_38200# 0.02fF
C14279 VP.n7144 a_400_38200# 0.24fF
C14280 VP.n7145 a_400_38200# 0.91fF
C14281 VP.n7146 a_400_38200# 0.05fF
C14282 VP.t195 a_400_38200# 34.79fF
C14283 VP.t881 a_400_38200# 0.02fF
C14284 VP.n7147 a_400_38200# 0.12fF
C14285 VP.n7148 a_400_38200# 0.14fF
C14286 VP.t782 a_400_38200# 0.02fF
C14287 VP.n7150 a_400_38200# 0.24fF
C14288 VP.n7151 a_400_38200# 0.91fF
C14289 VP.n7152 a_400_38200# 0.05fF
C14290 VP.t1061 a_400_38200# 0.02fF
C14291 VP.n7153 a_400_38200# 0.24fF
C14292 VP.n7154 a_400_38200# 0.35fF
C14293 VP.n7155 a_400_38200# 0.60fF
C14294 VP.n7156 a_400_38200# 0.04fF
C14295 VP.n7157 a_400_38200# 0.08fF
C14296 VP.n7158 a_400_38200# 0.72fF
C14297 VP.n7159 a_400_38200# 0.09fF
C14298 VP.n7160 a_400_38200# 0.00fF
C14299 VP.n7161 a_400_38200# 1.22fF
C14300 VP.n7162 a_400_38200# 0.19fF
C14301 VP.n7164 a_400_38200# 1.72fF
C14302 VP.n7165 a_400_38200# 1.96fF
C14303 VP.n7166 a_400_38200# 1.04fF
C14304 VP.n7167 a_400_38200# 0.05fF
C14305 VP.n7168 a_400_38200# 0.03fF
C14306 VP.n7169 a_400_38200# 0.06fF
C14307 VP.n7170 a_400_38200# 0.06fF
C14308 VP.n7171 a_400_38200# 0.06fF
C14309 VP.n7172 a_400_38200# 0.07fF
C14310 VP.n7173 a_400_38200# 0.03fF
C14311 VP.n7174 a_400_38200# 0.05fF
C14312 VP.n7175 a_400_38200# 0.07fF
C14313 VP.n7176 a_400_38200# 0.19fF
C14314 VP.n7177 a_400_38200# 0.60fF
C14315 VP.n7178 a_400_38200# 0.76fF
C14316 VP.n7179 a_400_38200# 0.40fF
C14317 VP.n7180 a_400_38200# 0.03fF
C14318 VP.n7181 a_400_38200# 0.01fF
C14319 VP.t603 a_400_38200# 0.02fF
C14320 VP.n7182 a_400_38200# 0.25fF
C14321 VP.t318 a_400_38200# 0.02fF
C14322 VP.n7183 a_400_38200# 0.95fF
C14323 VP.n7184 a_400_38200# 0.70fF
C14324 VP.n7185 a_400_38200# 1.93fF
C14325 VP.n7186 a_400_38200# 2.97fF
C14326 VP.n7187 a_400_38200# 2.27fF
C14327 VP.t535 a_400_38200# 0.02fF
C14328 VP.n7188 a_400_38200# 0.24fF
C14329 VP.n7189 a_400_38200# 0.35fF
C14330 VP.n7190 a_400_38200# 0.60fF
C14331 VP.n7191 a_400_38200# 0.12fF
C14332 VP.t1254 a_400_38200# 0.02fF
C14333 VP.n7192 a_400_38200# 0.14fF
C14334 VP.n7194 a_400_38200# 0.04fF
C14335 VP.n7195 a_400_38200# 0.02fF
C14336 VP.n7196 a_400_38200# 0.06fF
C14337 VP.n7197 a_400_38200# 0.30fF
C14338 VP.n7198 a_400_38200# 0.10fF
C14339 VP.n7199 a_400_38200# 0.28fF
C14340 VP.n7200 a_400_38200# 0.06fF
C14341 VP.n7201 a_400_38200# 0.06fF
C14342 VP.n7202 a_400_38200# 0.03fF
C14343 VP.n7203 a_400_38200# 0.15fF
C14344 VP.n7204 a_400_38200# 0.08fF
C14345 VP.n7205 a_400_38200# 0.14fF
C14346 VP.n7206 a_400_38200# 0.03fF
C14347 VP.n7207 a_400_38200# 0.06fF
C14348 VP.n7208 a_400_38200# 0.06fF
C14349 VP.n7209 a_400_38200# 0.06fF
C14350 VP.n7210 a_400_38200# 0.06fF
C14351 VP.n7211 a_400_38200# 0.03fF
C14352 VP.n7212 a_400_38200# 0.05fF
C14353 VP.n7213 a_400_38200# 0.07fF
C14354 VP.n7214 a_400_38200# 0.19fF
C14355 VP.n7215 a_400_38200# 0.59fF
C14356 VP.n7216 a_400_38200# 0.34fF
C14357 VP.n7217 a_400_38200# 1.88fF
C14358 VP.t968 a_400_38200# 0.02fF
C14359 VP.n7218 a_400_38200# 0.24fF
C14360 VP.n7219 a_400_38200# 0.91fF
C14361 VP.n7220 a_400_38200# 0.05fF
C14362 VP.t591 a_400_38200# 0.02fF
C14363 VP.n7221 a_400_38200# 0.12fF
C14364 VP.n7222 a_400_38200# 0.14fF
C14365 VP.n7224 a_400_38200# 0.19fF
C14366 VP.n7225 a_400_38200# 0.10fF
C14367 VP.n7226 a_400_38200# 0.10fF
C14368 VP.n7227 a_400_38200# 0.18fF
C14369 VP.n7228 a_400_38200# 0.09fF
C14370 VP.n7229 a_400_38200# 0.04fF
C14371 VP.n7230 a_400_38200# 0.19fF
C14372 VP.n7231 a_400_38200# 0.26fF
C14373 VP.n7232 a_400_38200# 1.17fF
C14374 VP.n7233 a_400_38200# 0.06fF
C14375 VP.n7234 a_400_38200# 0.44fF
C14376 VP.n7235 a_400_38200# 0.13fF
C14377 VP.n7236 a_400_38200# 0.02fF
C14378 VP.n7237 a_400_38200# 1.81fF
C14379 VP.n7238 a_400_38200# 0.12fF
C14380 VP.t810 a_400_38200# 0.02fF
C14381 VP.n7239 a_400_38200# 0.14fF
C14382 VP.t59 a_400_38200# 0.02fF
C14383 VP.n7241 a_400_38200# 0.24fF
C14384 VP.n7242 a_400_38200# 0.35fF
C14385 VP.n7243 a_400_38200# 0.60fF
C14386 VP.n7244 a_400_38200# 3.18fF
C14387 VP.n7245 a_400_38200# 2.06fF
C14388 VP.n7246 a_400_38200# 1.98fF
C14389 VP.t520 a_400_38200# 0.02fF
C14390 VP.n7247 a_400_38200# 0.24fF
C14391 VP.n7248 a_400_38200# 0.91fF
C14392 VP.n7249 a_400_38200# 0.05fF
C14393 VP.t909 a_400_38200# 0.02fF
C14394 VP.n7250 a_400_38200# 0.12fF
C14395 VP.n7251 a_400_38200# 0.14fF
C14396 VP.n7253 a_400_38200# 0.16fF
C14397 VP.n7254 a_400_38200# 0.19fF
C14398 VP.n7255 a_400_38200# 0.09fF
C14399 VP.n7256 a_400_38200# 0.04fF
C14400 VP.n7257 a_400_38200# 0.14fF
C14401 VP.n7258 a_400_38200# 0.64fF
C14402 VP.n7259 a_400_38200# 1.32fF
C14403 VP.n7260 a_400_38200# 1.81fF
C14404 VP.n7261 a_400_38200# 0.12fF
C14405 VP.t361 a_400_38200# 0.02fF
C14406 VP.n7262 a_400_38200# 0.14fF
C14407 VP.t944 a_400_38200# 0.02fF
C14408 VP.n7264 a_400_38200# 0.24fF
C14409 VP.n7265 a_400_38200# 0.35fF
C14410 VP.n7266 a_400_38200# 0.60fF
C14411 VP.n7267 a_400_38200# 2.97fF
C14412 VP.n7268 a_400_38200# 2.27fF
C14413 VP.n7269 a_400_38200# 2.00fF
C14414 VP.t40 a_400_38200# 0.02fF
C14415 VP.n7270 a_400_38200# 0.24fF
C14416 VP.n7271 a_400_38200# 0.91fF
C14417 VP.n7272 a_400_38200# 0.05fF
C14418 VP.t459 a_400_38200# 0.02fF
C14419 VP.n7273 a_400_38200# 0.12fF
C14420 VP.n7274 a_400_38200# 0.14fF
C14421 VP.n7276 a_400_38200# 0.24fF
C14422 VP.t485 a_400_38200# 0.02fF
C14423 VP.n7277 a_400_38200# 0.36fF
C14424 VP.n7278 a_400_38200# 0.36fF
C14425 VP.n7279 a_400_38200# 0.67fF
C14426 VP.n7280 a_400_38200# 0.16fF
C14427 VP.n7281 a_400_38200# 0.19fF
C14428 VP.n7282 a_400_38200# 0.09fF
C14429 VP.n7283 a_400_38200# 0.04fF
C14430 VP.n7284 a_400_38200# 0.14fF
C14431 VP.n7285 a_400_38200# 0.64fF
C14432 VP.n7286 a_400_38200# 1.32fF
C14433 VP.n7287 a_400_38200# 1.81fF
C14434 VP.n7288 a_400_38200# 2.97fF
C14435 VP.n7289 a_400_38200# 2.27fF
C14436 VP.n7290 a_400_38200# 0.75fF
C14437 VP.n7291 a_400_38200# 0.24fF
C14438 VP.t3 a_400_38200# 0.02fF
C14439 VP.n7292 a_400_38200# 0.35fF
C14440 VP.n7293 a_400_38200# 0.63fF
C14441 VP.n7294 a_400_38200# 0.40fF
C14442 VP.n7295 a_400_38200# 0.40fF
C14443 VP.n7296 a_400_38200# 0.12fF
C14444 VP.t767 a_400_38200# 0.02fF
C14445 VP.n7297 a_400_38200# 0.14fF
C14446 VP.t861 a_400_38200# 0.02fF
C14447 VP.n7299 a_400_38200# 0.12fF
C14448 VP.n7300 a_400_38200# 0.14fF
C14449 VP.n7302 a_400_38200# 0.16fF
C14450 VP.n7303 a_400_38200# 0.19fF
C14451 VP.n7304 a_400_38200# 0.09fF
C14452 VP.n7305 a_400_38200# 0.04fF
C14453 VP.n7306 a_400_38200# 0.14fF
C14454 VP.n7307 a_400_38200# 0.64fF
C14455 VP.n7308 a_400_38200# 1.32fF
C14456 VP.n7309 a_400_38200# 1.81fF
C14457 VP.n7310 a_400_38200# 0.12fF
C14458 VP.t1236 a_400_38200# 0.02fF
C14459 VP.n7311 a_400_38200# 0.14fF
C14460 VP.t455 a_400_38200# 0.02fF
C14461 VP.n7313 a_400_38200# 0.24fF
C14462 VP.n7314 a_400_38200# 0.35fF
C14463 VP.n7315 a_400_38200# 0.60fF
C14464 VP.n7316 a_400_38200# 2.97fF
C14465 VP.n7317 a_400_38200# 2.27fF
C14466 VP.n7318 a_400_38200# 2.00fF
C14467 VP.t882 a_400_38200# 0.02fF
C14468 VP.n7319 a_400_38200# 0.24fF
C14469 VP.n7320 a_400_38200# 0.91fF
C14470 VP.n7321 a_400_38200# 0.05fF
C14471 VP.t1270 a_400_38200# 0.02fF
C14472 VP.n7322 a_400_38200# 0.12fF
C14473 VP.n7323 a_400_38200# 0.14fF
C14474 VP.n7325 a_400_38200# 0.03fF
C14475 VP.n7326 a_400_38200# 0.19fF
C14476 VP.n7327 a_400_38200# 0.24fF
C14477 VP.n7328 a_400_38200# 0.98fF
C14478 VP.n7329 a_400_38200# 0.12fF
C14479 VP.n7330 a_400_38200# 0.19fF
C14480 VP.n7331 a_400_38200# 0.09fF
C14481 VP.n7332 a_400_38200# 0.18fF
C14482 VP.n7333 a_400_38200# 0.09fF
C14483 VP.n7334 a_400_38200# 0.08fF
C14484 VP.n7335 a_400_38200# 0.39fF
C14485 VP.n7336 a_400_38200# 0.24fF
C14486 VP.n7337 a_400_38200# 0.13fF
C14487 VP.n7338 a_400_38200# 0.02fF
C14488 VP.n7339 a_400_38200# 1.81fF
C14489 VP.n7340 a_400_38200# 0.12fF
C14490 VP.t345 a_400_38200# 0.02fF
C14491 VP.n7341 a_400_38200# 0.14fF
C14492 VP.t928 a_400_38200# 0.02fF
C14493 VP.n7343 a_400_38200# 0.24fF
C14494 VP.n7344 a_400_38200# 0.35fF
C14495 VP.n7345 a_400_38200# 0.60fF
C14496 VP.n7346 a_400_38200# 3.17fF
C14497 VP.n7347 a_400_38200# 2.27fF
C14498 VP.n7348 a_400_38200# 1.98fF
C14499 VP.t11 a_400_38200# 0.02fF
C14500 VP.n7349 a_400_38200# 0.24fF
C14501 VP.n7350 a_400_38200# 0.91fF
C14502 VP.n7351 a_400_38200# 0.05fF
C14503 VP.t374 a_400_38200# 0.02fF
C14504 VP.n7352 a_400_38200# 0.12fF
C14505 VP.n7353 a_400_38200# 0.14fF
C14506 VP.n7355 a_400_38200# 15.28fF
C14507 VP.n7356 a_400_38200# 0.10fF
C14508 VP.n7357 a_400_38200# 0.06fF
C14509 VP.n7358 a_400_38200# 0.06fF
C14510 VP.n7359 a_400_38200# 0.28fF
C14511 VP.n7360 a_400_38200# 0.03fF
C14512 VP.n7361 a_400_38200# 0.15fF
C14513 VP.n7362 a_400_38200# 0.08fF
C14514 VP.n7363 a_400_38200# 0.14fF
C14515 VP.n7364 a_400_38200# 0.03fF
C14516 VP.n7365 a_400_38200# 0.06fF
C14517 VP.n7366 a_400_38200# 0.06fF
C14518 VP.n7367 a_400_38200# 0.06fF
C14519 VP.n7368 a_400_38200# 0.06fF
C14520 VP.n7369 a_400_38200# 0.03fF
C14521 VP.n7370 a_400_38200# 0.05fF
C14522 VP.n7371 a_400_38200# 0.07fF
C14523 VP.n7372 a_400_38200# 0.19fF
C14524 VP.n7373 a_400_38200# 0.59fF
C14525 VP.n7374 a_400_38200# 0.34fF
C14526 VP.n7375 a_400_38200# 0.04fF
C14527 VP.n7376 a_400_38200# 0.02fF
C14528 VP.n7377 a_400_38200# 0.06fF
C14529 VP.n7378 a_400_38200# 0.30fF
C14530 VP.n7379 a_400_38200# 1.93fF
C14531 VP.n7380 a_400_38200# 0.12fF
C14532 VP.t135 a_400_38200# 0.02fF
C14533 VP.n7381 a_400_38200# 0.14fF
C14534 VP.t735 a_400_38200# 0.02fF
C14535 VP.n7383 a_400_38200# 0.24fF
C14536 VP.n7384 a_400_38200# 0.35fF
C14537 VP.n7385 a_400_38200# 0.60fF
C14538 VP.n7386 a_400_38200# 0.56fF
C14539 VP.n7387 a_400_38200# 1.24fF
C14540 VP.n7388 a_400_38200# 0.54fF
C14541 VP.n7389 a_400_38200# 0.22fF
C14542 VP.n7390 a_400_38200# 1.73fF
C14543 VP.t190 a_400_38200# 0.02fF
C14544 VP.n7391 a_400_38200# 0.12fF
C14545 VP.n7392 a_400_38200# 0.14fF
C14546 VP.t1161 a_400_38200# 0.02fF
C14547 VP.n7394 a_400_38200# 0.24fF
C14548 VP.n7395 a_400_38200# 0.91fF
C14549 VP.n7396 a_400_38200# 0.05fF
C14550 VP.n7397 a_400_38200# 0.10fF
C14551 VP.n7398 a_400_38200# 0.28fF
C14552 VP.n7399 a_400_38200# 0.06fF
C14553 VP.n7400 a_400_38200# 0.06fF
C14554 VP.n7401 a_400_38200# 0.03fF
C14555 VP.n7402 a_400_38200# 0.15fF
C14556 VP.n7403 a_400_38200# 0.08fF
C14557 VP.n7404 a_400_38200# 0.14fF
C14558 VP.n7405 a_400_38200# 0.03fF
C14559 VP.n7406 a_400_38200# 0.06fF
C14560 VP.n7407 a_400_38200# 0.06fF
C14561 VP.n7408 a_400_38200# 0.06fF
C14562 VP.n7409 a_400_38200# 0.06fF
C14563 VP.n7410 a_400_38200# 0.03fF
C14564 VP.n7411 a_400_38200# 0.05fF
C14565 VP.n7412 a_400_38200# 0.07fF
C14566 VP.n7413 a_400_38200# 0.19fF
C14567 VP.n7414 a_400_38200# 0.59fF
C14568 VP.n7415 a_400_38200# 0.34fF
C14569 VP.n7416 a_400_38200# 0.04fF
C14570 VP.n7417 a_400_38200# 0.02fF
C14571 VP.n7418 a_400_38200# 0.06fF
C14572 VP.n7419 a_400_38200# 0.30fF
C14573 VP.n7420 a_400_38200# 1.93fF
C14574 VP.n7421 a_400_38200# 0.12fF
C14575 VP.t1000 a_400_38200# 0.02fF
C14576 VP.n7422 a_400_38200# 0.14fF
C14577 VP.t283 a_400_38200# 0.02fF
C14578 VP.n7424 a_400_38200# 0.24fF
C14579 VP.n7425 a_400_38200# 0.35fF
C14580 VP.n7426 a_400_38200# 0.60fF
C14581 VP.n7427 a_400_38200# 0.71fF
C14582 VP.n7428 a_400_38200# 1.39fF
C14583 VP.n7429 a_400_38200# 0.54fF
C14584 VP.n7430 a_400_38200# 0.21fF
C14585 VP.n7431 a_400_38200# 1.73fF
C14586 VP.t1042 a_400_38200# 0.02fF
C14587 VP.n7432 a_400_38200# 0.12fF
C14588 VP.n7433 a_400_38200# 0.14fF
C14589 VP.t712 a_400_38200# 0.02fF
C14590 VP.n7435 a_400_38200# 0.24fF
C14591 VP.n7436 a_400_38200# 0.91fF
C14592 VP.n7437 a_400_38200# 0.05fF
C14593 VP.n7438 a_400_38200# 0.06fF
C14594 VP.n7439 a_400_38200# 0.06fF
C14595 VP.n7440 a_400_38200# 0.03fF
C14596 VP.n7441 a_400_38200# 0.10fF
C14597 VP.n7442 a_400_38200# 0.17fF
C14598 VP.n7443 a_400_38200# 0.10fF
C14599 VP.n7444 a_400_38200# 0.13fF
C14600 VP.n7445 a_400_38200# 0.02fF
C14601 VP.n7446 a_400_38200# 0.04fF
C14602 VP.n7447 a_400_38200# 0.06fF
C14603 VP.n7448 a_400_38200# 0.09fF
C14604 VP.n7449 a_400_38200# 0.10fF
C14605 VP.n7450 a_400_38200# 0.05fF
C14606 VP.n7451 a_400_38200# 0.19fF
C14607 VP.n7452 a_400_38200# 0.16fF
C14608 VP.n7453 a_400_38200# 0.04fF
C14609 VP.n7454 a_400_38200# 0.05fF
C14610 VP.n7455 a_400_38200# 0.04fF
C14611 VP.n7456 a_400_38200# 0.12fF
C14612 VP.n7457 a_400_38200# 0.09fF
C14613 VP.n7458 a_400_38200# 0.14fF
C14614 VP.n7459 a_400_38200# 0.56fF
C14615 VP.n7460 a_400_38200# 0.10fF
C14616 VP.n7461 a_400_38200# 1.93fF
C14617 VP.n7462 a_400_38200# 0.12fF
C14618 VP.t1214 a_400_38200# 0.02fF
C14619 VP.n7463 a_400_38200# 0.14fF
C14620 VP.t499 a_400_38200# 0.02fF
C14621 VP.n7465 a_400_38200# 0.24fF
C14622 VP.n7466 a_400_38200# 0.35fF
C14623 VP.n7467 a_400_38200# 0.60fF
C14624 VP.n7468 a_400_38200# 0.18fF
C14625 VP.n7469 a_400_38200# 0.45fF
C14626 VP.n7470 a_400_38200# 0.06fF
C14627 VP.n7471 a_400_38200# 0.01fF
C14628 VP.n7472 a_400_38200# 0.01fF
C14629 VP.n7473 a_400_38200# 0.04fF
C14630 VP.n7474 a_400_38200# 0.02fF
C14631 VP.n7475 a_400_38200# 0.07fF
C14632 VP.n7476 a_400_38200# 0.04fF
C14633 VP.n7477 a_400_38200# 0.14fF
C14634 VP.n7478 a_400_38200# 0.45fF
C14635 VP.n7479 a_400_38200# 1.46fF
C14636 VP.n7480 a_400_38200# 1.78fF
C14637 VP.t1308 a_400_38200# 0.02fF
C14638 VP.n7481 a_400_38200# 0.12fF
C14639 VP.n7482 a_400_38200# 0.14fF
C14640 VP.t930 a_400_38200# 0.02fF
C14641 VP.n7484 a_400_38200# 0.24fF
C14642 VP.n7485 a_400_38200# 0.91fF
C14643 VP.n7486 a_400_38200# 0.05fF
C14644 VP.n7487 a_400_38200# 1.93fF
C14645 VP.n7488 a_400_38200# 0.18fF
C14646 VP.n7489 a_400_38200# 0.45fF
C14647 VP.n7490 a_400_38200# 0.06fF
C14648 VP.n7491 a_400_38200# 0.01fF
C14649 VP.n7492 a_400_38200# 0.01fF
C14650 VP.n7493 a_400_38200# 0.04fF
C14651 VP.n7494 a_400_38200# 0.02fF
C14652 VP.n7495 a_400_38200# 0.07fF
C14653 VP.n7496 a_400_38200# 0.04fF
C14654 VP.n7497 a_400_38200# 0.14fF
C14655 VP.n7498 a_400_38200# 0.45fF
C14656 VP.n7499 a_400_38200# 1.46fF
C14657 VP.t906 a_400_38200# 0.02fF
C14658 VP.n7500 a_400_38200# 0.24fF
C14659 VP.n7501 a_400_38200# 0.35fF
C14660 VP.n7502 a_400_38200# 0.60fF
C14661 VP.n7503 a_400_38200# 0.12fF
C14662 VP.t314 a_400_38200# 0.02fF
C14663 VP.n7504 a_400_38200# 0.14fF
C14664 VP.n7506 a_400_38200# 0.10fF
C14665 VP.n7507 a_400_38200# 0.17fF
C14666 VP.n7508 a_400_38200# 0.06fF
C14667 VP.n7509 a_400_38200# 0.06fF
C14668 VP.n7510 a_400_38200# 0.03fF
C14669 VP.n7511 a_400_38200# 0.10fF
C14670 VP.n7512 a_400_38200# 0.13fF
C14671 VP.n7513 a_400_38200# 0.13fF
C14672 VP.n7514 a_400_38200# 0.04fF
C14673 VP.n7515 a_400_38200# 0.05fF
C14674 VP.n7516 a_400_38200# 0.04fF
C14675 VP.n7517 a_400_38200# 0.09fF
C14676 VP.n7518 a_400_38200# 0.09fF
C14677 VP.n7519 a_400_38200# 0.05fF
C14678 VP.n7520 a_400_38200# 0.19fF
C14679 VP.n7521 a_400_38200# 0.12fF
C14680 VP.n7522 a_400_38200# 0.09fF
C14681 VP.n7523 a_400_38200# 0.14fF
C14682 VP.n7524 a_400_38200# 0.04fF
C14683 VP.n7525 a_400_38200# 0.02fF
C14684 VP.n7526 a_400_38200# 0.06fF
C14685 VP.n7527 a_400_38200# 0.56fF
C14686 VP.n7528 a_400_38200# 0.10fF
C14687 VP.n7529 a_400_38200# 1.78fF
C14688 VP.t414 a_400_38200# 0.02fF
C14689 VP.n7530 a_400_38200# 0.12fF
C14690 VP.n7531 a_400_38200# 0.14fF
C14691 VP.t1333 a_400_38200# 0.02fF
C14692 VP.n7533 a_400_38200# 0.24fF
C14693 VP.n7534 a_400_38200# 0.91fF
C14694 VP.n7535 a_400_38200# 0.05fF
C14695 VP.n7536 a_400_38200# 1.93fF
C14696 VP.n7537 a_400_38200# 0.18fF
C14697 VP.n7538 a_400_38200# 0.45fF
C14698 VP.n7539 a_400_38200# 0.06fF
C14699 VP.n7540 a_400_38200# 0.01fF
C14700 VP.n7541 a_400_38200# 0.01fF
C14701 VP.n7542 a_400_38200# 0.04fF
C14702 VP.n7543 a_400_38200# 0.02fF
C14703 VP.n7544 a_400_38200# 0.07fF
C14704 VP.n7545 a_400_38200# 0.04fF
C14705 VP.n7546 a_400_38200# 0.14fF
C14706 VP.n7547 a_400_38200# 0.45fF
C14707 VP.n7548 a_400_38200# 1.46fF
C14708 VP.t37 a_400_38200# 0.02fF
C14709 VP.n7549 a_400_38200# 0.24fF
C14710 VP.n7550 a_400_38200# 0.35fF
C14711 VP.n7551 a_400_38200# 0.60fF
C14712 VP.n7552 a_400_38200# 0.12fF
C14713 VP.t791 a_400_38200# 0.02fF
C14714 VP.n7553 a_400_38200# 0.14fF
C14715 VP.n7555 a_400_38200# 0.10fF
C14716 VP.n7556 a_400_38200# 0.17fF
C14717 VP.n7557 a_400_38200# 0.06fF
C14718 VP.n7558 a_400_38200# 0.06fF
C14719 VP.n7559 a_400_38200# 0.03fF
C14720 VP.n7560 a_400_38200# 0.10fF
C14721 VP.n7561 a_400_38200# 0.13fF
C14722 VP.n7562 a_400_38200# 0.13fF
C14723 VP.n7563 a_400_38200# 0.04fF
C14724 VP.n7564 a_400_38200# 0.05fF
C14725 VP.n7565 a_400_38200# 0.04fF
C14726 VP.n7566 a_400_38200# 0.09fF
C14727 VP.n7567 a_400_38200# 0.09fF
C14728 VP.n7568 a_400_38200# 0.05fF
C14729 VP.n7569 a_400_38200# 0.19fF
C14730 VP.n7570 a_400_38200# 0.12fF
C14731 VP.n7571 a_400_38200# 0.09fF
C14732 VP.n7572 a_400_38200# 0.14fF
C14733 VP.n7573 a_400_38200# 0.04fF
C14734 VP.n7574 a_400_38200# 0.02fF
C14735 VP.n7575 a_400_38200# 0.06fF
C14736 VP.n7576 a_400_38200# 0.56fF
C14737 VP.n7577 a_400_38200# 0.10fF
C14738 VP.n7578 a_400_38200# 1.78fF
C14739 VP.t824 a_400_38200# 0.02fF
C14740 VP.n7579 a_400_38200# 0.12fF
C14741 VP.n7580 a_400_38200# 0.14fF
C14742 VP.t502 a_400_38200# 0.02fF
C14743 VP.n7582 a_400_38200# 0.24fF
C14744 VP.n7583 a_400_38200# 0.91fF
C14745 VP.n7584 a_400_38200# 0.05fF
C14746 VP.n7585 a_400_38200# 1.92fF
C14747 VP.n7586 a_400_38200# 2.51fF
C14748 VP.t1165 a_400_38200# 0.02fF
C14749 VP.n7587 a_400_38200# 0.24fF
C14750 VP.n7588 a_400_38200# 0.35fF
C14751 VP.n7589 a_400_38200# 0.60fF
C14752 VP.n7590 a_400_38200# 0.12fF
C14753 VP.t581 a_400_38200# 0.02fF
C14754 VP.n7591 a_400_38200# 0.14fF
C14755 VP.n7593 a_400_38200# 0.06fF
C14756 VP.n7594 a_400_38200# 0.30fF
C14757 VP.n7595 a_400_38200# 0.20fF
C14758 VP.n7596 a_400_38200# 0.09fF
C14759 VP.n7597 a_400_38200# 0.26fF
C14760 VP.n7598 a_400_38200# 0.22fF
C14761 VP.n7599 a_400_38200# 0.19fF
C14762 VP.n7600 a_400_38200# 0.05fF
C14763 VP.n7601 a_400_38200# 0.13fF
C14764 VP.n7602 a_400_38200# 0.09fF
C14765 VP.n7603 a_400_38200# 0.09fF
C14766 VP.n7604 a_400_38200# 0.07fF
C14767 VP.n7605 a_400_38200# 0.71fF
C14768 VP.n7606 a_400_38200# 0.24fF
C14769 VP.n7607 a_400_38200# 1.88fF
C14770 VP.t1230 a_400_38200# 0.02fF
C14771 VP.n7608 a_400_38200# 0.12fF
C14772 VP.n7609 a_400_38200# 0.14fF
C14773 VP.t295 a_400_38200# 0.02fF
C14774 VP.n7611 a_400_38200# 0.24fF
C14775 VP.n7612 a_400_38200# 0.91fF
C14776 VP.n7613 a_400_38200# 0.05fF
C14777 VP.t134 a_400_38200# 35.17fF
C14778 VP.t1188 a_400_38200# 0.02fF
C14779 VP.n7614 a_400_38200# 1.21fF
C14780 VP.n7615 a_400_38200# 0.25fF
C14781 VP.n7616 a_400_38200# 26.29fF
C14782 VP.n7617 a_400_38200# 26.29fF
C14783 VP.n7618 a_400_38200# 0.76fF
C14784 VP.n7619 a_400_38200# 0.27fF
C14785 VP.n7620 a_400_38200# 0.59fF
C14786 VP.n7621 a_400_38200# 0.10fF
C14787 VP.n7622 a_400_38200# 3.02fF
C14788 VP.t2 a_400_38200# 15.72fF
C14789 VP.n7623 a_400_38200# 1.15fF
C14790 VP.n7625 a_400_38200# 13.70fF
C14791 VP.n7627 a_400_38200# 1.99fF
C14792 VP.n7628 a_400_38200# 4.39fF
C14793 VP.n7629 a_400_38200# 0.03fF
C14794 VP.n7630 a_400_38200# 0.05fF
C14795 VP.n7631 a_400_38200# 0.07fF
C14796 VP.n7632 a_400_38200# 0.03fF
C14797 VP.n7633 a_400_38200# 0.06fF
C14798 VP.n7634 a_400_38200# 0.06fF
C14799 VP.n7635 a_400_38200# 0.06fF
C14800 VP.n7636 a_400_38200# 0.07fF
C14801 VP.n7637 a_400_38200# 0.57fF
C14802 VP.n7638 a_400_38200# 1.88fF
C14803 VP.n7639 a_400_38200# 0.92fF
C14804 VP.n7640 a_400_38200# 2.63fF
C14805 VP.n7641 a_400_38200# 0.10fF
C14806 VP.n7642 a_400_38200# 0.28fF
C14807 VP.n7643 a_400_38200# 0.15fF
C14808 VP.n7644 a_400_38200# 0.08fF
C14809 VP.n7645 a_400_38200# 0.14fF
C14810 VP.n7646 a_400_38200# 0.06fF
C14811 VP.n7647 a_400_38200# 0.06fF
C14812 VP.n7648 a_400_38200# 0.03fF
C14813 VP.n7649 a_400_38200# 0.05fF
C14814 VP.n7650 a_400_38200# 0.07fF
C14815 VP.n7651 a_400_38200# 0.19fF
C14816 VP.n7652 a_400_38200# 0.59fF
C14817 VP.n7653 a_400_38200# 0.34fF
C14818 VP.n7654 a_400_38200# 0.04fF
C14819 VP.n7655 a_400_38200# 0.02fF
C14820 VP.n7656 a_400_38200# 0.06fF
C14821 VP.n7657 a_400_38200# 0.30fF
C14822 VP.n7658 a_400_38200# 0.12fF
C14823 VP.t623 a_400_38200# 0.02fF
C14824 VP.n7659 a_400_38200# 0.14fF
C14825 VP.n7661 a_400_38200# 1.93fF
C14826 VP.t306 a_400_38200# 0.02fF
C14827 VP.n7662 a_400_38200# 0.24fF
C14828 VP.n7663 a_400_38200# 0.35fF
C14829 VP.n7664 a_400_38200# 0.60fF
C14830 VP.n7665 a_400_38200# 0.12fF
C14831 VP.t1014 a_400_38200# 0.02fF
C14832 VP.n7666 a_400_38200# 0.14fF
C14833 VP.n7668 a_400_38200# 0.04fF
C14834 VP.n7669 a_400_38200# 0.02fF
C14835 VP.n7670 a_400_38200# 0.06fF
C14836 VP.n7671 a_400_38200# 0.30fF
C14837 VP.n7672 a_400_38200# 0.10fF
C14838 VP.n7673 a_400_38200# 0.28fF
C14839 VP.n7674 a_400_38200# 0.15fF
C14840 VP.n7675 a_400_38200# 0.08fF
C14841 VP.n7676 a_400_38200# 0.14fF
C14842 VP.n7677 a_400_38200# 0.06fF
C14843 VP.n7678 a_400_38200# 0.06fF
C14844 VP.n7679 a_400_38200# 0.03fF
C14845 VP.n7680 a_400_38200# 0.05fF
C14846 VP.n7681 a_400_38200# 0.07fF
C14847 VP.n7682 a_400_38200# 0.19fF
C14848 VP.n7683 a_400_38200# 0.59fF
C14849 VP.n7684 a_400_38200# 0.34fF
C14850 VP.n7685 a_400_38200# 2.18fF
C14851 VP.t1327 a_400_38200# 0.02fF
C14852 VP.n7686 a_400_38200# 0.24fF
C14853 VP.n7687 a_400_38200# 0.91fF
C14854 VP.n7688 a_400_38200# 0.05fF
C14855 VP.t112 a_400_38200# 0.02fF
C14856 VP.n7689 a_400_38200# 0.12fF
C14857 VP.n7690 a_400_38200# 0.14fF
C14858 VP.n7692 a_400_38200# 0.10fF
C14859 VP.n7693 a_400_38200# 0.10fF
C14860 VP.n7694 a_400_38200# 0.18fF
C14861 VP.n7695 a_400_38200# 0.09fF
C14862 VP.n7696 a_400_38200# 0.04fF
C14863 VP.n7697 a_400_38200# 0.26fF
C14864 VP.n7698 a_400_38200# 1.17fF
C14865 VP.n7699 a_400_38200# 0.06fF
C14866 VP.n7700 a_400_38200# 0.44fF
C14867 VP.n7701 a_400_38200# 0.13fF
C14868 VP.n7702 a_400_38200# 0.02fF
C14869 VP.n7703 a_400_38200# 1.81fF
C14870 VP.n7704 a_400_38200# 0.12fF
C14871 VP.t1336 a_400_38200# 0.02fF
C14872 VP.n7705 a_400_38200# 0.14fF
C14873 VP.t553 a_400_38200# 0.02fF
C14874 VP.n7707 a_400_38200# 0.24fF
C14875 VP.n7708 a_400_38200# 0.35fF
C14876 VP.n7709 a_400_38200# 0.60fF
C14877 VP.n7710 a_400_38200# 2.28fF
C14878 VP.t266 a_400_38200# 0.02fF
C14879 VP.n7711 a_400_38200# 0.24fF
C14880 VP.n7712 a_400_38200# 0.91fF
C14881 VP.n7713 a_400_38200# 0.05fF
C14882 VP.t383 a_400_38200# 0.02fF
C14883 VP.n7714 a_400_38200# 0.12fF
C14884 VP.n7715 a_400_38200# 0.14fF
C14885 VP.n7717 a_400_38200# 0.06fF
C14886 VP.n7718 a_400_38200# 0.09fF
C14887 VP.n7719 a_400_38200# 0.09fF
C14888 VP.n7720 a_400_38200# 1.45fF
C14889 VP.n7721 a_400_38200# 0.14fF
C14890 VP.n7722 a_400_38200# 0.07fF
C14891 VP.n7723 a_400_38200# 0.72fF
C14892 VP.n7724 a_400_38200# 1.81fF
C14893 VP.n7725 a_400_38200# 0.12fF
C14894 VP.t886 a_400_38200# 0.02fF
C14895 VP.n7726 a_400_38200# 0.14fF
C14896 VP.t171 a_400_38200# 0.02fF
C14897 VP.n7728 a_400_38200# 0.24fF
C14898 VP.n7729 a_400_38200# 0.35fF
C14899 VP.n7730 a_400_38200# 0.60fF
C14900 VP.n7731 a_400_38200# 2.30fF
C14901 VP.t1195 a_400_38200# 0.02fF
C14902 VP.n7732 a_400_38200# 0.24fF
C14903 VP.n7733 a_400_38200# 0.91fF
C14904 VP.n7734 a_400_38200# 0.05fF
C14905 VP.t1239 a_400_38200# 0.02fF
C14906 VP.n7735 a_400_38200# 0.12fF
C14907 VP.n7736 a_400_38200# 0.14fF
C14908 VP.n7738 a_400_38200# 0.06fF
C14909 VP.n7739 a_400_38200# 0.25fF
C14910 VP.n7740 a_400_38200# 0.45fF
C14911 VP.n7741 a_400_38200# 0.03fF
C14912 VP.n7742 a_400_38200# 0.05fF
C14913 VP.n7743 a_400_38200# 0.07fF
C14914 VP.n7744 a_400_38200# 0.06fF
C14915 VP.n7745 a_400_38200# 0.06fF
C14916 VP.n7746 a_400_38200# 0.19fF
C14917 VP.n7747 a_400_38200# 0.59fF
C14918 VP.n7748 a_400_38200# 0.34fF
C14919 VP.n7749 a_400_38200# 0.05fF
C14920 VP.n7750 a_400_38200# 0.30fF
C14921 VP.n7751 a_400_38200# 1.93fF
C14922 VP.n7752 a_400_38200# 0.12fF
C14923 VP.t437 a_400_38200# 0.02fF
C14924 VP.n7753 a_400_38200# 0.14fF
C14925 VP.t1020 a_400_38200# 0.02fF
C14926 VP.n7755 a_400_38200# 0.24fF
C14927 VP.n7756 a_400_38200# 0.35fF
C14928 VP.n7757 a_400_38200# 0.60fF
C14929 VP.n7758 a_400_38200# 2.04fF
C14930 VP.t742 a_400_38200# 0.02fF
C14931 VP.n7759 a_400_38200# 0.24fF
C14932 VP.n7760 a_400_38200# 0.91fF
C14933 VP.n7761 a_400_38200# 0.05fF
C14934 VP.t794 a_400_38200# 0.02fF
C14935 VP.n7762 a_400_38200# 0.12fF
C14936 VP.n7763 a_400_38200# 0.14fF
C14937 VP.n7765 a_400_38200# 0.24fF
C14938 VP.t289 a_400_38200# 0.02fF
C14939 VP.n7766 a_400_38200# 0.36fF
C14940 VP.n7767 a_400_38200# 0.36fF
C14941 VP.n7768 a_400_38200# 0.67fF
C14942 VP.n7769 a_400_38200# 0.06fF
C14943 VP.n7770 a_400_38200# 0.09fF
C14944 VP.n7771 a_400_38200# 0.09fF
C14945 VP.n7772 a_400_38200# 1.45fF
C14946 VP.n7773 a_400_38200# 0.14fF
C14947 VP.n7774 a_400_38200# 0.07fF
C14948 VP.n7775 a_400_38200# 0.72fF
C14949 VP.n7776 a_400_38200# 1.81fF
C14950 VP.n7777 a_400_38200# 1.06fF
C14951 VP.n7778 a_400_38200# 0.24fF
C14952 VP.t573 a_400_38200# 0.02fF
C14953 VP.n7779 a_400_38200# 0.35fF
C14954 VP.n7780 a_400_38200# 0.63fF
C14955 VP.n7781 a_400_38200# 0.40fF
C14956 VP.n7782 a_400_38200# 0.40fF
C14957 VP.n7783 a_400_38200# 0.12fF
C14958 VP.t1291 a_400_38200# 0.02fF
C14959 VP.n7784 a_400_38200# 0.14fF
C14960 VP.t348 a_400_38200# 0.02fF
C14961 VP.n7786 a_400_38200# 0.12fF
C14962 VP.n7787 a_400_38200# 0.14fF
C14963 VP.n7789 a_400_38200# 1.93fF
C14964 VP.n7790 a_400_38200# 2.23fF
C14965 VP.t104 a_400_38200# 0.02fF
C14966 VP.n7791 a_400_38200# 0.24fF
C14967 VP.n7792 a_400_38200# 0.35fF
C14968 VP.n7793 a_400_38200# 0.60fF
C14969 VP.n7794 a_400_38200# 0.12fF
C14970 VP.t847 a_400_38200# 0.02fF
C14971 VP.n7795 a_400_38200# 0.14fF
C14972 VP.n7797 a_400_38200# 0.07fF
C14973 VP.n7798 a_400_38200# 0.30fF
C14974 VP.n7799 a_400_38200# 0.06fF
C14975 VP.n7800 a_400_38200# 0.25fF
C14976 VP.n7801 a_400_38200# 0.45fF
C14977 VP.n7802 a_400_38200# 0.06fF
C14978 VP.n7803 a_400_38200# 0.06fF
C14979 VP.n7804 a_400_38200# 0.03fF
C14980 VP.n7805 a_400_38200# 0.05fF
C14981 VP.n7806 a_400_38200# 0.07fF
C14982 VP.n7807 a_400_38200# 0.19fF
C14983 VP.n7808 a_400_38200# 0.59fF
C14984 VP.n7809 a_400_38200# 0.34fF
C14985 VP.n7810 a_400_38200# 2.04fF
C14986 VP.t1140 a_400_38200# 0.02fF
C14987 VP.n7811 a_400_38200# 0.24fF
C14988 VP.n7812 a_400_38200# 0.91fF
C14989 VP.n7813 a_400_38200# 0.05fF
C14990 VP.t1197 a_400_38200# 0.02fF
C14991 VP.n7814 a_400_38200# 0.12fF
C14992 VP.n7815 a_400_38200# 0.14fF
C14993 VP.n7817 a_400_38200# 0.06fF
C14994 VP.n7818 a_400_38200# 0.09fF
C14995 VP.n7819 a_400_38200# 0.09fF
C14996 VP.n7820 a_400_38200# 1.45fF
C14997 VP.n7821 a_400_38200# 0.14fF
C14998 VP.n7822 a_400_38200# 0.07fF
C14999 VP.n7823 a_400_38200# 0.72fF
C15000 VP.n7824 a_400_38200# 1.81fF
C15001 VP.n7825 a_400_38200# 0.12fF
C15002 VP.t397 a_400_38200# 0.02fF
C15003 VP.n7826 a_400_38200# 0.14fF
C15004 VP.t980 a_400_38200# 0.02fF
C15005 VP.n7828 a_400_38200# 0.24fF
C15006 VP.n7829 a_400_38200# 0.35fF
C15007 VP.n7830 a_400_38200# 0.60fF
C15008 VP.n7831 a_400_38200# 2.30fF
C15009 VP.t691 a_400_38200# 0.02fF
C15010 VP.n7832 a_400_38200# 0.24fF
C15011 VP.n7833 a_400_38200# 0.91fF
C15012 VP.n7834 a_400_38200# 0.05fF
C15013 VP.t745 a_400_38200# 0.02fF
C15014 VP.n7835 a_400_38200# 0.12fF
C15015 VP.n7836 a_400_38200# 0.14fF
C15016 VP.n7838 a_400_38200# 1.93fF
C15017 VP.n7839 a_400_38200# 2.23fF
C15018 VP.t533 a_400_38200# 0.02fF
C15019 VP.n7840 a_400_38200# 0.24fF
C15020 VP.n7841 a_400_38200# 0.35fF
C15021 VP.n7842 a_400_38200# 0.60fF
C15022 VP.n7843 a_400_38200# 0.12fF
C15023 VP.t1253 a_400_38200# 0.02fF
C15024 VP.n7844 a_400_38200# 0.14fF
C15025 VP.n7846 a_400_38200# 0.07fF
C15026 VP.n7847 a_400_38200# 0.30fF
C15027 VP.n7848 a_400_38200# 0.06fF
C15028 VP.n7849 a_400_38200# 0.25fF
C15029 VP.n7850 a_400_38200# 0.45fF
C15030 VP.n7851 a_400_38200# 0.06fF
C15031 VP.n7852 a_400_38200# 0.06fF
C15032 VP.n7853 a_400_38200# 0.03fF
C15033 VP.n7854 a_400_38200# 0.05fF
C15034 VP.n7855 a_400_38200# 0.07fF
C15035 VP.n7856 a_400_38200# 0.19fF
C15036 VP.n7857 a_400_38200# 0.59fF
C15037 VP.n7858 a_400_38200# 0.34fF
C15038 VP.n7859 a_400_38200# 2.04fF
C15039 VP.t247 a_400_38200# 0.02fF
C15040 VP.n7860 a_400_38200# 0.24fF
C15041 VP.n7861 a_400_38200# 0.91fF
C15042 VP.n7862 a_400_38200# 0.05fF
C15043 VP.t364 a_400_38200# 0.02fF
C15044 VP.n7863 a_400_38200# 0.12fF
C15045 VP.n7864 a_400_38200# 0.14fF
C15046 VP.n7866 a_400_38200# 0.06fF
C15047 VP.n7867 a_400_38200# 0.09fF
C15048 VP.n7868 a_400_38200# 0.09fF
C15049 VP.n7869 a_400_38200# 0.43fF
C15050 VP.n7870 a_400_38200# 0.69fF
C15051 VP.n7871 a_400_38200# 0.14fF
C15052 VP.n7872 a_400_38200# 0.07fF
C15053 VP.n7873 a_400_38200# 0.72fF
C15054 VP.n7874 a_400_38200# 1.81fF
C15055 VP.n7875 a_400_38200# 0.12fF
C15056 VP.t808 a_400_38200# 0.02fF
C15057 VP.n7876 a_400_38200# 0.14fF
C15058 VP.t56 a_400_38200# 0.02fF
C15059 VP.n7878 a_400_38200# 0.24fF
C15060 VP.n7879 a_400_38200# 0.35fF
C15061 VP.n7880 a_400_38200# 0.60fF
C15062 VP.n7881 a_400_38200# 2.30fF
C15063 VP.t1102 a_400_38200# 0.02fF
C15064 VP.n7882 a_400_38200# 0.24fF
C15065 VP.n7883 a_400_38200# 0.91fF
C15066 VP.n7884 a_400_38200# 0.05fF
C15067 VP.t1220 a_400_38200# 0.02fF
C15068 VP.n7885 a_400_38200# 0.12fF
C15069 VP.n7886 a_400_38200# 0.14fF
C15070 VP.n7888 a_400_38200# 0.31fF
C15071 VP.n7889 a_400_38200# 0.04fF
C15072 VP.n7890 a_400_38200# 0.88fF
C15073 VP.n7891 a_400_38200# 0.48fF
C15074 VP.n7892 a_400_38200# 0.88fF
C15075 VP.n7893 a_400_38200# 0.60fF
C15076 VP.n7894 a_400_38200# 2.33fF
C15077 VP.n7895 a_400_38200# 0.59fF
C15078 VP.n7896 a_400_38200# 0.02fF
C15079 VP.n7897 a_400_38200# 0.96fF
C15080 VP.t10 a_400_38200# 15.72fF
C15081 VP.n7898 a_400_38200# 15.42fF
C15082 VP.n7900 a_400_38200# 0.38fF
C15083 VP.n7901 a_400_38200# 0.23fF
C15084 VP.n7902 a_400_38200# 3.28fF
C15085 VP.n7903 a_400_38200# 1.41fF
C15086 VP.n7904 a_400_38200# 0.30fF
C15087 VP.t1192 a_400_38200# 0.02fF
C15088 VP.n7905 a_400_38200# 0.64fF
C15089 VP.n7906 a_400_38200# 0.60fF
C15090 VP.n7907 a_400_38200# 1.88fF
C15091 VP.n7908 a_400_38200# 4.64fF
C15092 VP.t912 a_400_38200# 0.02fF
C15093 VP.n7909 a_400_38200# 1.19fF
C15094 VP.n7910 a_400_38200# 0.05fF
C15095 VP.t1008 a_400_38200# 0.02fF
C15096 VP.n7911 a_400_38200# 0.01fF
C15097 VP.n7912 a_400_38200# 0.26fF
C15098 VP.n7914 a_400_38200# 15.28fF
C15099 VP.n7915 a_400_38200# 0.10fF
C15100 VP.n7916 a_400_38200# 0.28fF
C15101 VP.n7917 a_400_38200# 0.15fF
C15102 VP.n7918 a_400_38200# 0.08fF
C15103 VP.n7919 a_400_38200# 0.14fF
C15104 VP.n7920 a_400_38200# 0.06fF
C15105 VP.n7921 a_400_38200# 0.06fF
C15106 VP.n7922 a_400_38200# 0.03fF
C15107 VP.n7923 a_400_38200# 0.05fF
C15108 VP.n7924 a_400_38200# 0.07fF
C15109 VP.n7925 a_400_38200# 0.19fF
C15110 VP.n7926 a_400_38200# 0.59fF
C15111 VP.n7927 a_400_38200# 0.34fF
C15112 VP.n7928 a_400_38200# 0.04fF
C15113 VP.n7929 a_400_38200# 0.02fF
C15114 VP.n7930 a_400_38200# 0.06fF
C15115 VP.n7931 a_400_38200# 0.30fF
C15116 VP.n7932 a_400_38200# 1.93fF
C15117 VP.n7933 a_400_38200# 0.12fF
C15118 VP.t163 a_400_38200# 0.02fF
C15119 VP.n7934 a_400_38200# 0.14fF
C15120 VP.t758 a_400_38200# 0.02fF
C15121 VP.n7936 a_400_38200# 0.24fF
C15122 VP.n7937 a_400_38200# 0.35fF
C15123 VP.n7938 a_400_38200# 0.60fF
C15124 VP.n7939 a_400_38200# 2.39fF
C15125 VP.n7940 a_400_38200# 1.79fF
C15126 VP.t578 a_400_38200# 0.02fF
C15127 VP.n7941 a_400_38200# 0.12fF
C15128 VP.n7942 a_400_38200# 0.14fF
C15129 VP.t479 a_400_38200# 0.02fF
C15130 VP.n7944 a_400_38200# 0.24fF
C15131 VP.n7945 a_400_38200# 0.91fF
C15132 VP.n7946 a_400_38200# 0.05fF
C15133 VP.n7947 a_400_38200# 1.93fF
C15134 VP.n7948 a_400_38200# 2.72fF
C15135 VP.t943 a_400_38200# 0.02fF
C15136 VP.n7949 a_400_38200# 0.24fF
C15137 VP.n7950 a_400_38200# 0.35fF
C15138 VP.n7951 a_400_38200# 0.60fF
C15139 VP.n7952 a_400_38200# 0.12fF
C15140 VP.t359 a_400_38200# 0.02fF
C15141 VP.n7953 a_400_38200# 0.14fF
C15142 VP.n7955 a_400_38200# 0.02fF
C15143 VP.n7956 a_400_38200# 0.32fF
C15144 VP.n7957 a_400_38200# 0.04fF
C15145 VP.n7958 a_400_38200# 0.05fF
C15146 VP.n7959 a_400_38200# 0.04fF
C15147 VP.n7960 a_400_38200# 0.12fF
C15148 VP.n7961 a_400_38200# 0.09fF
C15149 VP.n7962 a_400_38200# 0.14fF
C15150 VP.n7963 a_400_38200# 0.08fF
C15151 VP.n7964 a_400_38200# 0.09fF
C15152 VP.n7965 a_400_38200# 0.07fF
C15153 VP.n7966 a_400_38200# 0.56fF
C15154 VP.n7967 a_400_38200# 0.20fF
C15155 VP.n7968 a_400_38200# 2.19fF
C15156 VP.t773 a_400_38200# 0.02fF
C15157 VP.n7969 a_400_38200# 0.12fF
C15158 VP.n7970 a_400_38200# 0.14fF
C15159 VP.t660 a_400_38200# 0.02fF
C15160 VP.n7972 a_400_38200# 0.24fF
C15161 VP.n7973 a_400_38200# 0.91fF
C15162 VP.n7974 a_400_38200# 0.05fF
C15163 VP.t111 a_400_38200# 34.79fF
C15164 VP.t1026 a_400_38200# 0.02fF
C15165 VP.n7975 a_400_38200# 0.12fF
C15166 VP.n7976 a_400_38200# 0.14fF
C15167 VP.t927 a_400_38200# 0.02fF
C15168 VP.n7978 a_400_38200# 0.24fF
C15169 VP.n7979 a_400_38200# 0.91fF
C15170 VP.n7980 a_400_38200# 0.05fF
C15171 VP.t1207 a_400_38200# 0.02fF
C15172 VP.n7981 a_400_38200# 0.24fF
C15173 VP.n7982 a_400_38200# 0.35fF
C15174 VP.n7983 a_400_38200# 0.60fF
C15175 VP.n7984 a_400_38200# 0.04fF
C15176 VP.n7985 a_400_38200# 0.08fF
C15177 VP.n7986 a_400_38200# 0.72fF
C15178 VP.n7987 a_400_38200# 0.09fF
C15179 VP.n7988 a_400_38200# 0.00fF
C15180 VP.n7989 a_400_38200# 1.22fF
C15181 VP.n7990 a_400_38200# 0.19fF
C15182 VP.n7992 a_400_38200# 1.72fF
C15183 VP.n7993 a_400_38200# 1.96fF
C15184 VP.n7994 a_400_38200# 1.04fF
C15185 VP.n7995 a_400_38200# 0.05fF
C15186 VP.n7996 a_400_38200# 0.03fF
C15187 VP.n7997 a_400_38200# 0.06fF
C15188 VP.n7998 a_400_38200# 0.06fF
C15189 VP.n7999 a_400_38200# 0.06fF
C15190 VP.n8000 a_400_38200# 0.07fF
C15191 VP.n8001 a_400_38200# 0.03fF
C15192 VP.n8002 a_400_38200# 0.05fF
C15193 VP.n8003 a_400_38200# 0.07fF
C15194 VP.n8004 a_400_38200# 0.19fF
C15195 VP.n8005 a_400_38200# 0.60fF
C15196 VP.n8006 a_400_38200# 0.76fF
C15197 VP.n8007 a_400_38200# 0.40fF
C15198 VP.n8008 a_400_38200# 0.03fF
C15199 VP.n8009 a_400_38200# 0.01fF
C15200 VP.t749 a_400_38200# 0.02fF
C15201 VP.n8010 a_400_38200# 0.25fF
C15202 VP.t470 a_400_38200# 0.02fF
C15203 VP.n8011 a_400_38200# 0.95fF
C15204 VP.n8012 a_400_38200# 0.70fF
C15205 VP.n8013 a_400_38200# 1.93fF
C15206 VP.n8014 a_400_38200# 2.97fF
C15207 VP.n8015 a_400_38200# 2.27fF
C15208 VP.t436 a_400_38200# 0.02fF
C15209 VP.n8016 a_400_38200# 0.24fF
C15210 VP.n8017 a_400_38200# 0.35fF
C15211 VP.n8018 a_400_38200# 0.60fF
C15212 VP.n8019 a_400_38200# 0.12fF
C15213 VP.t1145 a_400_38200# 0.02fF
C15214 VP.n8020 a_400_38200# 0.14fF
C15215 VP.n8022 a_400_38200# 0.04fF
C15216 VP.n8023 a_400_38200# 0.02fF
C15217 VP.n8024 a_400_38200# 0.06fF
C15218 VP.n8025 a_400_38200# 0.30fF
C15219 VP.n8026 a_400_38200# 0.10fF
C15220 VP.n8027 a_400_38200# 0.06fF
C15221 VP.n8028 a_400_38200# 0.06fF
C15222 VP.n8029 a_400_38200# 0.28fF
C15223 VP.n8030 a_400_38200# 0.03fF
C15224 VP.n8031 a_400_38200# 0.15fF
C15225 VP.n8032 a_400_38200# 0.08fF
C15226 VP.n8033 a_400_38200# 0.14fF
C15227 VP.n8034 a_400_38200# 0.03fF
C15228 VP.n8035 a_400_38200# 0.06fF
C15229 VP.n8036 a_400_38200# 0.06fF
C15230 VP.n8037 a_400_38200# 0.06fF
C15231 VP.n8038 a_400_38200# 0.06fF
C15232 VP.n8039 a_400_38200# 0.03fF
C15233 VP.n8040 a_400_38200# 0.05fF
C15234 VP.n8041 a_400_38200# 0.07fF
C15235 VP.n8042 a_400_38200# 0.19fF
C15236 VP.n8043 a_400_38200# 0.59fF
C15237 VP.n8044 a_400_38200# 0.34fF
C15238 VP.n8045 a_400_38200# 1.88fF
C15239 VP.t867 a_400_38200# 0.02fF
C15240 VP.n8046 a_400_38200# 0.24fF
C15241 VP.n8047 a_400_38200# 0.91fF
C15242 VP.n8048 a_400_38200# 0.05fF
C15243 VP.t1189 a_400_38200# 0.02fF
C15244 VP.n8049 a_400_38200# 0.12fF
C15245 VP.n8050 a_400_38200# 0.14fF
C15246 VP.n8052 a_400_38200# 0.19fF
C15247 VP.n8053 a_400_38200# 0.10fF
C15248 VP.n8054 a_400_38200# 0.10fF
C15249 VP.n8055 a_400_38200# 0.18fF
C15250 VP.n8056 a_400_38200# 0.09fF
C15251 VP.n8057 a_400_38200# 0.04fF
C15252 VP.n8058 a_400_38200# 0.19fF
C15253 VP.n8059 a_400_38200# 0.26fF
C15254 VP.n8060 a_400_38200# 1.17fF
C15255 VP.n8061 a_400_38200# 0.06fF
C15256 VP.n8062 a_400_38200# 0.44fF
C15257 VP.n8063 a_400_38200# 0.13fF
C15258 VP.n8064 a_400_38200# 0.02fF
C15259 VP.n8065 a_400_38200# 1.81fF
C15260 VP.n8066 a_400_38200# 0.12fF
C15261 VP.t71 a_400_38200# 0.02fF
C15262 VP.n8067 a_400_38200# 0.14fF
C15263 VP.t680 a_400_38200# 0.02fF
C15264 VP.n8069 a_400_38200# 0.24fF
C15265 VP.n8070 a_400_38200# 0.35fF
C15266 VP.n8071 a_400_38200# 0.60fF
C15267 VP.n8072 a_400_38200# 3.18fF
C15268 VP.n8073 a_400_38200# 2.06fF
C15269 VP.n8074 a_400_38200# 1.98fF
C15270 VP.t1111 a_400_38200# 0.02fF
C15271 VP.n8075 a_400_38200# 0.24fF
C15272 VP.n8076 a_400_38200# 0.91fF
C15273 VP.n8077 a_400_38200# 0.05fF
C15274 VP.t737 a_400_38200# 0.02fF
C15275 VP.n8078 a_400_38200# 0.12fF
C15276 VP.n8079 a_400_38200# 0.14fF
C15277 VP.n8081 a_400_38200# 0.16fF
C15278 VP.n8082 a_400_38200# 0.19fF
C15279 VP.n8083 a_400_38200# 0.09fF
C15280 VP.n8084 a_400_38200# 0.04fF
C15281 VP.n8085 a_400_38200# 0.14fF
C15282 VP.n8086 a_400_38200# 0.64fF
C15283 VP.n8087 a_400_38200# 1.32fF
C15284 VP.n8088 a_400_38200# 1.81fF
C15285 VP.n8089 a_400_38200# 0.12fF
C15286 VP.t954 a_400_38200# 0.02fF
C15287 VP.n8090 a_400_38200# 0.14fF
C15288 VP.t236 a_400_38200# 0.02fF
C15289 VP.n8092 a_400_38200# 0.24fF
C15290 VP.n8093 a_400_38200# 0.35fF
C15291 VP.n8094 a_400_38200# 0.60fF
C15292 VP.n8095 a_400_38200# 2.97fF
C15293 VP.n8096 a_400_38200# 2.27fF
C15294 VP.n8097 a_400_38200# 2.00fF
C15295 VP.t668 a_400_38200# 0.02fF
C15296 VP.n8098 a_400_38200# 0.24fF
C15297 VP.n8099 a_400_38200# 0.91fF
C15298 VP.n8100 a_400_38200# 0.05fF
C15299 VP.t1057 a_400_38200# 0.02fF
C15300 VP.n8101 a_400_38200# 0.12fF
C15301 VP.n8102 a_400_38200# 0.14fF
C15302 VP.n8104 a_400_38200# 0.24fF
C15303 VP.t1076 a_400_38200# 0.02fF
C15304 VP.n8105 a_400_38200# 0.36fF
C15305 VP.n8106 a_400_38200# 0.36fF
C15306 VP.n8107 a_400_38200# 0.67fF
C15307 VP.n8108 a_400_38200# 0.16fF
C15308 VP.n8109 a_400_38200# 0.19fF
C15309 VP.n8110 a_400_38200# 0.09fF
C15310 VP.n8111 a_400_38200# 0.04fF
C15311 VP.n8112 a_400_38200# 0.14fF
C15312 VP.n8113 a_400_38200# 0.64fF
C15313 VP.n8114 a_400_38200# 1.32fF
C15314 VP.n8115 a_400_38200# 1.81fF
C15315 VP.n8116 a_400_38200# 2.97fF
C15316 VP.n8117 a_400_38200# 2.27fF
C15317 VP.n8118 a_400_38200# 0.75fF
C15318 VP.n8119 a_400_38200# 0.24fF
C15319 VP.t649 a_400_38200# 0.02fF
C15320 VP.n8120 a_400_38200# 0.35fF
C15321 VP.n8121 a_400_38200# 0.63fF
C15322 VP.n8122 a_400_38200# 0.40fF
C15323 VP.n8123 a_400_38200# 0.40fF
C15324 VP.n8124 a_400_38200# 0.12fF
C15325 VP.t19 a_400_38200# 0.02fF
C15326 VP.n8125 a_400_38200# 0.14fF
C15327 VP.t145 a_400_38200# 0.02fF
C15328 VP.n8127 a_400_38200# 0.12fF
C15329 VP.n8128 a_400_38200# 0.14fF
C15330 VP.n8130 a_400_38200# 0.16fF
C15331 VP.n8131 a_400_38200# 0.19fF
C15332 VP.n8132 a_400_38200# 0.09fF
C15333 VP.n8133 a_400_38200# 0.04fF
C15334 VP.n8134 a_400_38200# 0.14fF
C15335 VP.n8135 a_400_38200# 0.64fF
C15336 VP.n8136 a_400_38200# 1.32fF
C15337 VP.n8137 a_400_38200# 1.81fF
C15338 VP.n8138 a_400_38200# 0.12fF
C15339 VP.t468 a_400_38200# 0.02fF
C15340 VP.n8139 a_400_38200# 0.14fF
C15341 VP.t1054 a_400_38200# 0.02fF
C15342 VP.n8141 a_400_38200# 0.24fF
C15343 VP.n8142 a_400_38200# 0.35fF
C15344 VP.n8143 a_400_38200# 0.60fF
C15345 VP.n8144 a_400_38200# 2.97fF
C15346 VP.n8145 a_400_38200# 2.27fF
C15347 VP.n8146 a_400_38200# 2.00fF
C15348 VP.t177 a_400_38200# 0.02fF
C15349 VP.n8147 a_400_38200# 0.24fF
C15350 VP.n8148 a_400_38200# 0.91fF
C15351 VP.n8149 a_400_38200# 0.05fF
C15352 VP.t560 a_400_38200# 0.02fF
C15353 VP.n8150 a_400_38200# 0.12fF
C15354 VP.n8151 a_400_38200# 0.14fF
C15355 VP.n8153 a_400_38200# 0.16fF
C15356 VP.n8154 a_400_38200# 0.19fF
C15357 VP.n8155 a_400_38200# 0.09fF
C15358 VP.n8156 a_400_38200# 0.04fF
C15359 VP.n8157 a_400_38200# 0.14fF
C15360 VP.n8158 a_400_38200# 0.64fF
C15361 VP.n8159 a_400_38200# 1.32fF
C15362 VP.n8160 a_400_38200# 1.81fF
C15363 VP.n8161 a_400_38200# 0.12fF
C15364 VP.t937 a_400_38200# 0.02fF
C15365 VP.n8162 a_400_38200# 0.14fF
C15366 VP.t219 a_400_38200# 0.02fF
C15367 VP.n8164 a_400_38200# 0.24fF
C15368 VP.n8165 a_400_38200# 0.35fF
C15369 VP.n8166 a_400_38200# 0.60fF
C15370 VP.n8167 a_400_38200# 2.97fF
C15371 VP.n8168 a_400_38200# 2.27fF
C15372 VP.n8169 a_400_38200# 2.00fF
C15373 VP.t652 a_400_38200# 0.02fF
C15374 VP.n8170 a_400_38200# 0.24fF
C15375 VP.n8171 a_400_38200# 0.91fF
C15376 VP.n8172 a_400_38200# 0.05fF
C15377 VP.t967 a_400_38200# 0.02fF
C15378 VP.n8173 a_400_38200# 0.12fF
C15379 VP.n8174 a_400_38200# 0.14fF
C15380 VP.n8176 a_400_38200# 0.09fF
C15381 VP.n8177 a_400_38200# 0.03fF
C15382 VP.n8178 a_400_38200# 0.04fF
C15383 VP.n8179 a_400_38200# 0.37fF
C15384 VP.n8180 a_400_38200# 0.11fF
C15385 VP.n8181 a_400_38200# 0.05fF
C15386 VP.n8182 a_400_38200# 0.08fF
C15387 VP.n8183 a_400_38200# 0.10fF
C15388 VP.n8184 a_400_38200# 0.06fF
C15389 VP.n8185 a_400_38200# 0.08fF
C15390 VP.n8186 a_400_38200# 0.19fF
C15391 VP.n8187 a_400_38200# 0.06fF
C15392 VP.n8188 a_400_38200# 0.15fF
C15393 VP.n8189 a_400_38200# 0.14fF
C15394 VP.n8190 a_400_38200# 0.13fF
C15395 VP.n8191 a_400_38200# 0.12fF
C15396 VP.n8192 a_400_38200# 0.05fF
C15397 VP.n8193 a_400_38200# 0.17fF
C15398 VP.n8194 a_400_38200# 0.26fF
C15399 VP.n8195 a_400_38200# 0.37fF
C15400 VP.n8196 a_400_38200# 0.27fF
C15401 VP.n8197 a_400_38200# 2.05fF
C15402 VP.n8198 a_400_38200# 0.12fF
C15403 VP.t726 a_400_38200# 0.02fF
C15404 VP.n8199 a_400_38200# 0.14fF
C15405 VP.t1318 a_400_38200# 0.02fF
C15406 VP.n8201 a_400_38200# 0.24fF
C15407 VP.n8202 a_400_38200# 0.35fF
C15408 VP.n8203 a_400_38200# 0.60fF
C15409 VP.n8204 a_400_38200# 2.87fF
C15410 VP.n8205 a_400_38200# 2.00fF
C15411 VP.t447 a_400_38200# 0.02fF
C15412 VP.n8206 a_400_38200# 0.24fF
C15413 VP.n8207 a_400_38200# 0.91fF
C15414 VP.n8208 a_400_38200# 0.05fF
C15415 VP.t39 a_400_38200# 0.02fF
C15416 VP.n8209 a_400_38200# 0.12fF
C15417 VP.n8210 a_400_38200# 0.14fF
C15418 VP.n8212 a_400_38200# 15.28fF
C15419 VP.n8213 a_400_38200# 0.10fF
C15420 VP.n8214 a_400_38200# 0.28fF
C15421 VP.n8215 a_400_38200# 0.06fF
C15422 VP.n8216 a_400_38200# 0.06fF
C15423 VP.n8217 a_400_38200# 0.03fF
C15424 VP.n8218 a_400_38200# 0.15fF
C15425 VP.n8219 a_400_38200# 0.08fF
C15426 VP.n8220 a_400_38200# 0.14fF
C15427 VP.n8221 a_400_38200# 0.03fF
C15428 VP.n8222 a_400_38200# 0.06fF
C15429 VP.n8223 a_400_38200# 0.06fF
C15430 VP.n8224 a_400_38200# 0.06fF
C15431 VP.n8225 a_400_38200# 0.06fF
C15432 VP.n8226 a_400_38200# 0.03fF
C15433 VP.n8227 a_400_38200# 0.05fF
C15434 VP.n8228 a_400_38200# 0.07fF
C15435 VP.n8229 a_400_38200# 0.19fF
C15436 VP.n8230 a_400_38200# 0.59fF
C15437 VP.n8231 a_400_38200# 0.34fF
C15438 VP.n8232 a_400_38200# 0.04fF
C15439 VP.n8233 a_400_38200# 0.02fF
C15440 VP.n8234 a_400_38200# 0.06fF
C15441 VP.n8235 a_400_38200# 0.30fF
C15442 VP.n8236 a_400_38200# 1.93fF
C15443 VP.n8237 a_400_38200# 0.12fF
C15444 VP.t294 a_400_38200# 0.02fF
C15445 VP.n8238 a_400_38200# 0.14fF
C15446 VP.t885 a_400_38200# 0.02fF
C15447 VP.n8240 a_400_38200# 0.24fF
C15448 VP.n8241 a_400_38200# 0.35fF
C15449 VP.n8242 a_400_38200# 0.60fF
C15450 VP.n8243 a_400_38200# 0.53fF
C15451 VP.n8244 a_400_38200# 1.39fF
C15452 VP.n8245 a_400_38200# 0.53fF
C15453 VP.n8246 a_400_38200# 0.21fF
C15454 VP.n8247 a_400_38200# 1.73fF
C15455 VP.t342 a_400_38200# 0.02fF
C15456 VP.n8248 a_400_38200# 0.12fF
C15457 VP.n8249 a_400_38200# 0.14fF
C15458 VP.t1316 a_400_38200# 0.02fF
C15459 VP.n8251 a_400_38200# 0.24fF
C15460 VP.n8252 a_400_38200# 0.91fF
C15461 VP.n8253 a_400_38200# 0.05fF
C15462 VP.n8254 a_400_38200# 0.06fF
C15463 VP.n8255 a_400_38200# 0.06fF
C15464 VP.n8256 a_400_38200# 0.03fF
C15465 VP.n8257 a_400_38200# 0.10fF
C15466 VP.n8258 a_400_38200# 0.17fF
C15467 VP.n8259 a_400_38200# 0.10fF
C15468 VP.n8260 a_400_38200# 0.13fF
C15469 VP.n8261 a_400_38200# 0.02fF
C15470 VP.n8262 a_400_38200# 0.04fF
C15471 VP.n8263 a_400_38200# 0.06fF
C15472 VP.n8264 a_400_38200# 0.09fF
C15473 VP.n8265 a_400_38200# 0.10fF
C15474 VP.n8266 a_400_38200# 0.05fF
C15475 VP.n8267 a_400_38200# 0.19fF
C15476 VP.n8268 a_400_38200# 0.16fF
C15477 VP.n8269 a_400_38200# 0.04fF
C15478 VP.n8270 a_400_38200# 0.05fF
C15479 VP.n8271 a_400_38200# 0.04fF
C15480 VP.n8272 a_400_38200# 0.12fF
C15481 VP.n8273 a_400_38200# 0.09fF
C15482 VP.n8274 a_400_38200# 0.14fF
C15483 VP.n8275 a_400_38200# 0.56fF
C15484 VP.n8276 a_400_38200# 0.10fF
C15485 VP.n8277 a_400_38200# 1.93fF
C15486 VP.n8278 a_400_38200# 0.12fF
C15487 VP.t508 a_400_38200# 0.02fF
C15488 VP.n8279 a_400_38200# 0.14fF
C15489 VP.t1091 a_400_38200# 0.02fF
C15490 VP.n8281 a_400_38200# 0.24fF
C15491 VP.n8282 a_400_38200# 0.35fF
C15492 VP.n8283 a_400_38200# 0.60fF
C15493 VP.n8284 a_400_38200# 2.23fF
C15494 VP.n8285 a_400_38200# 0.18fF
C15495 VP.n8286 a_400_38200# 0.45fF
C15496 VP.n8287 a_400_38200# 0.06fF
C15497 VP.n8288 a_400_38200# 0.01fF
C15498 VP.n8289 a_400_38200# 0.01fF
C15499 VP.n8290 a_400_38200# 0.04fF
C15500 VP.n8291 a_400_38200# 0.02fF
C15501 VP.n8292 a_400_38200# 0.07fF
C15502 VP.n8293 a_400_38200# 0.04fF
C15503 VP.n8294 a_400_38200# 0.14fF
C15504 VP.n8295 a_400_38200# 0.45fF
C15505 VP.n8296 a_400_38200# 1.46fF
C15506 VP.n8297 a_400_38200# 1.78fF
C15507 VP.t610 a_400_38200# 0.02fF
C15508 VP.n8298 a_400_38200# 0.12fF
C15509 VP.n8299 a_400_38200# 0.14fF
C15510 VP.t221 a_400_38200# 0.02fF
C15511 VP.n8301 a_400_38200# 0.24fF
C15512 VP.n8302 a_400_38200# 0.91fF
C15513 VP.n8303 a_400_38200# 0.05fF
C15514 VP.n8304 a_400_38200# 1.93fF
C15515 VP.n8305 a_400_38200# 0.18fF
C15516 VP.n8306 a_400_38200# 0.45fF
C15517 VP.n8307 a_400_38200# 0.06fF
C15518 VP.n8308 a_400_38200# 0.01fF
C15519 VP.n8309 a_400_38200# 0.01fF
C15520 VP.n8310 a_400_38200# 0.04fF
C15521 VP.n8311 a_400_38200# 0.02fF
C15522 VP.n8312 a_400_38200# 0.07fF
C15523 VP.n8313 a_400_38200# 0.04fF
C15524 VP.n8314 a_400_38200# 0.14fF
C15525 VP.n8315 a_400_38200# 0.45fF
C15526 VP.n8316 a_400_38200# 1.46fF
C15527 VP.t201 a_400_38200# 0.02fF
C15528 VP.n8317 a_400_38200# 0.24fF
C15529 VP.n8318 a_400_38200# 0.35fF
C15530 VP.n8319 a_400_38200# 0.60fF
C15531 VP.n8320 a_400_38200# 0.12fF
C15532 VP.t917 a_400_38200# 0.02fF
C15533 VP.n8321 a_400_38200# 0.14fF
C15534 VP.n8323 a_400_38200# 0.10fF
C15535 VP.n8324 a_400_38200# 0.17fF
C15536 VP.n8325 a_400_38200# 0.06fF
C15537 VP.n8326 a_400_38200# 0.06fF
C15538 VP.n8327 a_400_38200# 0.03fF
C15539 VP.n8328 a_400_38200# 0.10fF
C15540 VP.n8329 a_400_38200# 0.13fF
C15541 VP.n8330 a_400_38200# 0.13fF
C15542 VP.n8331 a_400_38200# 0.04fF
C15543 VP.n8332 a_400_38200# 0.05fF
C15544 VP.n8333 a_400_38200# 0.04fF
C15545 VP.n8334 a_400_38200# 0.09fF
C15546 VP.n8335 a_400_38200# 0.09fF
C15547 VP.n8336 a_400_38200# 0.05fF
C15548 VP.n8337 a_400_38200# 0.19fF
C15549 VP.n8338 a_400_38200# 0.12fF
C15550 VP.n8339 a_400_38200# 0.09fF
C15551 VP.n8340 a_400_38200# 0.14fF
C15552 VP.n8341 a_400_38200# 0.04fF
C15553 VP.n8342 a_400_38200# 0.02fF
C15554 VP.n8343 a_400_38200# 0.06fF
C15555 VP.n8344 a_400_38200# 0.56fF
C15556 VP.n8345 a_400_38200# 0.10fF
C15557 VP.n8346 a_400_38200# 1.78fF
C15558 VP.t1004 a_400_38200# 0.02fF
C15559 VP.n8347 a_400_38200# 0.12fF
C15560 VP.n8348 a_400_38200# 0.14fF
C15561 VP.t633 a_400_38200# 0.02fF
C15562 VP.n8350 a_400_38200# 0.24fF
C15563 VP.n8351 a_400_38200# 0.91fF
C15564 VP.n8352 a_400_38200# 0.05fF
C15565 VP.n8353 a_400_38200# 1.93fF
C15566 VP.n8354 a_400_38200# 0.18fF
C15567 VP.n8355 a_400_38200# 0.45fF
C15568 VP.n8356 a_400_38200# 0.06fF
C15569 VP.n8357 a_400_38200# 0.01fF
C15570 VP.n8358 a_400_38200# 0.01fF
C15571 VP.n8359 a_400_38200# 0.04fF
C15572 VP.n8360 a_400_38200# 0.02fF
C15573 VP.n8361 a_400_38200# 0.07fF
C15574 VP.n8362 a_400_38200# 0.04fF
C15575 VP.n8363 a_400_38200# 0.14fF
C15576 VP.n8364 a_400_38200# 0.45fF
C15577 VP.n8365 a_400_38200# 1.46fF
C15578 VP.t605 a_400_38200# 0.02fF
C15579 VP.n8366 a_400_38200# 0.24fF
C15580 VP.n8367 a_400_38200# 0.35fF
C15581 VP.n8368 a_400_38200# 0.60fF
C15582 VP.n8369 a_400_38200# 0.12fF
C15583 VP.t48 a_400_38200# 0.02fF
C15584 VP.n8370 a_400_38200# 0.14fF
C15585 VP.n8372 a_400_38200# 0.10fF
C15586 VP.n8373 a_400_38200# 0.17fF
C15587 VP.n8374 a_400_38200# 0.06fF
C15588 VP.n8375 a_400_38200# 0.06fF
C15589 VP.n8376 a_400_38200# 0.03fF
C15590 VP.n8377 a_400_38200# 0.10fF
C15591 VP.n8378 a_400_38200# 0.13fF
C15592 VP.n8379 a_400_38200# 0.13fF
C15593 VP.n8380 a_400_38200# 0.04fF
C15594 VP.n8381 a_400_38200# 0.05fF
C15595 VP.n8382 a_400_38200# 0.04fF
C15596 VP.n8383 a_400_38200# 0.09fF
C15597 VP.n8384 a_400_38200# 0.09fF
C15598 VP.n8385 a_400_38200# 0.05fF
C15599 VP.n8386 a_400_38200# 0.19fF
C15600 VP.n8387 a_400_38200# 0.12fF
C15601 VP.n8388 a_400_38200# 0.09fF
C15602 VP.n8389 a_400_38200# 0.14fF
C15603 VP.n8390 a_400_38200# 0.04fF
C15604 VP.n8391 a_400_38200# 0.02fF
C15605 VP.n8392 a_400_38200# 0.06fF
C15606 VP.n8393 a_400_38200# 0.56fF
C15607 VP.n8394 a_400_38200# 0.10fF
C15608 VP.n8395 a_400_38200# 1.78fF
C15609 VP.t89 a_400_38200# 0.02fF
C15610 VP.n8396 a_400_38200# 0.12fF
C15611 VP.n8397 a_400_38200# 0.14fF
C15612 VP.t1027 a_400_38200# 0.02fF
C15613 VP.n8399 a_400_38200# 0.24fF
C15614 VP.n8400 a_400_38200# 0.91fF
C15615 VP.n8401 a_400_38200# 0.05fF
C15616 VP.n8402 a_400_38200# 1.93fF
C15617 VP.n8403 a_400_38200# 0.18fF
C15618 VP.n8404 a_400_38200# 0.45fF
C15619 VP.n8405 a_400_38200# 0.06fF
C15620 VP.n8406 a_400_38200# 0.01fF
C15621 VP.n8407 a_400_38200# 0.01fF
C15622 VP.n8408 a_400_38200# 0.04fF
C15623 VP.n8409 a_400_38200# 0.02fF
C15624 VP.n8410 a_400_38200# 0.07fF
C15625 VP.n8411 a_400_38200# 0.04fF
C15626 VP.n8412 a_400_38200# 0.14fF
C15627 VP.n8413 a_400_38200# 0.53fF
C15628 VP.n8414 a_400_38200# 1.62fF
C15629 VP.t1074 a_400_38200# 0.02fF
C15630 VP.n8415 a_400_38200# 0.24fF
C15631 VP.n8416 a_400_38200# 0.35fF
C15632 VP.n8417 a_400_38200# 0.60fF
C15633 VP.n8418 a_400_38200# 0.12fF
C15634 VP.t491 a_400_38200# 0.02fF
C15635 VP.n8419 a_400_38200# 0.14fF
C15636 VP.n8421 a_400_38200# 0.10fF
C15637 VP.n8422 a_400_38200# 0.17fF
C15638 VP.n8423 a_400_38200# 0.06fF
C15639 VP.n8424 a_400_38200# 0.06fF
C15640 VP.n8425 a_400_38200# 0.03fF
C15641 VP.n8426 a_400_38200# 0.10fF
C15642 VP.n8427 a_400_38200# 0.13fF
C15643 VP.n8428 a_400_38200# 0.14fF
C15644 VP.n8429 a_400_38200# 0.04fF
C15645 VP.n8430 a_400_38200# 0.02fF
C15646 VP.n8431 a_400_38200# 0.03fF
C15647 VP.n8432 a_400_38200# 0.03fF
C15648 VP.n8433 a_400_38200# 0.05fF
C15649 VP.n8434 a_400_38200# 0.03fF
C15650 VP.n8435 a_400_38200# 0.04fF
C15651 VP.n8436 a_400_38200# 0.20fF
C15652 VP.n8437 a_400_38200# 0.14fF
C15653 VP.n8438 a_400_38200# 0.02fF
C15654 VP.n8439 a_400_38200# 0.07fF
C15655 VP.n8440 a_400_38200# 0.13fF
C15656 VP.n8441 a_400_38200# 0.04fF
C15657 VP.n8442 a_400_38200# 0.02fF
C15658 VP.n8443 a_400_38200# 0.06fF
C15659 VP.n8444 a_400_38200# 0.55fF
C15660 VP.n8445 a_400_38200# 0.10fF
C15661 VP.n8446 a_400_38200# 1.95fF
C15662 VP.t519 a_400_38200# 0.02fF
C15663 VP.n8447 a_400_38200# 0.12fF
C15664 VP.n8448 a_400_38200# 0.14fF
C15665 VP.t205 a_400_38200# 0.02fF
C15666 VP.n8450 a_400_38200# 0.24fF
C15667 VP.n8451 a_400_38200# 0.91fF
C15668 VP.n8452 a_400_38200# 0.05fF
C15669 VP.t18 a_400_38200# 35.17fF
C15670 VP.t1335 a_400_38200# 0.02fF
C15671 VP.n8453 a_400_38200# 1.21fF
C15672 VP.n8454 a_400_38200# 0.25fF
C15673 VP.n8455 a_400_38200# 26.29fF
C15674 VP.n8456 a_400_38200# 26.29fF
C15675 VP.n8457 a_400_38200# 0.76fF
C15676 VP.n8458 a_400_38200# 0.27fF
C15677 VP.n8459 a_400_38200# 0.59fF
C15678 VP.n8460 a_400_38200# 0.10fF
C15679 VP.n8461 a_400_38200# 3.02fF
C15680 VP.t200 a_400_38200# 15.72fF
C15681 VP.n8462 a_400_38200# 1.15fF
C15682 VP.n8464 a_400_38200# 13.70fF
C15683 VP.n8466 a_400_38200# 1.99fF
C15684 VP.n8467 a_400_38200# 4.39fF
C15685 VP.n8468 a_400_38200# 0.03fF
C15686 VP.n8469 a_400_38200# 0.05fF
C15687 VP.n8470 a_400_38200# 0.07fF
C15688 VP.n8471 a_400_38200# 0.03fF
C15689 VP.n8472 a_400_38200# 0.06fF
C15690 VP.n8473 a_400_38200# 0.06fF
C15691 VP.n8474 a_400_38200# 0.06fF
C15692 VP.n8475 a_400_38200# 0.07fF
C15693 VP.n8476 a_400_38200# 0.57fF
C15694 VP.n8477 a_400_38200# 1.88fF
C15695 VP.n8478 a_400_38200# 0.92fF
C15696 VP.n8479 a_400_38200# 2.63fF
C15697 VP.n8480 a_400_38200# 0.10fF
C15698 VP.n8481 a_400_38200# 0.28fF
C15699 VP.n8482 a_400_38200# 0.15fF
C15700 VP.n8483 a_400_38200# 0.08fF
C15701 VP.n8484 a_400_38200# 0.14fF
C15702 VP.n8485 a_400_38200# 0.06fF
C15703 VP.n8486 a_400_38200# 0.06fF
C15704 VP.n8487 a_400_38200# 0.03fF
C15705 VP.n8488 a_400_38200# 0.05fF
C15706 VP.n8489 a_400_38200# 0.07fF
C15707 VP.n8490 a_400_38200# 0.19fF
C15708 VP.n8491 a_400_38200# 0.59fF
C15709 VP.n8492 a_400_38200# 0.34fF
C15710 VP.n8493 a_400_38200# 0.04fF
C15711 VP.n8494 a_400_38200# 0.02fF
C15712 VP.n8495 a_400_38200# 0.06fF
C15713 VP.n8496 a_400_38200# 0.30fF
C15714 VP.n8497 a_400_38200# 0.12fF
C15715 VP.t771 a_400_38200# 0.02fF
C15716 VP.n8498 a_400_38200# 0.14fF
C15717 VP.n8500 a_400_38200# 1.93fF
C15718 VP.t907 a_400_38200# 0.02fF
C15719 VP.n8501 a_400_38200# 0.24fF
C15720 VP.n8502 a_400_38200# 0.35fF
C15721 VP.n8503 a_400_38200# 0.60fF
C15722 VP.n8504 a_400_38200# 0.12fF
C15723 VP.t319 a_400_38200# 0.02fF
C15724 VP.n8505 a_400_38200# 0.14fF
C15725 VP.n8507 a_400_38200# 0.04fF
C15726 VP.n8508 a_400_38200# 0.02fF
C15727 VP.n8509 a_400_38200# 0.06fF
C15728 VP.n8510 a_400_38200# 0.30fF
C15729 VP.n8511 a_400_38200# 0.10fF
C15730 VP.n8512 a_400_38200# 0.28fF
C15731 VP.n8513 a_400_38200# 0.15fF
C15732 VP.n8514 a_400_38200# 0.08fF
C15733 VP.n8515 a_400_38200# 0.14fF
C15734 VP.n8516 a_400_38200# 0.06fF
C15735 VP.n8517 a_400_38200# 0.06fF
C15736 VP.n8518 a_400_38200# 0.03fF
C15737 VP.n8519 a_400_38200# 0.05fF
C15738 VP.n8520 a_400_38200# 0.07fF
C15739 VP.n8521 a_400_38200# 0.19fF
C15740 VP.n8522 a_400_38200# 0.59fF
C15741 VP.n8523 a_400_38200# 0.34fF
C15742 VP.n8524 a_400_38200# 2.18fF
C15743 VP.t628 a_400_38200# 0.02fF
C15744 VP.n8525 a_400_38200# 0.24fF
C15745 VP.n8526 a_400_38200# 0.91fF
C15746 VP.n8527 a_400_38200# 0.05fF
C15747 VP.t721 a_400_38200# 0.02fF
C15748 VP.n8528 a_400_38200# 0.12fF
C15749 VP.n8529 a_400_38200# 0.14fF
C15750 VP.n8531 a_400_38200# 0.10fF
C15751 VP.n8532 a_400_38200# 0.10fF
C15752 VP.n8533 a_400_38200# 0.18fF
C15753 VP.n8534 a_400_38200# 0.09fF
C15754 VP.n8535 a_400_38200# 0.04fF
C15755 VP.n8536 a_400_38200# 0.26fF
C15756 VP.n8537 a_400_38200# 1.17fF
C15757 VP.n8538 a_400_38200# 0.06fF
C15758 VP.n8539 a_400_38200# 0.44fF
C15759 VP.n8540 a_400_38200# 0.13fF
C15760 VP.n8541 a_400_38200# 0.02fF
C15761 VP.n8542 a_400_38200# 1.81fF
C15762 VP.n8543 a_400_38200# 0.12fF
C15763 VP.t1162 a_400_38200# 0.02fF
C15764 VP.n8544 a_400_38200# 0.14fF
C15765 VP.t458 a_400_38200# 0.02fF
C15766 VP.n8546 a_400_38200# 0.24fF
C15767 VP.n8547 a_400_38200# 0.35fF
C15768 VP.n8548 a_400_38200# 0.60fF
C15769 VP.n8549 a_400_38200# 2.28fF
C15770 VP.t172 a_400_38200# 0.02fF
C15771 VP.n8550 a_400_38200# 0.24fF
C15772 VP.n8551 a_400_38200# 0.91fF
C15773 VP.n8552 a_400_38200# 0.05fF
C15774 VP.t274 a_400_38200# 0.02fF
C15775 VP.n8553 a_400_38200# 0.12fF
C15776 VP.n8554 a_400_38200# 0.14fF
C15777 VP.n8556 a_400_38200# 0.06fF
C15778 VP.n8557 a_400_38200# 0.09fF
C15779 VP.n8558 a_400_38200# 0.09fF
C15780 VP.n8559 a_400_38200# 1.45fF
C15781 VP.n8560 a_400_38200# 0.14fF
C15782 VP.n8561 a_400_38200# 0.07fF
C15783 VP.n8562 a_400_38200# 0.72fF
C15784 VP.n8563 a_400_38200# 1.81fF
C15785 VP.n8564 a_400_38200# 0.12fF
C15786 VP.t182 a_400_38200# 0.02fF
C15787 VP.n8565 a_400_38200# 0.14fF
C15788 VP.t695 a_400_38200# 0.02fF
C15789 VP.n8567 a_400_38200# 0.24fF
C15790 VP.n8568 a_400_38200# 0.35fF
C15791 VP.n8569 a_400_38200# 0.60fF
C15792 VP.n8570 a_400_38200# 2.30fF
C15793 VP.t421 a_400_38200# 0.02fF
C15794 VP.n8571 a_400_38200# 0.24fF
C15795 VP.n8572 a_400_38200# 0.91fF
C15796 VP.n8573 a_400_38200# 0.05fF
C15797 VP.t528 a_400_38200# 0.02fF
C15798 VP.n8574 a_400_38200# 0.12fF
C15799 VP.n8575 a_400_38200# 0.14fF
C15800 VP.n8577 a_400_38200# 0.06fF
C15801 VP.n8578 a_400_38200# 0.25fF
C15802 VP.n8579 a_400_38200# 0.45fF
C15803 VP.n8580 a_400_38200# 0.03fF
C15804 VP.n8581 a_400_38200# 0.05fF
C15805 VP.n8582 a_400_38200# 0.07fF
C15806 VP.n8583 a_400_38200# 0.06fF
C15807 VP.n8584 a_400_38200# 0.06fF
C15808 VP.n8585 a_400_38200# 0.19fF
C15809 VP.n8586 a_400_38200# 0.59fF
C15810 VP.n8587 a_400_38200# 0.34fF
C15811 VP.n8588 a_400_38200# 0.05fF
C15812 VP.n8589 a_400_38200# 0.30fF
C15813 VP.n8590 a_400_38200# 1.93fF
C15814 VP.n8591 a_400_38200# 0.12fF
C15815 VP.t1033 a_400_38200# 0.02fF
C15816 VP.n8592 a_400_38200# 0.14fF
C15817 VP.t325 a_400_38200# 0.02fF
C15818 VP.n8594 a_400_38200# 0.24fF
C15819 VP.n8595 a_400_38200# 0.35fF
C15820 VP.n8596 a_400_38200# 0.60fF
C15821 VP.n8597 a_400_38200# 2.04fF
C15822 VP.t1341 a_400_38200# 0.02fF
C15823 VP.n8598 a_400_38200# 0.24fF
C15824 VP.n8599 a_400_38200# 0.91fF
C15825 VP.n8600 a_400_38200# 0.05fF
C15826 VP.t51 a_400_38200# 0.02fF
C15827 VP.n8601 a_400_38200# 0.12fF
C15828 VP.n8602 a_400_38200# 0.14fF
C15829 VP.n8604 a_400_38200# 0.24fF
C15830 VP.t892 a_400_38200# 0.02fF
C15831 VP.n8605 a_400_38200# 0.36fF
C15832 VP.n8606 a_400_38200# 0.36fF
C15833 VP.n8607 a_400_38200# 0.67fF
C15834 VP.n8608 a_400_38200# 0.06fF
C15835 VP.n8609 a_400_38200# 0.09fF
C15836 VP.n8610 a_400_38200# 0.09fF
C15837 VP.n8611 a_400_38200# 1.45fF
C15838 VP.n8612 a_400_38200# 0.14fF
C15839 VP.n8613 a_400_38200# 0.07fF
C15840 VP.n8614 a_400_38200# 0.72fF
C15841 VP.n8615 a_400_38200# 1.81fF
C15842 VP.n8616 a_400_38200# 1.06fF
C15843 VP.n8617 a_400_38200# 0.24fF
C15844 VP.t1168 a_400_38200# 0.02fF
C15845 VP.n8618 a_400_38200# 0.35fF
C15846 VP.n8619 a_400_38200# 0.63fF
C15847 VP.n8620 a_400_38200# 0.40fF
C15848 VP.n8621 a_400_38200# 0.40fF
C15849 VP.n8622 a_400_38200# 0.12fF
C15850 VP.t585 a_400_38200# 0.02fF
C15851 VP.n8623 a_400_38200# 0.14fF
C15852 VP.t938 a_400_38200# 0.02fF
C15853 VP.n8625 a_400_38200# 0.12fF
C15854 VP.n8626 a_400_38200# 0.14fF
C15855 VP.n8628 a_400_38200# 1.93fF
C15856 VP.t716 a_400_38200# 0.02fF
C15857 VP.n8629 a_400_38200# 0.24fF
C15858 VP.n8630 a_400_38200# 0.35fF
C15859 VP.n8631 a_400_38200# 0.60fF
C15860 VP.n8632 a_400_38200# 0.12fF
C15861 VP.t118 a_400_38200# 0.02fF
C15862 VP.n8633 a_400_38200# 0.14fF
C15863 VP.n8635 a_400_38200# 0.07fF
C15864 VP.n8636 a_400_38200# 0.30fF
C15865 VP.n8637 a_400_38200# 0.06fF
C15866 VP.n8638 a_400_38200# 0.25fF
C15867 VP.n8639 a_400_38200# 0.45fF
C15868 VP.n8640 a_400_38200# 0.06fF
C15869 VP.n8641 a_400_38200# 0.06fF
C15870 VP.n8642 a_400_38200# 0.03fF
C15871 VP.n8643 a_400_38200# 0.05fF
C15872 VP.n8644 a_400_38200# 0.07fF
C15873 VP.n8645 a_400_38200# 0.19fF
C15874 VP.n8646 a_400_38200# 0.59fF
C15875 VP.n8647 a_400_38200# 0.34fF
C15876 VP.n8648 a_400_38200# 2.04fF
C15877 VP.t441 a_400_38200# 0.02fF
C15878 VP.n8649 a_400_38200# 0.24fF
C15879 VP.n8650 a_400_38200# 0.91fF
C15880 VP.n8651 a_400_38200# 0.05fF
C15881 VP.t493 a_400_38200# 0.02fF
C15882 VP.n8652 a_400_38200# 0.12fF
C15883 VP.n8653 a_400_38200# 0.14fF
C15884 VP.n8655 a_400_38200# 0.06fF
C15885 VP.n8656 a_400_38200# 0.09fF
C15886 VP.n8657 a_400_38200# 0.09fF
C15887 VP.n8658 a_400_38200# 1.45fF
C15888 VP.n8659 a_400_38200# 0.14fF
C15889 VP.n8660 a_400_38200# 0.07fF
C15890 VP.n8661 a_400_38200# 0.72fF
C15891 VP.n8662 a_400_38200# 1.81fF
C15892 VP.n8663 a_400_38200# 0.12fF
C15893 VP.t990 a_400_38200# 0.02fF
C15894 VP.n8664 a_400_38200# 0.14fF
C15895 VP.t270 a_400_38200# 0.02fF
C15896 VP.n8666 a_400_38200# 0.24fF
C15897 VP.n8667 a_400_38200# 0.35fF
C15898 VP.n8668 a_400_38200# 0.60fF
C15899 VP.n8669 a_400_38200# 2.30fF
C15900 VP.t1295 a_400_38200# 0.02fF
C15901 VP.n8670 a_400_38200# 0.24fF
C15902 VP.n8671 a_400_38200# 0.91fF
C15903 VP.n8672 a_400_38200# 0.05fF
C15904 VP.t1343 a_400_38200# 0.02fF
C15905 VP.n8673 a_400_38200# 0.12fF
C15906 VP.n8674 a_400_38200# 0.14fF
C15907 VP.n8676 a_400_38200# 1.93fF
C15908 VP.t1125 a_400_38200# 0.02fF
C15909 VP.n8677 a_400_38200# 0.24fF
C15910 VP.n8678 a_400_38200# 0.35fF
C15911 VP.n8679 a_400_38200# 0.60fF
C15912 VP.n8680 a_400_38200# 0.12fF
C15913 VP.t544 a_400_38200# 0.02fF
C15914 VP.n8681 a_400_38200# 0.14fF
C15915 VP.n8683 a_400_38200# 0.07fF
C15916 VP.n8684 a_400_38200# 0.30fF
C15917 VP.n8685 a_400_38200# 0.06fF
C15918 VP.n8686 a_400_38200# 0.25fF
C15919 VP.n8687 a_400_38200# 0.45fF
C15920 VP.n8688 a_400_38200# 0.06fF
C15921 VP.n8689 a_400_38200# 0.06fF
C15922 VP.n8690 a_400_38200# 0.03fF
C15923 VP.n8691 a_400_38200# 0.05fF
C15924 VP.n8692 a_400_38200# 0.07fF
C15925 VP.n8693 a_400_38200# 0.19fF
C15926 VP.n8694 a_400_38200# 0.59fF
C15927 VP.n8695 a_400_38200# 0.34fF
C15928 VP.n8696 a_400_38200# 2.04fF
C15929 VP.t849 a_400_38200# 0.02fF
C15930 VP.n8697 a_400_38200# 0.24fF
C15931 VP.n8698 a_400_38200# 0.91fF
C15932 VP.n8699 a_400_38200# 0.05fF
C15933 VP.t894 a_400_38200# 0.02fF
C15934 VP.n8700 a_400_38200# 0.12fF
C15935 VP.n8701 a_400_38200# 0.14fF
C15936 VP.n8703 a_400_38200# 0.06fF
C15937 VP.n8704 a_400_38200# 0.09fF
C15938 VP.n8705 a_400_38200# 0.09fF
C15939 VP.n8706 a_400_38200# 1.45fF
C15940 VP.n8707 a_400_38200# 0.14fF
C15941 VP.n8708 a_400_38200# 0.07fF
C15942 VP.n8709 a_400_38200# 0.72fF
C15943 VP.n8710 a_400_38200# 1.81fF
C15944 VP.n8711 a_400_38200# 0.12fF
C15945 VP.t67 a_400_38200# 0.02fF
C15946 VP.n8712 a_400_38200# 0.14fF
C15947 VP.t678 a_400_38200# 0.02fF
C15948 VP.n8714 a_400_38200# 0.24fF
C15949 VP.n8715 a_400_38200# 0.35fF
C15950 VP.n8716 a_400_38200# 0.60fF
C15951 VP.n8717 a_400_38200# 2.30fF
C15952 VP.t399 a_400_38200# 0.02fF
C15953 VP.n8718 a_400_38200# 0.24fF
C15954 VP.n8719 a_400_38200# 0.91fF
C15955 VP.n8720 a_400_38200# 0.05fF
C15956 VP.t511 a_400_38200# 0.02fF
C15957 VP.n8721 a_400_38200# 0.12fF
C15958 VP.n8722 a_400_38200# 0.14fF
C15959 VP.n8724 a_400_38200# 1.93fF
C15960 VP.t233 a_400_38200# 0.02fF
C15961 VP.n8725 a_400_38200# 0.24fF
C15962 VP.n8726 a_400_38200# 0.35fF
C15963 VP.n8727 a_400_38200# 0.60fF
C15964 VP.n8728 a_400_38200# 0.12fF
C15965 VP.t951 a_400_38200# 0.02fF
C15966 VP.n8729 a_400_38200# 0.14fF
C15967 VP.n8731 a_400_38200# 0.07fF
C15968 VP.n8732 a_400_38200# 0.30fF
C15969 VP.n8733 a_400_38200# 0.06fF
C15970 VP.n8734 a_400_38200# 0.25fF
C15971 VP.n8735 a_400_38200# 0.45fF
C15972 VP.n8736 a_400_38200# 0.06fF
C15973 VP.n8737 a_400_38200# 0.06fF
C15974 VP.n8738 a_400_38200# 0.03fF
C15975 VP.n8739 a_400_38200# 0.05fF
C15976 VP.n8740 a_400_38200# 0.07fF
C15977 VP.n8741 a_400_38200# 0.19fF
C15978 VP.n8742 a_400_38200# 0.59fF
C15979 VP.n8743 a_400_38200# 0.34fF
C15980 VP.n8744 a_400_38200# 2.04fF
C15981 VP.t1256 a_400_38200# 0.02fF
C15982 VP.n8745 a_400_38200# 0.24fF
C15983 VP.n8746 a_400_38200# 0.91fF
C15984 VP.n8747 a_400_38200# 0.05fF
C15985 VP.t29 a_400_38200# 0.02fF
C15986 VP.n8748 a_400_38200# 0.12fF
C15987 VP.n8749 a_400_38200# 0.14fF
C15988 VP.n8751 a_400_38200# 1.81fF
C15989 VP.t1088 a_400_38200# 0.02fF
C15990 VP.n8752 a_400_38200# 0.24fF
C15991 VP.n8753 a_400_38200# 0.35fF
C15992 VP.n8754 a_400_38200# 0.60fF
C15993 VP.n8755 a_400_38200# 0.12fF
C15994 VP.t505 a_400_38200# 0.02fF
C15995 VP.n8756 a_400_38200# 0.14fF
C15996 VP.n8758 a_400_38200# 0.03fF
C15997 VP.n8759 a_400_38200# 0.09fF
C15998 VP.n8760 a_400_38200# 0.09fF
C15999 VP.n8761 a_400_38200# 0.05fF
C16000 VP.n8762 a_400_38200# 0.11fF
C16001 VP.n8763 a_400_38200# 0.09fF
C16002 VP.n8764 a_400_38200# 0.02fF
C16003 VP.n8765 a_400_38200# 0.03fF
C16004 VP.n8766 a_400_38200# 0.11fF
C16005 VP.n8767 a_400_38200# 1.39fF
C16006 VP.n8768 a_400_38200# 0.06fF
C16007 VP.n8769 a_400_38200# 0.37fF
C16008 VP.n8770 a_400_38200# 2.30fF
C16009 VP.t812 a_400_38200# 0.02fF
C16010 VP.n8771 a_400_38200# 0.24fF
C16011 VP.n8772 a_400_38200# 0.91fF
C16012 VP.n8773 a_400_38200# 0.05fF
C16013 VP.t922 a_400_38200# 0.02fF
C16014 VP.n8774 a_400_38200# 0.12fF
C16015 VP.n8775 a_400_38200# 0.14fF
C16016 VP.n8777 a_400_38200# 0.88fF
C16017 VP.n8778 a_400_38200# 0.48fF
C16018 VP.n8779 a_400_38200# 0.88fF
C16019 VP.n8780 a_400_38200# 0.60fF
C16020 VP.n8781 a_400_38200# 2.33fF
C16021 VP.n8782 a_400_38200# 0.59fF
C16022 VP.n8783 a_400_38200# 0.02fF
C16023 VP.n8784 a_400_38200# 0.96fF
C16024 VP.t4 a_400_38200# 15.72fF
C16025 VP.n8785 a_400_38200# 15.42fF
C16026 VP.n8787 a_400_38200# 0.38fF
C16027 VP.n8788 a_400_38200# 0.23fF
C16028 VP.n8789 a_400_38200# 3.42fF
C16029 VP.n8790 a_400_38200# 0.21fF
C16030 VP.n8791 a_400_38200# 1.08fF
C16031 VP.n8792 a_400_38200# 0.03fF
C16032 VP.n8793 a_400_38200# 0.09fF
C16033 VP.n8794 a_400_38200# 0.43fF
C16034 VP.n8795 a_400_38200# 0.37fF
C16035 VP.t1339 a_400_38200# 0.02fF
C16036 VP.n8796 a_400_38200# 0.64fF
C16037 VP.n8797 a_400_38200# 0.60fF
C16038 VP.n8798 a_400_38200# 2.32fF
C16039 VP.n8799 a_400_38200# 4.93fF
C16040 VP.t1060 a_400_38200# 0.02fF
C16041 VP.n8800 a_400_38200# 1.19fF
C16042 VP.n8801 a_400_38200# 0.05fF
C16043 VP.t1153 a_400_38200# 0.02fF
C16044 VP.n8802 a_400_38200# 0.01fF
C16045 VP.n8803 a_400_38200# 0.26fF
C16046 VP.n8805 a_400_38200# 15.28fF
C16047 VP.t28 a_400_38200# 34.79fF
C16048 VP.t1174 a_400_38200# 0.02fF
C16049 VP.n8806 a_400_38200# 0.12fF
C16050 VP.n8807 a_400_38200# 0.14fF
C16051 VP.t1073 a_400_38200# 0.02fF
C16052 VP.n8809 a_400_38200# 0.24fF
C16053 VP.n8810 a_400_38200# 0.91fF
C16054 VP.n8811 a_400_38200# 0.05fF
C16055 VP.t5 a_400_38200# 0.02fF
C16056 VP.n8812 a_400_38200# 0.24fF
C16057 VP.n8813 a_400_38200# 0.35fF
C16058 VP.n8814 a_400_38200# 0.60fF
C16059 VP.n8815 a_400_38200# 0.02fF
C16060 VP.n8816 a_400_38200# 0.04fF
C16061 VP.n8817 a_400_38200# 0.06fF
C16062 VP.n8818 a_400_38200# 0.45fF
C16063 VP.n8819 a_400_38200# 0.10fF
C16064 VP.n8820 a_400_38200# 0.17fF
C16065 VP.n8821 a_400_38200# 0.10fF
C16066 VP.n8822 a_400_38200# 0.04fF
C16067 VP.n8823 a_400_38200# 0.09fF
C16068 VP.n8824 a_400_38200# 0.88fF
C16069 VP.n8825 a_400_38200# 0.10fF
C16070 VP.n8826 a_400_38200# 1.72fF
C16071 VP.n8827 a_400_38200# 1.93fF
C16072 VP.n8828 a_400_38200# 1.04fF
C16073 VP.n8829 a_400_38200# 0.05fF
C16074 VP.n8830 a_400_38200# 0.03fF
C16075 VP.n8831 a_400_38200# 0.06fF
C16076 VP.n8832 a_400_38200# 0.06fF
C16077 VP.n8833 a_400_38200# 0.06fF
C16078 VP.n8834 a_400_38200# 0.07fF
C16079 VP.n8835 a_400_38200# 0.03fF
C16080 VP.n8836 a_400_38200# 0.05fF
C16081 VP.n8837 a_400_38200# 0.07fF
C16082 VP.n8838 a_400_38200# 0.19fF
C16083 VP.n8839 a_400_38200# 0.60fF
C16084 VP.n8840 a_400_38200# 0.76fF
C16085 VP.n8841 a_400_38200# 0.40fF
C16086 VP.n8842 a_400_38200# 0.03fF
C16087 VP.n8843 a_400_38200# 0.01fF
C16088 VP.t898 a_400_38200# 0.02fF
C16089 VP.n8844 a_400_38200# 0.25fF
C16090 VP.t616 a_400_38200# 0.02fF
C16091 VP.n8845 a_400_38200# 0.95fF
C16092 VP.n8846 a_400_38200# 0.70fF
C16093 VP.n8847 a_400_38200# 1.92fF
C16094 VP.n8848 a_400_38200# 2.73fF
C16095 VP.n8849 a_400_38200# 0.19fF
C16096 VP.n8850 a_400_38200# 0.46fF
C16097 VP.n8851 a_400_38200# 0.11fF
C16098 VP.n8852 a_400_38200# 0.06fF
C16099 VP.n8853 a_400_38200# 0.01fF
C16100 VP.n8854 a_400_38200# 0.01fF
C16101 VP.n8855 a_400_38200# 0.04fF
C16102 VP.n8856 a_400_38200# 0.02fF
C16103 VP.n8857 a_400_38200# 0.07fF
C16104 VP.n8858 a_400_38200# 0.04fF
C16105 VP.n8859 a_400_38200# 0.14fF
C16106 VP.n8860 a_400_38200# 0.51fF
C16107 VP.n8861 a_400_38200# 1.62fF
C16108 VP.t1032 a_400_38200# 0.02fF
C16109 VP.n8862 a_400_38200# 0.24fF
C16110 VP.n8863 a_400_38200# 0.35fF
C16111 VP.n8864 a_400_38200# 0.60fF
C16112 VP.n8865 a_400_38200# 0.12fF
C16113 VP.t445 a_400_38200# 0.02fF
C16114 VP.n8866 a_400_38200# 0.14fF
C16115 VP.n8868 a_400_38200# 0.04fF
C16116 VP.n8869 a_400_38200# 0.02fF
C16117 VP.n8870 a_400_38200# 0.06fF
C16118 VP.n8871 a_400_38200# 0.30fF
C16119 VP.n8872 a_400_38200# 0.06fF
C16120 VP.n8873 a_400_38200# 0.33fF
C16121 VP.n8874 a_400_38200# 0.03fF
C16122 VP.n8875 a_400_38200# 0.15fF
C16123 VP.n8876 a_400_38200# 0.08fF
C16124 VP.n8877 a_400_38200# 0.14fF
C16125 VP.n8878 a_400_38200# 0.03fF
C16126 VP.n8879 a_400_38200# 0.06fF
C16127 VP.n8880 a_400_38200# 0.06fF
C16128 VP.n8881 a_400_38200# 0.06fF
C16129 VP.n8882 a_400_38200# 0.06fF
C16130 VP.n8883 a_400_38200# 0.03fF
C16131 VP.n8884 a_400_38200# 0.05fF
C16132 VP.n8885 a_400_38200# 0.07fF
C16133 VP.n8886 a_400_38200# 0.19fF
C16134 VP.n8887 a_400_38200# 0.59fF
C16135 VP.n8888 a_400_38200# 0.34fF
C16136 VP.n8889 a_400_38200# 1.94fF
C16137 VP.t154 a_400_38200# 0.02fF
C16138 VP.n8890 a_400_38200# 0.24fF
C16139 VP.n8891 a_400_38200# 0.91fF
C16140 VP.n8892 a_400_38200# 0.05fF
C16141 VP.t487 a_400_38200# 0.02fF
C16142 VP.n8893 a_400_38200# 0.12fF
C16143 VP.n8894 a_400_38200# 0.14fF
C16144 VP.n8896 a_400_38200# 0.19fF
C16145 VP.n8897 a_400_38200# 0.10fF
C16146 VP.n8898 a_400_38200# 0.10fF
C16147 VP.n8899 a_400_38200# 0.18fF
C16148 VP.n8900 a_400_38200# 0.09fF
C16149 VP.n8901 a_400_38200# 0.04fF
C16150 VP.n8902 a_400_38200# 0.19fF
C16151 VP.n8903 a_400_38200# 0.26fF
C16152 VP.n8904 a_400_38200# 1.17fF
C16153 VP.n8905 a_400_38200# 0.06fF
C16154 VP.n8906 a_400_38200# 0.44fF
C16155 VP.n8907 a_400_38200# 0.13fF
C16156 VP.n8908 a_400_38200# 0.02fF
C16157 VP.n8909 a_400_38200# 1.81fF
C16158 VP.n8910 a_400_38200# 0.12fF
C16159 VP.t1299 a_400_38200# 0.02fF
C16160 VP.n8911 a_400_38200# 0.14fF
C16161 VP.t584 a_400_38200# 0.02fF
C16162 VP.n8913 a_400_38200# 0.24fF
C16163 VP.n8914 a_400_38200# 0.35fF
C16164 VP.n8915 a_400_38200# 0.60fF
C16165 VP.n8916 a_400_38200# 3.18fF
C16166 VP.n8917 a_400_38200# 2.06fF
C16167 VP.n8918 a_400_38200# 1.98fF
C16168 VP.t1010 a_400_38200# 0.02fF
C16169 VP.n8919 a_400_38200# 0.24fF
C16170 VP.n8920 a_400_38200# 0.91fF
C16171 VP.n8921 a_400_38200# 0.05fF
C16172 VP.t1337 a_400_38200# 0.02fF
C16173 VP.n8922 a_400_38200# 0.12fF
C16174 VP.n8923 a_400_38200# 0.14fF
C16175 VP.n8925 a_400_38200# 0.16fF
C16176 VP.n8926 a_400_38200# 0.19fF
C16177 VP.n8927 a_400_38200# 0.09fF
C16178 VP.n8928 a_400_38200# 0.04fF
C16179 VP.n8929 a_400_38200# 0.14fF
C16180 VP.n8930 a_400_38200# 0.64fF
C16181 VP.n8931 a_400_38200# 1.32fF
C16182 VP.n8932 a_400_38200# 1.81fF
C16183 VP.n8933 a_400_38200# 0.12fF
C16184 VP.t241 a_400_38200# 0.02fF
C16185 VP.n8934 a_400_38200# 0.14fF
C16186 VP.t838 a_400_38200# 0.02fF
C16187 VP.n8936 a_400_38200# 0.24fF
C16188 VP.n8937 a_400_38200# 0.35fF
C16189 VP.n8938 a_400_38200# 0.60fF
C16190 VP.n8939 a_400_38200# 2.97fF
C16191 VP.n8940 a_400_38200# 2.27fF
C16192 VP.n8941 a_400_38200# 2.00fF
C16193 VP.t1266 a_400_38200# 0.02fF
C16194 VP.n8942 a_400_38200# 0.24fF
C16195 VP.n8943 a_400_38200# 0.91fF
C16196 VP.n8944 a_400_38200# 0.05fF
C16197 VP.t887 a_400_38200# 0.02fF
C16198 VP.n8945 a_400_38200# 0.12fF
C16199 VP.n8946 a_400_38200# 0.14fF
C16200 VP.n8948 a_400_38200# 0.24fF
C16201 VP.t371 a_400_38200# 0.02fF
C16202 VP.n8949 a_400_38200# 0.36fF
C16203 VP.n8950 a_400_38200# 0.36fF
C16204 VP.n8951 a_400_38200# 0.67fF
C16205 VP.n8952 a_400_38200# 0.16fF
C16206 VP.n8953 a_400_38200# 0.19fF
C16207 VP.n8954 a_400_38200# 0.09fF
C16208 VP.n8955 a_400_38200# 0.04fF
C16209 VP.n8956 a_400_38200# 0.14fF
C16210 VP.n8957 a_400_38200# 0.64fF
C16211 VP.n8958 a_400_38200# 1.32fF
C16212 VP.n8959 a_400_38200# 1.81fF
C16213 VP.n8960 a_400_38200# 2.97fF
C16214 VP.n8961 a_400_38200# 2.27fF
C16215 VP.n8962 a_400_38200# 0.75fF
C16216 VP.n8963 a_400_38200# 0.24fF
C16217 VP.t1243 a_400_38200# 0.02fF
C16218 VP.n8964 a_400_38200# 0.35fF
C16219 VP.n8965 a_400_38200# 0.63fF
C16220 VP.n8966 a_400_38200# 0.40fF
C16221 VP.n8967 a_400_38200# 0.40fF
C16222 VP.n8968 a_400_38200# 0.12fF
C16223 VP.t655 a_400_38200# 0.02fF
C16224 VP.n8969 a_400_38200# 0.14fF
C16225 VP.t755 a_400_38200# 0.02fF
C16226 VP.n8971 a_400_38200# 0.12fF
C16227 VP.n8972 a_400_38200# 0.14fF
C16228 VP.n8974 a_400_38200# 0.16fF
C16229 VP.n8975 a_400_38200# 0.19fF
C16230 VP.n8976 a_400_38200# 0.09fF
C16231 VP.n8977 a_400_38200# 0.04fF
C16232 VP.n8978 a_400_38200# 0.14fF
C16233 VP.n8979 a_400_38200# 0.64fF
C16234 VP.n8980 a_400_38200# 1.32fF
C16235 VP.n8981 a_400_38200# 1.81fF
C16236 VP.n8982 a_400_38200# 0.12fF
C16237 VP.t1062 a_400_38200# 0.02fF
C16238 VP.n8983 a_400_38200# 0.14fF
C16239 VP.t350 a_400_38200# 0.02fF
C16240 VP.n8985 a_400_38200# 0.24fF
C16241 VP.n8986 a_400_38200# 0.35fF
C16242 VP.n8987 a_400_38200# 0.60fF
C16243 VP.n8988 a_400_38200# 2.97fF
C16244 VP.n8989 a_400_38200# 2.27fF
C16245 VP.n8990 a_400_38200# 2.00fF
C16246 VP.t781 a_400_38200# 0.02fF
C16247 VP.n8991 a_400_38200# 0.24fF
C16248 VP.n8992 a_400_38200# 0.91fF
C16249 VP.n8993 a_400_38200# 0.05fF
C16250 VP.t1148 a_400_38200# 0.02fF
C16251 VP.n8994 a_400_38200# 0.12fF
C16252 VP.n8995 a_400_38200# 0.14fF
C16253 VP.n8997 a_400_38200# 0.16fF
C16254 VP.n8998 a_400_38200# 0.19fF
C16255 VP.n8999 a_400_38200# 0.09fF
C16256 VP.n9000 a_400_38200# 0.04fF
C16257 VP.n9001 a_400_38200# 0.14fF
C16258 VP.n9002 a_400_38200# 0.64fF
C16259 VP.n9003 a_400_38200# 1.32fF
C16260 VP.n9004 a_400_38200# 1.81fF
C16261 VP.n9005 a_400_38200# 0.12fF
C16262 VP.t226 a_400_38200# 0.02fF
C16263 VP.n9006 a_400_38200# 0.14fF
C16264 VP.t751 a_400_38200# 0.02fF
C16265 VP.n9008 a_400_38200# 0.24fF
C16266 VP.n9009 a_400_38200# 0.35fF
C16267 VP.n9010 a_400_38200# 0.60fF
C16268 VP.n9011 a_400_38200# 2.97fF
C16269 VP.n9012 a_400_38200# 2.27fF
C16270 VP.n9013 a_400_38200# 2.00fF
C16271 VP.t1176 a_400_38200# 0.02fF
C16272 VP.n9014 a_400_38200# 0.24fF
C16273 VP.n9015 a_400_38200# 0.91fF
C16274 VP.n9016 a_400_38200# 0.05fF
C16275 VP.t257 a_400_38200# 0.02fF
C16276 VP.n9017 a_400_38200# 0.12fF
C16277 VP.n9018 a_400_38200# 0.14fF
C16278 VP.n9020 a_400_38200# 0.03fF
C16279 VP.n9021 a_400_38200# 0.19fF
C16280 VP.n9022 a_400_38200# 0.24fF
C16281 VP.n9023 a_400_38200# 0.98fF
C16282 VP.n9024 a_400_38200# 0.12fF
C16283 VP.n9025 a_400_38200# 0.19fF
C16284 VP.n9026 a_400_38200# 0.09fF
C16285 VP.n9027 a_400_38200# 0.18fF
C16286 VP.n9028 a_400_38200# 0.09fF
C16287 VP.n9029 a_400_38200# 0.08fF
C16288 VP.n9030 a_400_38200# 0.39fF
C16289 VP.n9031 a_400_38200# 0.24fF
C16290 VP.n9032 a_400_38200# 0.13fF
C16291 VP.n9033 a_400_38200# 0.02fF
C16292 VP.n9034 a_400_38200# 1.81fF
C16293 VP.n9035 a_400_38200# 0.12fF
C16294 VP.t639 a_400_38200# 0.02fF
C16295 VP.n9036 a_400_38200# 0.14fF
C16296 VP.t1223 a_400_38200# 0.02fF
C16297 VP.n9038 a_400_38200# 0.24fF
C16298 VP.n9039 a_400_38200# 0.35fF
C16299 VP.n9040 a_400_38200# 0.60fF
C16300 VP.n9041 a_400_38200# 3.17fF
C16301 VP.n9042 a_400_38200# 2.27fF
C16302 VP.n9043 a_400_38200# 1.98fF
C16303 VP.t352 a_400_38200# 0.02fF
C16304 VP.n9044 a_400_38200# 0.24fF
C16305 VP.n9045 a_400_38200# 0.91fF
C16306 VP.n9046 a_400_38200# 0.05fF
C16307 VP.t666 a_400_38200# 0.02fF
C16308 VP.n9047 a_400_38200# 0.12fF
C16309 VP.n9048 a_400_38200# 0.14fF
C16310 VP.n9050 a_400_38200# 15.28fF
C16311 VP.n9051 a_400_38200# 0.06fF
C16312 VP.n9052 a_400_38200# 0.06fF
C16313 VP.n9053 a_400_38200# 0.03fF
C16314 VP.n9054 a_400_38200# 0.10fF
C16315 VP.n9055 a_400_38200# 0.17fF
C16316 VP.n9056 a_400_38200# 0.10fF
C16317 VP.n9057 a_400_38200# 0.13fF
C16318 VP.n9058 a_400_38200# 0.02fF
C16319 VP.n9059 a_400_38200# 0.04fF
C16320 VP.n9060 a_400_38200# 0.06fF
C16321 VP.n9061 a_400_38200# 0.09fF
C16322 VP.n9062 a_400_38200# 0.10fF
C16323 VP.n9063 a_400_38200# 0.05fF
C16324 VP.n9064 a_400_38200# 0.19fF
C16325 VP.n9065 a_400_38200# 0.16fF
C16326 VP.n9066 a_400_38200# 0.04fF
C16327 VP.n9067 a_400_38200# 0.05fF
C16328 VP.n9068 a_400_38200# 0.04fF
C16329 VP.n9069 a_400_38200# 0.12fF
C16330 VP.n9070 a_400_38200# 0.09fF
C16331 VP.n9071 a_400_38200# 0.14fF
C16332 VP.n9072 a_400_38200# 0.56fF
C16333 VP.n9073 a_400_38200# 0.10fF
C16334 VP.n9074 a_400_38200# 1.93fF
C16335 VP.n9075 a_400_38200# 0.12fF
C16336 VP.t1096 a_400_38200# 0.02fF
C16337 VP.n9076 a_400_38200# 0.14fF
C16338 VP.t387 a_400_38200# 0.02fF
C16339 VP.n9078 a_400_38200# 0.24fF
C16340 VP.n9079 a_400_38200# 0.35fF
C16341 VP.n9080 a_400_38200# 0.60fF
C16342 VP.n9081 a_400_38200# 2.23fF
C16343 VP.n9082 a_400_38200# 0.18fF
C16344 VP.n9083 a_400_38200# 0.45fF
C16345 VP.n9084 a_400_38200# 0.06fF
C16346 VP.n9085 a_400_38200# 0.01fF
C16347 VP.n9086 a_400_38200# 0.01fF
C16348 VP.n9087 a_400_38200# 0.04fF
C16349 VP.n9088 a_400_38200# 0.02fF
C16350 VP.n9089 a_400_38200# 0.07fF
C16351 VP.n9090 a_400_38200# 0.04fF
C16352 VP.n9091 a_400_38200# 0.14fF
C16353 VP.n9092 a_400_38200# 0.45fF
C16354 VP.n9093 a_400_38200# 1.46fF
C16355 VP.n9094 a_400_38200# 1.78fF
C16356 VP.t1203 a_400_38200# 0.02fF
C16357 VP.n9095 a_400_38200# 0.12fF
C16358 VP.n9096 a_400_38200# 0.14fF
C16359 VP.t822 a_400_38200# 0.02fF
C16360 VP.n9098 a_400_38200# 0.24fF
C16361 VP.n9099 a_400_38200# 0.91fF
C16362 VP.n9100 a_400_38200# 0.05fF
C16363 VP.n9101 a_400_38200# 1.93fF
C16364 VP.n9102 a_400_38200# 2.23fF
C16365 VP.n9103 a_400_38200# 0.18fF
C16366 VP.n9104 a_400_38200# 0.45fF
C16367 VP.n9105 a_400_38200# 0.06fF
C16368 VP.n9106 a_400_38200# 0.01fF
C16369 VP.n9107 a_400_38200# 0.01fF
C16370 VP.n9108 a_400_38200# 0.04fF
C16371 VP.n9109 a_400_38200# 0.02fF
C16372 VP.n9110 a_400_38200# 0.07fF
C16373 VP.n9111 a_400_38200# 0.04fF
C16374 VP.n9112 a_400_38200# 0.14fF
C16375 VP.n9113 a_400_38200# 0.45fF
C16376 VP.n9114 a_400_38200# 1.46fF
C16377 VP.t796 a_400_38200# 0.02fF
C16378 VP.n9115 a_400_38200# 0.24fF
C16379 VP.n9116 a_400_38200# 0.35fF
C16380 VP.n9117 a_400_38200# 0.60fF
C16381 VP.n9118 a_400_38200# 0.12fF
C16382 VP.t208 a_400_38200# 0.02fF
C16383 VP.n9119 a_400_38200# 0.14fF
C16384 VP.n9121 a_400_38200# 0.10fF
C16385 VP.n9122 a_400_38200# 0.17fF
C16386 VP.n9123 a_400_38200# 0.06fF
C16387 VP.n9124 a_400_38200# 0.06fF
C16388 VP.n9125 a_400_38200# 0.03fF
C16389 VP.n9126 a_400_38200# 0.10fF
C16390 VP.n9127 a_400_38200# 0.13fF
C16391 VP.n9128 a_400_38200# 0.13fF
C16392 VP.n9129 a_400_38200# 0.04fF
C16393 VP.n9130 a_400_38200# 0.05fF
C16394 VP.n9131 a_400_38200# 0.04fF
C16395 VP.n9132 a_400_38200# 0.09fF
C16396 VP.n9133 a_400_38200# 0.09fF
C16397 VP.n9134 a_400_38200# 0.05fF
C16398 VP.n9135 a_400_38200# 0.19fF
C16399 VP.n9136 a_400_38200# 0.12fF
C16400 VP.n9137 a_400_38200# 0.09fF
C16401 VP.n9138 a_400_38200# 0.14fF
C16402 VP.n9139 a_400_38200# 0.04fF
C16403 VP.n9140 a_400_38200# 0.02fF
C16404 VP.n9141 a_400_38200# 0.06fF
C16405 VP.n9142 a_400_38200# 0.56fF
C16406 VP.n9143 a_400_38200# 0.10fF
C16407 VP.n9144 a_400_38200# 1.78fF
C16408 VP.t301 a_400_38200# 0.02fF
C16409 VP.n9145 a_400_38200# 0.12fF
C16410 VP.n9146 a_400_38200# 0.14fF
C16411 VP.t1226 a_400_38200# 0.02fF
C16412 VP.n9148 a_400_38200# 0.24fF
C16413 VP.n9149 a_400_38200# 0.91fF
C16414 VP.n9150 a_400_38200# 0.05fF
C16415 VP.n9151 a_400_38200# 1.93fF
C16416 VP.n9152 a_400_38200# 2.23fF
C16417 VP.n9153 a_400_38200# 0.18fF
C16418 VP.n9154 a_400_38200# 0.45fF
C16419 VP.n9155 a_400_38200# 0.06fF
C16420 VP.n9156 a_400_38200# 0.01fF
C16421 VP.n9157 a_400_38200# 0.01fF
C16422 VP.n9158 a_400_38200# 0.04fF
C16423 VP.n9159 a_400_38200# 0.02fF
C16424 VP.n9160 a_400_38200# 0.07fF
C16425 VP.n9161 a_400_38200# 0.04fF
C16426 VP.n9162 a_400_38200# 0.14fF
C16427 VP.n9163 a_400_38200# 0.45fF
C16428 VP.n9164 a_400_38200# 1.46fF
C16429 VP.t1200 a_400_38200# 0.02fF
C16430 VP.n9165 a_400_38200# 0.24fF
C16431 VP.n9166 a_400_38200# 0.35fF
C16432 VP.n9167 a_400_38200# 0.60fF
C16433 VP.n9168 a_400_38200# 0.12fF
C16434 VP.t614 a_400_38200# 0.02fF
C16435 VP.n9169 a_400_38200# 0.14fF
C16436 VP.n9171 a_400_38200# 0.10fF
C16437 VP.n9172 a_400_38200# 0.17fF
C16438 VP.n9173 a_400_38200# 0.06fF
C16439 VP.n9174 a_400_38200# 0.06fF
C16440 VP.n9175 a_400_38200# 0.03fF
C16441 VP.n9176 a_400_38200# 0.10fF
C16442 VP.n9177 a_400_38200# 0.13fF
C16443 VP.n9178 a_400_38200# 0.13fF
C16444 VP.n9179 a_400_38200# 0.04fF
C16445 VP.n9180 a_400_38200# 0.05fF
C16446 VP.n9181 a_400_38200# 0.04fF
C16447 VP.n9182 a_400_38200# 0.09fF
C16448 VP.n9183 a_400_38200# 0.09fF
C16449 VP.n9184 a_400_38200# 0.05fF
C16450 VP.n9185 a_400_38200# 0.19fF
C16451 VP.n9186 a_400_38200# 0.12fF
C16452 VP.n9187 a_400_38200# 0.09fF
C16453 VP.n9188 a_400_38200# 0.14fF
C16454 VP.n9189 a_400_38200# 0.04fF
C16455 VP.n9190 a_400_38200# 0.02fF
C16456 VP.n9191 a_400_38200# 0.06fF
C16457 VP.n9192 a_400_38200# 0.56fF
C16458 VP.n9193 a_400_38200# 0.10fF
C16459 VP.n9194 a_400_38200# 1.78fF
C16460 VP.t700 a_400_38200# 0.02fF
C16461 VP.n9195 a_400_38200# 0.12fF
C16462 VP.n9196 a_400_38200# 0.14fF
C16463 VP.t332 a_400_38200# 0.02fF
C16464 VP.n9198 a_400_38200# 0.24fF
C16465 VP.n9199 a_400_38200# 0.91fF
C16466 VP.n9200 a_400_38200# 0.05fF
C16467 VP.n9201 a_400_38200# 1.93fF
C16468 VP.n9202 a_400_38200# 2.23fF
C16469 VP.n9203 a_400_38200# 0.18fF
C16470 VP.n9204 a_400_38200# 0.45fF
C16471 VP.n9205 a_400_38200# 0.06fF
C16472 VP.n9206 a_400_38200# 0.01fF
C16473 VP.n9207 a_400_38200# 0.01fF
C16474 VP.n9208 a_400_38200# 0.04fF
C16475 VP.n9209 a_400_38200# 0.02fF
C16476 VP.n9210 a_400_38200# 0.07fF
C16477 VP.n9211 a_400_38200# 0.04fF
C16478 VP.n9212 a_400_38200# 0.14fF
C16479 VP.n9213 a_400_38200# 0.45fF
C16480 VP.n9214 a_400_38200# 1.46fF
C16481 VP.t368 a_400_38200# 0.02fF
C16482 VP.n9215 a_400_38200# 0.24fF
C16483 VP.n9216 a_400_38200# 0.35fF
C16484 VP.n9217 a_400_38200# 0.60fF
C16485 VP.n9218 a_400_38200# 0.12fF
C16486 VP.t1082 a_400_38200# 0.02fF
C16487 VP.n9219 a_400_38200# 0.14fF
C16488 VP.n9221 a_400_38200# 0.10fF
C16489 VP.n9222 a_400_38200# 0.17fF
C16490 VP.n9223 a_400_38200# 0.06fF
C16491 VP.n9224 a_400_38200# 0.06fF
C16492 VP.n9225 a_400_38200# 0.03fF
C16493 VP.n9226 a_400_38200# 0.10fF
C16494 VP.n9227 a_400_38200# 0.13fF
C16495 VP.n9228 a_400_38200# 0.13fF
C16496 VP.n9229 a_400_38200# 0.04fF
C16497 VP.n9230 a_400_38200# 0.05fF
C16498 VP.n9231 a_400_38200# 0.04fF
C16499 VP.n9232 a_400_38200# 0.09fF
C16500 VP.n9233 a_400_38200# 0.09fF
C16501 VP.n9234 a_400_38200# 0.05fF
C16502 VP.n9235 a_400_38200# 0.19fF
C16503 VP.n9236 a_400_38200# 0.12fF
C16504 VP.n9237 a_400_38200# 0.09fF
C16505 VP.n9238 a_400_38200# 0.14fF
C16506 VP.n9239 a_400_38200# 0.04fF
C16507 VP.n9240 a_400_38200# 0.02fF
C16508 VP.n9241 a_400_38200# 0.06fF
C16509 VP.n9242 a_400_38200# 0.56fF
C16510 VP.n9243 a_400_38200# 0.10fF
C16511 VP.n9244 a_400_38200# 1.78fF
C16512 VP.t1110 a_400_38200# 0.02fF
C16513 VP.n9245 a_400_38200# 0.12fF
C16514 VP.n9246 a_400_38200# 0.14fF
C16515 VP.t800 a_400_38200# 0.02fF
C16516 VP.n9248 a_400_38200# 0.24fF
C16517 VP.n9249 a_400_38200# 0.91fF
C16518 VP.n9250 a_400_38200# 0.05fF
C16519 VP.n9251 a_400_38200# 1.92fF
C16520 VP.n9252 a_400_38200# 2.51fF
C16521 VP.t157 a_400_38200# 0.02fF
C16522 VP.n9253 a_400_38200# 0.24fF
C16523 VP.n9254 a_400_38200# 0.35fF
C16524 VP.n9255 a_400_38200# 0.60fF
C16525 VP.n9256 a_400_38200# 0.12fF
C16526 VP.t876 a_400_38200# 0.02fF
C16527 VP.n9257 a_400_38200# 0.14fF
C16528 VP.n9259 a_400_38200# 0.06fF
C16529 VP.n9260 a_400_38200# 0.30fF
C16530 VP.n9261 a_400_38200# 0.20fF
C16531 VP.n9262 a_400_38200# 0.09fF
C16532 VP.n9263 a_400_38200# 0.26fF
C16533 VP.n9264 a_400_38200# 0.22fF
C16534 VP.n9265 a_400_38200# 0.19fF
C16535 VP.n9266 a_400_38200# 0.05fF
C16536 VP.n9267 a_400_38200# 0.13fF
C16537 VP.n9268 a_400_38200# 0.09fF
C16538 VP.n9269 a_400_38200# 0.09fF
C16539 VP.n9270 a_400_38200# 0.07fF
C16540 VP.n9271 a_400_38200# 0.71fF
C16541 VP.n9272 a_400_38200# 0.24fF
C16542 VP.n9273 a_400_38200# 1.88fF
C16543 VP.t220 a_400_38200# 0.02fF
C16544 VP.n9274 a_400_38200# 0.12fF
C16545 VP.n9275 a_400_38200# 0.14fF
C16546 VP.t595 a_400_38200# 0.02fF
C16547 VP.n9277 a_400_38200# 0.24fF
C16548 VP.n9278 a_400_38200# 0.91fF
C16549 VP.n9279 a_400_38200# 0.05fF
C16550 VP.t207 a_400_38200# 35.17fF
C16551 VP.t180 a_400_38200# 0.02fF
C16552 VP.n9280 a_400_38200# 1.21fF
C16553 VP.n9281 a_400_38200# 0.25fF
C16554 VP.n9282 a_400_38200# 26.29fF
C16555 VP.n9283 a_400_38200# 26.29fF
C16556 VP.n9284 a_400_38200# 0.76fF
C16557 VP.n9285 a_400_38200# 0.27fF
C16558 VP.n9286 a_400_38200# 0.59fF
C16559 VP.n9287 a_400_38200# 0.10fF
C16560 VP.n9288 a_400_38200# 3.02fF
C16561 VP.t156 a_400_38200# 15.72fF
C16562 VP.n9289 a_400_38200# 1.15fF
C16563 VP.n9291 a_400_38200# 13.70fF
C16564 VP.n9293 a_400_38200# 1.99fF
C16565 VP.n9294 a_400_38200# 4.39fF
C16566 VP.n9295 a_400_38200# 0.03fF
C16567 VP.n9296 a_400_38200# 0.05fF
C16568 VP.n9297 a_400_38200# 0.07fF
C16569 VP.n9298 a_400_38200# 0.03fF
C16570 VP.n9299 a_400_38200# 0.06fF
C16571 VP.n9300 a_400_38200# 0.06fF
C16572 VP.n9301 a_400_38200# 0.06fF
C16573 VP.n9302 a_400_38200# 0.07fF
C16574 VP.n9303 a_400_38200# 0.57fF
C16575 VP.n9304 a_400_38200# 1.88fF
C16576 VP.n9305 a_400_38200# 0.91fF
C16577 VP.n9306 a_400_38200# 2.65fF
C16578 VP.n9307 a_400_38200# 0.07fF
C16579 VP.n9308 a_400_38200# 0.14fF
C16580 VP.n9309 a_400_38200# 0.13fF
C16581 VP.n9310 a_400_38200# 0.07fF
C16582 VP.n9311 a_400_38200# 0.22fF
C16583 VP.n9312 a_400_38200# 0.06fF
C16584 VP.n9313 a_400_38200# 0.05fF
C16585 VP.n9314 a_400_38200# 0.03fF
C16586 VP.n9315 a_400_38200# 0.08fF
C16587 VP.n9316 a_400_38200# 0.63fF
C16588 VP.n9317 a_400_38200# 0.72fF
C16589 VP.n9318 a_400_38200# 0.02fF
C16590 VP.n9319 a_400_38200# 0.11fF
C16591 VP.n9320 a_400_38200# 0.29fF
C16592 VP.n9321 a_400_38200# 0.12fF
C16593 VP.t1063 a_400_38200# 0.02fF
C16594 VP.n9322 a_400_38200# 0.14fF
C16595 VP.n9324 a_400_38200# 0.10fF
C16596 VP.n9325 a_400_38200# 0.10fF
C16597 VP.n9326 a_400_38200# 0.18fF
C16598 VP.n9327 a_400_38200# 0.09fF
C16599 VP.n9328 a_400_38200# 0.04fF
C16600 VP.n9329 a_400_38200# 0.26fF
C16601 VP.n9330 a_400_38200# 1.17fF
C16602 VP.n9331 a_400_38200# 0.06fF
C16603 VP.n9332 a_400_38200# 0.44fF
C16604 VP.n9333 a_400_38200# 0.13fF
C16605 VP.n9334 a_400_38200# 0.02fF
C16606 VP.n9335 a_400_38200# 1.81fF
C16607 VP.n9336 a_400_38200# 0.12fF
C16608 VP.t617 a_400_38200# 0.02fF
C16609 VP.n9337 a_400_38200# 0.14fF
C16610 VP.t1056 a_400_38200# 0.02fF
C16611 VP.n9339 a_400_38200# 0.24fF
C16612 VP.n9340 a_400_38200# 0.35fF
C16613 VP.n9341 a_400_38200# 0.60fF
C16614 VP.n9342 a_400_38200# 3.09fF
C16615 VP.n9343 a_400_38200# 2.28fF
C16616 VP.t776 a_400_38200# 0.02fF
C16617 VP.n9344 a_400_38200# 0.24fF
C16618 VP.n9345 a_400_38200# 0.91fF
C16619 VP.n9346 a_400_38200# 0.05fF
C16620 VP.t1016 a_400_38200# 0.02fF
C16621 VP.n9347 a_400_38200# 0.12fF
C16622 VP.n9348 a_400_38200# 0.14fF
C16623 VP.n9350 a_400_38200# 0.06fF
C16624 VP.n9351 a_400_38200# 0.09fF
C16625 VP.n9352 a_400_38200# 0.09fF
C16626 VP.n9353 a_400_38200# 1.45fF
C16627 VP.n9354 a_400_38200# 0.14fF
C16628 VP.n9355 a_400_38200# 0.07fF
C16629 VP.n9356 a_400_38200# 0.72fF
C16630 VP.n9357 a_400_38200# 1.81fF
C16631 VP.n9358 a_400_38200# 0.12fF
C16632 VP.t152 a_400_38200# 0.02fF
C16633 VP.n9359 a_400_38200# 0.14fF
C16634 VP.t609 a_400_38200# 0.02fF
C16635 VP.n9361 a_400_38200# 0.24fF
C16636 VP.n9362 a_400_38200# 0.35fF
C16637 VP.n9363 a_400_38200# 0.60fF
C16638 VP.n9364 a_400_38200# 2.97fF
C16639 VP.n9365 a_400_38200# 2.30fF
C16640 VP.t326 a_400_38200# 0.02fF
C16641 VP.n9366 a_400_38200# 0.24fF
C16642 VP.n9367 a_400_38200# 0.91fF
C16643 VP.n9368 a_400_38200# 0.05fF
C16644 VP.t571 a_400_38200# 0.02fF
C16645 VP.n9369 a_400_38200# 0.12fF
C16646 VP.n9370 a_400_38200# 0.14fF
C16647 VP.n9372 a_400_38200# 0.06fF
C16648 VP.n9373 a_400_38200# 0.25fF
C16649 VP.n9374 a_400_38200# 0.45fF
C16650 VP.n9375 a_400_38200# 0.03fF
C16651 VP.n9376 a_400_38200# 0.05fF
C16652 VP.n9377 a_400_38200# 0.07fF
C16653 VP.n9378 a_400_38200# 0.06fF
C16654 VP.n9379 a_400_38200# 0.06fF
C16655 VP.n9380 a_400_38200# 0.19fF
C16656 VP.n9381 a_400_38200# 0.59fF
C16657 VP.n9382 a_400_38200# 0.34fF
C16658 VP.n9383 a_400_38200# 0.09fF
C16659 VP.n9384 a_400_38200# 0.05fF
C16660 VP.n9385 a_400_38200# 0.30fF
C16661 VP.n9386 a_400_38200# 1.93fF
C16662 VP.n9387 a_400_38200# 0.12fF
C16663 VP.t482 a_400_38200# 0.02fF
C16664 VP.n9388 a_400_38200# 0.14fF
C16665 VP.t853 a_400_38200# 0.02fF
C16666 VP.n9390 a_400_38200# 0.24fF
C16667 VP.n9391 a_400_38200# 0.35fF
C16668 VP.n9392 a_400_38200# 0.60fF
C16669 VP.n9393 a_400_38200# 2.23fF
C16670 VP.n9394 a_400_38200# 2.04fF
C16671 VP.t566 a_400_38200# 0.02fF
C16672 VP.n9395 a_400_38200# 0.24fF
C16673 VP.n9396 a_400_38200# 0.91fF
C16674 VP.n9397 a_400_38200# 0.05fF
C16675 VP.t828 a_400_38200# 0.02fF
C16676 VP.n9398 a_400_38200# 0.12fF
C16677 VP.n9399 a_400_38200# 0.14fF
C16678 VP.n9401 a_400_38200# 0.24fF
C16679 VP.t189 a_400_38200# 0.02fF
C16680 VP.n9402 a_400_38200# 0.36fF
C16681 VP.n9403 a_400_38200# 0.36fF
C16682 VP.n9404 a_400_38200# 0.67fF
C16683 VP.n9405 a_400_38200# 0.06fF
C16684 VP.n9406 a_400_38200# 0.09fF
C16685 VP.n9407 a_400_38200# 0.09fF
C16686 VP.n9408 a_400_38200# 0.09fF
C16687 VP.n9409 a_400_38200# 1.45fF
C16688 VP.n9410 a_400_38200# 0.14fF
C16689 VP.n9411 a_400_38200# 0.07fF
C16690 VP.n9412 a_400_38200# 0.72fF
C16691 VP.n9413 a_400_38200# 1.81fF
C16692 VP.n9414 a_400_38200# 2.97fF
C16693 VP.n9415 a_400_38200# 1.06fF
C16694 VP.n9416 a_400_38200# 0.24fF
C16695 VP.t474 a_400_38200# 0.02fF
C16696 VP.n9417 a_400_38200# 0.35fF
C16697 VP.n9418 a_400_38200# 0.63fF
C16698 VP.n9419 a_400_38200# 0.40fF
C16699 VP.n9420 a_400_38200# 0.40fF
C16700 VP.n9421 a_400_38200# 0.12fF
C16701 VP.t1329 a_400_38200# 0.02fF
C16702 VP.n9422 a_400_38200# 0.14fF
C16703 VP.t378 a_400_38200# 0.02fF
C16704 VP.n9424 a_400_38200# 0.12fF
C16705 VP.n9425 a_400_38200# 0.14fF
C16706 VP.n9427 a_400_38200# 1.93fF
C16707 VP.n9428 a_400_38200# 2.23fF
C16708 VP.t1322 a_400_38200# 0.02fF
C16709 VP.n9429 a_400_38200# 0.24fF
C16710 VP.n9430 a_400_38200# 0.35fF
C16711 VP.n9431 a_400_38200# 0.60fF
C16712 VP.n9432 a_400_38200# 0.12fF
C16713 VP.t880 a_400_38200# 0.02fF
C16714 VP.n9433 a_400_38200# 0.14fF
C16715 VP.n9435 a_400_38200# 0.09fF
C16716 VP.n9436 a_400_38200# 0.07fF
C16717 VP.n9437 a_400_38200# 0.30fF
C16718 VP.n9438 a_400_38200# 0.06fF
C16719 VP.n9439 a_400_38200# 0.25fF
C16720 VP.n9440 a_400_38200# 0.45fF
C16721 VP.n9441 a_400_38200# 0.06fF
C16722 VP.n9442 a_400_38200# 0.06fF
C16723 VP.n9443 a_400_38200# 0.03fF
C16724 VP.n9444 a_400_38200# 0.05fF
C16725 VP.n9445 a_400_38200# 0.07fF
C16726 VP.n9446 a_400_38200# 0.19fF
C16727 VP.n9447 a_400_38200# 0.59fF
C16728 VP.n9448 a_400_38200# 0.34fF
C16729 VP.n9449 a_400_38200# 2.04fF
C16730 VP.t1039 a_400_38200# 0.02fF
C16731 VP.n9450 a_400_38200# 0.24fF
C16732 VP.n9451 a_400_38200# 0.91fF
C16733 VP.n9452 a_400_38200# 0.05fF
C16734 VP.t1234 a_400_38200# 0.02fF
C16735 VP.n9453 a_400_38200# 0.12fF
C16736 VP.n9454 a_400_38200# 0.14fF
C16737 VP.n9456 a_400_38200# 0.06fF
C16738 VP.n9457 a_400_38200# 0.09fF
C16739 VP.n9458 a_400_38200# 0.09fF
C16740 VP.n9459 a_400_38200# 1.45fF
C16741 VP.n9460 a_400_38200# 0.14fF
C16742 VP.n9461 a_400_38200# 0.07fF
C16743 VP.n9462 a_400_38200# 0.72fF
C16744 VP.n9463 a_400_38200# 1.81fF
C16745 VP.n9464 a_400_38200# 0.12fF
C16746 VP.t431 a_400_38200# 0.02fF
C16747 VP.n9465 a_400_38200# 0.14fF
C16748 VP.t871 a_400_38200# 0.02fF
C16749 VP.n9467 a_400_38200# 0.24fF
C16750 VP.n9468 a_400_38200# 0.35fF
C16751 VP.n9469 a_400_38200# 0.60fF
C16752 VP.n9470 a_400_38200# 2.97fF
C16753 VP.n9471 a_400_38200# 2.30fF
C16754 VP.t589 a_400_38200# 0.02fF
C16755 VP.n9472 a_400_38200# 0.24fF
C16756 VP.n9473 a_400_38200# 0.91fF
C16757 VP.n9474 a_400_38200# 0.05fF
C16758 VP.t788 a_400_38200# 0.02fF
C16759 VP.n9475 a_400_38200# 0.12fF
C16760 VP.n9476 a_400_38200# 0.14fF
C16761 VP.n9478 a_400_38200# 1.93fF
C16762 VP.n9479 a_400_38200# 2.23fF
C16763 VP.t425 a_400_38200# 0.02fF
C16764 VP.n9480 a_400_38200# 0.24fF
C16765 VP.n9481 a_400_38200# 0.35fF
C16766 VP.n9482 a_400_38200# 0.60fF
C16767 VP.n9483 a_400_38200# 0.12fF
C16768 VP.t1286 a_400_38200# 0.02fF
C16769 VP.n9484 a_400_38200# 0.14fF
C16770 VP.n9486 a_400_38200# 0.09fF
C16771 VP.n9487 a_400_38200# 0.07fF
C16772 VP.n9488 a_400_38200# 0.30fF
C16773 VP.n9489 a_400_38200# 0.06fF
C16774 VP.n9490 a_400_38200# 0.25fF
C16775 VP.n9491 a_400_38200# 0.45fF
C16776 VP.n9492 a_400_38200# 0.06fF
C16777 VP.n9493 a_400_38200# 0.06fF
C16778 VP.n9494 a_400_38200# 0.03fF
C16779 VP.n9495 a_400_38200# 0.05fF
C16780 VP.n9496 a_400_38200# 0.07fF
C16781 VP.n9497 a_400_38200# 0.19fF
C16782 VP.n9498 a_400_38200# 0.59fF
C16783 VP.n9499 a_400_38200# 0.34fF
C16784 VP.n9500 a_400_38200# 2.04fF
C16785 VP.t121 a_400_38200# 0.02fF
C16786 VP.n9501 a_400_38200# 0.24fF
C16787 VP.n9502 a_400_38200# 0.91fF
C16788 VP.n9503 a_400_38200# 0.05fF
C16789 VP.t341 a_400_38200# 0.02fF
C16790 VP.n9504 a_400_38200# 0.12fF
C16791 VP.n9505 a_400_38200# 0.14fF
C16792 VP.n9507 a_400_38200# 0.06fF
C16793 VP.n9508 a_400_38200# 0.09fF
C16794 VP.n9509 a_400_38200# 0.09fF
C16795 VP.n9510 a_400_38200# 1.45fF
C16796 VP.n9511 a_400_38200# 0.14fF
C16797 VP.n9512 a_400_38200# 0.07fF
C16798 VP.n9513 a_400_38200# 0.72fF
C16799 VP.n9514 a_400_38200# 1.81fF
C16800 VP.n9515 a_400_38200# 0.12fF
C16801 VP.t842 a_400_38200# 0.02fF
C16802 VP.n9516 a_400_38200# 0.14fF
C16803 VP.t1279 a_400_38200# 0.02fF
C16804 VP.n9518 a_400_38200# 0.24fF
C16805 VP.n9519 a_400_38200# 0.35fF
C16806 VP.n9520 a_400_38200# 0.60fF
C16807 VP.n9521 a_400_38200# 2.97fF
C16808 VP.n9522 a_400_38200# 2.30fF
C16809 VP.t993 a_400_38200# 0.02fF
C16810 VP.n9523 a_400_38200# 0.24fF
C16811 VP.n9524 a_400_38200# 0.91fF
C16812 VP.n9525 a_400_38200# 0.05fF
C16813 VP.t1187 a_400_38200# 0.02fF
C16814 VP.n9526 a_400_38200# 0.12fF
C16815 VP.n9527 a_400_38200# 0.14fF
C16816 VP.n9529 a_400_38200# 1.93fF
C16817 VP.n9530 a_400_38200# 2.23fF
C16818 VP.t835 a_400_38200# 0.02fF
C16819 VP.n9531 a_400_38200# 0.24fF
C16820 VP.n9532 a_400_38200# 0.35fF
C16821 VP.n9533 a_400_38200# 0.60fF
C16822 VP.n9534 a_400_38200# 0.12fF
C16823 VP.t390 a_400_38200# 0.02fF
C16824 VP.n9535 a_400_38200# 0.14fF
C16825 VP.n9537 a_400_38200# 0.09fF
C16826 VP.n9538 a_400_38200# 0.07fF
C16827 VP.n9539 a_400_38200# 0.30fF
C16828 VP.n9540 a_400_38200# 0.06fF
C16829 VP.n9541 a_400_38200# 0.25fF
C16830 VP.n9542 a_400_38200# 0.45fF
C16831 VP.n9543 a_400_38200# 0.06fF
C16832 VP.n9544 a_400_38200# 0.06fF
C16833 VP.n9545 a_400_38200# 0.03fF
C16834 VP.n9546 a_400_38200# 0.05fF
C16835 VP.n9547 a_400_38200# 0.07fF
C16836 VP.n9548 a_400_38200# 0.19fF
C16837 VP.n9549 a_400_38200# 0.59fF
C16838 VP.n9550 a_400_38200# 0.34fF
C16839 VP.n9551 a_400_38200# 2.04fF
C16840 VP.t548 a_400_38200# 0.02fF
C16841 VP.n9552 a_400_38200# 0.24fF
C16842 VP.n9553 a_400_38200# 0.91fF
C16843 VP.n9554 a_400_38200# 0.05fF
C16844 VP.t809 a_400_38200# 0.02fF
C16845 VP.n9555 a_400_38200# 0.12fF
C16846 VP.n9556 a_400_38200# 0.14fF
C16847 VP.n9558 a_400_38200# 0.06fF
C16848 VP.n9559 a_400_38200# 0.09fF
C16849 VP.n9560 a_400_38200# 0.09fF
C16850 VP.n9561 a_400_38200# 0.43fF
C16851 VP.n9562 a_400_38200# 0.69fF
C16852 VP.n9563 a_400_38200# 0.14fF
C16853 VP.n9564 a_400_38200# 0.07fF
C16854 VP.n9565 a_400_38200# 0.72fF
C16855 VP.n9566 a_400_38200# 1.81fF
C16856 VP.n9567 a_400_38200# 0.12fF
C16857 VP.t1247 a_400_38200# 0.02fF
C16858 VP.n9568 a_400_38200# 0.14fF
C16859 VP.t384 a_400_38200# 0.02fF
C16860 VP.n9570 a_400_38200# 0.24fF
C16861 VP.n9571 a_400_38200# 0.35fF
C16862 VP.n9572 a_400_38200# 0.60fF
C16863 VP.n9573 a_400_38200# 2.97fF
C16864 VP.n9574 a_400_38200# 2.30fF
C16865 VP.t74 a_400_38200# 0.02fF
C16866 VP.n9575 a_400_38200# 0.24fF
C16867 VP.n9576 a_400_38200# 0.91fF
C16868 VP.n9577 a_400_38200# 0.05fF
C16869 VP.t360 a_400_38200# 0.02fF
C16870 VP.n9578 a_400_38200# 0.12fF
C16871 VP.n9579 a_400_38200# 0.14fF
C16872 VP.n9581 a_400_38200# 0.88fF
C16873 VP.n9582 a_400_38200# 0.48fF
C16874 VP.n9583 a_400_38200# 0.88fF
C16875 VP.n9584 a_400_38200# 0.60fF
C16876 VP.n9585 a_400_38200# 2.33fF
C16877 VP.n9586 a_400_38200# 0.59fF
C16878 VP.n9587 a_400_38200# 0.02fF
C16879 VP.n9588 a_400_38200# 0.96fF
C16880 VP.t153 a_400_38200# 15.72fF
C16881 VP.n9589 a_400_38200# 15.42fF
C16882 VP.n9591 a_400_38200# 0.38fF
C16883 VP.n9592 a_400_38200# 0.23fF
C16884 VP.n9593 a_400_38200# 3.42fF
C16885 VP.n9594 a_400_38200# 0.10fF
C16886 VP.n9595 a_400_38200# 0.10fF
C16887 VP.n9596 a_400_38200# 0.06fF
C16888 VP.n9597 a_400_38200# 0.21fF
C16889 VP.n9598 a_400_38200# 1.08fF
C16890 VP.n9599 a_400_38200# 0.03fF
C16891 VP.n9600 a_400_38200# 0.56fF
C16892 VP.n9601 a_400_38200# 0.17fF
C16893 VP.t185 a_400_38200# 0.02fF
C16894 VP.n9602 a_400_38200# 0.64fF
C16895 VP.n9603 a_400_38200# 0.60fF
C16896 VP.n9604 a_400_38200# 2.32fF
C16897 VP.n9605 a_400_38200# 4.93fF
C16898 VP.t1205 a_400_38200# 0.02fF
C16899 VP.n9606 a_400_38200# 1.19fF
C16900 VP.n9607 a_400_38200# 0.05fF
C16901 VP.t144 a_400_38200# 0.02fF
C16902 VP.n9608 a_400_38200# 0.01fF
C16903 VP.n9609 a_400_38200# 0.26fF
C16904 VP.n9611 a_400_38200# 15.28fF
C16905 VP.n9612 a_400_38200# 1.93fF
C16906 VP.n9613 a_400_38200# 2.96fF
C16907 VP.t1240 a_400_38200# 0.02fF
C16908 VP.n9614 a_400_38200# 0.24fF
C16909 VP.n9615 a_400_38200# 0.35fF
C16910 VP.n9616 a_400_38200# 0.60fF
C16911 VP.n9617 a_400_38200# 0.12fF
C16912 VP.t802 a_400_38200# 0.02fF
C16913 VP.n9618 a_400_38200# 0.14fF
C16914 VP.n9620 a_400_38200# 0.02fF
C16915 VP.n9621 a_400_38200# 0.32fF
C16916 VP.n9622 a_400_38200# 0.04fF
C16917 VP.n9623 a_400_38200# 0.05fF
C16918 VP.n9624 a_400_38200# 0.04fF
C16919 VP.n9625 a_400_38200# 0.12fF
C16920 VP.n9626 a_400_38200# 0.09fF
C16921 VP.n9627 a_400_38200# 0.14fF
C16922 VP.n9628 a_400_38200# 0.08fF
C16923 VP.n9629 a_400_38200# 0.09fF
C16924 VP.n9630 a_400_38200# 0.07fF
C16925 VP.n9631 a_400_38200# 0.56fF
C16926 VP.n9632 a_400_38200# 0.20fF
C16927 VP.n9633 a_400_38200# 2.19fF
C16928 VP.t1213 a_400_38200# 0.02fF
C16929 VP.n9634 a_400_38200# 0.12fF
C16930 VP.n9635 a_400_38200# 0.14fF
C16931 VP.t956 a_400_38200# 0.02fF
C16932 VP.n9637 a_400_38200# 0.24fF
C16933 VP.n9638 a_400_38200# 0.91fF
C16934 VP.n9639 a_400_38200# 0.05fF
C16935 VP.t143 a_400_38200# 34.79fF
C16936 VP.t165 a_400_38200# 0.02fF
C16937 VP.n9640 a_400_38200# 0.12fF
C16938 VP.n9641 a_400_38200# 0.14fF
C16939 VP.t1222 a_400_38200# 0.02fF
C16940 VP.n9643 a_400_38200# 0.24fF
C16941 VP.n9644 a_400_38200# 0.91fF
C16942 VP.n9645 a_400_38200# 0.05fF
C16943 VP.t204 a_400_38200# 0.02fF
C16944 VP.n9646 a_400_38200# 0.24fF
C16945 VP.n9647 a_400_38200# 0.35fF
C16946 VP.n9648 a_400_38200# 0.60fF
C16947 VP.n9649 a_400_38200# 0.02fF
C16948 VP.n9650 a_400_38200# 0.04fF
C16949 VP.n9651 a_400_38200# 0.06fF
C16950 VP.n9652 a_400_38200# 0.45fF
C16951 VP.n9653 a_400_38200# 0.10fF
C16952 VP.n9654 a_400_38200# 0.17fF
C16953 VP.n9655 a_400_38200# 0.10fF
C16954 VP.n9656 a_400_38200# 0.04fF
C16955 VP.n9657 a_400_38200# 0.09fF
C16956 VP.n9658 a_400_38200# 0.10fF
C16957 VP.n9659 a_400_38200# 1.82fF
C16958 VP.n9660 a_400_38200# 2.21fF
C16959 VP.n9661 a_400_38200# 26.29fF
C16960 VP.n9662 a_400_38200# 26.29fF
C16961 VP.n9663 a_400_38200# 0.76fF
C16962 VP.n9664 a_400_38200# 0.27fF
C16963 VP.n9665 a_400_38200# 0.59fF
C16964 VP.n9666 a_400_38200# 0.10fF
C16965 VP.n9667 a_400_38200# 3.02fF
C16966 VP.t31 a_400_38200# 15.72fF
C16967 VP.n9668 a_400_38200# 1.15fF
C16968 VP.n9670 a_400_38200# 13.70fF
C16969 VP.n9672 a_400_38200# 1.99fF
C16970 VP.n9673 a_400_38200# 4.39fF
C16971 VP.n9674 a_400_38200# 0.03fF
C16972 VP.n9675 a_400_38200# 0.05fF
C16973 VP.n9676 a_400_38200# 0.07fF
C16974 VP.n9677 a_400_38200# 0.03fF
C16975 VP.n9678 a_400_38200# 0.06fF
C16976 VP.n9679 a_400_38200# 0.06fF
C16977 VP.n9680 a_400_38200# 0.06fF
C16978 VP.n9681 a_400_38200# 0.07fF
C16979 VP.n9682 a_400_38200# 0.57fF
C16980 VP.n9683 a_400_38200# 1.88fF
C16981 VP.n9684 a_400_38200# 0.01fF
C16982 VP.t1044 a_400_38200# 0.02fF
C16983 VP.n9685 a_400_38200# 0.25fF
C16984 VP.t911 a_400_38200# 0.02fF
C16985 VP.n9686 a_400_38200# 0.95fF
C16986 VP.n9687 a_400_38200# 0.70fF
C16987 VP.n9688 a_400_38200# 0.10fF
C16988 VP.n9689 a_400_38200# 0.18fF
C16989 VP.n9690 a_400_38200# 0.09fF
C16990 VP.n9691 a_400_38200# 0.04fF
C16991 VP.n9692 a_400_38200# 0.19fF
C16992 VP.n9693 a_400_38200# 0.26fF
C16993 VP.n9694 a_400_38200# 1.17fF
C16994 VP.n9695 a_400_38200# 0.26fF
C16995 VP.n9696 a_400_38200# 0.05fF
C16996 VP.n9697 a_400_38200# 0.44fF
C16997 VP.n9698 a_400_38200# 0.13fF
C16998 VP.n9699 a_400_38200# 0.02fF
C16999 VP.n9700 a_400_38200# 1.82fF
C17000 VP.n9701 a_400_38200# 0.12fF
C17001 VP.t593 a_400_38200# 0.02fF
C17002 VP.n9702 a_400_38200# 0.14fF
C17003 VP.t1181 a_400_38200# 0.02fF
C17004 VP.n9704 a_400_38200# 0.24fF
C17005 VP.n9705 a_400_38200# 0.35fF
C17006 VP.n9706 a_400_38200# 0.60fF
C17007 VP.n9707 a_400_38200# 0.19fF
C17008 VP.n9708 a_400_38200# 0.11fF
C17009 VP.n9709 a_400_38200# 0.06fF
C17010 VP.n9710 a_400_38200# 0.07fF
C17011 VP.n9711 a_400_38200# 0.10fF
C17012 VP.n9712 a_400_38200# 0.04fF
C17013 VP.n9713 a_400_38200# 0.01fF
C17014 VP.n9714 a_400_38200# 0.01fF
C17015 VP.n9715 a_400_38200# 0.02fF
C17016 VP.n9716 a_400_38200# 0.15fF
C17017 VP.n9717 a_400_38200# 0.37fF
C17018 VP.n9718 a_400_38200# 1.57fF
C17019 VP.n9719 a_400_38200# 2.00fF
C17020 VP.t461 a_400_38200# 0.02fF
C17021 VP.n9720 a_400_38200# 0.24fF
C17022 VP.n9721 a_400_38200# 0.91fF
C17023 VP.n9722 a_400_38200# 0.05fF
C17024 VP.t636 a_400_38200# 0.02fF
C17025 VP.n9723 a_400_38200# 0.12fF
C17026 VP.n9724 a_400_38200# 0.14fF
C17027 VP.n9726 a_400_38200# 0.16fF
C17028 VP.n9727 a_400_38200# 0.19fF
C17029 VP.n9728 a_400_38200# 0.09fF
C17030 VP.n9729 a_400_38200# 0.04fF
C17031 VP.n9730 a_400_38200# 0.14fF
C17032 VP.n9731 a_400_38200# 0.64fF
C17033 VP.n9732 a_400_38200# 1.32fF
C17034 VP.n9733 a_400_38200# 1.81fF
C17035 VP.n9734 a_400_38200# 0.12fF
C17036 VP.t127 a_400_38200# 0.02fF
C17037 VP.n9735 a_400_38200# 0.14fF
C17038 VP.t729 a_400_38200# 0.02fF
C17039 VP.n9737 a_400_38200# 0.24fF
C17040 VP.n9738 a_400_38200# 0.35fF
C17041 VP.n9739 a_400_38200# 0.60fF
C17042 VP.n9740 a_400_38200# 2.27fF
C17043 VP.n9741 a_400_38200# 2.00fF
C17044 VP.t1310 a_400_38200# 0.02fF
C17045 VP.n9742 a_400_38200# 0.24fF
C17046 VP.n9743 a_400_38200# 0.91fF
C17047 VP.n9744 a_400_38200# 0.05fF
C17048 VP.t183 a_400_38200# 0.02fF
C17049 VP.n9745 a_400_38200# 0.12fF
C17050 VP.n9746 a_400_38200# 0.14fF
C17051 VP.n9748 a_400_38200# 0.16fF
C17052 VP.n9749 a_400_38200# 0.19fF
C17053 VP.n9750 a_400_38200# 0.09fF
C17054 VP.n9751 a_400_38200# 0.04fF
C17055 VP.n9752 a_400_38200# 0.14fF
C17056 VP.n9753 a_400_38200# 0.64fF
C17057 VP.n9754 a_400_38200# 1.43fF
C17058 VP.n9755 a_400_38200# 1.81fF
C17059 VP.n9756 a_400_38200# 0.12fF
C17060 VP.t355 a_400_38200# 0.02fF
C17061 VP.n9757 a_400_38200# 0.14fF
C17062 VP.t941 a_400_38200# 0.02fF
C17063 VP.n9759 a_400_38200# 0.24fF
C17064 VP.n9760 a_400_38200# 0.35fF
C17065 VP.n9761 a_400_38200# 0.60fF
C17066 VP.n9762 a_400_38200# 2.27fF
C17067 VP.n9763 a_400_38200# 2.00fF
C17068 VP.t217 a_400_38200# 0.02fF
C17069 VP.n9764 a_400_38200# 0.24fF
C17070 VP.n9765 a_400_38200# 0.91fF
C17071 VP.n9766 a_400_38200# 0.05fF
C17072 VP.t453 a_400_38200# 0.02fF
C17073 VP.n9767 a_400_38200# 0.12fF
C17074 VP.n9768 a_400_38200# 0.14fF
C17075 VP.n9770 a_400_38200# 0.16fF
C17076 VP.n9771 a_400_38200# 0.19fF
C17077 VP.n9772 a_400_38200# 0.09fF
C17078 VP.n9773 a_400_38200# 0.04fF
C17079 VP.n9774 a_400_38200# 0.14fF
C17080 VP.n9775 a_400_38200# 0.64fF
C17081 VP.n9776 a_400_38200# 1.43fF
C17082 VP.n9777 a_400_38200# 1.81fF
C17083 VP.n9778 a_400_38200# 0.12fF
C17084 VP.t759 a_400_38200# 0.02fF
C17085 VP.n9779 a_400_38200# 0.14fF
C17086 VP.t1347 a_400_38200# 0.02fF
C17087 VP.n9781 a_400_38200# 0.24fF
C17088 VP.n9782 a_400_38200# 0.35fF
C17089 VP.n9783 a_400_38200# 0.60fF
C17090 VP.n9784 a_400_38200# 2.27fF
C17091 VP.n9785 a_400_38200# 2.00fF
C17092 VP.t624 a_400_38200# 0.02fF
C17093 VP.n9786 a_400_38200# 0.24fF
C17094 VP.n9787 a_400_38200# 0.91fF
C17095 VP.n9788 a_400_38200# 0.05fF
C17096 VP.t856 a_400_38200# 0.02fF
C17097 VP.n9789 a_400_38200# 0.12fF
C17098 VP.n9790 a_400_38200# 0.14fF
C17099 VP.n9792 a_400_38200# 0.16fF
C17100 VP.n9793 a_400_38200# 0.19fF
C17101 VP.n9794 a_400_38200# 0.09fF
C17102 VP.n9795 a_400_38200# 0.04fF
C17103 VP.n9796 a_400_38200# 0.14fF
C17104 VP.n9797 a_400_38200# 0.64fF
C17105 VP.n9798 a_400_38200# 1.43fF
C17106 VP.n9799 a_400_38200# 1.81fF
C17107 VP.n9800 a_400_38200# 0.12fF
C17108 VP.t1233 a_400_38200# 0.02fF
C17109 VP.n9801 a_400_38200# 0.14fF
C17110 VP.t514 a_400_38200# 0.02fF
C17111 VP.n9803 a_400_38200# 0.24fF
C17112 VP.n9804 a_400_38200# 0.35fF
C17113 VP.n9805 a_400_38200# 0.60fF
C17114 VP.n9806 a_400_38200# 2.27fF
C17115 VP.n9807 a_400_38200# 2.00fF
C17116 VP.t1089 a_400_38200# 0.02fF
C17117 VP.n9808 a_400_38200# 0.24fF
C17118 VP.n9809 a_400_38200# 0.91fF
C17119 VP.n9810 a_400_38200# 0.05fF
C17120 VP.t1263 a_400_38200# 0.02fF
C17121 VP.n9811 a_400_38200# 0.12fF
C17122 VP.n9812 a_400_38200# 0.14fF
C17123 VP.n9814 a_400_38200# 15.28fF
C17124 VP.n9815 a_400_38200# 0.06fF
C17125 VP.n9816 a_400_38200# 0.06fF
C17126 VP.n9817 a_400_38200# 0.03fF
C17127 VP.n9818 a_400_38200# 0.10fF
C17128 VP.n9819 a_400_38200# 0.17fF
C17129 VP.n9820 a_400_38200# 0.10fF
C17130 VP.n9821 a_400_38200# 0.13fF
C17131 VP.n9822 a_400_38200# 0.02fF
C17132 VP.n9823 a_400_38200# 0.04fF
C17133 VP.n9824 a_400_38200# 0.06fF
C17134 VP.n9825 a_400_38200# 0.10fF
C17135 VP.n9826 a_400_38200# 0.05fF
C17136 VP.n9827 a_400_38200# 0.19fF
C17137 VP.n9828 a_400_38200# 0.16fF
C17138 VP.n9829 a_400_38200# 0.04fF
C17139 VP.n9830 a_400_38200# 0.05fF
C17140 VP.n9831 a_400_38200# 0.04fF
C17141 VP.n9832 a_400_38200# 0.12fF
C17142 VP.n9833 a_400_38200# 0.09fF
C17143 VP.n9834 a_400_38200# 0.14fF
C17144 VP.n9835 a_400_38200# 0.56fF
C17145 VP.n9836 a_400_38200# 0.10fF
C17146 VP.n9837 a_400_38200# 1.93fF
C17147 VP.n9838 a_400_38200# 0.12fF
C17148 VP.t393 a_400_38200# 0.02fF
C17149 VP.n9839 a_400_38200# 0.14fF
C17150 VP.t979 a_400_38200# 0.02fF
C17151 VP.n9841 a_400_38200# 0.24fF
C17152 VP.n9842 a_400_38200# 0.35fF
C17153 VP.n9843 a_400_38200# 0.60fF
C17154 VP.n9844 a_400_38200# 0.18fF
C17155 VP.n9845 a_400_38200# 0.45fF
C17156 VP.n9846 a_400_38200# 0.06fF
C17157 VP.n9847 a_400_38200# 0.01fF
C17158 VP.n9848 a_400_38200# 0.01fF
C17159 VP.n9849 a_400_38200# 0.04fF
C17160 VP.n9850 a_400_38200# 0.02fF
C17161 VP.n9851 a_400_38200# 0.07fF
C17162 VP.n9852 a_400_38200# 0.04fF
C17163 VP.n9853 a_400_38200# 0.14fF
C17164 VP.n9854 a_400_38200# 0.45fF
C17165 VP.n9855 a_400_38200# 1.46fF
C17166 VP.n9856 a_400_38200# 1.78fF
C17167 VP.t1034 a_400_38200# 0.02fF
C17168 VP.n9857 a_400_38200# 0.12fF
C17169 VP.n9858 a_400_38200# 0.14fF
C17170 VP.t253 a_400_38200# 0.02fF
C17171 VP.n9860 a_400_38200# 0.24fF
C17172 VP.n9861 a_400_38200# 0.91fF
C17173 VP.n9862 a_400_38200# 0.05fF
C17174 VP.n9863 a_400_38200# 1.93fF
C17175 VP.n9864 a_400_38200# 0.18fF
C17176 VP.n9865 a_400_38200# 0.45fF
C17177 VP.n9866 a_400_38200# 0.06fF
C17178 VP.n9867 a_400_38200# 0.01fF
C17179 VP.n9868 a_400_38200# 0.01fF
C17180 VP.n9869 a_400_38200# 0.04fF
C17181 VP.n9870 a_400_38200# 0.02fF
C17182 VP.n9871 a_400_38200# 0.07fF
C17183 VP.n9872 a_400_38200# 0.04fF
C17184 VP.n9873 a_400_38200# 0.14fF
C17185 VP.n9874 a_400_38200# 0.45fF
C17186 VP.n9875 a_400_38200# 1.46fF
C17187 VP.t52 a_400_38200# 0.02fF
C17188 VP.n9876 a_400_38200# 0.24fF
C17189 VP.n9877 a_400_38200# 0.35fF
C17190 VP.n9878 a_400_38200# 0.60fF
C17191 VP.n9879 a_400_38200# 0.12fF
C17192 VP.t804 a_400_38200# 0.02fF
C17193 VP.n9880 a_400_38200# 0.14fF
C17194 VP.n9882 a_400_38200# 0.10fF
C17195 VP.n9883 a_400_38200# 0.17fF
C17196 VP.n9884 a_400_38200# 0.06fF
C17197 VP.n9885 a_400_38200# 0.06fF
C17198 VP.n9886 a_400_38200# 0.03fF
C17199 VP.n9887 a_400_38200# 0.10fF
C17200 VP.n9888 a_400_38200# 0.13fF
C17201 VP.n9889 a_400_38200# 0.13fF
C17202 VP.n9890 a_400_38200# 0.04fF
C17203 VP.n9891 a_400_38200# 0.05fF
C17204 VP.n9892 a_400_38200# 0.04fF
C17205 VP.n9893 a_400_38200# 0.09fF
C17206 VP.n9894 a_400_38200# 0.05fF
C17207 VP.n9895 a_400_38200# 0.19fF
C17208 VP.n9896 a_400_38200# 0.12fF
C17209 VP.n9897 a_400_38200# 0.09fF
C17210 VP.n9898 a_400_38200# 0.14fF
C17211 VP.n9899 a_400_38200# 0.04fF
C17212 VP.n9900 a_400_38200# 0.02fF
C17213 VP.n9901 a_400_38200# 0.06fF
C17214 VP.n9902 a_400_38200# 0.56fF
C17215 VP.n9903 a_400_38200# 0.10fF
C17216 VP.n9904 a_400_38200# 1.78fF
C17217 VP.t905 a_400_38200# 0.02fF
C17218 VP.n9905 a_400_38200# 0.12fF
C17219 VP.n9906 a_400_38200# 0.14fF
C17220 VP.t664 a_400_38200# 0.02fF
C17221 VP.n9908 a_400_38200# 0.24fF
C17222 VP.n9909 a_400_38200# 0.91fF
C17223 VP.n9910 a_400_38200# 0.05fF
C17224 VP.n9911 a_400_38200# 1.93fF
C17225 VP.n9912 a_400_38200# 0.18fF
C17226 VP.n9913 a_400_38200# 0.45fF
C17227 VP.n9914 a_400_38200# 0.06fF
C17228 VP.n9915 a_400_38200# 0.01fF
C17229 VP.n9916 a_400_38200# 0.01fF
C17230 VP.n9917 a_400_38200# 0.04fF
C17231 VP.n9918 a_400_38200# 0.02fF
C17232 VP.n9919 a_400_38200# 0.07fF
C17233 VP.n9920 a_400_38200# 0.04fF
C17234 VP.n9921 a_400_38200# 0.14fF
C17235 VP.n9922 a_400_38200# 0.45fF
C17236 VP.n9923 a_400_38200# 1.46fF
C17237 VP.t496 a_400_38200# 0.02fF
C17238 VP.n9924 a_400_38200# 0.24fF
C17239 VP.n9925 a_400_38200# 0.35fF
C17240 VP.n9926 a_400_38200# 0.60fF
C17241 VP.n9927 a_400_38200# 0.12fF
C17242 VP.t1208 a_400_38200# 0.02fF
C17243 VP.n9928 a_400_38200# 0.14fF
C17244 VP.n9930 a_400_38200# 0.10fF
C17245 VP.n9931 a_400_38200# 0.17fF
C17246 VP.n9932 a_400_38200# 0.06fF
C17247 VP.n9933 a_400_38200# 0.06fF
C17248 VP.n9934 a_400_38200# 0.03fF
C17249 VP.n9935 a_400_38200# 0.10fF
C17250 VP.n9936 a_400_38200# 0.13fF
C17251 VP.n9937 a_400_38200# 0.13fF
C17252 VP.n9938 a_400_38200# 0.04fF
C17253 VP.n9939 a_400_38200# 0.05fF
C17254 VP.n9940 a_400_38200# 0.04fF
C17255 VP.n9941 a_400_38200# 0.09fF
C17256 VP.n9942 a_400_38200# 0.05fF
C17257 VP.n9943 a_400_38200# 0.19fF
C17258 VP.n9944 a_400_38200# 0.12fF
C17259 VP.n9945 a_400_38200# 0.09fF
C17260 VP.n9946 a_400_38200# 0.14fF
C17261 VP.n9947 a_400_38200# 0.04fF
C17262 VP.n9948 a_400_38200# 0.02fF
C17263 VP.n9949 a_400_38200# 0.06fF
C17264 VP.n9950 a_400_38200# 0.56fF
C17265 VP.n9951 a_400_38200# 0.10fF
C17266 VP.n9952 a_400_38200# 1.78fF
C17267 VP.t1303 a_400_38200# 0.02fF
C17268 VP.n9953 a_400_38200# 0.12fF
C17269 VP.n9954 a_400_38200# 0.14fF
C17270 VP.t1070 a_400_38200# 0.02fF
C17271 VP.n9956 a_400_38200# 0.24fF
C17272 VP.n9957 a_400_38200# 0.91fF
C17273 VP.n9958 a_400_38200# 0.05fF
C17274 VP.n9959 a_400_38200# 1.93fF
C17275 VP.n9960 a_400_38200# 0.18fF
C17276 VP.n9961 a_400_38200# 0.45fF
C17277 VP.n9962 a_400_38200# 0.06fF
C17278 VP.n9963 a_400_38200# 0.01fF
C17279 VP.n9964 a_400_38200# 0.01fF
C17280 VP.n9965 a_400_38200# 0.04fF
C17281 VP.n9966 a_400_38200# 0.02fF
C17282 VP.n9967 a_400_38200# 0.07fF
C17283 VP.n9968 a_400_38200# 0.04fF
C17284 VP.n9969 a_400_38200# 0.14fF
C17285 VP.n9970 a_400_38200# 0.45fF
C17286 VP.n9971 a_400_38200# 1.46fF
C17287 VP.t900 a_400_38200# 0.02fF
C17288 VP.n9972 a_400_38200# 0.24fF
C17289 VP.n9973 a_400_38200# 0.35fF
C17290 VP.n9974 a_400_38200# 0.60fF
C17291 VP.n9975 a_400_38200# 0.12fF
C17292 VP.t376 a_400_38200# 0.02fF
C17293 VP.n9976 a_400_38200# 0.14fF
C17294 VP.n9978 a_400_38200# 0.10fF
C17295 VP.n9979 a_400_38200# 0.17fF
C17296 VP.n9980 a_400_38200# 0.06fF
C17297 VP.n9981 a_400_38200# 0.06fF
C17298 VP.n9982 a_400_38200# 0.03fF
C17299 VP.n9983 a_400_38200# 0.10fF
C17300 VP.n9984 a_400_38200# 0.13fF
C17301 VP.n9985 a_400_38200# 0.13fF
C17302 VP.n9986 a_400_38200# 0.04fF
C17303 VP.n9987 a_400_38200# 0.05fF
C17304 VP.n9988 a_400_38200# 0.04fF
C17305 VP.n9989 a_400_38200# 0.09fF
C17306 VP.n9990 a_400_38200# 0.05fF
C17307 VP.n9991 a_400_38200# 0.19fF
C17308 VP.n9992 a_400_38200# 0.12fF
C17309 VP.n9993 a_400_38200# 0.09fF
C17310 VP.n9994 a_400_38200# 0.14fF
C17311 VP.n9995 a_400_38200# 0.04fF
C17312 VP.n9996 a_400_38200# 0.02fF
C17313 VP.n9997 a_400_38200# 0.06fF
C17314 VP.n9998 a_400_38200# 0.56fF
C17315 VP.n9999 a_400_38200# 0.10fF
C17316 VP.n10000 a_400_38200# 1.78fF
C17317 VP.t409 a_400_38200# 0.02fF
C17318 VP.n10001 a_400_38200# 0.12fF
C17319 VP.n10002 a_400_38200# 0.14fF
C17320 VP.t168 a_400_38200# 0.02fF
C17321 VP.n10004 a_400_38200# 0.24fF
C17322 VP.n10005 a_400_38200# 0.91fF
C17323 VP.n10006 a_400_38200# 0.05fF
C17324 VP.n10007 a_400_38200# 1.93fF
C17325 VP.n10008 a_400_38200# 2.27fF
C17326 VP.t32 a_400_38200# 0.02fF
C17327 VP.n10009 a_400_38200# 0.24fF
C17328 VP.n10010 a_400_38200# 0.35fF
C17329 VP.n10011 a_400_38200# 0.60fF
C17330 VP.n10012 a_400_38200# 0.12fF
C17331 VP.t787 a_400_38200# 0.02fF
C17332 VP.n10013 a_400_38200# 0.14fF
C17333 VP.n10015 a_400_38200# 0.10fF
C17334 VP.n10016 a_400_38200# 0.17fF
C17335 VP.n10017 a_400_38200# 0.06fF
C17336 VP.n10018 a_400_38200# 0.06fF
C17337 VP.n10019 a_400_38200# 0.03fF
C17338 VP.n10020 a_400_38200# 0.10fF
C17339 VP.n10021 a_400_38200# 0.13fF
C17340 VP.n10022 a_400_38200# 0.14fF
C17341 VP.n10023 a_400_38200# 0.04fF
C17342 VP.n10024 a_400_38200# 0.02fF
C17343 VP.n10025 a_400_38200# 0.03fF
C17344 VP.n10026 a_400_38200# 0.03fF
C17345 VP.n10027 a_400_38200# 0.05fF
C17346 VP.n10028 a_400_38200# 0.03fF
C17347 VP.n10029 a_400_38200# 0.04fF
C17348 VP.n10030 a_400_38200# 0.20fF
C17349 VP.n10031 a_400_38200# 0.14fF
C17350 VP.n10032 a_400_38200# 0.02fF
C17351 VP.n10033 a_400_38200# 0.07fF
C17352 VP.n10034 a_400_38200# 0.13fF
C17353 VP.n10035 a_400_38200# 0.04fF
C17354 VP.n10036 a_400_38200# 0.02fF
C17355 VP.n10037 a_400_38200# 0.06fF
C17356 VP.n10038 a_400_38200# 0.55fF
C17357 VP.n10039 a_400_38200# 0.10fF
C17358 VP.n10040 a_400_38200# 1.89fF
C17359 VP.t819 a_400_38200# 0.02fF
C17360 VP.n10041 a_400_38200# 0.12fF
C17361 VP.n10042 a_400_38200# 0.14fF
C17362 VP.t646 a_400_38200# 0.02fF
C17363 VP.n10044 a_400_38200# 0.24fF
C17364 VP.n10045 a_400_38200# 0.91fF
C17365 VP.n10046 a_400_38200# 0.05fF
C17366 VP.n10047 a_400_38200# 1.92fF
C17367 VP.n10048 a_400_38200# 2.51fF
C17368 VP.t312 a_400_38200# 0.02fF
C17369 VP.n10049 a_400_38200# 0.24fF
C17370 VP.n10050 a_400_38200# 0.35fF
C17371 VP.n10051 a_400_38200# 0.60fF
C17372 VP.n10052 a_400_38200# 0.12fF
C17373 VP.t1022 a_400_38200# 0.02fF
C17374 VP.n10053 a_400_38200# 0.14fF
C17375 VP.n10055 a_400_38200# 0.04fF
C17376 VP.n10056 a_400_38200# 0.02fF
C17377 VP.n10057 a_400_38200# 0.06fF
C17378 VP.n10058 a_400_38200# 0.30fF
C17379 VP.n10059 a_400_38200# 0.10fF
C17380 VP.n10060 a_400_38200# 0.28fF
C17381 VP.n10061 a_400_38200# 0.06fF
C17382 VP.n10062 a_400_38200# 0.06fF
C17383 VP.n10063 a_400_38200# 0.03fF
C17384 VP.n10064 a_400_38200# 0.15fF
C17385 VP.n10065 a_400_38200# 0.08fF
C17386 VP.n10066 a_400_38200# 0.14fF
C17387 VP.n10067 a_400_38200# 0.17fF
C17388 VP.n10068 a_400_38200# 0.22fF
C17389 VP.n10069 a_400_38200# 0.64fF
C17390 VP.n10070 a_400_38200# 0.34fF
C17391 VP.n10071 a_400_38200# 1.88fF
C17392 VP.t369 a_400_38200# 0.02fF
C17393 VP.n10072 a_400_38200# 0.12fF
C17394 VP.n10073 a_400_38200# 0.14fF
C17395 VP.t891 a_400_38200# 0.02fF
C17396 VP.n10075 a_400_38200# 0.24fF
C17397 VP.n10076 a_400_38200# 0.91fF
C17398 VP.n10077 a_400_38200# 0.05fF
C17399 VP.n10078 a_400_38200# 0.12fF
C17400 VP.t1249 a_400_38200# 0.02fF
C17401 VP.n10079 a_400_38200# 0.14fF
C17402 VP.t1350 a_400_38200# 0.02fF
C17403 VP.n10080 a_400_38200# 0.12fF
C17404 VP.n10081 a_400_38200# 0.14fF
C17405 VP.n10082 a_400_38200# 2.27fF
C17406 VP.n10083 a_400_38200# 1.81fF
C17407 VP.n10084 a_400_38200# 0.89fF
C17408 VP.n10085 a_400_38200# 0.15fF
C17409 VP.n10086 a_400_38200# 0.16fF
C17410 VP.n10087 a_400_38200# 0.16fF
C17411 VP.n10088 a_400_38200# 0.04fF
C17412 VP.n10089 a_400_38200# 0.15fF
C17413 VP.n10090 a_400_38200# 0.36fF
C17414 VP.n10091 a_400_38200# 0.55fF
C17415 VP.n10092 a_400_38200# 0.38fF
C17416 VP.n10093 a_400_38200# 0.24fF
C17417 VP.t531 a_400_38200# 0.02fF
C17418 VP.n10094 a_400_38200# 0.35fF
C17419 VP.n10095 a_400_38200# 0.60fF
C17420 VP.n10096 a_400_38200# 2.00fF
C17421 VP.n10097 a_400_38200# 0.24fF
C17422 VP.t1107 a_400_38200# 0.02fF
C17423 VP.n10098 a_400_38200# 0.91fF
C17424 VP.n10099 a_400_38200# 0.05fF
C17425 VP.t126 a_400_38200# 35.17fF
C17426 VP.t335 a_400_38200# 0.02fF
C17427 VP.n10100 a_400_38200# 1.21fF
C17428 VP.n10101 a_400_38200# 0.25fF
C17429 VP.n10102 a_400_38200# 0.40fF
C17430 VP.n10103 a_400_38200# 0.03fF
C17431 VP.n10104 a_400_38200# 1.04fF
C17432 VP.n10105 a_400_38200# 0.05fF
C17433 VP.n10106 a_400_38200# 0.06fF
C17434 VP.n10107 a_400_38200# 0.09fF
C17435 VP.n10108 a_400_38200# 0.12fF
C17436 VP.n10109 a_400_38200# 0.20fF
C17437 VP.n10110 a_400_38200# 0.60fF
C17438 VP.n10111 a_400_38200# 0.76fF
C17439 VP.n10112 a_400_38200# 0.92fF
C17440 VP.n10113 a_400_38200# 2.46fF
C17441 VP.n10114 a_400_38200# 1.04fF
C17442 VP.n10115 a_400_38200# 0.49fF
C17443 VP.n10116 a_400_38200# 0.10fF
C17444 VP.n10117 a_400_38200# 0.06fF
C17445 VP.n10118 a_400_38200# 0.07fF
C17446 VP.n10119 a_400_38200# 0.20fF
C17447 VP.n10120 a_400_38200# 0.65fF
C17448 VP.n10121 a_400_38200# 0.32fF
C17449 VP.n10122 a_400_38200# 0.36fF
C17450 VP.n10123 a_400_38200# 0.03fF
C17451 VP.n10124 a_400_38200# 0.01fF
C17452 VP.t1191 a_400_38200# 0.02fF
C17453 VP.n10125 a_400_38200# 0.25fF
C17454 VP.t1059 a_400_38200# 0.02fF
C17455 VP.n10126 a_400_38200# 0.95fF
C17456 VP.n10127 a_400_38200# 0.70fF
C17457 VP.n10128 a_400_38200# 0.06fF
C17458 VP.n10129 a_400_38200# 0.07fF
C17459 VP.n10130 a_400_38200# 0.03fF
C17460 VP.n10131 a_400_38200# 0.05fF
C17461 VP.n10132 a_400_38200# 0.07fF
C17462 VP.n10133 a_400_38200# 0.56fF
C17463 VP.n10134 a_400_38200# 1.86fF
C17464 VP.n10135 a_400_38200# 1.79fF
C17465 VP.n10136 a_400_38200# 1.78fF
C17466 VP.n10137 a_400_38200# 0.12fF
C17467 VP.t739 a_400_38200# 0.02fF
C17468 VP.n10138 a_400_38200# 0.14fF
C17469 VP.t1331 a_400_38200# 0.02fF
C17470 VP.n10140 a_400_38200# 0.24fF
C17471 VP.n10141 a_400_38200# 0.35fF
C17472 VP.n10142 a_400_38200# 0.60fF
C17473 VP.n10143 a_400_38200# 2.11fF
C17474 VP.n10144 a_400_38200# 2.11fF
C17475 VP.t612 a_400_38200# 0.02fF
C17476 VP.n10145 a_400_38200# 0.24fF
C17477 VP.n10146 a_400_38200# 0.91fF
C17478 VP.n10147 a_400_38200# 0.05fF
C17479 VP.t784 a_400_38200# 0.02fF
C17480 VP.n10148 a_400_38200# 0.12fF
C17481 VP.n10149 a_400_38200# 0.14fF
C17482 VP.n10151 a_400_38200# 0.24fF
C17483 VP.t405 a_400_38200# 0.02fF
C17484 VP.n10152 a_400_38200# 0.36fF
C17485 VP.n10153 a_400_38200# 0.36fF
C17486 VP.n10154 a_400_38200# 0.67fF
C17487 VP.n10155 a_400_38200# 2.24fF
C17488 VP.n10156 a_400_38200# 2.59fF
C17489 VP.n10157 a_400_38200# 2.21fF
C17490 VP.n10158 a_400_38200# 2.11fF
C17491 VP.n10159 a_400_38200# 0.74fF
C17492 VP.n10160 a_400_38200# 0.24fF
C17493 VP.t1123 a_400_38200# 0.02fF
C17494 VP.n10161 a_400_38200# 0.35fF
C17495 VP.n10162 a_400_38200# 0.63fF
C17496 VP.n10163 a_400_38200# 0.40fF
C17497 VP.n10164 a_400_38200# 0.40fF
C17498 VP.n10165 a_400_38200# 0.12fF
C17499 VP.t539 a_400_38200# 0.02fF
C17500 VP.n10166 a_400_38200# 0.14fF
C17501 VP.t1182 a_400_38200# 0.02fF
C17502 VP.n10168 a_400_38200# 0.12fF
C17503 VP.n10169 a_400_38200# 0.14fF
C17504 VP.n10171 a_400_38200# 26.29fF
C17505 VP.n10172 a_400_38200# 4.40fF
C17506 VP.n10173 a_400_38200# 3.82fF
C17507 VP.n10174 a_400_38200# 119.55fF
C17508 VP.n10175 a_400_38200# 26.29fF
C17509 VP.n10176 a_400_38200# 5.85fF
C17510 VP.n10177 a_400_38200# 2.59fF
C17511 VP.n10178 a_400_38200# 0.33fF
C17512 VP.n10179 a_400_38200# 6.03fF
C17513 VP.n10180 a_400_38200# 1.02fF
C17514 VP.n10181 a_400_38200# 0.33fF
C17515 VP.n10182 a_400_38200# 2.74fF
C17516 VP.n10183 a_400_38200# 0.72fF
C17517 VP.n10184 a_400_38200# 0.27fF
C17518 VP.n10185 a_400_38200# 1.25fF
C17519 VP.n10186 a_400_38200# 0.49fF
C17520 VP.n10187 a_400_38200# 1.25fF
C17521 VP.n10188 a_400_38200# 0.48fF
C17522 VP.n10189 a_400_38200# 0.91fF
C17523 VP.n10190 a_400_38200# 0.26fF
C17524 VP.t913 a_400_38200# 0.02fF
C17525 VP.n10191 a_400_38200# 0.89fF
C17526 VP.t1317 a_400_38200# 0.02fF
C17527 VP.n10192 a_400_38200# 0.89fF
C17528 VP.n10193 a_400_38200# 2.77fF
C17529 VP.n10194 a_400_38200# 0.06fF
C17530 VP.n10195 a_400_38200# 0.27fF
C17531 VP.n10196 a_400_38200# 0.70fF
C17532 VP.n10197 a_400_38200# 94.45fF
C17533 VP.n10198 a_400_38200# 26.29fF
C17534 VP.n10199 a_400_38200# 94.45fF
C17535 VP.n10200 a_400_38200# 26.29fF
C17536 VP.n10201 a_400_38200# 6.07fF
C17537 VP.n10202 a_400_38200# 1.66fF
C17538 VP.n10203 a_400_38200# 0.02fF
C17539 VP.t197 a_400_38200# 0.02fF
C17540 VP.n10204 a_400_38200# 0.37fF
C17541 VP.n10205 a_400_38200# 0.02fF
C17542 VP.t1050 a_400_38200# 0.02fF
C17543 VP.n10206 a_400_38200# 0.37fF
C17544 VP.n10207 a_400_38200# 1.25fF
C17545 VP.n10208 a_400_38200# 0.48fF
C17546 VP.n10209 a_400_38200# 0.91fF
C17547 VP.n10210 a_400_38200# 0.26fF
C17548 VP.t778 a_400_38200# 0.02fF
C17549 VP.n10211 a_400_38200# 0.89fF
C17550 VP.t1113 a_400_38200# 0.02fF
C17551 VP.n10212 a_400_38200# 0.89fF
C17552 VP.n10213 a_400_38200# 2.77fF
C17553 VP.n10214 a_400_38200# 26.29fF
C17554 VP.n10215 a_400_38200# 26.29fF
C17555 VP.n10216 a_400_38200# 5.98fF
C17556 VP.n10217 a_400_38200# 0.06fF
C17557 VP.n10218 a_400_38200# 0.27fF
C17558 VP.n10219 a_400_38200# 0.70fF
C17559 VP.n10220 a_400_38200# 1.66fF
C17560 VP.n10221 a_400_38200# 0.02fF
C17561 VP.t1292 a_400_38200# 0.02fF
C17562 VP.n10222 a_400_38200# 0.37fF
C17563 VP.n10223 a_400_38200# 1.25fF
C17564 VP.n10224 a_400_38200# 0.48fF
C17565 VP.n10225 a_400_38200# 0.91fF
C17566 VP.n10226 a_400_38200# 0.26fF
C17567 VP.t329 a_400_38200# 0.02fF
C17568 VP.n10227 a_400_38200# 0.89fF
C17569 VP.t669 a_400_38200# 0.02fF
C17570 VP.n10228 a_400_38200# 0.89fF
C17571 VP.n10229 a_400_38200# 26.29fF
C17572 VP.n10230 a_400_38200# 26.29fF
C17573 VP.n10231 a_400_38200# 5.88fF
C17574 VP.n10232 a_400_38200# 2.84fF
C17575 VP.n10233 a_400_38200# 0.02fF
C17576 VP.t919 a_400_38200# 0.02fF
C17577 VP.n10234 a_400_38200# 0.37fF
C17578 VP.n10235 a_400_38200# 1.25fF
C17579 VP.n10236 a_400_38200# 0.48fF
C17580 VP.n10237 a_400_38200# 0.91fF
C17581 VP.n10238 a_400_38200# 0.26fF
C17582 VP.t1173 a_400_38200# 0.02fF
C17583 VP.n10239 a_400_38200# 0.89fF
C17584 VP.t222 a_400_38200# 0.02fF
C17585 VP.n10240 a_400_38200# 0.89fF
C17586 VP.n10241 a_400_38200# 2.77fF
C17587 VP.n10242 a_400_38200# 26.29fF
C17588 VP.n10243 a_400_38200# 26.29fF
C17589 VP.n10244 a_400_38200# 5.98fF
C17590 VP.n10245 a_400_38200# 0.06fF
C17591 VP.n10246 a_400_38200# 0.27fF
C17592 VP.n10247 a_400_38200# 0.70fF
C17593 VP.n10248 a_400_38200# 1.66fF
C17594 VP.n10249 a_400_38200# 0.02fF
C17595 VP.t469 a_400_38200# 0.02fF
C17596 VP.n10250 a_400_38200# 0.37fF
C17597 VP.n10251 a_400_38200# 1.25fF
C17598 VP.n10252 a_400_38200# 0.48fF
C17599 VP.n10253 a_400_38200# 0.91fF
C17600 VP.n10254 a_400_38200# 0.26fF
C17601 VP.t720 a_400_38200# 0.02fF
C17602 VP.n10255 a_400_38200# 0.89fF
C17603 VP.t1077 a_400_38200# 0.02fF
C17604 VP.n10256 a_400_38200# 0.89fF
C17605 VP.n10257 a_400_38200# 26.29fF
C17606 VP.n10258 a_400_38200# 26.29fF
C17607 VP.n10259 a_400_38200# 5.88fF
C17608 VP.n10260 a_400_38200# 2.84fF
C17609 VP.n10261 a_400_38200# 0.02fF
C17610 VP.t1315 a_400_38200# 0.02fF
C17611 VP.n10262 a_400_38200# 0.37fF
C17612 VP.n10263 a_400_38200# 1.25fF
C17613 VP.n10264 a_400_38200# 0.48fF
C17614 VP.n10265 a_400_38200# 0.91fF
C17615 VP.n10266 a_400_38200# 0.26fF
C17616 VP.t273 a_400_38200# 0.02fF
C17617 VP.n10267 a_400_38200# 0.89fF
C17618 VP.t635 a_400_38200# 0.02fF
C17619 VP.n10268 a_400_38200# 0.89fF
C17620 VP.n10269 a_400_38200# 2.77fF
C17621 VP.n10270 a_400_38200# 26.29fF
C17622 VP.n10271 a_400_38200# 26.29fF
C17623 VP.n10272 a_400_38200# 5.98fF
C17624 VP.n10273 a_400_38200# 0.06fF
C17625 VP.n10274 a_400_38200# 0.27fF
C17626 VP.n10275 a_400_38200# 0.70fF
C17627 VP.n10276 a_400_38200# 1.66fF
C17628 VP.n10277 a_400_38200# 0.02fF
C17629 VP.t866 a_400_38200# 0.02fF
C17630 VP.n10278 a_400_38200# 0.37fF
C17631 VP.n10279 a_400_38200# 1.25fF
C17632 VP.n10280 a_400_38200# 0.48fF
C17633 VP.n10281 a_400_38200# 0.91fF
C17634 VP.n10282 a_400_38200# 0.26fF
C17635 VP.t1129 a_400_38200# 0.02fF
C17636 VP.n10283 a_400_38200# 0.89fF
C17637 VP.t181 a_400_38200# 0.02fF
C17638 VP.n10284 a_400_38200# 0.89fF
C17639 VP.n10285 a_400_38200# 26.29fF
C17640 VP.n10286 a_400_38200# 26.29fF
C17641 VP.n10287 a_400_38200# 5.88fF
C17642 VP.n10288 a_400_38200# 2.84fF
C17643 VP.n10289 a_400_38200# 0.02fF
C17644 VP.t419 a_400_38200# 0.02fF
C17645 VP.n10290 a_400_38200# 0.37fF
C17646 VP.n10291 a_400_38200# 1.25fF
C17647 VP.n10292 a_400_38200# 0.48fF
C17648 VP.n10293 a_400_38200# 0.91fF
C17649 VP.n10294 a_400_38200# 0.26fF
C17650 VP.t682 a_400_38200# 0.02fF
C17651 VP.n10295 a_400_38200# 0.89fF
C17652 VP.t1095 a_400_38200# 0.02fF
C17653 VP.n10296 a_400_38200# 0.89fF
C17654 VP.n10297 a_400_38200# 2.77fF
C17655 VP.n10298 a_400_38200# 26.29fF
C17656 VP.n10299 a_400_38200# 26.29fF
C17657 VP.n10300 a_400_38200# 5.98fF
C17658 VP.n10301 a_400_38200# 0.06fF
C17659 VP.n10302 a_400_38200# 0.27fF
C17660 VP.n10303 a_400_38200# 0.70fF
C17661 VP.n10304 a_400_38200# 1.66fF
C17662 VP.n10305 a_400_38200# 0.02fF
C17663 VP.t1276 a_400_38200# 0.02fF
C17664 VP.n10306 a_400_38200# 0.37fF
C17665 VP.n10307 a_400_38200# 1.13fF
C17666 VP.n10308 a_400_38200# 0.48fF
C17667 VP.n10309 a_400_38200# 0.91fF
C17668 VP.n10310 a_400_38200# 0.26fF
C17669 VP.t237 a_400_38200# 0.02fF
C17670 VP.n10311 a_400_38200# 0.89fF
C17671 VP.t654 a_400_38200# 0.02fF
C17672 VP.n10312 a_400_38200# 0.89fF
C17673 VP.n10313 a_400_38200# 2.77fF
C17674 VP.n10314 a_400_38200# 37.85fF
C17675 VP.n10315 a_400_38200# 26.29fF
C17676 VP.n10316 a_400_38200# 37.85fF
C17677 VP.n10317 a_400_38200# 26.29fF
C17678 VP.n10318 a_400_38200# 5.98fF
C17679 VP.n10319 a_400_38200# 0.06fF
C17680 VP.n10320 a_400_38200# 0.27fF
C17681 VP.n10321 a_400_38200# 0.70fF
C17682 VP.n10322 a_400_38200# 1.66fF
C17683 VP.n10323 a_400_38200# 0.02fF
C17684 VP.t831 a_400_38200# 0.02fF
C17685 VP.n10324 a_400_38200# 0.37fF
C17686 VP.n10325 a_400_38200# 6.13fF
C17687 VP.n10326 a_400_38200# 1.93fF
C17688 VP.t1092 a_400_38200# 0.02fF
C17689 VP.n10327 a_400_38200# 0.89fF
C17690 VP.t206 a_400_38200# 0.02fF
C17691 VP.n10328 a_400_38200# 0.89fF
C17692 VP.n10329 a_400_38200# 2.61fF
C17693 VP.n10330 a_400_38200# 1.07fF
C17694 VP.n10331 a_400_38200# 0.31fF
C17695 VP.n10332 a_400_38200# 1.02fF
C17696 VP.n10333 a_400_38200# 0.24fF
C17697 VP.n10334 a_400_38200# 0.46fF
C17698 VP.n10335 a_400_38200# 0.02fF
C17699 VP.t379 a_400_38200# 0.02fF
C17700 VP.n10336 a_400_38200# 0.37fF
C17701 VP.t471 a_400_38200# 0.02fF
C17702 VP.n10337 a_400_38200# 0.89fF
C17703 VP.n10338 a_400_38200# 0.02fF
C17704 VP.t645 a_400_38200# 0.02fF
C17705 VP.n10339 a_400_38200# 0.37fF
C17706 VP.t9 a_400_38200# 0.02fF
C17707 VP.n10340 a_400_38200# 0.89fF
C17708 VP.t451 a_400_38200# 0.02fF
C17709 VP.n10341 a_400_38200# 0.44fF
C17710 VP.t631 a_400_38200# 0.02fF
C17711 VP.n10342 a_400_38200# 1.30fF
C17712 VP.n10343 a_400_38200# 1.59fF
C17713 VP.n10344 a_400_38200# 12.08fF
C17714 VP.n10345 a_400_38200# 0.88fF
C17715 VP.n10346 a_400_38200# 43.82fF
C17716 VP.n10347 a_400_38200# 0.52fF
C17717 VP.n10348 a_400_38200# 3.57fF
C17718 VP.n10349 a_400_38200# 1.77fF
C17719 VP.n10350 a_400_38200# 0.50fF
C17720 VP.n10351 a_400_38200# 6.23fF
C17721 VP.n10352 a_400_38200# 0.25fF
C17722 VP.t462 a_400_38200# 0.02fF
C17723 VP.n10353 a_400_38200# 0.89fF
C17724 VP.t868 a_400_38200# 0.02fF
C17725 VP.n10354 a_400_38200# 0.89fF
C17726 VP.n10355 a_400_38200# 0.91fF
C17727 VP.n10356 a_400_38200# 0.26fF
C17728 VP.n10357 a_400_38200# 1.25fF
C17729 VP.n10358 a_400_38200# 0.48fF
C17730 VP.t8 a_400_38200# 78.13fF
C17731 VP.n10359 a_400_38200# 2.59fF
C17732 VP.n10360 a_400_38200# 2.21fF
C17733 VP.n10361 a_400_38200# 2.11fF
C17734 VP.t231 a_400_38200# 0.02fF
C17735 VP.n10362 a_400_38200# 0.24fF
C17736 VP.n10363 a_400_38200# 0.35fF
C17737 VP.n10364 a_400_38200# 0.60fF
C17738 VP.n10365 a_400_38200# 0.12fF
C17739 VP.t948 a_400_38200# 0.02fF
C17740 VP.n10366 a_400_38200# 0.14fF
C17741 VP.n10368 a_400_38200# 2.02fF
C17742 VP.n10369 a_400_38200# 1.98fF
C17743 VP.t816 a_400_38200# 0.02fF
C17744 VP.n10370 a_400_38200# 0.24fF
C17745 VP.n10371 a_400_38200# 0.91fF
C17746 VP.n10372 a_400_38200# 0.05fF
C17747 VP.t1051 a_400_38200# 0.02fF
C17748 VP.n10373 a_400_38200# 0.12fF
C17749 VP.n10374 a_400_38200# 0.14fF
C17750 VP.n10376 a_400_38200# 2.59fF
C17751 VP.n10377 a_400_38200# 2.21fF
C17752 VP.n10378 a_400_38200# 2.11fF
C17753 VP.t643 a_400_38200# 0.02fF
C17754 VP.n10379 a_400_38200# 0.24fF
C17755 VP.n10380 a_400_38200# 0.35fF
C17756 VP.n10381 a_400_38200# 0.60fF
C17757 VP.n10382 a_400_38200# 0.12fF
C17758 VP.t7 a_400_38200# 0.02fF
C17759 VP.n10383 a_400_38200# 0.14fF
C17760 VP.n10385 a_400_38200# 2.02fF
C17761 VP.n10386 a_400_38200# 1.98fF
C17762 VP.t1219 a_400_38200# 0.02fF
C17763 VP.n10387 a_400_38200# 0.24fF
C17764 VP.n10388 a_400_38200# 0.91fF
C17765 VP.n10389 a_400_38200# 0.05fF
C17766 VP.t133 a_400_38200# 0.02fF
C17767 VP.n10390 a_400_38200# 0.12fF
C17768 VP.n10391 a_400_38200# 0.14fF
C17769 VP.n10393 a_400_38200# 2.59fF
C17770 VP.n10394 a_400_38200# 2.21fF
C17771 VP.n10395 a_400_38200# 2.11fF
C17772 VP.t1045 a_400_38200# 0.02fF
C17773 VP.n10396 a_400_38200# 0.24fF
C17774 VP.n10397 a_400_38200# 0.35fF
C17775 VP.n10398 a_400_38200# 0.60fF
C17776 VP.n10399 a_400_38200# 0.12fF
C17777 VP.t521 a_400_38200# 0.02fF
C17778 VP.n10400 a_400_38200# 0.14fF
C17779 VP.n10402 a_400_38200# 2.02fF
C17780 VP.n10403 a_400_38200# 1.98fF
C17781 VP.t324 a_400_38200# 0.02fF
C17782 VP.n10404 a_400_38200# 0.24fF
C17783 VP.n10405 a_400_38200# 0.91fF
C17784 VP.n10406 a_400_38200# 0.05fF
C17785 VP.t554 a_400_38200# 0.02fF
C17786 VP.n10407 a_400_38200# 0.12fF
C17787 VP.n10408 a_400_38200# 0.14fF
C17788 VP.n10410 a_400_38200# 1.39fF
C17789 VP.n10411 a_400_38200# 0.06fF
C17790 VP.n10412 a_400_38200# 0.19fF
C17791 VP.n10413 a_400_38200# 0.10fF
C17792 VP.n10414 a_400_38200# 0.10fF
C17793 VP.n10415 a_400_38200# 0.18fF
C17794 VP.n10416 a_400_38200# 0.09fF
C17795 VP.n10417 a_400_38200# 0.04fF
C17796 VP.n10418 a_400_38200# 0.46fF
C17797 VP.n10419 a_400_38200# 0.13fF
C17798 VP.n10420 a_400_38200# 0.02fF
C17799 VP.n10421 a_400_38200# 2.43fF
C17800 VP.n10422 a_400_38200# 0.12fF
C17801 VP.t1170 a_400_38200# 0.02fF
C17802 VP.n10423 a_400_38200# 0.14fF
C17803 VP.t465 a_400_38200# 0.02fF
C17804 VP.n10425 a_400_38200# 0.24fF
C17805 VP.n10426 a_400_38200# 0.35fF
C17806 VP.n10427 a_400_38200# 0.60fF
C17807 VP.n10428 a_400_38200# 3.13fF
C17808 VP.n10429 a_400_38200# 1.80fF
C17809 VP.t1037 a_400_38200# 0.02fF
C17810 VP.n10430 a_400_38200# 0.24fF
C17811 VP.n10431 a_400_38200# 0.91fF
C17812 VP.n10432 a_400_38200# 0.05fF
C17813 VP.t515 a_400_38200# 0.02fF
C17814 VP.n10433 a_400_38200# 0.12fF
C17815 VP.n10434 a_400_38200# 0.14fF
C17816 VP.t147 a_400_38200# 17.67fF
C17817 VP.n10436 a_400_38200# 15.28fF
C17818 VP.n10437 a_400_38200# 0.11fF
C17819 VP.n10438 a_400_38200# 0.32fF
C17820 VP.n10439 a_400_38200# 0.11fF
C17821 VP.n10440 a_400_38200# 0.12fF
C17822 VP.n10441 a_400_38200# 0.08fF
C17823 VP.n10442 a_400_38200# 0.08fF
C17824 VP.n10443 a_400_38200# 0.06fF
C17825 VP.n10444 a_400_38200# 0.10fF
C17826 VP.n10445 a_400_38200# 0.05fF
C17827 VP.n10446 a_400_38200# 0.19fF
C17828 VP.n10447 a_400_38200# 0.16fF
C17829 VP.n10448 a_400_38200# 0.04fF
C17830 VP.n10449 a_400_38200# 0.05fF
C17831 VP.n10450 a_400_38200# 0.04fF
C17832 VP.n10451 a_400_38200# 0.12fF
C17833 VP.n10452 a_400_38200# 0.09fF
C17834 VP.n10453 a_400_38200# 0.14fF
C17835 VP.n10454 a_400_38200# 0.56fF
C17836 VP.n10455 a_400_38200# 0.15fF
C17837 VP.n10456 a_400_38200# 1.96fF
C17838 VP.n10457 a_400_38200# 0.12fF
C17839 VP.t287 a_400_38200# 0.02fF
C17840 VP.n10458 a_400_38200# 0.14fF
C17841 VP.t879 a_400_38200# 0.02fF
C17842 VP.n10460 a_400_38200# 0.24fF
C17843 VP.n10461 a_400_38200# 0.35fF
C17844 VP.n10462 a_400_38200# 0.60fF
C17845 VP.n10463 a_400_38200# 2.00fF
C17846 VP.n10464 a_400_38200# 1.89fF
C17847 VP.t336 a_400_38200# 0.02fF
C17848 VP.n10465 a_400_38200# 0.12fF
C17849 VP.n10466 a_400_38200# 0.14fF
C17850 VP.t148 a_400_38200# 0.02fF
C17851 VP.n10468 a_400_38200# 0.24fF
C17852 VP.n10469 a_400_38200# 0.91fF
C17853 VP.n10470 a_400_38200# 0.05fF
C17854 VP.n10471 a_400_38200# 1.96fF
C17855 VP.n10472 a_400_38200# 2.00fF
C17856 VP.t676 a_400_38200# 0.02fF
C17857 VP.n10473 a_400_38200# 0.24fF
C17858 VP.n10474 a_400_38200# 0.35fF
C17859 VP.n10475 a_400_38200# 0.60fF
C17860 VP.n10476 a_400_38200# 0.12fF
C17861 VP.t63 a_400_38200# 0.02fF
C17862 VP.n10477 a_400_38200# 0.14fF
C17863 VP.n10479 a_400_38200# 0.11fF
C17864 VP.n10480 a_400_38200# 0.12fF
C17865 VP.n10481 a_400_38200# 0.08fF
C17866 VP.n10482 a_400_38200# 0.08fF
C17867 VP.n10483 a_400_38200# 0.06fF
C17868 VP.n10484 a_400_38200# 0.12fF
C17869 VP.n10485 a_400_38200# 0.11fF
C17870 VP.n10486 a_400_38200# 0.32fF
C17871 VP.n10487 a_400_38200# 0.18fF
C17872 VP.n10488 a_400_38200# 0.03fF
C17873 VP.n10489 a_400_38200# 0.05fF
C17874 VP.n10490 a_400_38200# 0.04fF
C17875 VP.n10491 a_400_38200# 0.11fF
C17876 VP.n10492 a_400_38200# 0.06fF
C17877 VP.n10493 a_400_38200# 0.06fF
C17878 VP.n10494 a_400_38200# 0.07fF
C17879 VP.n10495 a_400_38200# 0.12fF
C17880 VP.n10496 a_400_38200# 0.22fF
C17881 VP.n10497 a_400_38200# 0.48fF
C17882 VP.n10498 a_400_38200# 0.21fF
C17883 VP.n10499 a_400_38200# 1.88fF
C17884 VP.t198 a_400_38200# 0.02fF
C17885 VP.n10500 a_400_38200# 0.12fF
C17886 VP.n10501 a_400_38200# 0.14fF
C17887 VP.t1261 a_400_38200# 0.02fF
C17888 VP.n10503 a_400_38200# 0.24fF
C17889 VP.n10504 a_400_38200# 0.91fF
C17890 VP.n10505 a_400_38200# 0.05fF
C17891 VP.n10506 a_400_38200# 1.96fF
C17892 VP.n10507 a_400_38200# 2.00fF
C17893 VP.t1086 a_400_38200# 0.02fF
C17894 VP.n10508 a_400_38200# 0.24fF
C17895 VP.n10509 a_400_38200# 0.35fF
C17896 VP.n10510 a_400_38200# 0.60fF
C17897 VP.n10511 a_400_38200# 0.12fF
C17898 VP.t500 a_400_38200# 0.02fF
C17899 VP.n10512 a_400_38200# 0.14fF
C17900 VP.n10514 a_400_38200# 0.11fF
C17901 VP.n10515 a_400_38200# 0.12fF
C17902 VP.n10516 a_400_38200# 0.08fF
C17903 VP.n10517 a_400_38200# 0.08fF
C17904 VP.n10518 a_400_38200# 0.06fF
C17905 VP.n10519 a_400_38200# 0.12fF
C17906 VP.n10520 a_400_38200# 0.11fF
C17907 VP.n10521 a_400_38200# 0.32fF
C17908 VP.n10522 a_400_38200# 0.18fF
C17909 VP.n10523 a_400_38200# 0.03fF
C17910 VP.n10524 a_400_38200# 0.05fF
C17911 VP.n10525 a_400_38200# 0.04fF
C17912 VP.n10526 a_400_38200# 0.11fF
C17913 VP.n10527 a_400_38200# 0.06fF
C17914 VP.n10528 a_400_38200# 0.06fF
C17915 VP.n10529 a_400_38200# 0.07fF
C17916 VP.n10530 a_400_38200# 0.12fF
C17917 VP.n10531 a_400_38200# 0.22fF
C17918 VP.n10532 a_400_38200# 0.48fF
C17919 VP.n10533 a_400_38200# 0.21fF
C17920 VP.n10534 a_400_38200# 1.88fF
C17921 VP.t601 a_400_38200# 0.02fF
C17922 VP.n10535 a_400_38200# 0.12fF
C17923 VP.n10536 a_400_38200# 0.14fF
C17924 VP.t365 a_400_38200# 0.02fF
C17925 VP.n10538 a_400_38200# 0.24fF
C17926 VP.n10539 a_400_38200# 0.91fF
C17927 VP.n10540 a_400_38200# 0.05fF
C17928 VP.n10541 a_400_38200# 1.96fF
C17929 VP.n10542 a_400_38200# 2.00fF
C17930 VP.t193 a_400_38200# 0.02fF
C17931 VP.n10543 a_400_38200# 0.24fF
C17932 VP.n10544 a_400_38200# 0.35fF
C17933 VP.n10545 a_400_38200# 0.60fF
C17934 VP.n10546 a_400_38200# 0.12fF
C17935 VP.t908 a_400_38200# 0.02fF
C17936 VP.n10547 a_400_38200# 0.14fF
C17937 VP.n10549 a_400_38200# 0.11fF
C17938 VP.n10550 a_400_38200# 0.12fF
C17939 VP.n10551 a_400_38200# 0.08fF
C17940 VP.n10552 a_400_38200# 0.08fF
C17941 VP.n10553 a_400_38200# 0.06fF
C17942 VP.n10554 a_400_38200# 0.12fF
C17943 VP.n10555 a_400_38200# 0.11fF
C17944 VP.n10556 a_400_38200# 0.32fF
C17945 VP.n10557 a_400_38200# 0.18fF
C17946 VP.n10558 a_400_38200# 0.03fF
C17947 VP.n10559 a_400_38200# 0.05fF
C17948 VP.n10560 a_400_38200# 0.04fF
C17949 VP.n10561 a_400_38200# 0.11fF
C17950 VP.n10562 a_400_38200# 0.06fF
C17951 VP.n10563 a_400_38200# 0.06fF
C17952 VP.n10564 a_400_38200# 0.07fF
C17953 VP.n10565 a_400_38200# 0.12fF
C17954 VP.n10566 a_400_38200# 0.22fF
C17955 VP.n10567 a_400_38200# 0.48fF
C17956 VP.n10568 a_400_38200# 0.21fF
C17957 VP.n10569 a_400_38200# 1.88fF
C17958 VP.t999 a_400_38200# 0.02fF
C17959 VP.n10570 a_400_38200# 0.12fF
C17960 VP.n10571 a_400_38200# 0.14fF
C17961 VP.t775 a_400_38200# 0.02fF
C17962 VP.n10573 a_400_38200# 0.24fF
C17963 VP.n10574 a_400_38200# 0.91fF
C17964 VP.n10575 a_400_38200# 0.05fF
C17965 VP.n10576 a_400_38200# 1.96fF
C17966 VP.n10577 a_400_38200# 2.09fF
C17967 VP.t662 a_400_38200# 0.02fF
C17968 VP.n10578 a_400_38200# 0.24fF
C17969 VP.n10579 a_400_38200# 0.35fF
C17970 VP.n10580 a_400_38200# 0.60fF
C17971 VP.n10581 a_400_38200# 0.12fF
C17972 VP.t42 a_400_38200# 0.02fF
C17973 VP.n10582 a_400_38200# 0.14fF
C17974 VP.n10584 a_400_38200# 0.11fF
C17975 VP.n10585 a_400_38200# 0.12fF
C17976 VP.n10586 a_400_38200# 0.08fF
C17977 VP.n10587 a_400_38200# 0.08fF
C17978 VP.n10588 a_400_38200# 0.06fF
C17979 VP.n10589 a_400_38200# 0.12fF
C17980 VP.n10590 a_400_38200# 0.11fF
C17981 VP.n10591 a_400_38200# 0.32fF
C17982 VP.n10592 a_400_38200# 0.18fF
C17983 VP.n10593 a_400_38200# 0.03fF
C17984 VP.n10594 a_400_38200# 0.05fF
C17985 VP.n10595 a_400_38200# 0.04fF
C17986 VP.n10596 a_400_38200# 0.11fF
C17987 VP.n10597 a_400_38200# 0.06fF
C17988 VP.n10598 a_400_38200# 0.06fF
C17989 VP.n10599 a_400_38200# 0.07fF
C17990 VP.n10600 a_400_38200# 0.12fF
C17991 VP.n10601 a_400_38200# 0.22fF
C17992 VP.n10602 a_400_38200# 0.48fF
C17993 VP.n10603 a_400_38200# 0.21fF
C17994 VP.n10604 a_400_38200# 1.88fF
C17995 VP.t82 a_400_38200# 0.02fF
C17996 VP.n10605 a_400_38200# 0.12fF
C17997 VP.n10606 a_400_38200# 0.14fF
C17998 VP.t1241 a_400_38200# 0.02fF
C17999 VP.n10608 a_400_38200# 0.24fF
C18000 VP.n10609 a_400_38200# 0.91fF
C18001 VP.n10610 a_400_38200# 0.05fF
C18002 VP.n10611 a_400_38200# 1.96fF
C18003 VP.n10612 a_400_38200# 0.22fF
C18004 VP.n10613 a_400_38200# 0.56fF
C18005 VP.n10614 a_400_38200# 1.22fF
C18006 VP.n10615 a_400_38200# 0.55fF
C18007 VP.t214 a_400_38200# 0.02fF
C18008 VP.n10616 a_400_38200# 0.24fF
C18009 VP.n10617 a_400_38200# 0.35fF
C18010 VP.n10618 a_400_38200# 0.60fF
C18011 VP.n10619 a_400_38200# 0.12fF
C18012 VP.t931 a_400_38200# 0.02fF
C18013 VP.n10620 a_400_38200# 0.14fF
C18014 VP.n10622 a_400_38200# 0.11fF
C18015 VP.n10623 a_400_38200# 0.12fF
C18016 VP.n10624 a_400_38200# 0.08fF
C18017 VP.n10625 a_400_38200# 0.08fF
C18018 VP.n10626 a_400_38200# 0.06fF
C18019 VP.n10627 a_400_38200# 0.30fF
C18020 VP.n10628 a_400_38200# 0.11fF
C18021 VP.n10629 a_400_38200# 0.40fF
C18022 VP.n10630 a_400_38200# 0.23fF
C18023 VP.n10631 a_400_38200# 0.06fF
C18024 VP.n10632 a_400_38200# 0.04fF
C18025 VP.n10633 a_400_38200# 0.04fF
C18026 VP.n10634 a_400_38200# 0.05fF
C18027 VP.n10635 a_400_38200# 0.03fF
C18028 VP.n10636 a_400_38200# 0.05fF
C18029 VP.n10637 a_400_38200# 0.04fF
C18030 VP.n10638 a_400_38200# 0.05fF
C18031 VP.n10639 a_400_38200# 0.20fF
C18032 VP.n10640 a_400_38200# 0.54fF
C18033 VP.n10641 a_400_38200# 0.34fF
C18034 VP.n10642 a_400_38200# 1.73fF
C18035 VP.t962 a_400_38200# 0.02fF
C18036 VP.n10643 a_400_38200# 0.12fF
C18037 VP.n10644 a_400_38200# 0.14fF
C18038 VP.t795 a_400_38200# 0.02fF
C18039 VP.n10646 a_400_38200# 0.24fF
C18040 VP.n10647 a_400_38200# 0.91fF
C18041 VP.n10648 a_400_38200# 0.05fF
C18042 VP.t6 a_400_38200# 35.17fF
C18043 VP.t481 a_400_38200# 0.02fF
C18044 VP.n10649 a_400_38200# 1.21fF
C18045 VP.n10650 a_400_38200# 0.25fF
C18046 VP.n10651 a_400_38200# 0.03fF
C18047 VP.n10652 a_400_38200# 0.06fF
C18048 VP.n10653 a_400_38200# 0.06fF
C18049 VP.n10654 a_400_38200# 0.06fF
C18050 VP.n10655 a_400_38200# 0.07fF
C18051 VP.n10656 a_400_38200# 0.03fF
C18052 VP.n10657 a_400_38200# 0.05fF
C18053 VP.n10658 a_400_38200# 0.07fF
C18054 VP.n10659 a_400_38200# 0.57fF
C18055 VP.n10660 a_400_38200# 82.60fF
C18056 VP.n10661 a_400_38200# 82.60fF
C18057 VP.n10662 a_400_38200# 0.88fF
C18058 VP.n10663 a_400_38200# 0.26fF
C18059 VP.n10664 a_400_38200# 1.35fF
C18060 VP.n10665 a_400_38200# 0.88fF
C18061 VP.n10666 a_400_38200# 0.10fF
C18062 VP.n10667 a_400_38200# 3.02fF
C18063 VP.t0 a_400_38200# 15.72fF
C18064 VP.n10668 a_400_38200# 1.15fF
C18065 VP.n10670 a_400_38200# 13.70fF
C18066 VP.n10672 a_400_38200# 1.99fF
C18067 VP.n10673 a_400_38200# 4.39fF
C18068 VP.n10674 a_400_38200# 1.88fF
C18069 VP.n10675 a_400_38200# 0.92fF
C18070 VP.n10676 a_400_38200# 0.11fF
C18071 VP.n10677 a_400_38200# 0.24fF
C18072 VP.n10678 a_400_38200# 0.13fF
C18073 VP.n10679 a_400_38200# 0.13fF
C18074 VP.n10680 a_400_38200# 0.24fF
C18075 VP.n10681 a_400_38200# 0.44fF
C18076 VP.n10682 a_400_38200# 0.10fF
C18077 VP.n10683 a_400_38200# 0.12fF
C18078 VP.n10684 a_400_38200# 0.08fF
C18079 VP.n10685 a_400_38200# 0.08fF
C18080 VP.n10686 a_400_38200# 0.06fF
C18081 VP.n10687 a_400_38200# 0.51fF
C18082 VP.n10688 a_400_38200# 0.12fF
C18083 VP.t1209 a_400_38200# 0.02fF
C18084 VP.n10689 a_400_38200# 0.14fF
C18085 VP.n10691 a_400_38200# 0.09fF
C18086 VP.n10692 a_400_38200# 0.06fF
C18087 VP.n10693 a_400_38200# 0.06fF
C18088 VP.n10694 a_400_38200# 0.03fF
C18089 VP.n10696 a_400_38200# 1.45fF
C18090 VP.n10697 a_400_38200# 0.19fF
C18091 VP.n10698 a_400_38200# 0.04fF
C18092 VP.n10699 a_400_38200# 0.02fF
C18093 VP.n10700 a_400_38200# 0.06fF
C18094 VP.n10701 a_400_38200# 0.72fF
C18095 VP.n10702 a_400_38200# 1.81fF
C18096 VP.n10703 a_400_38200# 0.12fF
C18097 VP.t762 a_400_38200# 0.02fF
C18098 VP.n10704 a_400_38200# 0.14fF
C18099 VP.t1349 a_400_38200# 0.02fF
C18100 VP.n10706 a_400_38200# 0.24fF
C18101 VP.n10707 a_400_38200# 0.35fF
C18102 VP.n10708 a_400_38200# 0.60fF
C18103 VP.n10709 a_400_38200# 2.97fF
C18104 VP.n10710 a_400_38200# 2.30fF
C18105 VP.t924 a_400_38200# 0.02fF
C18106 VP.n10711 a_400_38200# 0.24fF
C18107 VP.n10712 a_400_38200# 0.91fF
C18108 VP.n10713 a_400_38200# 0.05fF
C18109 VP.t1164 a_400_38200# 0.02fF
C18110 VP.n10714 a_400_38200# 0.12fF
C18111 VP.n10715 a_400_38200# 0.14fF
C18112 VP.n10717 a_400_38200# 0.06fF
C18113 VP.n10718 a_400_38200# 0.25fF
C18114 VP.n10719 a_400_38200# 0.45fF
C18115 VP.n10720 a_400_38200# 0.03fF
C18116 VP.n10721 a_400_38200# 0.05fF
C18117 VP.n10722 a_400_38200# 0.07fF
C18118 VP.n10723 a_400_38200# 0.06fF
C18119 VP.n10724 a_400_38200# 0.06fF
C18120 VP.n10725 a_400_38200# 0.19fF
C18121 VP.n10726 a_400_38200# 0.59fF
C18122 VP.n10727 a_400_38200# 0.34fF
C18123 VP.n10728 a_400_38200# 0.09fF
C18124 VP.n10729 a_400_38200# 0.05fF
C18125 VP.n10730 a_400_38200# 0.30fF
C18126 VP.n10731 a_400_38200# 1.93fF
C18127 VP.n10732 a_400_38200# 0.12fF
C18128 VP.t309 a_400_38200# 0.02fF
C18129 VP.n10733 a_400_38200# 0.14fF
C18130 VP.t903 a_400_38200# 0.02fF
C18131 VP.n10735 a_400_38200# 0.24fF
C18132 VP.n10736 a_400_38200# 0.35fF
C18133 VP.n10737 a_400_38200# 0.60fF
C18134 VP.n10738 a_400_38200# 2.18fF
C18135 VP.n10739 a_400_38200# 2.04fF
C18136 VP.t475 a_400_38200# 0.02fF
C18137 VP.n10740 a_400_38200# 0.24fF
C18138 VP.n10741 a_400_38200# 0.91fF
C18139 VP.n10742 a_400_38200# 0.05fF
C18140 VP.t714 a_400_38200# 0.02fF
C18141 VP.n10743 a_400_38200# 0.12fF
C18142 VP.n10744 a_400_38200# 0.14fF
C18143 VP.n10746 a_400_38200# 0.24fF
C18144 VP.t707 a_400_38200# 0.02fF
C18145 VP.n10747 a_400_38200# 0.36fF
C18146 VP.n10748 a_400_38200# 0.36fF
C18147 VP.n10749 a_400_38200# 0.67fF
C18148 VP.n10750 a_400_38200# 1.82fF
C18149 VP.n10751 a_400_38200# 2.85fF
C18150 VP.n10752 a_400_38200# 2.97fF
C18151 VP.n10753 a_400_38200# 1.52fF
C18152 VP.n10754 a_400_38200# 0.24fF
C18153 VP.t1138 a_400_38200# 0.02fF
C18154 VP.n10755 a_400_38200# 0.35fF
C18155 VP.n10756 a_400_38200# 0.63fF
C18156 VP.n10757 a_400_38200# 0.40fF
C18157 VP.n10758 a_400_38200# 0.40fF
C18158 VP.n10759 a_400_38200# 0.12fF
C18159 VP.t629 a_400_38200# 0.02fF
C18160 VP.n10760 a_400_38200# 0.14fF
C18161 VP.t971 a_400_38200# 0.02fF
C18162 VP.n10762 a_400_38200# 0.12fF
C18163 VP.n10763 a_400_38200# 0.14fF
C18164 VP.n10765 a_400_38200# 1.93fF
C18165 VP.n10766 a_400_38200# 2.18fF
C18166 VP.t769 a_400_38200# 0.02fF
C18167 VP.n10767 a_400_38200# 0.24fF
C18168 VP.n10768 a_400_38200# 0.35fF
C18169 VP.n10769 a_400_38200# 0.60fF
C18170 VP.n10770 a_400_38200# 0.12fF
C18171 VP.t175 a_400_38200# 0.02fF
C18172 VP.n10771 a_400_38200# 0.14fF
C18173 VP.n10773 a_400_38200# 0.04fF
C18174 VP.n10774 a_400_38200# 0.02fF
C18175 VP.n10775 a_400_38200# 0.06fF
C18176 VP.n10776 a_400_38200# 0.30fF
C18177 VP.n10777 a_400_38200# 0.11fF
C18178 VP.n10778 a_400_38200# 0.05fF
C18179 VP.n10779 a_400_38200# 0.28fF
C18180 VP.n10780 a_400_38200# 0.06fF
C18181 VP.n10781 a_400_38200# 0.03fF
C18182 VP.n10782 a_400_38200# 0.15fF
C18183 VP.n10783 a_400_38200# 0.08fF
C18184 VP.n10784 a_400_38200# 0.14fF
C18185 VP.n10785 a_400_38200# 0.06fF
C18186 VP.n10786 a_400_38200# 0.06fF
C18187 VP.n10787 a_400_38200# 0.03fF
C18188 VP.n10788 a_400_38200# 0.05fF
C18189 VP.n10789 a_400_38200# 0.07fF
C18190 VP.n10790 a_400_38200# 0.19fF
C18191 VP.n10791 a_400_38200# 0.59fF
C18192 VP.n10792 a_400_38200# 0.34fF
C18193 VP.n10793 a_400_38200# 2.04fF
C18194 VP.t340 a_400_38200# 0.02fF
C18195 VP.n10794 a_400_38200# 0.24fF
C18196 VP.n10795 a_400_38200# 0.91fF
C18197 VP.n10796 a_400_38200# 0.05fF
C18198 VP.t523 a_400_38200# 0.02fF
C18199 VP.n10797 a_400_38200# 0.12fF
C18200 VP.n10798 a_400_38200# 0.14fF
C18201 VP.n10800 a_400_38200# 3.10fF
C18202 VP.n10801 a_400_38200# 1.82fF
C18203 VP.n10802 a_400_38200# 0.12fF
C18204 VP.t1025 a_400_38200# 0.02fF
C18205 VP.n10803 a_400_38200# 0.14fF
C18206 VP.t316 a_400_38200# 0.02fF
C18207 VP.n10805 a_400_38200# 0.24fF
C18208 VP.n10806 a_400_38200# 0.35fF
C18209 VP.n10807 a_400_38200# 0.60fF
C18210 VP.n10808 a_400_38200# 2.97fF
C18211 VP.n10809 a_400_38200# 2.76fF
C18212 VP.t1186 a_400_38200# 0.02fF
C18213 VP.n10810 a_400_38200# 0.24fF
C18214 VP.n10811 a_400_38200# 0.91fF
C18215 VP.n10812 a_400_38200# 0.05fF
C18216 VP.t43 a_400_38200# 0.02fF
C18217 VP.n10813 a_400_38200# 0.12fF
C18218 VP.n10814 a_400_38200# 0.14fF
C18219 VP.n10816 a_400_38200# 1.93fF
C18220 VP.n10817 a_400_38200# 2.18fF
C18221 VP.t1159 a_400_38200# 0.02fF
C18222 VP.n10818 a_400_38200# 0.24fF
C18223 VP.n10819 a_400_38200# 0.35fF
C18224 VP.n10820 a_400_38200# 0.60fF
C18225 VP.n10821 a_400_38200# 0.12fF
C18226 VP.t577 a_400_38200# 0.02fF
C18227 VP.n10822 a_400_38200# 0.14fF
C18228 VP.n10824 a_400_38200# 0.04fF
C18229 VP.n10825 a_400_38200# 0.02fF
C18230 VP.n10826 a_400_38200# 0.06fF
C18231 VP.n10827 a_400_38200# 0.30fF
C18232 VP.n10828 a_400_38200# 0.11fF
C18233 VP.n10829 a_400_38200# 0.05fF
C18234 VP.n10830 a_400_38200# 0.28fF
C18235 VP.n10831 a_400_38200# 0.06fF
C18236 VP.n10832 a_400_38200# 0.03fF
C18237 VP.n10833 a_400_38200# 0.15fF
C18238 VP.n10834 a_400_38200# 0.08fF
C18239 VP.n10835 a_400_38200# 0.14fF
C18240 VP.n10836 a_400_38200# 0.06fF
C18241 VP.n10837 a_400_38200# 0.06fF
C18242 VP.n10838 a_400_38200# 0.03fF
C18243 VP.n10839 a_400_38200# 0.05fF
C18244 VP.n10840 a_400_38200# 0.07fF
C18245 VP.n10841 a_400_38200# 0.19fF
C18246 VP.n10842 a_400_38200# 0.59fF
C18247 VP.n10843 a_400_38200# 0.34fF
C18248 VP.n10844 a_400_38200# 2.04fF
C18249 VP.t734 a_400_38200# 0.02fF
C18250 VP.n10845 a_400_38200# 0.24fF
C18251 VP.n10846 a_400_38200# 0.91fF
C18252 VP.n10847 a_400_38200# 0.05fF
C18253 VP.t932 a_400_38200# 0.02fF
C18254 VP.n10848 a_400_38200# 0.12fF
C18255 VP.n10849 a_400_38200# 0.14fF
C18256 VP.n10851 a_400_38200# 3.10fF
C18257 VP.n10852 a_400_38200# 1.82fF
C18258 VP.n10853 a_400_38200# 0.12fF
C18259 VP.t110 a_400_38200# 0.02fF
C18260 VP.n10854 a_400_38200# 0.14fF
C18261 VP.t710 a_400_38200# 0.02fF
C18262 VP.n10856 a_400_38200# 0.24fF
C18263 VP.n10857 a_400_38200# 0.35fF
C18264 VP.n10858 a_400_38200# 0.60fF
C18265 VP.n10859 a_400_38200# 2.97fF
C18266 VP.n10860 a_400_38200# 2.76fF
C18267 VP.t282 a_400_38200# 0.02fF
C18268 VP.n10861 a_400_38200# 0.24fF
C18269 VP.n10862 a_400_38200# 0.91fF
C18270 VP.n10863 a_400_38200# 0.05fF
C18271 VP.t486 a_400_38200# 0.02fF
C18272 VP.n10864 a_400_38200# 0.12fF
C18273 VP.n10865 a_400_38200# 0.14fF
C18274 VP.n10867 a_400_38200# 1.93fF
C18275 VP.n10868 a_400_38200# 2.18fF
C18276 VP.t264 a_400_38200# 0.02fF
C18277 VP.n10869 a_400_38200# 0.24fF
C18278 VP.n10870 a_400_38200# 0.35fF
C18279 VP.n10871 a_400_38200# 0.60fF
C18280 VP.n10872 a_400_38200# 0.12fF
C18281 VP.t984 a_400_38200# 0.02fF
C18282 VP.n10873 a_400_38200# 0.14fF
C18283 VP.n10875 a_400_38200# 0.04fF
C18284 VP.n10876 a_400_38200# 0.02fF
C18285 VP.n10877 a_400_38200# 0.06fF
C18286 VP.n10878 a_400_38200# 0.30fF
C18287 VP.n10879 a_400_38200# 0.11fF
C18288 VP.n10880 a_400_38200# 0.05fF
C18289 VP.n10881 a_400_38200# 0.28fF
C18290 VP.n10882 a_400_38200# 0.06fF
C18291 VP.n10883 a_400_38200# 0.03fF
C18292 VP.n10884 a_400_38200# 0.15fF
C18293 VP.n10885 a_400_38200# 0.08fF
C18294 VP.n10886 a_400_38200# 0.14fF
C18295 VP.n10887 a_400_38200# 0.06fF
C18296 VP.n10888 a_400_38200# 0.06fF
C18297 VP.n10889 a_400_38200# 0.03fF
C18298 VP.n10890 a_400_38200# 0.05fF
C18299 VP.n10891 a_400_38200# 0.07fF
C18300 VP.n10892 a_400_38200# 0.19fF
C18301 VP.n10893 a_400_38200# 0.59fF
C18302 VP.n10894 a_400_38200# 0.34fF
C18303 VP.n10895 a_400_38200# 2.04fF
C18304 VP.t1136 a_400_38200# 0.02fF
C18305 VP.n10896 a_400_38200# 0.24fF
C18306 VP.n10897 a_400_38200# 0.91fF
C18307 VP.n10898 a_400_38200# 0.05fF
C18308 VP.t1334 a_400_38200# 0.02fF
C18309 VP.n10899 a_400_38200# 0.12fF
C18310 VP.n10900 a_400_38200# 0.14fF
C18311 VP.n10902 a_400_38200# 3.10fF
C18312 VP.n10903 a_400_38200# 1.82fF
C18313 VP.n10904 a_400_38200# 0.12fF
C18314 VP.t536 a_400_38200# 0.02fF
C18315 VP.n10905 a_400_38200# 0.14fF
C18316 VP.t1119 a_400_38200# 0.02fF
C18317 VP.n10907 a_400_38200# 0.24fF
C18318 VP.n10908 a_400_38200# 0.35fF
C18319 VP.n10909 a_400_38200# 0.60fF
C18320 VP.n10910 a_400_38200# 2.97fF
C18321 VP.n10911 a_400_38200# 2.76fF
C18322 VP.t687 a_400_38200# 0.02fF
C18323 VP.n10912 a_400_38200# 0.24fF
C18324 VP.n10913 a_400_38200# 0.91fF
C18325 VP.n10914 a_400_38200# 0.05fF
C18326 VP.t953 a_400_38200# 0.02fF
C18327 VP.n10915 a_400_38200# 0.12fF
C18328 VP.n10916 a_400_38200# 0.14fF
C18329 VP.n10918 a_400_38200# 1.93fF
C18330 VP.n10919 a_400_38200# 2.97fF
C18331 VP.t674 a_400_38200# 0.02fF
C18332 VP.n10920 a_400_38200# 0.24fF
C18333 VP.n10921 a_400_38200# 0.35fF
C18334 VP.n10922 a_400_38200# 0.60fF
C18335 VP.n10923 a_400_38200# 0.12fF
C18336 VP.t62 a_400_38200# 0.02fF
C18337 VP.n10924 a_400_38200# 0.14fF
C18338 VP.n10926 a_400_38200# 0.04fF
C18339 VP.n10927 a_400_38200# 0.02fF
C18340 VP.n10928 a_400_38200# 0.06fF
C18341 VP.n10929 a_400_38200# 0.30fF
C18342 VP.n10930 a_400_38200# 0.11fF
C18343 VP.n10931 a_400_38200# 0.05fF
C18344 VP.n10932 a_400_38200# 0.28fF
C18345 VP.n10933 a_400_38200# 0.06fF
C18346 VP.n10934 a_400_38200# 0.03fF
C18347 VP.n10935 a_400_38200# 0.15fF
C18348 VP.n10936 a_400_38200# 0.08fF
C18349 VP.n10937 a_400_38200# 0.14fF
C18350 VP.n10938 a_400_38200# 0.06fF
C18351 VP.n10939 a_400_38200# 0.06fF
C18352 VP.n10940 a_400_38200# 0.03fF
C18353 VP.n10941 a_400_38200# 0.05fF
C18354 VP.n10942 a_400_38200# 0.07fF
C18355 VP.n10943 a_400_38200# 0.19fF
C18356 VP.n10944 a_400_38200# 0.59fF
C18357 VP.n10945 a_400_38200# 0.34fF
C18358 VP.n10946 a_400_38200# 2.20fF
C18359 VP.t243 a_400_38200# 0.02fF
C18360 VP.n10947 a_400_38200# 0.24fF
C18361 VP.n10948 a_400_38200# 0.91fF
C18362 VP.n10949 a_400_38200# 0.05fF
C18363 VP.t507 a_400_38200# 0.02fF
C18364 VP.n10950 a_400_38200# 0.12fF
C18365 VP.n10951 a_400_38200# 0.14fF
C18366 VP.n10953 a_400_38200# 1.88fF
C18367 VP.t483 a_400_38200# 0.02fF
C18368 VP.n10954 a_400_38200# 0.64fF
C18369 VP.n10955 a_400_38200# 0.60fF
C18370 VP.n10956 a_400_38200# 0.88fF
C18371 VP.n10957 a_400_38200# 0.48fF
C18372 VP.n10958 a_400_38200# 0.88fF
C18373 VP.n10959 a_400_38200# 0.60fF
C18374 VP.n10960 a_400_38200# 2.33fF
C18375 VP.n10961 a_400_38200# 0.59fF
C18376 VP.n10962 a_400_38200# 0.02fF
C18377 VP.n10963 a_400_38200# 0.96fF
C18378 VP.t167 a_400_38200# 15.72fF
C18379 VP.n10964 a_400_38200# 15.42fF
C18380 VP.n10966 a_400_38200# 0.38fF
C18381 VP.n10967 a_400_38200# 0.23fF
C18382 VP.n10968 a_400_38200# 3.40fF
C18383 VP.n10969 a_400_38200# 1.98fF
C18384 VP.n10970 a_400_38200# 4.90fF
C18385 VP.t1 a_400_38200# 0.02fF
C18386 VP.n10971 a_400_38200# 1.19fF
C18387 VP.n10972 a_400_38200# 0.05fF
C18388 VP.t300 a_400_38200# 0.02fF
C18389 VP.n10973 a_400_38200# 0.01fF
C18390 VP.n10974 a_400_38200# 0.26fF
C18391 VP.n10976 a_400_38200# 15.28fF
C18392 VP.n10977 a_400_38200# 1.93fF
C18393 VP.n10978 a_400_38200# 2.62fF
C18394 VP.t228 a_400_38200# 0.02fF
C18395 VP.n10979 a_400_38200# 0.24fF
C18396 VP.n10980 a_400_38200# 0.35fF
C18397 VP.n10981 a_400_38200# 0.60fF
C18398 VP.n10982 a_400_38200# 0.12fF
C18399 VP.t945 a_400_38200# 0.02fF
C18400 VP.n10983 a_400_38200# 0.14fF
C18401 VP.n10985 a_400_38200# 0.04fF
C18402 VP.n10986 a_400_38200# 0.02fF
C18403 VP.n10987 a_400_38200# 0.06fF
C18404 VP.n10988 a_400_38200# 0.30fF
C18405 VP.n10989 a_400_38200# 0.07fF
C18406 VP.n10990 a_400_38200# 0.05fF
C18407 VP.n10991 a_400_38200# 0.26fF
C18408 VP.n10992 a_400_38200# 0.06fF
C18409 VP.n10993 a_400_38200# 0.03fF
C18410 VP.n10994 a_400_38200# 0.15fF
C18411 VP.n10995 a_400_38200# 0.08fF
C18412 VP.n10996 a_400_38200# 0.14fF
C18413 VP.n10997 a_400_38200# 0.06fF
C18414 VP.n10998 a_400_38200# 0.06fF
C18415 VP.n10999 a_400_38200# 0.03fF
C18416 VP.n11000 a_400_38200# 0.05fF
C18417 VP.n11001 a_400_38200# 0.07fF
C18418 VP.n11002 a_400_38200# 0.19fF
C18419 VP.n11003 a_400_38200# 0.59fF
C18420 VP.n11004 a_400_38200# 0.34fF
C18421 VP.n11005 a_400_38200# 2.18fF
C18422 VP.t17 a_400_38200# 0.02fF
C18423 VP.n11006 a_400_38200# 0.12fF
C18424 VP.n11007 a_400_38200# 0.14fF
C18425 VP.t1097 a_400_38200# 0.02fF
C18426 VP.n11009 a_400_38200# 0.24fF
C18427 VP.n11010 a_400_38200# 0.91fF
C18428 VP.n11011 a_400_38200# 0.05fF
C18429 VP.t16 a_400_38200# 34.79fF
C18430 VP.t322 a_400_38200# 0.02fF
C18431 VP.n11012 a_400_38200# 0.12fF
C18432 VP.n11013 a_400_38200# 0.14fF
C18433 VP.t30 a_400_38200# 0.02fF
C18434 VP.n11015 a_400_38200# 0.24fF
C18435 VP.n11016 a_400_38200# 0.91fF
C18436 VP.n11017 a_400_38200# 0.05fF
C18437 VP.t498 a_400_38200# 0.02fF
C18438 VP.n11018 a_400_38200# 0.24fF
C18439 VP.n11019 a_400_38200# 0.35fF
C18440 VP.n11020 a_400_38200# 0.60fF
C18441 VP.n11021 a_400_38200# 0.04fF
C18442 VP.n11022 a_400_38200# 0.02fF
C18443 VP.n11023 a_400_38200# 0.06fF
C18444 VP.n11024 a_400_38200# 0.45fF
C18445 VP.n11025 a_400_38200# 0.10fF
C18446 VP.n11026 a_400_38200# 0.17fF
C18447 VP.n11027 a_400_38200# 0.10fF
C18448 VP.n11028 a_400_38200# 0.04fF
C18449 VP.n11029 a_400_38200# 0.09fF
C18450 VP.n11030 a_400_38200# 0.45fF
C18451 VP.n11031 a_400_38200# 0.10fF
C18452 VP.n11032 a_400_38200# 1.65fF
C18453 VP.n11033 a_400_38200# 2.24fF
C18454 VP.n11034 a_400_38200# 2.43fF
C18455 VP.n11035 a_400_38200# 40.92fF
C18456 VP.n11036 a_400_38200# 26.56fF
C18457 VP.n11037 a_400_38200# 26.56fF
C18458 VP.n11038 a_400_38200# 26.56fF
C18459 VP.n11039 a_400_38200# 26.56fF
C18460 VP.n11040 a_400_38200# 26.56fF
C18461 VP.n11041 a_400_38200# 26.56fF
C18462 VP.n11042 a_400_38200# 26.56fF
C18463 VP.n11043 a_400_38200# 26.56fF
C18464 VP.n11044 a_400_38200# 26.56fF
C18465 VP.n11045 a_400_38200# 26.56fF
C18466 VP.n11046 a_400_38200# 95.01fF
C18467 VP.n11047 a_400_38200# 81.17fF
C18468 VP.n11048 a_400_38200# 26.68fF
C18469 VP.n11049 a_400_38200# 26.70fF
C18470 VP.n11050 a_400_38200# 26.68fF
C18471 VP.n11051 a_400_38200# 26.68fF
C18472 VP.n11052 a_400_38200# 26.68fF
C18473 VP.n11053 a_400_38200# 26.68fF
C18474 VP.n11054 a_400_38200# 26.68fF
C18475 VP.n11055 a_400_38200# 26.68fF
C18476 VP.n11056 a_400_38200# 26.68fF
C18477 VP.n11057 a_400_38200# 26.68fF
C18478 VP.n11058 a_400_38200# 25.05fF
.ends

