magic
tech sky130A
timestamp 1675433101
<< error_p >>
rect 507 607 610 663
rect 497 586 1575 607
rect 48 553 1575 586
rect 48 550 81 553
rect 345 550 385 553
rect 497 550 1575 553
rect 81 517 519 550
rect 775 517 1075 550
rect -36 469 0 502
rect -36 205 -3 469
rect 0 205 33 469
rect 156 447 160 517
rect -36 165 33 205
rect -36 43 -3 165
rect 0 160 33 165
rect 0 156 156 160
rect 0 43 160 156
rect -113 29 160 43
rect -113 0 519 29
rect 775 0 1075 33
rect -113 -2 552 0
rect -113 -113 43 -2
rect 48 -33 552 -2
rect 742 -33 1108 0
<< nwell >>
rect 0 0 1175 550
<< mvpmos >>
rect 81 500 519 550
rect 0 31 50 469
<< mvpdiff >>
rect 81 550 519 553
rect 81 494 519 500
rect 81 477 87 494
rect 513 477 519 494
rect 81 471 519 477
rect 81 469 114 471
rect -3 31 0 469
rect 50 463 114 469
rect 50 37 56 463
rect 73 436 114 463
rect 73 64 79 436
rect 73 37 114 64
rect 50 31 114 37
rect 81 29 114 31
rect 81 23 519 29
rect 81 6 87 23
rect 513 6 519 23
rect 81 0 519 6
<< mvpdiffc >>
rect 87 477 513 494
rect 56 37 73 463
rect 87 6 513 23
<< mvnsubdiff >>
rect 775 19 787 550
rect 1063 19 1075 550
rect 775 0 1075 19
<< mvnsubdiffcont >>
rect 787 19 1063 550
<< poly >>
rect 0 542 81 550
rect 0 508 8 542
rect 42 508 81 542
rect 0 500 81 508
rect 519 542 600 550
rect 519 508 558 542
rect 592 508 600 542
rect 519 500 600 508
rect 0 469 50 500
rect 0 0 50 31
rect 550 0 600 500
<< polycont >>
rect 8 508 42 542
rect 558 508 592 542
<< locali >>
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 79 477 87 494
rect 513 477 521 494
rect 79 471 114 477
rect 56 463 114 471
rect 73 436 114 463
rect 73 37 114 64
rect 56 29 114 37
rect 79 23 114 29
rect 79 6 87 23
rect 513 6 521 23
rect 775 19 787 550
rect 1063 19 1075 550
rect 775 0 1075 19
<< viali >>
rect 8 508 42 542
rect 558 508 592 542
rect 87 477 513 494
rect 56 37 73 463
rect 87 6 513 23
rect 787 19 1063 550
<< metal1 >>
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 81 494 519 497
rect 81 477 87 494
rect 513 477 519 494
rect 81 474 519 477
rect 76 469 524 474
rect 53 463 524 469
rect 53 37 56 463
rect 73 415 524 463
rect 73 85 135 415
rect 465 85 524 415
rect 73 37 524 85
rect 53 31 524 37
rect 76 26 524 31
rect 81 23 519 26
rect 81 6 87 23
rect 513 6 519 23
rect 81 3 519 6
rect 775 19 787 550
rect 1063 19 1075 550
rect 775 0 1075 19
<< via1 >>
rect 8 508 42 542
rect 558 508 592 542
rect 135 85 465 415
<< metal2 >>
rect 0 542 775 550
rect 0 508 8 542
rect 42 508 558 542
rect 592 508 775 542
rect 0 500 775 508
rect 0 0 50 500
rect 125 415 475 425
rect 125 85 135 415
rect 465 85 475 415
rect 125 75 475 85
rect 550 0 775 500
<< via2 >>
rect 240 190 360 310
<< metal3 >>
rect 0 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 1575 550
rect 0 412 266 510
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 1575 510
rect 0 324 364 412
tri 0 226 98 324 ne
rect 98 314 364 324
tri 364 314 462 412 sw
rect 98 310 1075 314
rect 98 226 240 310
tri 0 186 40 226 sw
tri 98 186 138 226 ne
rect 138 190 240 226
rect 360 190 1075 310
rect 138 186 1075 190
rect 0 88 40 186
tri 40 88 138 186 sw
tri 138 88 236 186 ne
rect 236 88 1075 186
rect 0 0 138 88
tri 138 0 226 88 sw
tri 236 0 324 88 ne
rect 324 0 1075 88
<< via3 >>
rect 240 190 360 310
<< metal4 >>
rect 0 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 1575 550
rect 0 412 266 510
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 1575 510
rect 0 324 364 412
tri 0 226 98 324 ne
rect 98 314 364 324
tri 364 314 462 412 sw
rect 98 310 1075 314
rect 98 226 240 310
tri 0 186 40 226 sw
tri 98 186 138 226 ne
rect 138 190 240 226
rect 360 190 1075 310
rect 138 186 1075 190
rect 0 88 40 186
tri 40 88 138 186 sw
tri 138 88 236 186 ne
rect 236 88 1075 186
rect 0 0 138 88
tri 138 0 226 88 sw
tri 236 0 324 88 ne
rect 324 0 1075 88
<< via4 >>
rect 240 190 360 310
<< metal5 >>
rect 0 447 156 550
tri 156 447 259 550 sw
tri 394 447 497 550 ne
rect 497 447 1575 550
rect 0 394 259 447
tri 0 156 238 394 ne
rect 238 310 259 394
tri 259 310 396 447 sw
rect 238 190 240 310
rect 360 208 396 310
tri 396 208 498 310 sw
rect 360 190 1075 208
rect 238 156 1075 190
tri 0 0 156 156 sw
tri 238 0 394 156 ne
rect 394 0 1075 156
<< end >>
