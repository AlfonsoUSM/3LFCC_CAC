**.subckt postlayout_cap_pmos
.include pmos_flat_12x12.spice
VG VP GND PULSE(0 {VGS} 20n 0 0 100n 120n)
.save i(vg)
VSS VSS GND 0
.save i(vss)
R1 G VP 100 m=1
VG1 VP2 GND {VGS}
.save i(vg1)
VX PW GND 0
XU1 G VP2 VSS PW pmos_flat_12x12
**** begin user architecture code


.param VGS = 5
.option temp=70
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.control
compose voltage values (2.5) 5
foreach volt $&voltage
alterparam VGS=$volt
reset
save v(G)
tran 50f 120n
wrdata SPICE_files/PMOS/POSTLAYOUT_CAP/PMOS_cap_calc_POSTLAYOUT.txt v(G)
set appendwrite
end

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
.control
quit
.endc