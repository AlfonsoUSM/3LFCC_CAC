magic
tech sky130A
timestamp 1674760439
<< pwell >>
rect -1125 -1175 1175 1125
<< mvnmos >>
rect 0 31 50 469
rect -469 -50 -31 0
rect 81 -50 519 0
rect 0 -519 50 -81
<< mvndiff >>
rect 79 469 521 471
rect -29 463 0 469
rect -29 64 -23 463
rect -64 37 -23 64
rect -6 37 0 463
rect -64 31 0 37
rect 50 463 521 469
rect 50 37 56 463
rect 73 415 521 463
rect 73 85 135 415
rect 465 85 521 415
rect 73 37 521 85
rect 50 31 521 37
rect -64 29 -31 31
rect -469 23 -31 29
rect -469 6 -463 23
rect -37 6 -31 23
rect -469 0 -31 6
rect 79 29 521 31
rect 81 23 519 29
rect 81 6 87 23
rect 513 6 519 23
rect 81 0 519 6
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 81 -56 519 -50
rect 81 -73 87 -56
rect 513 -73 519 -56
rect 81 -79 519 -73
rect 81 -81 114 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 50 -87 114 -81
rect 50 -513 56 -87
rect 73 -114 114 -87
rect 73 -513 79 -114
rect 50 -519 79 -513
rect -471 -521 -29 -519
<< mvndiffc >>
rect -23 37 -6 463
rect 56 37 73 463
rect -463 6 -37 23
rect 87 6 513 23
rect -463 -73 -37 -56
rect 87 -73 513 -56
rect -23 -513 -6 -87
rect 56 -513 73 -87
<< mvpsubdiff >>
rect -1025 1013 1075 1025
rect -1025 17 -1013 1013
rect -19 737 0 1013
rect -737 725 787 737
rect -737 17 -725 725
rect -1025 0 -725 17
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect 135 403 465 415
rect 135 97 147 403
rect 453 97 465 403
rect 135 85 465 97
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 775 17 787 725
rect 1063 17 1075 1013
rect 775 0 1075 17
rect 775 -775 787 0
rect -737 -787 787 -775
rect -17 -1063 0 -787
rect 1063 -1063 1075 0
rect -1025 -1075 1075 -1063
<< mvpsubdiffcont >>
rect -1013 737 -19 1013
rect 0 737 1063 1013
rect -1013 17 -737 737
rect -1013 -787 -737 0
rect 147 97 453 403
rect -403 -453 -97 -147
rect 787 17 1063 737
rect 787 -787 1063 0
rect -1013 -1063 -17 -787
rect 0 -1063 1063 -787
<< poly >>
rect -550 542 600 550
rect -550 508 -542 542
rect -508 508 8 542
rect 42 508 558 542
rect 592 508 600 542
rect -550 500 600 508
rect -550 0 -500 500
rect 0 469 50 500
rect 0 0 50 31
rect 550 0 600 500
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -8 81 0
rect -31 -42 8 -8
rect 42 -42 81 -8
rect -31 -50 81 -42
rect 519 -8 600 0
rect 519 -42 558 -8
rect 592 -42 600 -8
rect 519 -50 600 -42
rect -550 -550 -500 -50
rect 0 -81 50 -50
rect 0 -550 50 -519
rect 550 -550 600 -50
rect -550 -558 600 -550
rect -550 -592 -542 -558
rect -508 -592 8 -558
rect 42 -592 558 -558
rect 592 -592 600 -558
rect -550 -600 600 -592
<< polycont >>
rect -542 508 -508 542
rect 8 508 42 542
rect 558 508 592 542
rect -542 -42 -508 -8
rect 8 -42 42 -8
rect 558 -42 592 -8
rect -542 -592 -508 -558
rect 8 -592 42 -558
rect 558 -592 592 -558
<< locali >>
rect -1025 1013 1075 1025
rect -1025 17 -1013 1013
rect -19 737 0 1013
rect -737 725 787 737
rect -737 17 -725 725
rect -550 542 -500 550
rect -550 508 -542 542
rect -508 508 -500 542
rect -550 500 -500 508
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 73 471 527 477
rect -23 463 -6 471
rect -64 37 -23 64
rect -64 29 -6 37
rect 56 463 527 471
rect 73 415 527 463
rect 73 85 135 415
rect 465 85 527 415
rect 73 37 527 85
rect 56 29 527 37
rect -64 23 -29 29
rect 73 23 527 29
rect -1025 0 -725 17
rect -471 6 -463 23
rect -37 6 -29 23
rect 79 6 87 23
rect 513 6 521 23
rect 775 17 787 725
rect 1063 17 1075 1013
rect 775 0 1075 17
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 0 -8 50 0
rect 0 -42 8 -8
rect 42 -42 50 -8
rect 0 -50 50 -42
rect 550 -8 600 0
rect 550 -42 558 -8
rect 592 -42 600 -8
rect 550 -50 600 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 79 -73 87 -56
rect 513 -73 521 -56
rect -477 -79 -23 -73
rect 79 -79 114 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 56 -87 114 -79
rect 73 -114 114 -87
rect 56 -521 73 -513
rect -477 -527 -23 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 0 -558 50 -550
rect 0 -592 8 -558
rect 42 -592 50 -558
rect 0 -600 50 -592
rect 550 -558 600 -550
rect 550 -592 558 -558
rect 592 -592 600 -558
rect 550 -600 600 -592
rect 775 -775 787 0
rect -737 -787 787 -775
rect -17 -1063 0 -787
rect 1063 -1063 1075 0
rect -1025 -1075 1075 -1063
<< viali >>
rect -1013 737 -19 1013
rect 0 737 1063 1013
rect -1013 19 -737 737
rect -542 508 -508 542
rect 8 508 42 542
rect 558 508 592 542
rect -23 37 -6 463
rect 56 37 73 463
rect 135 403 465 415
rect 135 97 147 403
rect 147 97 453 403
rect 453 97 465 403
rect 135 85 465 97
rect -463 6 -37 23
rect 87 6 513 23
rect 787 19 1063 737
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 8 -42 42 -8
rect 558 -42 592 -8
rect -463 -73 -37 -56
rect 87 -73 513 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 56 -513 73 -87
rect -542 -592 -508 -558
rect 8 -592 42 -558
rect 558 -592 592 -558
rect 787 -787 1063 0
rect -1013 -1063 -19 -787
rect 0 -1063 1063 -787
<< metal1 >>
rect -1025 1013 1075 1025
rect -1025 19 -1013 1013
rect -19 737 0 1013
rect -737 725 787 737
rect -737 19 -725 725
rect -550 542 -500 550
rect -550 508 -542 542
rect -508 508 -500 542
rect -550 500 -500 508
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect -474 469 -26 474
rect 76 469 524 474
rect -474 463 -3 469
rect -474 415 -23 463
rect -474 85 -415 415
rect -85 85 -23 415
rect -474 37 -23 85
rect -6 37 -3 463
rect -474 31 -3 37
rect 53 463 524 469
rect 53 37 56 463
rect 73 415 524 463
rect 73 85 135 415
rect 465 85 524 415
rect 73 37 524 85
rect 53 31 524 37
rect -474 26 -26 31
rect 76 26 524 31
rect -1025 0 -725 19
rect -469 23 -31 26
rect -469 6 -463 23
rect -37 6 -31 23
rect -469 3 -31 6
rect 81 23 519 26
rect 81 6 87 23
rect 513 6 519 23
rect 81 3 519 6
rect 775 19 787 725
rect 1063 19 1075 1013
rect 775 0 1075 19
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 0 -8 50 0
rect 0 -42 8 -8
rect 42 -42 50 -8
rect 0 -50 50 -42
rect 550 -8 600 0
rect 550 -42 558 -8
rect 592 -42 600 -8
rect 550 -50 600 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 81 -56 519 -53
rect 81 -73 87 -56
rect 513 -73 519 -56
rect 81 -76 519 -73
rect -474 -81 -26 -76
rect 76 -81 524 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 53 -87 524 -81
rect 53 -513 56 -87
rect 73 -135 524 -87
rect 73 -465 135 -135
rect 465 -465 524 -135
rect 73 -513 524 -465
rect 53 -519 524 -513
rect -474 -524 -26 -519
rect 76 -524 524 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 0 -558 50 -550
rect 0 -592 8 -558
rect 42 -592 50 -558
rect 0 -600 50 -592
rect 550 -558 600 -550
rect 550 -592 558 -558
rect 592 -592 600 -558
rect 550 -600 600 -592
rect 775 -775 787 0
rect -737 -787 787 -775
rect -19 -1063 0 -787
rect 1063 -1063 1075 0
rect -1025 -1075 1075 -1063
<< via1 >>
rect 88 825 188 925
rect -542 508 -508 542
rect 8 508 42 542
rect 558 508 592 542
rect -415 85 -85 415
rect 135 85 465 415
rect 875 38 975 138
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 8 -42 42 -8
rect 558 -42 592 -8
rect -415 -465 -85 -135
rect 135 -465 465 -135
rect -542 -592 -508 -558
rect 8 -592 42 -558
rect 558 -592 592 -558
rect -138 -975 -38 -875
<< metal2 >>
rect 78 925 198 935
rect 78 825 88 925
rect 188 825 198 925
rect 78 815 198 825
rect -725 542 775 725
rect -725 508 -542 542
rect -508 508 8 542
rect 42 508 558 542
rect 592 508 775 542
rect -725 500 775 508
rect -725 0 -500 500
rect -425 415 -75 425
rect -425 85 -415 415
rect -85 85 -75 415
rect -425 75 -75 85
rect 0 0 50 500
rect 125 415 475 425
rect 125 85 135 415
rect 465 85 475 415
rect 125 75 475 85
rect 550 0 775 500
rect 865 138 985 148
rect 865 38 875 138
rect 975 38 985 138
rect 865 28 985 38
rect -725 -8 775 0
rect -725 -42 -542 -8
rect -508 -42 8 -8
rect 42 -42 558 -8
rect 592 -42 775 -8
rect -725 -50 775 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 0 -550 50 -50
rect 125 -135 475 -125
rect 125 -465 135 -135
rect 465 -465 475 -135
rect 125 -475 475 -465
rect 550 -550 775 -50
rect -725 -558 775 -550
rect -725 -592 -542 -558
rect -508 -592 8 -558
rect 42 -592 558 -558
rect 592 -592 775 -558
rect -725 -775 775 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
<< via2 >>
rect 88 825 188 925
rect -310 190 -190 310
rect 240 190 360 310
rect 875 38 975 138
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 240 -360 360 -240
rect -138 -975 -38 -875
<< metal3 >>
rect -638 638 -186 1525
rect -1525 314 -186 638
rect -88 925 364 1025
rect -88 825 88 925
rect 188 825 364 925
rect -88 412 364 825
tri -186 314 -88 412 sw
tri -88 314 10 412 ne
rect 10 314 364 412
tri 364 314 462 412 sw
rect -1525 310 -88 314
rect -1525 190 -310 310
rect -190 226 -88 310
tri -88 226 0 314 sw
tri 10 226 98 314 ne
rect 98 310 1575 314
rect 98 226 240 310
rect -190 190 0 226
rect -1525 186 0 190
tri -412 88 -314 186 ne
rect -314 138 0 186
tri 0 138 88 226 sw
tri 98 138 186 226 ne
rect 186 190 240 226
rect 360 190 1575 310
rect 186 138 1575 190
rect -314 88 88 138
rect -1025 0 -412 88
tri -412 0 -324 88 sw
tri -314 0 -226 88 ne
rect -226 58 88 88
tri 88 58 168 138 sw
tri 186 58 266 138 ne
rect 266 58 875 138
rect -226 0 168 58
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 168 0
tri 168 -40 266 58 sw
tri 266 -40 364 58 ne
rect 364 38 875 58
rect 975 38 1575 138
rect 364 -40 1575 38
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 266 -40
tri 266 -138 364 -40 sw
tri 364 -138 462 -40 ne
rect 462 -138 1575 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -236 10 -138 ne
rect 10 -236 364 -138
tri 364 -236 462 -138 sw
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
tri 10 -324 98 -236 ne
rect 98 -240 1075 -236
rect 98 -324 240 -240
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri 0 -364 40 -324 sw
tri 98 -364 138 -324 ne
rect 138 -360 240 -324
rect 360 -360 1075 -240
rect 138 -364 1075 -360
tri -412 -462 -314 -364 ne
rect -314 -462 40 -364
tri 40 -462 138 -364 sw
tri 138 -462 236 -364 ne
rect -314 -875 138 -462
rect -314 -975 -138 -875
rect -38 -975 138 -875
rect -314 -1575 138 -975
rect 236 -688 1075 -364
rect 236 -1075 688 -688
<< via3 >>
rect 88 825 188 925
rect -310 190 -190 310
rect 240 190 360 310
rect 875 38 975 138
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 240 -360 360 -240
rect -138 -975 -38 -875
<< metal4 >>
rect -638 638 -186 1525
rect -1525 314 -186 638
rect -88 925 364 1025
rect -88 825 88 925
rect 188 825 364 925
rect -88 412 364 825
tri -186 314 -88 412 sw
tri -88 314 10 412 ne
rect 10 314 364 412
tri 364 314 462 412 sw
rect -1525 310 -88 314
rect -1525 190 -310 310
rect -190 226 -88 310
tri -88 226 0 314 sw
tri 10 226 98 314 ne
rect 98 310 1575 314
rect 98 226 240 310
rect -190 190 0 226
rect -1525 186 0 190
tri -412 88 -314 186 ne
rect -314 138 0 186
tri 0 138 88 226 sw
tri 98 138 186 226 ne
rect 186 190 240 226
rect 360 190 1575 310
rect 186 138 1575 190
rect -314 88 88 138
rect -1025 0 -412 88
tri -412 0 -324 88 sw
tri -314 0 -226 88 ne
rect -226 58 88 88
tri 88 58 168 138 sw
tri 186 58 266 138 ne
rect 266 58 875 138
rect -226 0 168 58
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 168 0
tri 168 -40 266 58 sw
tri 266 -40 364 58 ne
rect 364 38 875 58
rect 975 38 1575 138
rect 364 -40 1575 38
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 266 -40
tri 266 -138 364 -40 sw
tri 364 -138 462 -40 ne
rect 462 -138 1575 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -236 10 -138 ne
rect 10 -236 364 -138
tri 364 -236 462 -138 sw
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
tri 10 -324 98 -236 ne
rect 98 -240 1075 -236
rect 98 -324 240 -240
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri 0 -364 40 -324 sw
tri 98 -364 138 -324 ne
rect 138 -360 240 -324
rect 360 -360 1075 -240
rect 138 -364 1075 -360
tri -412 -462 -314 -364 ne
rect -314 -462 40 -364
tri 40 -462 138 -364 sw
tri 138 -462 236 -364 ne
rect -314 -875 138 -462
rect -314 -975 -138 -875
rect -38 -975 138 -875
rect -314 -1575 138 -975
rect 236 -688 1075 -364
rect 236 -1075 688 -688
<< via4 >>
rect -310 190 -190 310
rect 240 190 360 310
rect -310 -360 -190 -240
rect 240 -360 360 -240
<< metal5 >>
rect -603 603 -292 1525
rect -1525 310 -292 603
tri -292 310 -154 448 sw
rect -53 447 258 1025
tri -53 310 84 447 ne
rect 84 310 258 447
tri 258 310 396 448 sw
rect -1525 292 -310 310
tri -448 190 -346 292 ne
rect -346 190 -310 292
rect -190 190 -154 310
rect -1025 0 -447 53
tri -447 0 -394 53 sw
tri -346 0 -156 190 ne
rect -156 156 -154 190
tri -154 156 0 310 sw
tri 84 156 238 310 ne
rect 238 190 240 310
rect 360 208 396 310
tri 396 208 498 310 sw
rect 360 190 1575 208
rect 238 156 1575 190
rect -156 0 0 156
tri 0 0 156 156 sw
tri 238 0 394 156 ne
rect 394 0 1575 156
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 156 0
tri 156 -103 259 0 sw
tri 394 -103 497 0 ne
rect 497 -103 1575 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -240 84 -103 ne
rect 84 -240 259 -103
tri 259 -240 396 -103 sw
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
tri 84 -394 238 -240 ne
rect 238 -360 240 -240
rect 360 -342 396 -240
tri 396 -342 498 -240 sw
rect 360 -360 1075 -342
rect 238 -394 1075 -360
rect -208 -497 0 -394
tri 0 -497 103 -394 sw
rect -208 -1575 103 -497
tri 238 -498 342 -394 ne
rect 342 -653 1075 -394
rect 342 -1075 653 -653
<< end >>
