* NGSPICE file created from nmos_18x18_flat.ext - technology: sky130A

.subckt nmos_18x18_flat
X0 D.t611 G S.t638 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1 D.t610 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 S.t636 G D.t609 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D.t608 G S.t635 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 S.t634 G D.t607 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 D.t606 G S.t633 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 D.t605 G S.t632 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 D.t604 G S.t630 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 D.t603 G S.t631 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 S.t629 G D.t602 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 D.t601 G S.t628 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 D.t600 G S.t627 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 S.t625 G D.t599 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D.t598 G S.t626 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 S.t624 G D.t597 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D.t596 G S.t623 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 S.t622 G D.t595 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 S.t492 G D.t594 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 S.t621 G D.t593 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 D.t592 G S.t572 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 S.t620 G D.t591 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 S.t619 G D.t590 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 D.t589 G S.t618 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D.t588 G S.t617 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 D.t587 G S.t614 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 S.t616 G D.t586 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 S.t615 G D.t585 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 S.t613 G D.t584 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 S.t612 G D.t583 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 D.t582 G S.t611 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 S.t610 G D.t581 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 D.t580 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 S.t609 G D.t579 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 S.t607 G D.t578 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 D.t577 G S.t606 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 D.t576 G S.t487 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 S.t491 G D.t575 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t605 G D.t574 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 D.t573 G S.t577 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 D.t572 G S.t604 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D.t571 G S.t603 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 S.t602 G D.t570 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 S.t597 G D.t569 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 D.t568 G S.t598 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 D.t567 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 S.t600 G D.t566 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 D.t565 G S.t599 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 D.t564 G S.t596 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 S.t595 G D.t563 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 D.t562 G S.t594 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 D.t561 G S.t592 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 S.t593 G D.t560 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 D.t559 G S.t591 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 S.t590 G D.t558 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 D.t557 G S.t589 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 S.t488 G D.t556 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 S.t0 G D.t555 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 S.t494 G D.t554 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 S.t587 G D.t553 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D.t552 G S.t586 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 S.t585 G D.t551 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 D.t550 G S.t584 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 S.t580 G D.t549 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 D.t548 G S.t583 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 D.t547 G S.t582 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 S.t581 G D.t546 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 D.t545 G S.t579 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 D.t544 G S.t578 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 S.t574 G D.t543 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 D.t542 G S.t576 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 D.t541 G S.t575 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 S.t573 G D.t540 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 D.t539 G S.t571 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 S.t493 G D.t538 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 D.t537 G S.t495 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 D.t536 G S.t496 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 S.t0 G D.t535 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 D.t534 G S.t570 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 D.t533 G S.t569 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 S.t568 G D.t532 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 S.t563 G D.t531 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 S.t565 G D.t530 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 D.t529 G S.t567 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 S.t566 G D.t528 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 S.t564 G D.t527 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 S.t562 G D.t526 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 S.t554 G D.t525 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 S.t561 G D.t524 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 D.t523 G S.t560 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 S.t559 G D.t522 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D.t521 G S.t553 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 S.t558 G D.t520 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 S.t557 G D.t519 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 D.t518 G S.t556 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 S.t555 G D.t517 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 S.t552 G D.t516 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D.t515 G S.t551 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 D.t514 G S.t548 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 D.t513 G S.t549 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 S.t550 G D.t512 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 S.t547 G D.t511 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 D.t510 G S.t546 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 D.t509 G S.t545 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 D.t508 G S.t544 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 D.t507 G S.t543 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 D.t506 G S.t535 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 S.t542 G D.t505 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 D.t504 G S.t541 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 D.t503 G S.t540 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 S.t539 G D.t502 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D.t501 G S.t534 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 D.t500 G S.t538 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t537 G D.t499 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 D.t498 G S.t536 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 S.t533 G D.t497 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 S.t532 G D.t496 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 D.t495 G S.t530 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 D.t494 G S.t531 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 S.t529 G D.t493 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 D.t492 G S.t528 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 D.t491 G S.t527 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 D.t490 G S.t515 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 S.t526 G D.t489 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 S.t0 G D.t488 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 S.t516 G D.t487 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 D.t486 G S.t524 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 S.t523 G D.t485 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 S.t522 G D.t484 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 S.t0 G D.t483 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 S.t518 G D.t482 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 S.t521 G D.t481 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 D.t480 G S.t520 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 D.t479 G S.t519 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t514 G D.t478 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 S.t513 G D.t477 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 D.t476 G S.t512 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 S.t511 G D.t475 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 S.t510 G D.t474 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 S.t509 G D.t473 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 S.t508 G D.t472 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 D.t471 G S.t507 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 D.t470 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 S.t505 G D.t469 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 D.t468 G S.t490 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 D.t467 G S.t504 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 S.t503 G D.t466 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 D.t465 G S.t502 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 D.t464 G S.t501 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 S.t489 G D.t463 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 D.t462 G S.t500 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 D.t461 G S.t499 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 D.t460 G S.t498 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 D.t459 G S.t486 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 D.t458 G S.t485 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 S.t482 G D.t457 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 D.t456 G S.t483 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 D.t455 G S.t484 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 S.t481 G D.t454 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 D.t453 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 D.t452 G S.t479 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 D.t451 G S.t478 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 S.t477 G D.t450 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 S.t476 G D.t449 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 S.t475 G D.t448 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 D.t447 G S.t474 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 S.t472 G D.t446 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 D.t445 G S.t473 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 D.t444 G S.t471 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 S.t470 G D.t443 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 S.t469 G D.t442 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 D.t441 G S.t339 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 S.t468 G D.t440 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 D.t439 G S.t340 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 S.t0 G D.t438 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 S.t466 G D.t437 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 D.t436 G S.t465 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 S.t0 G D.t435 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 D.t434 G S.t460 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 S.t463 G D.t433 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 D.t432 G S.t462 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 S.t461 G D.t431 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 D.t430 G S.t459 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 D.t429 G S.t458 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 S.t455 G D.t428 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 D.t427 G S.t457 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 D.t426 G S.t456 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 S.t454 G D.t425 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 S.t453 G D.t424 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 D.t423 G S.t452 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 D.t422 G S.t418 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 S.t419 G D.t421 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 S.t420 G D.t420 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 S.t451 G D.t419 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 D.t418 G S.t450 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 D.t417 G S.t449 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 S.t446 G D.t416 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 D.t415 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 D.t414 G S.t448 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 S.t445 G D.t413 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 D.t412 G S.t444 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 S.t443 G D.t411 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 D.t410 G S.t442 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 D.t409 G S.t441 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 D.t408 G S.t440 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 S.t439 G D.t407 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 D.t406 G S.t438 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 S.t437 G D.t405 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 D.t404 G S.t436 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 D.t403 G S.t336 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 S.t417 G D.t402 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 D.t401 G S.t421 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 S.t435 G D.t400 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 S.t434 G D.t399 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 D.t398 G S.t433 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 S.t429 G D.t397 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 S.t430 G D.t396 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 D.t395 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 S.t431 G D.t394 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 S.t428 G D.t393 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 D.t392 G S.t427 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 S.t426 G D.t391 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 D.t390 G S.t425 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 S.t424 G D.t389 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 S.t423 G D.t388 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 D.t387 G S.t422 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 D.t386 G S.t416 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 S.t415 G D.t385 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 D.t384 G S.t338 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 D.t383 G S.t334 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 S.t343 G D.t382 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 D.t381 G S.t414 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 D.t380 G S.t413 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 S.t412 G D.t379 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 D.t378 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 D.t377 G S.t410 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 D.t376 G S.t411 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 S.t409 G D.t375 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 S.t408 G D.t374 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 D.t373 G S.t397 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 D.t372 G S.t399 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 D.t371 G S.t407 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 D.t370 G S.t406 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 S.t405 G D.t369 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 S.t400 G D.t368 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 D.t367 G S.t401 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 D.t366 G S.t404 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 D.t365 G S.t403 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 D.t364 G S.t402 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 S.t0 G D.t363 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 S.t395 G D.t362 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 S.t392 G D.t361 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 D.t360 G S.t393 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 S.t394 G D.t359 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 S.t391 G D.t358 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 D.t357 G S.t390 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 S.t389 G D.t356 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 D.t355 G S.t388 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 S.t387 G D.t354 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 S.t378 G D.t353 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 D.t352 G S.t386 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 S.t385 G D.t351 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 D.t350 G S.t384 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 S.t379 G D.t349 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 D.t348 G S.t380 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 S.t383 G D.t347 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 D.t346 G S.t382 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 D.t345 G S.t381 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 D.t344 G S.t377 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 D.t343 G S.t376 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 S.t373 G D.t342 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 S.t374 G D.t341 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 D.t340 G S.t375 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 S.t372 G D.t339 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 S.t371 G D.t338 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 D.t337 G S.t360 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 S.t370 G D.t336 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 S.t359 G D.t335 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 D.t334 G S.t362 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 S.t369 G D.t333 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 S.t368 G D.t332 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 D.t331 G S.t367 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 S.t363 G D.t330 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 S.t366 G D.t329 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D.t328 G S.t365 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 D.t327 G S.t364 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 S.t361 G D.t326 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 S.t358 G D.t325 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 S.t357 G D.t324 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 D.t323 G S.t356 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 D.t322 G S.t355 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 D.t321 G S.t354 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 S.t353 G D.t320 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 D.t319 G S.t352 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 D.t318 G S.t335 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 D.t317 G S.t341 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 D.t316 G S.t337 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 D.t315 G S.t345 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 S.t351 G D.t314 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 D.t313 G S.t350 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 D.t312 G S.t349 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 D.t311 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 S.t344 G D.t310 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 D.t309 G S.t347 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 S.t346 G D.t308 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 D.t307 G S.t342 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 S.t333 G D.t306 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 S.t332 G D.t305 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 S.t329 G D.t304 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 D.t303 G S.t330 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 S.t331 G D.t302 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 S.t328 G D.t301 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 S.t327 G D.t300 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 D.t299 G S.t326 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 D.t298 G S.t324 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 S.t325 G D.t297 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 D.t296 G S.t323 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 D.t295 G S.t322 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 S.t319 G D.t294 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 D.t293 G S.t320 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 S.t321 G D.t292 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 S.t318 G D.t291 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 D.t290 G S.t317 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 S.t316 G D.t289 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 D.t288 G S.t182 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 S.t185 G D.t287 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 S.t304 G D.t286 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 D.t285 G S.t315 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 S.t314 G D.t284 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 S.t313 G D.t283 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 D.t282 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 D.t281 G S.t311 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 S.t312 G D.t280 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 D.t279 G S.t309 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 S.t308 G D.t278 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 D.t277 G S.t307 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 D.t276 G S.t306 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 D.t275 G S.t302 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 D.t274 G S.t303 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 S.t305 G D.t273 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 D.t272 G S.t301 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 D.t271 G S.t300 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 D.t270 G S.t187 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 S.t299 G D.t269 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 D.t268 G S.t298 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 D.t267 G S.t191 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 D.t266 G S.t297 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 S.t296 G D.t265 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 S.t295 G D.t264 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 S.t290 G D.t263 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t0 G D.t262 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 S.t293 G D.t261 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 D.t260 G S.t292 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 S.t291 G D.t259 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 S.t289 G D.t258 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 S.t288 G D.t257 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 D.t256 G S.t287 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 S.t285 G D.t255 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 S.t286 G D.t254 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 S.t0 G D.t253 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 S.t283 G D.t252 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 S.t282 G D.t251 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 S.t281 G D.t250 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 D.t249 G S.t280 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 S.t0 G D.t248 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 S.t279 G D.t247 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 D.t246 G S.t278 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 S.t0 G D.t245 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 D.t244 G S.t276 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 S.t272 G D.t243 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 D.t242 G S.t275 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 S.t274 G D.t241 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 S.t273 G D.t240 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 D.t239 G S.t271 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 D.t238 G S.t270 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 D.t237 G S.t267 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 S.t269 G D.t236 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 D.t235 G S.t268 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 D.t234 G S.t266 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 S.t265 G D.t233 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 S.t264 G D.t232 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 S.t189 G D.t231 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 D.t230 G S.t186 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 D.t229 G S.t219 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 S.t263 G D.t228 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 D.t227 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 S.t261 G D.t226 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 D.t225 G S.t260 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 S.t246 G D.t224 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 S.t259 G D.t223 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 D.t222 G S.t258 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 S.t257 G D.t221 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 D.t220 G S.t256 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 D.t219 G S.t247 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 S.t255 G D.t218 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 S.t254 G D.t217 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 D.t216 G S.t253 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 S.t248 G D.t215 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 D.t214 G S.t249 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 S.t252 G D.t213 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 D.t212 G S.t251 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 D.t211 G S.t250 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 S.t245 G D.t210 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 S.t244 G D.t209 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 D.t208 G S.t243 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 S.t0 G D.t207 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 S.t241 G D.t206 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 D.t205 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 S.t239 G D.t204 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 S.t237 G D.t203 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 S.t238 G D.t202 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 D.t201 G S.t236 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 S.t227 G D.t200 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 S.t235 G D.t199 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 S.t234 G D.t198 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 D.t197 G S.t233 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 S.t232 G D.t196 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 D.t195 G S.t228 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 D.t194 G S.t231 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 S.t230 G D.t193 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 S.t229 G D.t192 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 D.t191 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 D.t190 G S.t225 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 D.t189 G S.t224 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 D.t188 G S.t223 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 S.t222 G D.t187 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 D.t186 G S.t221 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 D.t185 G S.t220 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 D.t184 G S.t218 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 S.t217 G D.t183 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 D.t182 G S.t216 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 S.t207 G D.t181 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 D.t180 G S.t215 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 D.t179 G S.t214 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 D.t178 G S.t213 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 S.t0 G D.t177 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 S.t211 G D.t176 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 S.t210 G D.t175 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 D.t174 G S.t209 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 D.t173 G S.t208 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 S.t206 G D.t172 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 S.t205 G D.t171 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 D.t170 G S.t202 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 D.t169 G S.t203 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 S.t204 G D.t168 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 D.t167 G S.t201 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 S.t200 G D.t166 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 S.t199 G D.t165 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 S.t183 G D.t164 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 D.t163 G S.t188 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 S.t190 G D.t162 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 D.t161 G S.t198 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 S.t197 G D.t160 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 S.t196 G D.t159 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 S.t195 G D.t158 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 S.t184 G D.t157 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 S.t194 G D.t156 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 D.t155 G S.t193 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 S.t192 G D.t154 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 S.t180 G D.t153 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 D.t152 G S.t179 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 D.t151 G S.t178 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 D.t150 G S.t177 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 D.t149 G S.t176 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t175 G D.t148 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 D.t147 G S.t174 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 S.t171 G D.t146 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 S.t173 G D.t145 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 D.t144 G S.t172 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 S.t170 G D.t143 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 S.t169 G D.t142 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 D.t141 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 D.t140 G S.t168 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 S.t166 G D.t139 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 S.t165 G D.t138 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 D.t137 G S.t164 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 S.t163 G D.t136 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 S.t162 G D.t135 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 D.t134 G S.t142 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 S.t145 G D.t133 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 S.t0 G D.t132 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 S.t160 G D.t131 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 S.t159 G D.t130 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 D.t129 G S.t158 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 D.t128 G S.t154 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 D.t127 G S.t157 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 S.t156 G D.t126 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 D.t125 G S.t155 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 D.t124 G S.t153 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 D.t123 G S.t152 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 S.t151 G D.t122 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 D.t121 G S.t149 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 D.t120 G S.t150 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 D.t119 G S.t148 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 S.t147 G D.t118 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t146 G D.t117 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 D.t116 G S.t143 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 D.t115 G S.t141 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 D.t114 G S.t3 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 D.t113 G S.t140 S.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 S.t138 G D.t112 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 D.t111 G S.t137 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 D.t110 G S.t136 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 S.t135 G D.t109 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 S.t134 G D.t108 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 S.t133 G D.t107 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 D.t106 G S.t132 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 S.t131 G D.t105 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 S.t130 G D.t104 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 S.t129 G D.t103 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 S.t127 G D.t102 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t128 G D.t101 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 D.t100 G S.t126 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 S.t125 G D.t99 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 S.t124 G D.t98 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 S.t6 G D.t97 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 D.t96 G S.t105 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 S.t111 G D.t95 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 S.t123 G D.t94 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 D.t93 G S.t122 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 D.t92 G S.t121 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 D.t91 G S.t115 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 S.t120 G D.t90 S.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 S.t118 G D.t89 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 D.t88 G S.t117 S.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 D.t87 G S.t116 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 S.t114 G D.t86 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 S.t113 G D.t85 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 S.t110 G D.t84 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 D.t83 G S.t112 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 S.t109 G D.t82 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 S.t108 G D.t81 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D.t80 G S.t107 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 D.t79 G S.t106 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 D.t78 G S.t104 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 D.t77 G S.t103 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 D.t76 G S.t8 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 D.t75 G S.t102 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 D.t74 G S.t101 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 D.t73 G S.t100 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 D.t72 G S.t95 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 D.t71 G S.t98 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 S.t97 G D.t70 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 S.t0 G D.t69 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 S.t93 G D.t68 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 D.t67 G S.t92 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t82 G D.t66 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 S.t91 G D.t65 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 D.t64 G S.t90 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 S.t89 G D.t63 S.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 S.t83 G D.t62 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 S.t87 G D.t61 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 S.t86 G D.t60 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 S.t85 G D.t59 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 D.t58 G S.t84 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 S.t81 G D.t57 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 S.t0 G D.t56 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 S.t79 G D.t55 S.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 D.t54 G S.t77 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 S.t76 G D.t53 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 D.t52 G S.t75 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 S.t74 G D.t51 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 D.t50 G S.t63 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 D.t49 G S.t68 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 D.t48 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 S.t73 G D.t47 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 D.t46 G S.t72 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 D.t45 G S.t71 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 S.t70 G D.t44 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 D.t43 G S.t62 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 D.t42 G S.t67 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 S.t66 G D.t41 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 D.t40 G S.t65 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 D.t39 G S.t64 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 S.t61 G D.t38 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 D.t37 G S.t60 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 D.t36 G S.t59 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 S.t57 G D.t35 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 D.t34 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 D.t33 G S.t56 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 S.t54 G D.t32 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 S.t53 G D.t31 S.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 S.t51 G D.t30 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 S.t37 G D.t29 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 D.t28 G S.t38 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 D.t27 G S.t50 S.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 S.t48 G D.t26 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 D.t25 G S.t46 S.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 S.t39 G D.t24 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 D.t23 G S.t40 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 D.t22 G S.t44 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 S.t43 G D.t21 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 D.t20 G S.t42 S.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 S.t0 G D.t19 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 S.t35 G D.t18 S.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 D.t17 G S.t33 S.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 S.t30 G D.t16 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 S.t0 G D.t15 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 D.t14 G S.t29 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 D.t13 G S.t28 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 S.t11 G D.t12 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 S.t27 G D.t11 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D.t10 G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 S.t21 G D.t9 S.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 D.t8 G S.t26 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 S.t24 G D.t7 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 S.t22 G D.t6 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 D.t5 G S.t4 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 S.t19 G D.t4 S.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 D.t3 G S.t17 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 S.t15 G D.t2 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 S.t13 G D.t1 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 D.t0 G S.t1 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 S.n60 S.n171 169.035
R1 S.n62 S.n338 169.035
R2 S.n64 S.n475 169.035
R3 S.n66 S.n603 169.035
R4 S.n9 S.n741 169.035
R5 S.n3 S.n265 169.035
R6 S.n59 S.n172 137.94
R7 S.n61 S.n339 137.94
R8 S.n63 S.n476 137.94
R9 S.n65 S.n604 137.94
R10 S.n682 S.n681 129.201
R11 S.n670 S.n669 129.201
R12 S.n538 S.n537 129.201
R13 S.n404 S.n403 129.201
R14 S.n264 S.n263 129.201
R15 S.n9 S.t12 95.334
R16 S.n3 S.t7 95.333
R17 S.n59 S.t23 95.333
R18 S.n4 S.t119 95.333
R19 S.n61 S.t88 95.333
R20 S.n5 S.t20 95.333
R21 S.n63 S.t5 95.333
R22 S.n6 S.t16 95.333
R23 S.n65 S.t25 95.333
R24 S.n7 S.t10 95.333
R25 S.t14 S.n211 91.963
R26 S.t144 S.n323 91.963
R27 S.t99 S.n381 91.963
R28 S.t18 S.n452 91.963
R29 S.t139 S.n512 91.963
R30 S.t78 S.n577 91.963
R31 S.t41 S.n632 91.963
R32 S.t49 S.n709 91.963
R33 S.t55 S.n763 91.963
R34 S.t34 S.n992 91.963
R35 S.t45 S.n961 91.519
R36 S.t34 S.n1091 91.519
R37 S.t14 S.n173 91.519
R38 S.t41 S.n605 91.519
R39 S.t55 S.n742 91.519
R40 S.t47 S.n1006 91.519
R41 S.t32 S.n813 91.519
R42 S.t99 S.n340 91.519
R43 S.t139 S.n477 91.519
R44 S.t94 S.n257 91.519
R45 S.t144 S.n399 91.519
R46 S.t18 S.n531 91.519
R47 S.t78 S.n663 91.519
R48 S.t49 S.n797 91.519
R49 S.t52 S.n906 91.519
R50 S.t0 S.n970 87.091
R51 S.t0 S.n964 87.091
R52 S.t2 S.n135 87.091
R53 S.t2 S.n123 87.091
R54 S.t2 S.n137 87.091
R55 S.t2 S.n126 87.091
R56 S.t2 S.n130 87.091
R57 S.t2 S.n134 87.091
R58 S.t2 S.n118 87.091
R59 S.t2 S.n136 87.091
R60 S.t0 S.n965 87.091
R61 S.t0 S.n966 87.091
R62 S.t0 S.n967 87.091
R63 S.t0 S.n968 87.091
R64 S.t0 S.n969 87.091
R65 S.t0 S.n963 87.091
R66 S.t14 S.t536 3.838
R67 S.t99 S.t388 3.838
R68 S.t139 S.t258 3.838
R69 S.t41 S.t153 3.838
R70 S.t55 S.t638 3.838
R71 S.t32 S.t356 3.838
R72 S.t45 S.t311 3.838
R73 S.t47 S.t490 3.838
R74 S.t55 S.t191 3.773
R75 S.t55 S.n738 3.773
R76 S.t55 S.n739 3.773
R77 S.t55 S.t74 3.773
R78 S.n10 S.t499 3.773
R79 S.t0 S.t496 3.773
R80 S.n11 S.t286 3.773
R81 S.t45 S.t401 3.773
R82 S.n910 S.t244 3.773
R83 S.t0 S.t72 3.773
R84 S.n962 S.t101 3.773
R85 S.t34 S.t520 3.773
R86 S.t47 S.n1019 3.773
R87 S.t47 S.t165 3.773
R88 S.t47 S.t452 3.773
R89 S.t47 S.n1027 3.773
R90 S.n1026 S.t479 3.773
R91 S.n1026 S.n1025 3.773
R92 S.n1020 S.n1021 3.773
R93 S.n1020 S.t129 3.773
R94 S.t52 S.n861 3.773
R95 S.t52 S.t255 3.773
R96 S.t52 S.t462 3.773
R97 S.t52 S.n866 3.773
R98 S.n865 S.t406 3.773
R99 S.n865 S.n864 3.773
R100 S.n862 S.n863 3.773
R101 S.n862 S.t199 3.773
R102 S.t0 S.t178 3.773
R103 S.n23 S.t522 3.773
R104 S.n22 S.t103 3.773
R105 S.t45 S.n920 3.773
R106 S.t45 S.t265 3.773
R107 S.t45 S.t339 3.773
R108 S.t45 S.n923 3.773
R109 S.n922 S.t416 3.773
R110 S.n922 S.n921 3.773
R111 S.n918 S.n919 3.773
R112 S.n918 S.t207 3.773
R113 S.t32 S.n860 3.773
R114 S.t32 S.t263 3.773
R115 S.t32 S.t465 3.773
R116 S.t32 S.n859 3.773
R117 S.n858 S.t413 3.773
R118 S.n858 S.n857 3.773
R119 S.n811 S.n812 3.773
R120 S.n811 S.t205 3.773
R121 S.t14 S.t264 3.773
R122 S.n170 S.t461 3.773
R123 S.t94 S.n251 3.773
R124 S.t94 S.t113 3.773
R125 S.t94 S.t326 3.773
R126 S.t94 S.n250 3.773
R127 S.n256 S.t386 3.773
R128 S.n256 S.n255 3.773
R129 S.n252 S.n253 3.773
R130 S.n252 S.t316 3.773
R131 S.t2 S.t166 3.773
R132 S.n29 S.t494 3.773
R133 S.n30 S.t177 3.773
R134 S.t2 S.t563 3.773
R135 S.n39 S.t616 3.773
R136 S.n38 S.t221 3.773
R137 S.t94 S.n155 3.773
R138 S.t94 S.t622 3.773
R139 S.t94 S.t320 3.773
R140 S.t94 S.n160 3.773
R141 S.n159 S.t157 3.773
R142 S.n159 S.n158 3.773
R143 S.n156 S.n157 3.773
R144 S.n156 S.t493 3.773
R145 S.t14 S.n186 3.773
R146 S.t14 S.t259 3.773
R147 S.t14 S.t436 3.773
R148 S.t14 S.n191 3.773
R149 S.n190 S.t486 3.773
R150 S.n190 S.n189 3.773
R151 S.n187 S.n188 3.773
R152 S.n187 S.t426 3.773
R153 S.n57 S.n349 3.773
R154 S.n57 S.t511 3.773
R155 S.t99 S.t100 3.773
R156 S.t99 S.n354 3.773
R157 S.n353 S.t148 3.773
R158 S.n353 S.n352 3.773
R159 S.n347 S.n348 3.773
R160 S.n347 S.t89 3.773
R161 S.t139 S.n480 3.773
R162 S.t139 S.t163 3.773
R163 S.t139 S.t384 3.773
R164 S.t139 S.n485 3.773
R165 S.n484 S.t444 3.773
R166 S.n484 S.n483 3.773
R167 S.n478 S.n479 3.773
R168 S.n478 S.t372 3.773
R169 S.t41 S.t518 3.773
R170 S.n602 S.t93 3.773
R171 S.t78 S.n581 3.773
R172 S.t78 S.t304 3.773
R173 S.t78 S.t531 3.773
R174 S.t78 S.n586 3.773
R175 S.n588 S.t583 3.773
R176 S.n588 S.n587 3.773
R177 S.n578 S.n579 3.773
R178 S.n578 S.t564 3.773
R179 S.n77 S.n413 3.773
R180 S.n77 S.t19 3.773
R181 S.t18 S.t249 3.773
R182 S.t18 S.n418 3.773
R183 S.n417 S.t307 3.773
R184 S.n417 S.n416 3.773
R185 S.n410 S.n411 3.773
R186 S.n410 S.t239 3.773
R187 S.t2 S.t134 3.773
R188 S.t2 S.t184 3.773
R189 S.n26 S.t397 3.773
R190 S.t94 S.n163 3.773
R191 S.t94 S.t200 3.773
R192 S.t94 S.t414 3.773
R193 S.t94 S.n168 3.773
R194 S.n167 S.t355 3.773
R195 S.n167 S.n166 3.773
R196 S.n164 S.n165 3.773
R197 S.n164 S.t138 3.773
R198 S.t14 S.n192 3.773
R199 S.t14 S.t206 3.773
R200 S.t14 S.t422 3.773
R201 S.t14 S.n198 3.773
R202 S.n197 S.t364 3.773
R203 S.n197 S.n196 3.773
R204 S.n193 S.n194 3.773
R205 S.n193 S.t146 3.773
R206 S.t55 S.t370 3.773
R207 S.n740 S.t565 3.773
R208 S.t49 S.n712 3.773
R209 S.t49 S.t227 3.773
R210 S.t49 S.t442 3.773
R211 S.t49 S.n715 3.773
R212 S.n717 S.t504 3.773
R213 S.n717 S.n716 3.773
R214 S.n713 S.n714 3.773
R215 S.n713 S.t434 3.773
R216 S.t41 S.n606 3.773
R217 S.t41 S.t85 3.773
R218 S.t41 S.t301 3.773
R219 S.t41 S.n611 3.773
R220 S.n610 S.t335 3.773
R221 S.n610 S.n609 3.773
R222 S.n607 S.n608 3.773
R223 S.n607 S.t293 3.773
R224 S.t78 S.n546 3.773
R225 S.t78 S.t514 3.773
R226 S.t78 S.t102 3.773
R227 S.t78 S.n551 3.773
R228 S.n550 S.t152 3.773
R229 S.n550 S.n549 3.773
R230 S.n547 S.n548 3.773
R231 S.n547 S.t130 3.773
R232 S.t139 S.n486 3.773
R233 S.t139 S.t363 3.773
R234 S.t139 S.t576 3.773
R235 S.t139 S.n491 3.773
R236 S.n490 S.t632 3.773
R237 S.n490 S.n489 3.773
R238 S.n487 S.n488 3.773
R239 S.n487 S.t562 3.773
R240 S.t18 S.n421 3.773
R241 S.t18 S.t232 3.773
R242 S.t18 S.t438 3.773
R243 S.t18 S.n426 3.773
R244 S.n425 S.t500 3.773
R245 S.n425 S.n424 3.773
R246 S.n422 S.n423 3.773
R247 S.n422 S.t431 3.773
R248 S.t99 S.n355 3.773
R249 S.t99 S.t108 3.773
R250 S.t99 S.t298 3.773
R251 S.t99 S.n360 3.773
R252 S.n359 S.t345 3.773
R253 S.n359 S.n358 3.773
R254 S.n356 S.n357 3.773
R255 S.n356 S.t288 3.773
R256 S.t144 S.n291 3.773
R257 S.t144 S.t217 3.773
R258 S.t144 S.t174 3.773
R259 S.t144 S.n298 3.773
R260 S.n297 S.t362 3.773
R261 S.n297 S.n296 3.773
R262 S.n292 S.n293 3.773
R263 S.n292 S.t156 3.773
R264 S.t14 S.n169 3.773
R265 S.t14 S.t392 3.773
R266 S.t14 S.t577 3.773
R267 S.t14 S.n218 3.773
R268 S.n220 S.t556 3.773
R269 S.n220 S.n219 3.773
R270 S.n221 S.n222 3.773
R271 S.n221 S.t351 3.773
R272 S.t94 S.n223 3.773
R273 S.t94 S.t394 3.773
R274 S.t94 S.t598 3.773
R275 S.t94 S.n229 3.773
R276 S.n228 S.t549 3.773
R277 S.n228 S.n227 3.773
R278 S.n224 S.n225 3.773
R279 S.n224 S.t344 3.773
R280 S.t2 S.t333 3.773
R281 S.n36 S.t385 3.773
R282 S.n35 S.t592 3.773
R283 S.t144 S.n301 3.773
R284 S.t144 S.t405 3.773
R285 S.t144 S.t611 3.773
R286 S.t144 S.n305 3.773
R287 S.n304 S.t560 3.773
R288 S.n304 S.n303 3.773
R289 S.n299 S.n300 3.773
R290 S.n299 S.t353 3.773
R291 S.t99 S.n363 3.773
R292 S.t99 S.t412 3.773
R293 S.t99 S.t572 3.773
R294 S.t99 S.n368 3.773
R295 S.n367 S.t567 3.773
R296 S.n367 S.n366 3.773
R297 S.n361 S.n362 3.773
R298 S.n361 S.t358 3.773
R299 S.t18 S.n430 3.773
R300 S.t18 S.t415 3.773
R301 S.t18 S.t28 3.773
R302 S.t18 S.n435 3.773
R303 S.n434 S.t495 3.773
R304 S.n434 S.n433 3.773
R305 S.n427 S.n428 3.773
R306 S.n427 S.t369 3.773
R307 S.t139 S.n494 3.773
R308 S.t139 S.t585 3.773
R309 S.t139 S.t140 3.773
R310 S.t139 S.n499 3.773
R311 S.n498 S.t213 3.773
R312 S.n498 S.n497 3.773
R313 S.n492 S.n493 3.773
R314 S.n492 S.t128 3.773
R315 S.t78 S.n555 3.773
R316 S.t78 S.t79 3.773
R317 S.t78 S.t187 3.773
R318 S.t78 S.n560 3.773
R319 S.n559 S.t341 3.773
R320 S.n559 S.n558 3.773
R321 S.n552 S.n553 3.773
R322 S.n552 S.t328 3.773
R323 S.t41 S.n614 3.773
R324 S.t41 S.t282 3.773
R325 S.t41 S.t485 3.773
R326 S.t41 S.n619 3.773
R327 S.n618 S.t544 3.773
R328 S.n618 S.n617 3.773
R329 S.n612 S.n613 3.773
R330 S.n612 S.t472 3.773
R331 S.n74 S.n687 3.773
R332 S.n74 S.t424 3.773
R333 S.t49 S.t628 3.773
R334 S.t49 S.n692 3.773
R335 S.n691 S.t71 3.773
R336 S.n691 S.n690 3.773
R337 S.n684 S.n685 3.773
R338 S.n684 S.t613 3.773
R339 S.n88 S.n745 3.773
R340 S.n88 S.t559 3.773
R341 S.t55 S.t143 3.773
R342 S.t55 S.n750 3.773
R343 S.n749 S.t223 3.773
R344 S.n749 S.n748 3.773
R345 S.n743 S.n744 3.773
R346 S.n743 S.t133 3.773
R347 S.t34 S.n996 3.773
R348 S.t34 S.t87 3.773
R349 S.t34 S.t302 3.773
R350 S.t34 S.n1001 3.773
R351 S.n1003 S.t354 3.773
R352 S.n1003 S.n1002 3.773
R353 S.n993 S.n994 3.773
R354 S.n993 S.t290 3.773
R355 S.t47 S.t237 3.773
R356 S.n1005 S.t435 3.773
R357 S.t144 S.n306 3.773
R358 S.t144 S.t590 3.773
R359 S.t144 S.t193 3.773
R360 S.t144 S.n313 3.773
R361 S.n312 S.t126 3.773
R362 S.n312 S.n311 3.773
R363 S.n307 S.n308 3.773
R364 S.n307 S.t547 3.773
R365 S.t14 S.n199 3.773
R366 S.t14 S.t587 3.773
R367 S.t14 S.t176 3.773
R368 S.t14 S.n204 3.773
R369 S.n203 S.t105 3.773
R370 S.n203 S.n202 3.773
R371 S.n200 S.n201 3.773
R372 S.n200 S.t542 3.773
R373 S.t94 S.n231 3.773
R374 S.t94 S.t580 3.773
R375 S.t94 S.t172 3.773
R376 S.t94 S.n239 3.773
R377 S.n238 S.t121 3.773
R378 S.n238 S.n237 3.773
R379 S.n232 S.n233 3.773
R380 S.n232 S.t539 3.773
R381 S.t2 S.t533 3.773
R382 S.n34 S.t574 3.773
R383 S.n33 S.t164 3.773
R384 S.t32 S.t91 3.773
R385 S.n103 S.t296 3.773
R386 S.t52 S.n869 3.773
R387 S.t52 S.t554 3.773
R388 S.t52 S.t149 3.773
R389 S.t52 S.n871 3.773
R390 S.n873 S.t224 3.773
R391 S.n873 S.n872 3.773
R392 S.n867 S.n868 3.773
R393 S.n867 S.t135 3.773
R394 S.t47 S.n1009 3.773
R395 S.t47 S.t428 3.773
R396 S.t47 S.t630 3.773
R397 S.t47 S.n1012 3.773
R398 S.n1011 S.t68 3.773
R399 S.n1011 S.n1010 3.773
R400 S.n1007 S.n1008 3.773
R401 S.n1007 S.t619 3.773
R402 S.t34 S.n980 3.773
R403 S.t34 S.t285 3.773
R404 S.t34 S.t498 3.773
R405 S.t34 S.n983 3.773
R406 S.n982 S.t546 3.773
R407 S.n982 S.n981 3.773
R408 S.n978 S.n979 3.773
R409 S.n978 S.t475 3.773
R410 S.t55 S.n753 3.773
R411 S.t55 S.t125 3.773
R412 S.t55 S.t350 3.773
R413 S.t55 S.n756 3.773
R414 S.n755 S.t407 3.773
R415 S.n755 S.n754 3.773
R416 S.n751 S.n752 3.773
R417 S.n751 S.t332 3.773
R418 S.t49 S.n697 3.773
R419 S.t49 S.t491 3.773
R420 S.t49 S.t209 3.773
R421 S.t49 S.n700 3.773
R422 S.n699 S.t267 3.773
R423 S.n699 S.n698 3.773
R424 S.n695 S.n696 3.773
R425 S.n695 S.t195 3.773
R426 S.t41 S.n622 3.773
R427 S.t41 S.t505 3.773
R428 S.t41 S.t64 3.773
R429 S.t41 S.n625 3.773
R430 S.n624 S.t116 3.773
R431 S.n624 S.n623 3.773
R432 S.n620 S.n621 3.773
R433 S.n620 S.t37 3.773
R434 S.t78 S.n565 3.773
R435 S.t78 S.t620 3.773
R436 S.t78 S.t524 3.773
R437 S.t78 S.n568 3.773
R438 S.n567 S.t155 3.773
R439 S.n567 S.n566 3.773
R440 S.n563 S.n564 3.773
R441 S.n563 S.t39 3.773
R442 S.t139 S.n502 3.773
R443 S.t139 S.t609 3.773
R444 S.t139 S.t215 3.773
R445 S.t139 S.n505 3.773
R446 S.n504 S.t141 3.773
R447 S.n504 S.n503 3.773
R448 S.n500 S.n501 3.773
R449 S.n500 S.t566 3.773
R450 S.t18 S.n440 3.773
R451 S.t18 S.t602 3.773
R452 S.t18 S.t202 3.773
R453 S.t18 S.n443 3.773
R454 S.n442 S.t137 3.773
R455 S.n442 S.n441 3.773
R456 S.n438 S.n439 3.773
R457 S.n438 S.t558 3.773
R458 S.t99 S.n371 3.773
R459 S.t99 S.t600 3.773
R460 S.t99 S.t188 3.773
R461 S.t99 S.n374 3.773
R462 S.n373 S.t132 3.773
R463 S.n373 S.n372 3.773
R464 S.n369 S.n370 3.773
R465 S.n369 S.t555 3.773
R466 S.t2 S.t329 3.773
R467 S.n32 S.t30 3.773
R468 S.n31 S.t367 3.773
R469 S.t94 S.n244 3.773
R470 S.t94 S.t151 3.773
R471 S.t94 S.t375 3.773
R472 S.t94 S.n249 3.773
R473 S.n248 S.t182 3.773
R474 S.n248 S.n247 3.773
R475 S.n245 S.n246 3.773
R476 S.n245 S.t109 3.773
R477 S.t14 S.n205 3.773
R478 S.t14 S.t159 3.773
R479 S.t14 S.t376 3.773
R480 S.t14 S.n210 3.773
R481 S.n209 S.t322 3.773
R482 S.n209 S.n208 3.773
R483 S.n206 S.n207 3.773
R484 S.n206 S.t110 3.773
R485 S.t45 S.n924 3.773
R486 S.t45 S.t430 3.773
R487 S.t45 S.t633 3.773
R488 S.t45 S.n927 3.773
R489 S.n929 S.t75 3.773
R490 S.n929 S.n928 3.773
R491 S.n925 S.n926 3.773
R492 S.n925 S.t492 3.773
R493 S.t32 S.n814 3.773
R494 S.t32 S.t291 3.773
R495 S.t32 S.t501 3.773
R496 S.t32 S.n819 3.773
R497 S.n818 S.t548 3.773
R498 S.n818 S.n817 3.773
R499 S.n815 S.n816 3.773
R500 S.n815 S.t477 3.773
R501 S.t52 S.n805 3.773
R502 S.t52 S.t127 3.773
R503 S.t52 S.t337 3.773
R504 S.t52 S.n810 3.773
R505 S.n809 S.t411 3.773
R506 S.n809 S.n808 3.773
R507 S.n806 S.n807 3.773
R508 S.n806 S.t346 3.773
R509 S.t47 S.n1013 3.773
R510 S.t47 S.t607 3.773
R511 S.t47 S.t214 3.773
R512 S.t47 S.n1018 3.773
R513 S.n1017 S.t270 3.773
R514 S.n1017 S.n1016 3.773
R515 S.n1014 S.n1015 3.773
R516 S.n1014 S.t196 3.773
R517 S.t34 S.n986 3.773
R518 S.t34 S.t468 3.773
R519 S.t34 S.t65 3.773
R520 S.t34 S.n991 3.773
R521 S.n990 S.t115 3.773
R522 S.n990 S.n989 3.773
R523 S.n987 S.n988 3.773
R524 S.n987 S.t51 3.773
R525 S.t55 S.n757 3.773
R526 S.t55 S.t357 3.773
R527 S.t55 S.t541 3.773
R528 S.t55 S.n762 3.773
R529 S.n761 S.t594 3.773
R530 S.n761 S.n760 3.773
R531 S.n758 S.n759 3.773
R532 S.n758 S.t532 3.773
R533 S.t49 S.n703 3.773
R534 S.t49 S.t312 3.773
R535 S.t49 S.t421 3.773
R536 S.t49 S.n708 3.773
R537 S.n707 S.t459 3.773
R538 S.n707 S.n706 3.773
R539 S.n704 S.n705 3.773
R540 S.n704 S.t261 3.773
R541 S.n89 S.n626 3.773
R542 S.n89 S.t305 3.773
R543 S.t41 S.t519 3.773
R544 S.t41 S.n631 3.773
R545 S.n630 S.t418 3.773
R546 S.n630 S.n629 3.773
R547 S.n627 S.n628 3.773
R548 S.n627 S.t254 3.773
R549 S.n68 S.n571 3.773
R550 S.n68 S.t197 3.773
R551 S.t78 S.t410 3.773
R552 S.t78 S.n576 3.773
R553 S.n575 S.t352 3.773
R554 S.n575 S.n574 3.773
R555 S.n572 S.n573 3.773
R556 S.n572 S.t252 3.773
R557 S.t139 S.n506 3.773
R558 S.t139 S.t180 3.773
R559 S.t139 S.t404 3.773
R560 S.t139 S.n511 3.773
R561 S.n510 S.t349 3.773
R562 S.n510 S.n509 3.773
R563 S.n507 S.n508 3.773
R564 S.n507 S.t131 3.773
R565 S.t18 S.n446 3.773
R566 S.t18 S.t175 3.773
R567 S.t18 S.t393 3.773
R568 S.t18 S.n451 3.773
R569 S.n450 S.t347 3.773
R570 S.n450 S.n449 3.773
R571 S.n447 S.n448 3.773
R572 S.n447 S.t124 3.773
R573 S.t99 S.n375 3.773
R574 S.t99 S.t170 3.773
R575 S.t99 S.t390 3.773
R576 S.t99 S.n380 3.773
R577 S.n379 S.t330 3.773
R578 S.n379 S.n378 3.773
R579 S.n376 S.n377 3.773
R580 S.n376 S.t111 3.773
R581 S.t144 S.n317 3.773
R582 S.t144 S.t162 3.773
R583 S.t144 S.t380 3.773
R584 S.t144 S.n322 3.773
R585 S.n321 S.t324 3.773
R586 S.n321 S.n320 3.773
R587 S.n318 S.n319 3.773
R588 S.n318 S.t120 3.773
R589 S.t144 S.n280 3.773
R590 S.t144 S.t361 3.773
R591 S.t144 S.t571 3.773
R592 S.t144 S.n287 3.773
R593 S.n286 S.t631 3.773
R594 S.n286 S.n285 3.773
R595 S.n281 S.n282 3.773
R596 S.n281 S.t561 3.773
R597 S.t2 S.t368 3.773
R598 S.n42 S.t160 3.773
R599 S.n41 S.t377 3.773
R600 S.t94 S.n141 3.773
R601 S.t94 S.t313 3.773
R602 S.t94 S.t527 3.773
R603 S.t94 S.n146 3.773
R604 S.n145 S.t578 3.773
R605 S.n145 S.n144 3.773
R606 S.n142 S.n143 3.773
R607 S.n142 S.t521 3.773
R608 S.t14 S.n174 3.773
R609 S.t14 S.t419 3.773
R610 S.t14 S.t40 3.773
R611 S.t14 S.n179 3.773
R612 S.n178 S.t8 3.773
R613 S.n178 S.n177 3.773
R614 S.n175 S.n176 3.773
R615 S.n175 S.t24 3.773
R616 S.t99 S.t114 3.773
R617 S.n337 S.t321 3.773
R618 S.t2 S.t557 3.773
R619 S.n27 S.t389 3.773
R620 S.n28 S.t570 3.773
R621 S.t94 S.n149 3.773
R622 S.t94 S.t510 3.773
R623 S.t94 S.t95 3.773
R624 S.t94 S.n154 3.773
R625 S.n153 S.t3 3.773
R626 S.n153 S.n152 3.773
R627 S.n150 S.n151 3.773
R628 S.n150 S.t86 3.773
R629 S.t14 S.n180 3.773
R630 S.t14 S.t15 3.773
R631 S.t14 S.t251 3.773
R632 S.t14 S.n185 3.773
R633 S.n184 S.t303 3.773
R634 S.n184 S.n183 3.773
R635 S.n181 S.n182 3.773
R636 S.n181 S.t238 3.773
R637 S.t139 S.t593 3.773
R638 S.n474 S.t171 3.773
R639 S.t18 S.n455 3.773
R640 S.t18 S.t454 3.773
R641 S.t18 S.t38 3.773
R642 S.t18 S.n458 3.773
R643 S.n460 S.t104 3.773
R644 S.n460 S.n459 3.773
R645 S.n456 S.n457 3.773
R646 S.n456 S.t21 3.773
R647 S.t99 S.n341 3.773
R648 S.t99 S.t314 3.773
R649 S.t99 S.t528 3.773
R650 S.t99 S.n346 3.773
R651 S.n345 S.t579 3.773
R652 S.n345 S.n344 3.773
R653 S.n342 S.n343 3.773
R654 S.n342 S.t523 3.773
R655 S.t144 S.n270 3.773
R656 S.t144 S.t145 3.773
R657 S.t144 S.t382 3.773
R658 S.t144 S.n277 3.773
R659 S.n276 S.t441 3.773
R660 S.n276 S.n275 3.773
R661 S.n271 S.n272 3.773
R662 S.n271 S.t359 3.773
R663 S.t144 S.n328 3.773
R664 S.t144 S.t488 3.773
R665 S.t144 S.t179 3.773
R666 S.t144 S.n333 3.773
R667 S.n335 S.t247 3.773
R668 S.n335 S.n334 3.773
R669 S.n329 S.n330 3.773
R670 S.n329 S.t169 3.773
R671 S.t2 S.t395 3.773
R672 S.n138 S.t595 3.773
R673 S.t94 S.t323 3.773
R674 S.n258 S.t617 3.773
R675 S.n259 S.t550 3.773
R676 S.t14 S.n212 3.773
R677 S.t14 S.t597 3.773
R678 S.t14 S.t569 3.773
R679 S.t14 S.n215 3.773
R680 S.n217 S.t603 3.773
R681 S.n217 S.n216 3.773
R682 S.n213 S.n214 3.773
R683 S.n213 S.t274 3.773
R684 S.t144 S.n393 3.773
R685 S.t144 S.t366 3.773
R686 S.t144 S.t575 3.773
R687 S.t144 S.n396 3.773
R688 S.n398 S.t515 3.773
R689 S.n398 S.n397 3.773
R690 S.n394 S.n395 3.773
R691 S.n394 S.t185 3.773
R692 S.t99 S.n336 3.773
R693 S.t99 S.t371 3.773
R694 S.t99 S.t582 3.773
R695 S.t99 S.n388 3.773
R696 S.n390 S.t530 3.773
R697 S.n390 S.n389 3.773
R698 S.n391 S.n392 3.773
R699 S.n391 S.t319 3.773
R700 S.t18 S.n467 3.773
R701 S.t18 S.t373 3.773
R702 S.t18 S.t586 3.773
R703 S.t18 S.n470 3.773
R704 S.n472 S.t534 3.773
R705 S.n472 S.n471 3.773
R706 S.n468 S.n469 3.773
R707 S.n468 S.t325 3.773
R708 S.n78 S.n461 3.773
R709 S.n78 S.t383 3.773
R710 S.n78 S.t589 3.773
R711 S.n78 S.n462 3.773
R712 S.n464 S.t540 3.773
R713 S.n464 S.n463 3.773
R714 S.n465 S.n466 3.773
R715 S.n465 S.t331 3.773
R716 S.t78 S.n589 3.773
R717 S.t78 S.t387 3.773
R718 S.t78 S.t599 3.773
R719 S.t78 S.n592 3.773
R720 S.n594 S.t545 3.773
R721 S.n594 S.n593 3.773
R722 S.n590 S.n591 3.773
R723 S.n590 S.t437 3.773
R724 S.t41 S.n633 3.773
R725 S.t41 S.t482 3.773
R726 S.t41 S.t84 3.773
R727 S.t41 S.n636 3.773
R728 S.n638 S.t17 3.773
R729 S.n638 S.n637 3.773
R730 S.n634 S.n635 3.773
R731 S.n634 S.t443 3.773
R732 S.t49 S.n718 3.773
R733 S.t49 S.t503 3.773
R734 S.t49 S.t92 3.773
R735 S.t49 S.n721 3.773
R736 S.n723 S.t26 3.773
R737 S.n723 S.n722 3.773
R738 S.n719 S.n720 3.773
R739 S.n719 S.t446 3.773
R740 S.t55 S.n764 3.773
R741 S.t55 S.t508 3.773
R742 S.t55 S.t98 3.773
R743 S.t55 S.n767 3.773
R744 S.n769 S.t29 3.773
R745 S.n769 S.n768 3.773
R746 S.n765 S.n766 3.773
R747 S.n765 S.t451 3.773
R748 S.t34 S.n1053 3.773
R749 S.t34 S.t513 3.773
R750 S.t34 S.t297 3.773
R751 S.t34 S.n1056 3.773
R752 S.n1058 S.t44 3.773
R753 S.n1058 S.n1057 3.773
R754 S.n1054 S.n1055 3.773
R755 S.n1054 S.t455 3.773
R756 S.t47 S.n1004 3.773
R757 S.t47 S.t229 3.773
R758 S.t47 S.t402 3.773
R759 S.t47 S.n1048 3.773
R760 S.n1050 S.t458 3.773
R761 S.n1050 S.n1049 3.773
R762 S.n1051 S.n1052 3.773
R763 S.n1051 S.t378 3.773
R764 S.t52 S.n874 3.773
R765 S.t52 S.t327 3.773
R766 S.t52 S.t543 3.773
R767 S.t52 S.n877 3.773
R768 S.n879 S.t596 3.773
R769 S.n879 S.n878 3.773
R770 S.n875 S.n876 3.773
R771 S.n875 S.t537 3.773
R772 S.t32 S.n827 3.773
R773 S.t32 S.t469 3.773
R774 S.t32 S.t62 3.773
R775 S.t32 S.n830 3.773
R776 S.n832 S.t122 3.773
R777 S.n832 S.n831 3.773
R778 S.n828 S.n829 3.773
R779 S.n828 S.t54 3.773
R780 S.n67 S.n930 3.773
R781 S.n67 S.t610 3.773
R782 S.t45 S.t216 3.773
R783 S.t45 S.n934 3.773
R784 S.n936 S.t275 3.773
R785 S.n936 S.n935 3.773
R786 S.n931 S.n932 3.773
R787 S.n931 S.t190 3.773
R788 S.t0 S.t483 3.773
R789 S.n20 S.t615 3.773
R790 S.n21 S.t220 3.773
R791 S.t34 S.n1061 3.773
R792 S.t34 S.t81 3.773
R793 S.t34 S.t300 3.773
R794 S.t34 S.n1068 3.773
R795 S.n1070 S.t250 3.773
R796 S.n1070 S.n1069 3.773
R797 S.n1059 S.n1060 3.773
R798 S.n1059 S.t22 3.773
R799 S.n90 S.n1067 3.773
R800 S.n90 S.t82 3.773
R801 S.n90 S.t309 3.773
R802 S.n90 S.n1066 3.773
R803 S.n1065 S.t253 3.773
R804 S.n1065 S.n1064 3.773
R805 S.n1062 S.n1063 3.773
R806 S.n1062 S.t27 3.773
R807 S.t32 S.n835 3.773
R808 S.t32 S.t76 3.773
R809 S.t32 S.t266 3.773
R810 S.t32 S.n836 3.773
R811 S.n838 S.t317 3.773
R812 S.n838 S.n837 3.773
R813 S.n833 S.n834 3.773
R814 S.n833 S.t257 3.773
R815 S.t0 S.t60 3.773
R816 S.n18 S.t194 3.773
R817 S.n19 S.t399 3.773
R818 S.t45 S.n939 3.773
R819 S.t45 S.t192 3.773
R820 S.t45 S.t403 3.773
R821 S.t45 S.n940 3.773
R822 S.n942 S.t460 3.773
R823 S.n942 S.n941 3.773
R824 S.n937 S.n938 3.773
R825 S.n937 S.t391 3.773
R826 S.t52 S.n882 3.773
R827 S.t52 S.t97 3.773
R828 S.t52 S.t136 3.773
R829 S.t52 S.n883 3.773
R830 S.n885 S.t260 3.773
R831 S.n885 S.n884 3.773
R832 S.n880 S.n881 3.773
R833 S.n880 S.t43 3.773
R834 S.t49 S.n724 3.773
R835 S.t49 S.t70 3.773
R836 S.t49 S.t292 3.773
R837 S.t49 S.n727 3.773
R838 S.n729 S.t236 3.773
R839 S.n729 S.n728 3.773
R840 S.n725 S.n726 3.773
R841 S.n725 S.t636 3.773
R842 S.t41 S.n639 3.773
R843 S.t41 S.t61 3.773
R844 S.t41 S.t280 3.773
R845 S.t41 S.n642 3.773
R846 S.n644 S.t228 3.773
R847 S.n644 S.n643 3.773
R848 S.n640 S.n641 3.773
R849 S.n640 S.t629 3.773
R850 S.t78 S.n595 3.773
R851 S.t78 S.t581 3.773
R852 S.t78 S.t168 3.773
R853 S.t78 S.n598 3.773
R854 S.n600 S.t117 3.773
R855 S.n600 S.n599 3.773
R856 S.n596 S.n597 3.773
R857 S.n596 S.t624 3.773
R858 S.t139 S.n473 3.773
R859 S.t139 S.t573 3.773
R860 S.t139 S.t142 3.773
R861 S.t139 S.n520 3.773
R862 S.n522 S.t112 3.773
R863 S.n522 S.n521 3.773
R864 S.n523 S.n524 3.773
R865 S.n523 S.t529 3.773
R866 S.t18 S.n525 3.773
R867 S.t18 S.t568 3.773
R868 S.t18 S.t154 3.773
R869 S.t18 S.n528 3.773
R870 S.n530 S.t107 3.773
R871 S.n530 S.n529 3.773
R872 S.n526 S.n527 3.773
R873 S.n526 S.t526 3.773
R874 S.t99 S.n382 3.773
R875 S.t99 S.t552 3.773
R876 S.t99 S.t150 3.773
R877 S.t99 S.n385 3.773
R878 S.n387 S.t535 3.773
R879 S.n387 S.n386 3.773
R880 S.n383 S.n384 3.773
R881 S.n383 S.t183 3.773
R882 S.t144 S.t276 3.773
R883 S.n400 S.t474 3.773
R884 S.n401 S.t409 3.773
R885 S.t18 S.t231 3.773
R886 S.n532 S.t342 3.773
R887 S.n533 S.t273 3.773
R888 S.t139 S.n513 3.773
R889 S.t139 S.t509 3.773
R890 S.t139 S.t365 3.773
R891 S.t139 S.n517 3.773
R892 S.n519 S.t471 3.773
R893 S.n519 S.n518 3.773
R894 S.n515 S.n516 3.773
R895 S.n515 S.t6 3.773
R896 S.t78 S.n657 3.773
R897 S.t78 S.t147 3.773
R898 S.t78 S.t360 3.773
R899 S.t78 S.n660 3.773
R900 S.n662 S.t315 3.773
R901 S.n662 S.n661 3.773
R902 S.n658 S.n659 3.773
R903 S.n658 S.t204 3.773
R904 S.t0 S.t219 3.773
R905 S.n16 S.t379 3.773
R906 S.n17 S.t591 3.773
R907 S.t45 S.n943 3.773
R908 S.t45 S.t308 3.773
R909 S.t45 S.t626 3.773
R910 S.t45 S.n946 3.773
R911 S.n948 S.t457 3.773
R912 S.n948 S.n947 3.773
R913 S.n944 S.n945 3.773
R914 S.n944 S.t246 3.773
R915 S.t32 S.n839 3.773
R916 S.t32 S.t299 3.773
R917 S.t32 S.t512 3.773
R918 S.t32 S.n842 3.773
R919 S.n844 S.t450 3.773
R920 S.n844 S.n843 3.773
R921 S.n840 S.n841 3.773
R922 S.n840 S.t248 3.773
R923 S.t52 S.n886 3.773
R924 S.t52 S.t295 3.773
R925 S.t52 S.t507 3.773
R926 S.t52 S.n889 3.773
R927 S.n891 S.t448 3.773
R928 S.n891 S.n890 3.773
R929 S.n887 S.n888 3.773
R930 S.n887 S.t245 3.773
R931 S.t47 S.n1028 3.773
R932 S.t47 S.t289 3.773
R933 S.t47 S.t502 3.773
R934 S.t47 S.n1031 3.773
R935 S.n1033 S.t440 3.773
R936 S.n1033 S.n1032 3.773
R937 S.n1029 S.n1030 3.773
R938 S.n1029 S.t241 3.773
R939 S.n83 S.n1071 3.773
R940 S.n83 S.t279 3.773
R941 S.t34 S.t484 3.773
R942 S.t34 S.n1074 3.773
R943 S.n1076 S.t336 3.773
R944 S.n1076 S.n1075 3.773
R945 S.n1072 S.n1073 3.773
R946 S.n1072 S.t234 3.773
R947 S.t55 S.n770 3.773
R948 S.t55 S.t272 3.773
R949 S.t55 S.t478 3.773
R950 S.t55 S.n773 3.773
R951 S.n775 S.t433 3.773
R952 S.n775 S.n774 3.773
R953 S.n771 S.n772 3.773
R954 S.n771 S.t230 3.773
R955 S.t49 S.n730 3.773
R956 S.t49 S.t269 3.773
R957 S.t49 S.t473 3.773
R958 S.t49 S.n733 3.773
R959 S.n735 S.t425 3.773
R960 S.n735 S.n734 3.773
R961 S.n731 S.n732 3.773
R962 S.n731 S.t222 3.773
R963 S.t41 S.n601 3.773
R964 S.t41 S.t189 3.773
R965 S.t41 S.t340 3.773
R966 S.t41 S.n652 3.773
R967 S.n654 S.t334 3.773
R968 S.n654 S.n653 3.773
R969 S.n655 S.n656 3.773
R970 S.n655 S.t210 3.773
R971 S.t78 S.t158 3.773
R972 S.n664 S.t198 3.773
R973 S.n665 S.t173 3.773
R974 S.t41 S.n645 3.773
R975 S.t41 S.t283 3.773
R976 S.t41 S.t42 3.773
R977 S.t41 S.n649 3.773
R978 S.n651 S.t618 3.773
R979 S.n651 S.n650 3.773
R980 S.n647 S.n648 3.773
R981 S.n647 S.t281 3.773
R982 S.t49 S.n791 3.773
R983 S.t49 S.t453 3.773
R984 S.t49 S.t50 3.773
R985 S.t49 S.n794 3.773
R986 S.n796 S.t487 3.773
R987 S.n796 S.n795 3.773
R988 S.n792 S.n793 3.773
R989 S.n792 S.t408 3.773
R990 S.t0 S.t427 3.773
R991 S.n14 S.t123 3.773
R992 S.n15 S.t203 3.773
R993 S.t45 S.n949 3.773
R994 S.t45 S.t489 3.773
R995 S.t45 S.t90 3.773
R996 S.t45 S.n952 3.773
R997 S.n954 S.t4 3.773
R998 S.n954 S.n953 3.773
R999 S.n950 S.n951 3.773
R1000 S.n950 S.t445 3.773
R1001 S.t32 S.n845 3.773
R1002 S.t32 S.t481 3.773
R1003 S.t32 S.t77 3.773
R1004 S.t32 S.n848 3.773
R1005 S.n850 S.t1 3.773
R1006 S.n850 S.n849 3.773
R1007 S.n846 S.n847 3.773
R1008 S.n846 S.t439 3.773
R1009 S.t52 S.n892 3.773
R1010 S.t52 S.t476 3.773
R1011 S.t52 S.t63 3.773
R1012 S.t52 S.n895 3.773
R1013 S.n897 S.t635 3.773
R1014 S.n897 S.n896 3.773
R1015 S.n893 S.n894 3.773
R1016 S.n893 S.t417 3.773
R1017 S.t47 S.n1034 3.773
R1018 S.t47 S.t470 3.773
R1019 S.t47 S.t67 3.773
R1020 S.t47 S.n1037 3.773
R1021 S.n1039 S.t627 3.773
R1022 S.n1039 S.n1038 3.773
R1023 S.n1035 S.n1036 3.773
R1024 S.n1035 S.t429 3.773
R1025 S.t34 S.n1077 3.773
R1026 S.t34 S.t466 3.773
R1027 S.t34 S.t59 3.773
R1028 S.t34 S.n1080 3.773
R1029 S.n1082 S.t623 3.773
R1030 S.n1082 S.n1081 3.773
R1031 S.n1078 S.n1079 3.773
R1032 S.n1078 S.t423 3.773
R1033 S.t55 S.n736 3.773
R1034 S.t55 S.t463 3.773
R1035 S.t55 S.t56 3.773
R1036 S.t55 S.n786 3.773
R1037 S.n788 S.t614 3.773
R1038 S.n788 S.n787 3.773
R1039 S.n789 S.n790 3.773
R1040 S.n789 S.t343 3.773
R1041 S.t0 S.t606 3.773
R1042 S.n12 S.t318 3.773
R1043 S.n13 S.t538 3.773
R1044 S.t45 S.n955 3.773
R1045 S.t45 S.t66 3.773
R1046 S.t45 S.t287 3.773
R1047 S.t45 S.n958 3.773
R1048 S.n960 S.t233 3.773
R1049 S.n960 S.n959 3.773
R1050 S.n956 S.n957 3.773
R1051 S.n956 S.t634 3.773
R1052 S.t32 S.n851 3.773
R1053 S.t32 S.t57 3.773
R1054 S.t32 S.t278 3.773
R1055 S.t32 S.n854 3.773
R1056 S.n856 S.t225 3.773
R1057 S.n856 S.n855 3.773
R1058 S.n852 S.n853 3.773
R1059 S.n852 S.t625 3.773
R1060 S.t52 S.n900 3.773
R1061 S.t52 S.t53 3.773
R1062 S.t52 S.t271 3.773
R1063 S.t52 S.n903 3.773
R1064 S.n905 S.t218 3.773
R1065 S.n905 S.n904 3.773
R1066 S.n901 S.n902 3.773
R1067 S.n901 S.t621 3.773
R1068 S.t47 S.n1042 3.773
R1069 S.t47 S.t48 3.773
R1070 S.t47 S.t268 3.773
R1071 S.t47 S.n1045 3.773
R1072 S.n1047 S.t208 3.773
R1073 S.n1047 S.n1046 3.773
R1074 S.n1043 S.n1044 3.773
R1075 S.n1043 S.t612 3.773
R1076 S.t34 S.n1085 3.773
R1077 S.t34 S.t35 3.773
R1078 S.t34 S.t186 3.773
R1079 S.t34 S.n1088 3.773
R1080 S.n1090 S.t201 3.773
R1081 S.n1090 S.n1089 3.773
R1082 S.n1086 S.n1087 3.773
R1083 S.n1086 S.t605 3.773
R1084 S.t55 S.n778 3.773
R1085 S.t55 S.t235 3.773
R1086 S.t55 S.t256 3.773
R1087 S.t55 S.n782 3.773
R1088 S.n784 S.t551 3.773
R1089 S.n784 S.n783 3.773
R1090 S.n779 S.n780 3.773
R1091 S.n779 S.t211 3.773
R1092 S.t49 S.t553 3.773
R1093 S.n798 S.t106 3.773
R1094 S.n799 S.t11 3.773
R1095 S.t0 S.t381 3.773
R1096 S.n25 S.t83 3.773
R1097 S.n24 S.t306 3.773
R1098 S.t45 S.n914 3.773
R1099 S.t45 S.t420 3.773
R1100 S.t45 S.t46 3.773
R1101 S.t45 S.n917 3.773
R1102 S.n916 S.t604 3.773
R1103 S.n916 S.n915 3.773
R1104 S.n911 S.n912 3.773
R1105 S.n911 S.t400 3.773
R1106 S.t32 S.n823 3.773
R1107 S.t32 S.t118 3.773
R1108 S.t32 S.t33 3.773
R1109 S.t32 S.n826 3.773
R1110 S.n825 S.t338 3.773
R1111 S.n825 S.n824 3.773
R1112 S.n821 S.n822 3.773
R1113 S.n821 S.t73 3.773
R1114 S.t52 S.t456 3.773
R1115 S.n907 S.t449 3.773
R1116 S.n908 S.t374 3.773
R1117 S.n1092 S.t516 3.773
R1118 S.n1093 S.t584 3.773
R1119 S.n86 S.t243 3.773
R1120 S.n86 S.n737 3.773
R1121 S.n85 S.n785 3.773
R1122 S.n85 S.t13 3.773
R1123 S.n3 S.n264 2.502
R1124 S.n4 S.n404 2.502
R1125 S.n5 S.n538 2.502
R1126 S.n6 S.n670 2.502
R1127 S.n7 S.n682 2.502
R1128 S.n71 S.n678 0.176
R1129 S.n51 S.n802 0.176
R1130 S.t2 S 0.176
R1131 S.n140 S.n262 0.171
R1132 S.n7 S.n683 0.157
R1133 S.t52 S.n909 0.152
R1134 S.t14 S.n195 0.145
R1135 S.n971 S.t0 0.141
R1136 S.t41 S.n65 0.132
R1137 S.t139 S.n63 0.132
R1138 S.t14 S.n59 0.132
R1139 S.t99 S.n61 0.131
R1140 S.t49 S.n7 0.129
R1141 S.t144 S.n310 0.127
R1142 S.t18 S.n436 0.127
R1143 S.t78 S.n561 0.127
R1144 S.t49 S.n693 0.127
R1145 S.t34 S.n976 0.127
R1146 S.n972 S.t52 0.124
R1147 S.t94 S.n230 0.123
R1148 S.n3 S.n266 0.117
R1149 S.n4 S.n405 0.117
R1150 S.n5 S.n539 0.117
R1151 S.n6 S.n671 0.117
R1152 S.n1098 S.t144 0.112
R1153 S.n1099 S.t94 0.111
R1154 S.n1097 S.t18 0.111
R1155 S.n1096 S.t78 0.111
R1156 S.n1095 S.t49 0.111
R1157 S.n1094 S.t34 0.11
R1158 S.n971 S.t45 0.11
R1159 S.t34 S.n94 0.108
R1160 S.t49 S.n93 0.108
R1161 S.t78 S.n95 0.108
R1162 S.t18 S.n92 0.108
R1163 S.t144 S.n91 0.108
R1164 S.n974 S.n973 0.101
R1165 S.n56 S.n1023 0.099
R1166 S.n974 S.n975 0.095
R1167 S.t2 S.n122 0.111
R1168 S.t45 S.n913 0.092
R1169 S.t45 S.n104 0.092
R1170 S.n53 S.n236 0.088
R1171 S.t99 S.n101 0.085
R1172 S.t139 S.n100 0.085
R1173 S.t41 S.n99 0.085
R1174 S.t55 S.n98 0.085
R1175 S.t47 S.n97 0.085
R1176 S.t139 S.n514 0.082
R1177 S.t41 S.n646 0.082
R1178 S.t32 S.n820 0.082
R1179 S.n542 S.n543 0.079
R1180 S.n673 S.n675 0.079
R1181 S.t55 S.n9 0.132
R1182 S.n666 S.n6 0.121
R1183 S.n534 S.n5 0.121
R1184 S.n406 S.n4 0.121
R1185 S.n140 S.n3 0.121
R1186 S.t18 S.n412 0.077
R1187 S.t18 S.n429 0.077
R1188 S.t78 S.n554 0.077
R1189 S.t49 S.n686 0.077
R1190 S.t78 S.n580 0.077
R1191 S.t34 S.n995 0.077
R1192 S.n235 S.n234 0.077
R1193 S.n680 S.n679 0.077
R1194 S.n69 S.n680 0.075
R1195 S.t144 S.n294 0.075
R1196 S.t144 S.n273 0.073
R1197 S.t144 S.n283 0.073
R1198 S.t18 S.n408 0.073
R1199 S.t18 S.n542 0.073
R1200 S.t78 S.n673 0.073
R1201 S.n76 S.n710 0.072
R1202 S.n81 S.n453 0.072
R1203 S.t94 S.n0 0.072
R1204 S.t144 S.n302 0.071
R1205 S.t94 S.n254 0.071
R1206 S.t34 S.n977 0.071
R1207 S.n75 S.n694 0.071
R1208 S.t78 S.n562 0.071
R1209 S.n80 S.n437 0.071
R1210 S.t144 S.n309 0.071
R1211 S.t144 S.n269 0.069
R1212 S.t144 S.n290 0.069
R1213 S.t144 S.n316 0.069
R1214 S.n71 S.n676 0.068
R1215 S.n51 S.n800 0.068
R1216 S.n541 S.n540 0.068
R1217 S.n1023 S.n1022 0.068
R1218 S.n121 S.n119 0.067
R1219 S.n133 S.n131 0.067
R1220 S.n133 S.n132 0.067
R1221 S.n129 S.n128 0.067
R1222 S.n129 S.n127 0.067
R1223 S.n122 S.n124 0.067
R1224 S.n122 S.n125 0.067
R1225 S.n108 S.n107 0.067
R1226 S.n108 S.n106 0.067
R1227 S.n121 S.n120 0.067
R1228 S.n117 S.n115 0.067
R1229 S.n111 S.n110 0.067
R1230 S.n111 S.n109 0.067
R1231 S.n117 S.n116 0.067
R1232 S.n114 S.n112 0.067
R1233 S.n114 S.n113 0.067
R1234 S.n140 S.n261 0.067
R1235 S.n140 S.n260 0.067
R1236 S.n406 S.n407 0.067
R1237 S.n534 S.n536 0.067
R1238 S.n534 S.n535 0.067
R1239 S.n666 S.n668 0.067
R1240 S.n666 S.n667 0.067
R1241 S.n406 S.n402 0.067
R1242 S.n542 S.n541 0.065
R1243 S.n673 S.n672 0.065
R1244 S.t94 S.n242 0.065
R1245 S.t144 S.n331 0.063
R1246 S.t18 S.n534 0.063
R1247 S.t78 S.n666 0.063
R1248 S.t99 S.n350 0.063
R1249 S.t18 S.n414 0.063
R1250 S.t139 S.n481 0.063
R1251 S.t78 S.n544 0.063
R1252 S.t18 S.n419 0.063
R1253 S.t144 S.n288 0.063
R1254 S.t52 S.n803 0.063
R1255 S.t34 S.n984 0.063
R1256 S.t49 S.n701 0.063
R1257 S.t78 S.n569 0.063
R1258 S.t18 S.n444 0.063
R1259 S.t144 S.n314 0.063
R1260 S.t94 S.n240 0.063
R1261 S.t99 S.n364 0.063
R1262 S.t18 S.n431 0.063
R1263 S.t139 S.n495 0.063
R1264 S.t78 S.n556 0.063
R1265 S.t41 S.n615 0.063
R1266 S.t49 S.n688 0.063
R1267 S.t55 S.n746 0.063
R1268 S.t94 S.n161 0.063
R1269 S.t144 S.n278 0.063
R1270 S.t144 S.n267 0.063
R1271 S.t94 S.n147 0.063
R1272 S.t52 S.n898 0.063
R1273 S.t47 S.n1040 0.063
R1274 S.t34 S.n1083 0.063
R1275 S.t55 S.n776 0.063
R1276 S.t55 S.n781 0.062
R1277 S.t2 S.n129 0.062
R1278 S.t2 S.n121 0.062
R1279 S.t2 S.n117 0.062
R1280 S.t2 S.n133 0.06
R1281 S.t2 S.n108 0.06
R1282 S.t2 S.n111 0.06
R1283 S.t2 S.n114 0.06
R1284 S.t45 S.n933 0.059
R1285 S.t144 S.n332 0.059
R1286 S.t52 S.n870 0.059
R1287 S.t144 S.n406 0.058
R1288 S.t52 S.n105 0.056
R1289 S.n56 S.n1024 0.056
R1290 S.t94 S.t14 0.055
R1291 S.t32 S.n103 0.055
R1292 S.t2 S.n138 0.055
R1293 S.t45 S.n910 0.054
R1294 S.t14 S.n170 0.054
R1295 S.t41 S.n602 0.054
R1296 S.t55 S.n740 0.054
R1297 S.t47 S.n1005 0.054
R1298 S.t99 S.n337 0.054
R1299 S.t139 S.n474 0.054
R1300 S.t94 S.n258 0.054
R1301 S.t144 S.n400 0.054
R1302 S.t18 S.n532 0.054
R1303 S.t78 S.n664 0.054
R1304 S.t49 S.n798 0.054
R1305 S.t52 S.n907 0.054
R1306 S.t34 S.n1093 0.054
R1307 S.t94 S.n96 0.053
R1308 S.t94 S.n102 0.053
R1309 S S.n1099 0.053
R1310 S.t47 S.n1026 0.053
R1311 S.t52 S.n865 0.053
R1312 S.t45 S.n922 0.053
R1313 S.t32 S.n858 0.053
R1314 S.t94 S.n256 0.053
R1315 S.t94 S.n159 0.053
R1316 S.t14 S.n190 0.053
R1317 S.t99 S.n353 0.053
R1318 S.t139 S.n484 0.053
R1319 S.t78 S.n588 0.053
R1320 S.t18 S.n417 0.053
R1321 S.t94 S.n167 0.053
R1322 S.t14 S.n197 0.053
R1323 S.t49 S.n717 0.053
R1324 S.t41 S.n610 0.053
R1325 S.t78 S.n550 0.053
R1326 S.t139 S.n490 0.053
R1327 S.t18 S.n425 0.053
R1328 S.t99 S.n359 0.053
R1329 S.t144 S.n297 0.053
R1330 S.t14 S.n220 0.053
R1331 S.t94 S.n228 0.053
R1332 S.t144 S.n304 0.053
R1333 S.t99 S.n367 0.053
R1334 S.t18 S.n434 0.053
R1335 S.t139 S.n498 0.053
R1336 S.t78 S.n559 0.053
R1337 S.t41 S.n618 0.053
R1338 S.t49 S.n691 0.053
R1339 S.t55 S.n749 0.053
R1340 S.t34 S.n1003 0.053
R1341 S.t144 S.n312 0.053
R1342 S.t14 S.n203 0.053
R1343 S.t94 S.n238 0.053
R1344 S.t52 S.n873 0.053
R1345 S.t47 S.n1011 0.053
R1346 S.t34 S.n982 0.053
R1347 S.t55 S.n755 0.053
R1348 S.t49 S.n699 0.053
R1349 S.t41 S.n624 0.053
R1350 S.t78 S.n567 0.053
R1351 S.t139 S.n504 0.053
R1352 S.t18 S.n442 0.053
R1353 S.t99 S.n373 0.053
R1354 S.t94 S.n248 0.053
R1355 S.t14 S.n209 0.053
R1356 S.t45 S.n929 0.053
R1357 S.t32 S.n818 0.053
R1358 S.t52 S.n809 0.053
R1359 S.t47 S.n1017 0.053
R1360 S.t34 S.n990 0.053
R1361 S.t55 S.n761 0.053
R1362 S.t49 S.n707 0.053
R1363 S.t41 S.n630 0.053
R1364 S.t78 S.n575 0.053
R1365 S.t139 S.n510 0.053
R1366 S.t18 S.n450 0.053
R1367 S.t99 S.n379 0.053
R1368 S.t144 S.n321 0.053
R1369 S.t144 S.n286 0.053
R1370 S.t94 S.n145 0.053
R1371 S.t14 S.n178 0.053
R1372 S.t94 S.n153 0.053
R1373 S.t14 S.n184 0.053
R1374 S.t18 S.n460 0.053
R1375 S.t99 S.n345 0.053
R1376 S.t144 S.n276 0.053
R1377 S.t144 S.n335 0.053
R1378 S.t14 S.n217 0.053
R1379 S.t144 S.n398 0.053
R1380 S.t99 S.n390 0.053
R1381 S.t18 S.n472 0.053
R1382 S.n78 S.n464 0.053
R1383 S.t78 S.n594 0.053
R1384 S.t41 S.n638 0.053
R1385 S.t49 S.n723 0.053
R1386 S.t55 S.n769 0.053
R1387 S.t34 S.n1058 0.053
R1388 S.t47 S.n1050 0.053
R1389 S.t52 S.n879 0.053
R1390 S.t32 S.n832 0.053
R1391 S.t45 S.n936 0.053
R1392 S.t34 S.n1070 0.053
R1393 S.n90 S.n1065 0.053
R1394 S.t32 S.n838 0.053
R1395 S.t45 S.n942 0.053
R1396 S.t52 S.n885 0.053
R1397 S.t49 S.n729 0.053
R1398 S.t41 S.n644 0.053
R1399 S.t78 S.n600 0.053
R1400 S.t139 S.n522 0.053
R1401 S.t18 S.n530 0.053
R1402 S.t99 S.n387 0.053
R1403 S.t139 S.n519 0.053
R1404 S.t78 S.n662 0.053
R1405 S.t45 S.n948 0.053
R1406 S.t32 S.n844 0.053
R1407 S.t52 S.n891 0.053
R1408 S.t47 S.n1033 0.053
R1409 S.t34 S.n1076 0.053
R1410 S.t55 S.n775 0.053
R1411 S.t49 S.n735 0.053
R1412 S.t41 S.n654 0.053
R1413 S.t41 S.n651 0.053
R1414 S.t49 S.n796 0.053
R1415 S.t45 S.n954 0.053
R1416 S.t32 S.n850 0.053
R1417 S.t52 S.n897 0.053
R1418 S.t47 S.n1039 0.053
R1419 S.t34 S.n1082 0.053
R1420 S.t55 S.n788 0.053
R1421 S.t45 S.n960 0.053
R1422 S.t32 S.n856 0.053
R1423 S.t52 S.n905 0.053
R1424 S.t47 S.n1047 0.053
R1425 S.t34 S.n1090 0.053
R1426 S.t55 S.n784 0.053
R1427 S.t45 S.n916 0.053
R1428 S.t32 S.n825 0.053
R1429 S.n675 S.n674 0.052
R1430 S.t0 S.n962 0.052
R1431 S.t94 S.n226 0.052
R1432 S.t94 S.n142 0.051
R1433 S.t94 S.n150 0.051
R1434 S.t94 S.n156 0.051
R1435 S.t94 S.n164 0.051
R1436 S.t14 S.n175 0.051
R1437 S.t14 S.n181 0.051
R1438 S.t14 S.n187 0.051
R1439 S.t14 S.n193 0.051
R1440 S.t14 S.n200 0.051
R1441 S.t14 S.n206 0.051
R1442 S.t14 S.n213 0.051
R1443 S.t14 S.n221 0.051
R1444 S.t94 S.n224 0.051
R1445 S.t94 S.n232 0.051
R1446 S.t94 S.n245 0.051
R1447 S.t94 S.n252 0.051
R1448 S.t94 S.n259 0.051
R1449 S.t144 S.n271 0.051
R1450 S.t144 S.n281 0.051
R1451 S.t144 S.n292 0.051
R1452 S.t144 S.n299 0.051
R1453 S.t144 S.n307 0.051
R1454 S.t144 S.n318 0.051
R1455 S.t144 S.n329 0.051
R1456 S.t99 S.n342 0.051
R1457 S.t99 S.n347 0.051
R1458 S.t99 S.n356 0.051
R1459 S.t99 S.n361 0.051
R1460 S.t99 S.n369 0.051
R1461 S.t99 S.n376 0.051
R1462 S.t99 S.n383 0.051
R1463 S.t99 S.n391 0.051
R1464 S.t144 S.n394 0.051
R1465 S.t144 S.n401 0.051
R1466 S.t18 S.n410 0.051
R1467 S.t18 S.n422 0.051
R1468 S.t18 S.n427 0.051
R1469 S.t18 S.n438 0.051
R1470 S.t18 S.n447 0.051
R1471 S.t18 S.n456 0.051
R1472 S.n78 S.n465 0.051
R1473 S.t18 S.n468 0.051
R1474 S.t139 S.n478 0.051
R1475 S.t139 S.n487 0.051
R1476 S.t139 S.n492 0.051
R1477 S.t139 S.n500 0.051
R1478 S.t139 S.n507 0.051
R1479 S.t139 S.n515 0.051
R1480 S.t139 S.n523 0.051
R1481 S.t18 S.n526 0.051
R1482 S.t18 S.n533 0.051
R1483 S.t78 S.n547 0.051
R1484 S.t78 S.n552 0.051
R1485 S.t78 S.n563 0.051
R1486 S.t78 S.n572 0.051
R1487 S.t78 S.n578 0.051
R1488 S.t78 S.n590 0.051
R1489 S.t78 S.n596 0.051
R1490 S.t41 S.n607 0.051
R1491 S.t41 S.n612 0.051
R1492 S.t41 S.n620 0.051
R1493 S.t41 S.n627 0.051
R1494 S.t41 S.n634 0.051
R1495 S.t41 S.n640 0.051
R1496 S.t41 S.n647 0.051
R1497 S.t41 S.n655 0.051
R1498 S.t78 S.n658 0.051
R1499 S.t78 S.n665 0.051
R1500 S.t49 S.n684 0.051
R1501 S.t49 S.n695 0.051
R1502 S.t49 S.n704 0.051
R1503 S.t49 S.n713 0.051
R1504 S.t49 S.n719 0.051
R1505 S.t49 S.n725 0.051
R1506 S.t49 S.n731 0.051
R1507 S.t55 S.n743 0.051
R1508 S.t55 S.n751 0.051
R1509 S.t55 S.n758 0.051
R1510 S.t55 S.n765 0.051
R1511 S.t55 S.n771 0.051
R1512 S.t55 S.n779 0.051
R1513 S.t55 S.n789 0.051
R1514 S.t49 S.n792 0.051
R1515 S.t49 S.n799 0.051
R1516 S.t52 S.n806 0.051
R1517 S.t32 S.n811 0.051
R1518 S.t32 S.n815 0.051
R1519 S.t32 S.n821 0.051
R1520 S.t32 S.n828 0.051
R1521 S.t32 S.n833 0.051
R1522 S.t32 S.n840 0.051
R1523 S.t32 S.n846 0.051
R1524 S.t32 S.n852 0.051
R1525 S.t52 S.n862 0.051
R1526 S.t52 S.n867 0.051
R1527 S.t52 S.n875 0.051
R1528 S.t52 S.n880 0.051
R1529 S.t52 S.n887 0.051
R1530 S.t52 S.n893 0.051
R1531 S.t52 S.n901 0.051
R1532 S.t52 S.n908 0.051
R1533 S.t45 S.n911 0.051
R1534 S.t45 S.n918 0.051
R1535 S.t45 S.n925 0.051
R1536 S.t45 S.n931 0.051
R1537 S.t45 S.n937 0.051
R1538 S.t45 S.n944 0.051
R1539 S.t45 S.n950 0.051
R1540 S.t45 S.n956 0.051
R1541 S.t34 S.n978 0.051
R1542 S.t34 S.n987 0.051
R1543 S.t34 S.n993 0.051
R1544 S.t47 S.n1007 0.051
R1545 S.t47 S.n1014 0.051
R1546 S.t47 S.n1020 0.051
R1547 S.t47 S.n1029 0.051
R1548 S.t47 S.n1035 0.051
R1549 S.t47 S.n1043 0.051
R1550 S.t47 S.n1051 0.051
R1551 S.t34 S.n1054 0.051
R1552 S.t34 S.n1059 0.051
R1553 S.n90 S.n1062 0.051
R1554 S.t34 S.n1072 0.051
R1555 S.t34 S.n1078 0.051
R1556 S.t34 S.n1086 0.051
R1557 S.t34 S.n1092 0.051
R1558 S.t55 S.n85 0.051
R1559 S.t55 S.n86 0.051
R1560 S.n583 S.n584 0.051
R1561 S.n998 S.n999 0.051
R1562 S.n324 S.n325 0.051
R1563 S.t78 S.n47 0.05
R1564 S.t49 S.n76 0.05
R1565 S.t34 S.n46 0.05
R1566 S.t18 S.n81 0.05
R1567 S.t144 S.n2 0.05
R1568 S.t34 S.n45 0.048
R1569 S.t34 S.n44 0.048
R1570 S.t2 S.n37 0.046
R1571 S.t2 S.n40 0.046
R1572 S.t18 S.n78 0.046
R1573 S.t18 S.t139 0.046
R1574 S.t2 S.n43 0.045
R1575 S.t78 S.t41 0.044
R1576 S.t49 S.t55 0.044
R1577 S.t78 S.n49 0.044
R1578 S.t49 S.n73 0.044
R1579 S.t52 S.n50 0.044
R1580 S.t49 S.n70 0.044
R1581 S.n139 S.t2 0.08
R1582 S.t49 S.n71 0.038
R1583 S.t18 S.n80 0.037
R1584 S.t49 S.n75 0.037
R1585 S.n53 S.n235 0.035
R1586 S.t55 S.n87 0.034
R1587 S.t18 S.n82 0.034
R1588 S.t0 S.n11 0.034
R1589 S.t0 S.n22 0.034
R1590 S.t0 S.n23 0.034
R1591 S.t2 S.n30 0.034
R1592 S.t2 S.n29 0.034
R1593 S.t2 S.n38 0.034
R1594 S.t2 S.n39 0.034
R1595 S.t2 S.n35 0.034
R1596 S.t2 S.n36 0.034
R1597 S.t2 S.n33 0.034
R1598 S.t2 S.n34 0.034
R1599 S.t2 S.n31 0.034
R1600 S.t2 S.n32 0.034
R1601 S.t2 S.n41 0.034
R1602 S.t2 S.n42 0.034
R1603 S.t2 S.n28 0.034
R1604 S.t2 S.n27 0.034
R1605 S.t0 S.n21 0.034
R1606 S.t0 S.n20 0.034
R1607 S.t0 S.n19 0.034
R1608 S.t0 S.n18 0.034
R1609 S.t0 S.n17 0.034
R1610 S.t0 S.n16 0.034
R1611 S.t0 S.n15 0.034
R1612 S.t0 S.n14 0.034
R1613 S.t0 S.n13 0.034
R1614 S.t0 S.n12 0.034
R1615 S.t0 S.n24 0.034
R1616 S.t0 S.n25 0.034
R1617 S.t49 S.n69 0.032
R1618 S.t18 S.n79 0.032
R1619 S.t49 S.n72 0.032
R1620 S.n1099 S.n1098 0.031
R1621 S.n1098 S.n1097 0.031
R1622 S.n1097 S.n1096 0.031
R1623 S.n1096 S.n1095 0.031
R1624 S.n1095 S.n1094 0.031
R1625 S.n1094 S.n972 0.031
R1626 S.n972 S.n971 0.031
R1627 S.n583 S.n585 0.022
R1628 S.n998 S.n1000 0.022
R1629 S.n324 S.n326 0.022
R1630 S.n47 S.n583 0.021
R1631 S.n240 S.n241 0.021
R1632 S.n46 S.n998 0.021
R1633 S.n161 S.n162 0.021
R1634 S.n2 S.n324 0.021
R1635 S.n147 S.n148 0.021
R1636 S.n242 S.n243 0.02
R1637 S.n47 S.n582 0.02
R1638 S.n76 S.n711 0.02
R1639 S.n46 S.n997 0.02
R1640 S.n81 S.n454 0.02
R1641 S.n2 S.n327 0.02
R1642 S.n408 S.n409 0.015
R1643 S.n283 S.n284 0.015
R1644 S.n294 S.n295 0.015
R1645 S.n273 S.n274 0.015
R1646 S.n676 S.n677 0.014
R1647 S.n800 S.n801 0.014
R1648 S.n350 S.n351 0.008
R1649 S.n414 S.n415 0.008
R1650 S.n481 S.n482 0.008
R1651 S.n544 S.n545 0.008
R1652 S.n419 S.n420 0.008
R1653 S.n288 S.n289 0.008
R1654 S.n803 S.n804 0.008
R1655 S.n984 S.n985 0.008
R1656 S.n701 S.n702 0.008
R1657 S.n569 S.n570 0.008
R1658 S.n444 S.n445 0.008
R1659 S.n314 S.n315 0.008
R1660 S.n364 S.n365 0.008
R1661 S.n431 S.n432 0.008
R1662 S.n495 S.n496 0.008
R1663 S.n556 S.n557 0.008
R1664 S.n615 S.n616 0.008
R1665 S.n688 S.n689 0.008
R1666 S.n746 S.n747 0.008
R1667 S.n278 S.n279 0.008
R1668 S.n267 S.n268 0.008
R1669 S.n898 S.n899 0.008
R1670 S.n1040 S.n1041 0.008
R1671 S.n1083 S.n1084 0.008
R1672 S.n776 S.n777 0.008
R1673 S.t34 S.n974 0.097
R1674 S.t52 S.t32 0.085
R1675 S.t34 S.t47 0.083
R1676 S.t144 S.t99 0.083
R1677 S.t78 S.n48 0.081
R1678 S.n9 S.n8 0.077
R1679 S.t52 S.n51 0.073
R1680 S.t0 S.n10 0.071
R1681 S.t94 S.n1 0.07
R1682 S.t139 S.n54 0.069
R1683 S.t32 S.n58 0.069
R1684 S.t2 S.n26 0.068
R1685 S.n65 S.n66 0.067
R1686 S.n63 S.n64 0.067
R1687 S.n61 S.n62 0.067
R1688 S.n59 S.n60 0.067
R1689 S.t2 S.n55 0.065
R1690 S.t144 S.n52 0.064
R1691 S.t99 S.n57 0.063
R1692 S.t94 S.n140 0.062
R1693 S.t45 S.n67 0.062
R1694 S.t49 S.n74 0.061
R1695 S.t78 S.n68 0.061
R1696 S.t18 S.n77 0.06
R1697 S.t34 S.n83 0.059
R1698 S.t94 S.n53 0.058
R1699 S.t52 S.n84 0.058
R1700 S.t47 S.n56 0.058
R1701 S.t55 S.n88 0.055
R1702 S.t34 S.n90 0.054
R1703 S.t41 S.n89 0.053
R1704 D.n1136 D.n1135 41.943
R1705 D.n1135 D.n1134 8.553
R1706 D.n1123 D.t89 4.386
R1707 D.n1078 D.t299 4.386
R1708 D.n1061 D.t491 4.386
R1709 D.n1059 D.t85 4.386
R1710 D.n1103 D.t253 4.386
R1711 D.n1760 D.t569 4.386
R1712 D.n1774 D.t120 4.386
R1713 D.n1772 D.t338 4.386
R1714 D.n1794 D.t134 4.386
R1715 D.n1792 D.t347 4.386
R1716 D.n1814 D.t249 4.386
R1717 D.n1812 D.t457 4.386
R1718 D.n1834 D.t267 4.386
R1719 D.n1832 D.t472 4.386
R1720 D.n1854 D.t279 4.386
R1721 D.n1852 D.t192 4.386
R1722 D.n1874 D.t234 4.386
R1723 D.n1872 D.t442 4.386
R1724 D.n1893 D.t470 4.386
R1725 D.n1891 D.t69 4.386
R1726 D.n1883 D.t365 4.386
R1727 D.n1880 D.t581 4.386
R1728 D.n1864 D.t110 4.386
R1729 D.n1861 D.t300 4.386
R1730 D.n1844 D.t271 4.386
R1731 D.n1841 D.t477 4.386
R1732 D.n1824 D.t260 4.386
R1733 D.n1821 D.t466 4.386
R1734 D.n1804 D.t140 4.386
R1735 D.n1801 D.t354 4.386
R1736 D.n1784 D.t128 4.386
R1737 D.n1781 D.t342 4.386
R1738 D.n1754 D.t244 4.386
R1739 D.n1751 D.t329 4.386
R1740 D.n1591 D.t516 4.386
R1741 D.n1615 D.t328 4.386
R1742 D.n1613 D.t540 4.386
R1743 D.n1635 D.t439 4.386
R1744 D.n1633 D.t38 4.386
R1745 D.n1655 D.t451 4.386
R1746 D.n1653 D.t51 4.386
R1747 D.n1675 D.t465 4.386
R1748 D.n1673 D.t66 4.386
R1749 D.n1695 D.t476 4.386
R1750 D.n1693 D.t53 4.386
R1751 D.n1715 D.t48 4.386
R1752 D.n1713 D.t262 4.386
R1753 D.n1704 D.t598 4.386
R1754 D.n1701 D.t154 4.386
R1755 D.n1684 D.t471 4.386
R1756 D.n1681 D.t70 4.386
R1757 D.n1664 D.t455 4.386
R1758 D.n1661 D.t57 4.386
R1759 D.n1644 D.t445 4.386
R1760 D.n1641 D.t44 4.386
R1761 D.n1624 D.t337 4.386
R1762 D.n1621 D.t546 4.386
R1763 D.n1604 D.t194 4.386
R1764 D.n1601 D.t532 4.386
R1765 D.n1467 D.t473 4.386
R1766 D.n1481 D.t20 4.386
R1767 D.n1479 D.t231 4.386
R1768 D.n1501 D.t33 4.386
R1769 D.n1499 D.t243 4.386
R1770 D.n1521 D.t42 4.386
R1771 D.n1519 D.t258 4.386
R1772 D.n1541 D.t54 4.386
R1773 D.n1539 D.t269 4.386
R1774 D.n1560 D.t453 4.386
R1775 D.n1558 D.t483 4.386
R1776 D.n1550 D.t64 4.386
R1777 D.n1547 D.t278 4.386
R1778 D.n1531 D.t50 4.386
R1779 D.n1528 D.t264 4.386
R1780 D.n1511 D.t36 4.386
R1781 D.n1508 D.t247 4.386
R1782 D.n1491 D.t27 4.386
R1783 D.n1488 D.t236 4.386
R1784 D.n1461 D.t129 4.386
R1785 D.n1458 D.t118 4.386
R1786 D.n1338 D.t252 4.386
R1787 D.n1362 D.t220 4.386
R1788 D.n1360 D.t433 4.386
R1789 D.n1382 D.t235 4.386
R1790 D.n1380 D.t443 4.386
R1791 D.n1402 D.t246 4.386
R1792 D.n1400 D.t454 4.386
R1793 D.n1422 D.t34 4.386
R1794 D.n1420 D.t245 4.386
R1795 D.n1411 D.t256 4.386
R1796 D.n1408 D.t463 4.386
R1797 D.n1391 D.t239 4.386
R1798 D.n1388 D.t449 4.386
R1799 D.n1371 D.t230 4.386
R1800 D.n1368 D.t437 4.386
R1801 D.n1351 D.t521 4.386
R1802 D.n1348 D.t424 4.386
R1803 D.n1254 D.t199 4.386
R1804 D.n1268 D.t423 4.386
R1805 D.n1266 D.t26 4.386
R1806 D.n1288 D.t436 4.386
R1807 D.n1286 D.t35 4.386
R1808 D.n1307 D.t227 4.386
R1809 D.n1305 D.t435 4.386
R1810 D.n1297 D.t441 4.386
R1811 D.n1294 D.t41 4.386
R1812 D.n1278 D.t432 4.386
R1813 D.n1275 D.t31 4.386
R1814 D.n1248 D.t480 4.386
R1815 D.n1245 D.t18 4.386
R1816 D.n1165 D.t138 4.386
R1817 D.n1189 D.t17 4.386
R1818 D.n1187 D.t228 4.386
R1819 D.n1209 D.t415 4.386
R1820 D.n1207 D.t15 4.386
R1821 D.n1198 D.t25 4.386
R1822 D.n1195 D.t233 4.386
R1823 D.n1178 D.t426 4.386
R1824 D.n1175 D.t218 4.386
R1825 D.n16 D.t533 4.386
R1826 D.n14 D.t130 4.386
R1827 D.n36 D.t547 4.386
R1828 D.n34 D.t143 4.386
R1829 D.n56 D.t557 4.386
R1830 D.n54 D.t153 4.386
R1831 D.n76 D.t58 4.386
R1832 D.n74 D.t273 4.386
R1833 D.n96 D.t71 4.386
R1834 D.n94 D.t324 4.386
R1835 D.n116 D.t364 4.386
R1836 D.n114 D.t578 4.386
R1837 D.n136 D.t43 4.386
R1838 D.n134 D.t259 4.386
R1839 D.n172 D.t282 4.386
R1840 D.n169 D.t488 4.386
R1841 D.n147 D.t182 4.386
R1842 D.n144 D.t396 4.386
R1843 D.n126 D.t507 4.386
R1844 D.n123 D.t102 4.386
R1845 D.n106 D.t266 4.386
R1846 D.n103 D.t440 4.386
R1847 D.n86 D.t67 4.386
R1848 D.n83 D.t280 4.386
R1849 D.n66 D.t565 4.386
R1850 D.n63 D.t160 4.386
R1851 D.n46 D.t552 4.386
R1852 D.n43 D.t148 4.386
R1853 D.n26 D.t541 4.386
R1854 D.n23 D.t135 4.386
R1855 D.n4 D.t296 4.386
R1856 D.n1 D.t122 4.386
R1857 D.n232 D.t343 4.386
R1858 D.n230 D.t553 4.386
R1859 D.n411 D.t606 4.386
R1860 D.n400 D.t464 4.386
R1861 D.n398 D.t65 4.386
R1862 D.n386 D.t316 4.386
R1863 D.n384 D.t525 4.386
R1864 D.n372 D.t179 4.386
R1865 D.n370 D.t393 4.386
R1866 D.n358 D.t40 4.386
R1867 D.n356 D.t255 4.386
R1868 D.n344 D.t504 4.386
R1869 D.n342 D.t99 4.386
R1870 D.n330 D.t401 4.386
R1871 D.n328 D.t575 4.386
R1872 D.n316 D.t479 4.386
R1873 D.n314 D.t469 4.386
R1874 D.n302 D.t377 4.386
R1875 D.n300 D.t591 4.386
R1876 D.n288 D.t366 4.386
R1877 D.n286 D.t579 4.386
R1878 D.n274 D.t360 4.386
R1879 D.n272 D.t570 4.386
R1880 D.n260 D.t357 4.386
R1881 D.n258 D.t566 4.386
R1882 D.n246 D.t348 4.386
R1883 D.n244 D.t558 4.386
R1884 D.n220 D.t340 4.386
R1885 D.n218 D.t549 4.386
R1886 D.n443 D.t149 4.386
R1887 D.n441 D.t361 4.386
R1888 D.n594 D.t121 4.386
R1889 D.n583 D.t604 4.386
R1890 D.n581 D.t203 4.386
R1891 D.n569 D.t460 4.386
R1892 D.n567 D.t61 4.386
R1893 D.n555 D.t313 4.386
R1894 D.n553 D.t522 4.386
R1895 D.n541 D.t174 4.386
R1896 D.n539 D.t389 4.386
R1897 D.n527 D.t39 4.386
R1898 D.n525 D.t251 4.386
R1899 D.n513 D.t486 4.386
R1900 D.n511 D.t55 4.386
R1901 D.n499 D.t180 4.386
R1902 D.n497 D.t551 4.386
R1903 D.n485 D.t170 4.386
R1904 D.n483 D.t385 4.386
R1905 D.n471 D.t163 4.386
R1906 D.n469 D.t379 4.386
R1907 D.n457 D.t155 4.386
R1908 D.n455 D.t369 4.386
R1909 D.n431 D.t144 4.386
R1910 D.n429 D.t359 4.386
R1911 D.n623 D.t573 4.386
R1912 D.n621 D.t172 4.386
R1913 D.n746 D.t275 4.386
R1914 D.n735 D.t116 4.386
R1915 D.n733 D.t336 4.386
R1916 D.n721 D.t601 4.386
R1917 D.n719 D.t200 4.386
R1918 D.n707 D.t458 4.386
R1919 D.n705 D.t59 4.386
R1920 D.n693 D.t270 4.386
R1921 D.n691 D.t478 4.386
R1922 D.n679 D.t113 4.386
R1923 D.n677 D.t330 4.386
R1924 D.n665 D.t13 4.386
R1925 D.n663 D.t196 4.386
R1926 D.n651 D.t592 4.386
R1927 D.n649 D.t81 4.386
R1928 D.n637 D.t582 4.386
R1929 D.n635 D.t183 4.386
R1930 D.n611 D.t568 4.386
R1931 D.n609 D.t166 4.386
R1932 D.n775 D.t387 4.386
R1933 D.n773 D.t223 4.386
R1934 D.n870 D.t410 4.386
R1935 D.n859 D.t272 4.386
R1936 D.n857 D.t482 4.386
R1937 D.n845 D.t75 4.386
R1938 D.n843 D.t286 4.386
R1939 D.n831 D.t542 4.386
R1940 D.n829 D.t136 4.386
R1941 D.n817 D.t406 4.386
R1942 D.n815 D.t4 4.386
R1943 D.n803 D.t268 4.386
R1944 D.n801 D.t475 4.386
R1945 D.n789 D.t147 4.386
R1946 D.n787 D.t326 4.386
R1947 D.n763 D.t381 4.386
R1948 D.n761 D.t595 4.386
R1949 D.n899 D.t404 4.386
R1950 D.n897 D.t2 4.386
R1951 D.n966 D.t494 4.386
R1952 D.n955 D.t350 4.386
R1953 D.n953 D.t560 4.386
R1954 D.n941 D.t214 4.386
R1955 D.n939 D.t425 4.386
R1956 D.n927 D.t73 4.386
R1957 D.n925 D.t284 4.386
R1958 D.n913 D.t539 4.386
R1959 D.n911 D.t133 4.386
R1960 D.n887 D.t293 4.386
R1961 D.n885 D.t474 4.386
R1962 D.n995 D.t212 4.386
R1963 D.n993 D.t421 4.386
R1964 D.n1036 D.t28 4.386
R1965 D.n1023 D.t492 4.386
R1966 D.n1021 D.t86 4.386
R1967 D.n1009 D.t346 4.386
R1968 D.n1007 D.t556 4.386
R1969 D.n983 D.t72 4.386
R1970 D.n981 D.t283 4.386
R1971 D.n1046 D.t152 4.386
R1972 D.n1070 D.t23 4.386
R1973 D.n1067 D.t232 4.386
R1974 D.n1117 D.t367 4.386
R1975 D.n1114 D.t420 4.386
R1976 D.n1133 D.t207 4.386
R1977 D.n1139 D.t610 4.386
R1978 D.n1154 D.t132 4.327
R1979 D.n1062 D.t139 4.327
R1980 D.n1058 D.t76 4.327
R1981 D.n1100 D.t535 4.327
R1982 D.n1775 D.t287 4.327
R1983 D.n1771 D.t80 4.327
R1984 D.n1795 D.t297 4.327
R1985 D.n1791 D.t88 4.327
R1986 D.n1815 D.t405 4.327
R1987 D.n1811 D.t201 4.327
R1988 D.n1835 D.t416 4.327
R1989 D.n1831 D.t211 4.327
R1990 D.n1855 D.t428 4.327
R1991 D.n1851 D.t225 4.327
R1992 D.n1875 D.t499 4.327
R1993 D.n1871 D.t434 4.327
R1994 D.n1894 D.t162 4.327
R1995 D.n1890 D.t37 4.327
R1996 D.n1911 D.t248 4.327
R1997 D.n1884 D.t32 4.327
R1998 D.n1881 D.t567 4.327
R1999 D.n1865 D.t353 4.327
R2000 D.n1862 D.t290 4.327
R2001 D.n1845 D.t419 4.327
R2002 D.n1842 D.t216 4.327
R2003 D.n1825 D.t411 4.327
R2004 D.n1822 D.t208 4.327
R2005 D.n1805 D.t302 4.327
R2006 D.n1802 D.t195 4.327
R2007 D.n1785 D.t294 4.327
R2008 D.n1782 D.t83 4.327
R2009 D.n1755 D.t241 4.327
R2010 D.n1752 D.t506 4.327
R2011 D.n1616 D.t489 4.327
R2012 D.n1612 D.t285 4.327
R2013 D.n1636 D.t597 4.327
R2014 D.n1632 D.t390 4.327
R2015 D.n1656 D.t609 4.327
R2016 D.n1652 D.t403 4.327
R2017 D.n1676 D.t6 4.327
R2018 D.n1672 D.t414 4.327
R2019 D.n1696 D.t21 4.327
R2020 D.n1692 D.t427 4.327
R2021 D.n1716 D.t358 4.327
R2022 D.n1712 D.t229 4.327
R2023 D.n1732 D.t438 4.327
R2024 D.n1705 D.t221 4.327
R2025 D.n1702 D.t141 4.327
R2026 D.n1685 D.t11 4.327
R2027 D.n1682 D.t418 4.327
R2028 D.n1665 D.t1 4.327
R2029 D.n1662 D.t408 4.327
R2030 D.n1645 D.t602 4.327
R2031 D.n1642 D.t398 4.327
R2032 D.n1625 D.t493 4.327
R2033 D.n1622 D.t383 4.327
R2034 D.n1605 D.t164 4.327
R2035 D.n1602 D.t444 4.327
R2036 D.n1482 D.t168 4.327
R2037 D.n1478 D.t576 4.327
R2038 D.n1502 D.t187 4.327
R2039 D.n1498 D.t596 4.327
R2040 D.n1522 D.t198 4.327
R2041 D.n1518 D.t608 4.327
R2042 D.n1542 D.t210 4.327
R2043 D.n1538 D.t5 4.327
R2044 D.n1561 D.t224 4.327
R2045 D.n1557 D.t392 4.327
R2046 D.n1577 D.t19 4.327
R2047 D.n1551 D.t215 4.327
R2048 D.n1548 D.t10 4.327
R2049 D.n1532 D.t206 4.327
R2050 D.n1529 D.t0 4.327
R2051 D.n1512 D.t193 4.327
R2052 D.n1509 D.t600 4.327
R2053 D.n1492 D.t175 4.327
R2054 D.n1489 D.t587 4.327
R2055 D.n1462 D.t97 4.327
R2056 D.n1459 D.t589 4.327
R2057 D.n1363 D.t374 4.327
R2058 D.n1359 D.t167 4.327
R2059 D.n1383 D.t388 4.327
R2060 D.n1379 D.t184 4.327
R2061 D.n1403 D.t402 4.327
R2062 D.n1399 D.t197 4.327
R2063 D.n1423 D.t413 4.327
R2064 D.n1419 D.t577 4.327
R2065 D.n1439 D.t177 4.327
R2066 D.n1412 D.t407 4.327
R2067 D.n1409 D.t205 4.327
R2068 D.n1392 D.t397 4.327
R2069 D.n1389 D.t190 4.327
R2070 D.n1372 D.t382 4.327
R2071 D.n1369 D.t173 4.327
R2072 D.n1352 D.t250 4.327
R2073 D.n1349 D.t515 4.327
R2074 D.n1269 D.t574 4.327
R2075 D.n1265 D.t370 4.327
R2076 D.n1289 D.t593 4.327
R2077 D.n1285 D.t386 4.327
R2078 D.n1308 D.t607 4.327
R2079 D.n1304 D.t151 4.327
R2080 D.n1324 D.t363 4.327
R2081 D.n1298 D.t599 4.327
R2082 D.n1295 D.t395 4.327
R2083 D.n1279 D.t583 4.327
R2084 D.n1276 D.t380 4.327
R2085 D.n1249 D.t176 4.327
R2086 D.n1246 D.t452 4.327
R2087 D.n1190 D.t165 4.327
R2088 D.n1186 D.t572 4.327
R2089 D.n1210 D.t181 4.327
R2090 D.n1206 D.t345 4.327
R2091 D.n1226 D.t555 4.327
R2092 D.n1199 D.t171 4.327
R2093 D.n1196 D.t580 4.327
R2094 D.n1179 D.t103 4.327
R2095 D.n1176 D.t384 4.327
R2096 D.n17 D.t82 4.327
R2097 D.n13 D.t490 4.327
R2098 D.n37 D.t90 4.327
R2099 D.n33 D.t501 4.327
R2100 D.n57 D.t98 4.327
R2101 D.n53 D.t509 4.327
R2102 D.n77 D.t213 4.327
R2103 D.n73 D.t8 4.327
R2104 D.n97 D.t226 4.327
R2105 D.n93 D.t22 4.327
R2106 D.n117 D.t30 4.327
R2107 D.n113 D.t564 4.327
R2108 D.n137 D.t308 4.327
R2109 D.n133 D.t242 4.327
R2110 D.n173 D.t594 4.327
R2111 D.n170 D.t456 4.327
R2112 D.n148 D.t450 4.327
R2113 D.n145 D.t378 4.327
R2114 D.n127 D.t159 4.327
R2115 D.n124 D.t93 4.327
R2116 D.n107 D.t496 4.327
R2117 D.n104 D.t429 4.327
R2118 D.n87 D.t217 4.327
R2119 D.n84 D.t14 4.327
R2120 D.n67 D.t105 4.327
R2121 D.n64 D.t3 4.327
R2122 D.n47 D.t95 4.327
R2123 D.n44 D.t503 4.327
R2124 D.n27 D.t84 4.327
R2125 D.n24 D.t495 4.327
R2126 D.n5 D.t304 4.327
R2127 D.n2 D.t571 4.327
R2128 D.n212 D.t288 4.327
R2129 D.n233 D.t502 4.327
R2130 D.n229 D.t298 4.327
R2131 D.n401 D.t109 4.327
R2132 D.n397 D.t52 4.327
R2133 D.n387 D.t590 4.327
R2134 D.n383 D.t514 4.327
R2135 D.n373 D.t448 4.327
R2136 D.n369 D.t376 4.327
R2137 D.n359 D.t305 4.327
R2138 D.n355 D.t238 4.327
R2139 D.n345 D.t158 4.327
R2140 D.n341 D.t91 4.327
R2141 D.n331 D.t29 4.327
R2142 D.n327 D.t562 4.327
R2143 D.n317 D.t24 4.327
R2144 D.n313 D.t430 4.327
R2145 D.n303 D.t528 4.327
R2146 D.n299 D.t422 4.327
R2147 D.n289 D.t520 4.327
R2148 D.n285 D.t319 4.327
R2149 D.n275 D.t517 4.327
R2150 D.n271 D.t312 4.327
R2151 D.n261 D.t511 4.327
R2152 D.n257 D.t309 4.327
R2153 D.n247 D.t505 4.327
R2154 D.n243 D.t303 4.327
R2155 D.n221 D.t497 4.327
R2156 D.n217 D.t295 4.327
R2157 D.n423 D.t92 4.327
R2158 D.n444 D.t310 4.327
R2159 D.n440 D.t100 4.327
R2160 D.n584 D.t263 4.327
R2161 D.n580 D.t189 4.327
R2162 D.n570 D.t107 4.327
R2163 D.n566 D.t49 4.327
R2164 D.n556 D.t584 4.327
R2165 D.n552 D.t510 4.327
R2166 D.n542 D.t446 4.327
R2167 D.n538 D.t371 4.327
R2168 D.n528 D.t301 4.327
R2169 D.n524 D.t237 4.327
R2170 D.n514 D.t101 4.327
R2171 D.n510 D.t87 4.327
R2172 D.n500 D.t333 4.327
R2173 D.n496 D.t125 4.327
R2174 D.n486 D.t325 4.327
R2175 D.n482 D.t115 4.327
R2176 D.n472 D.t320 4.327
R2177 D.n468 D.t111 4.327
R2178 D.n458 D.t314 4.327
R2179 D.n454 D.t106 4.327
R2180 D.n432 D.t306 4.327
R2181 D.n428 D.t96 4.327
R2182 D.n603 D.t513 4.327
R2183 D.n624 D.t112 4.327
R2184 D.n620 D.t523 4.327
R2185 D.n736 D.t399 4.327
R2186 D.n732 D.t321 4.327
R2187 D.n722 D.t261 4.327
R2188 D.n718 D.t188 4.327
R2189 D.n708 D.t104 4.327
R2190 D.n704 D.t45 4.327
R2191 D.n694 D.t526 4.327
R2192 D.n690 D.t508 4.327
R2193 D.n680 D.t394 4.327
R2194 D.n676 D.t317 4.327
R2195 D.n666 D.t257 4.327
R2196 D.n662 D.t178 4.327
R2197 D.n652 D.t126 4.327
R2198 D.n648 D.t537 4.327
R2199 D.n638 D.t117 4.327
R2200 D.n634 D.t529 4.327
R2201 D.n612 D.t108 4.327
R2202 D.n608 D.t518 4.327
R2203 D.n755 D.t322 4.327
R2204 D.n776 D.t538 4.327
R2205 D.n772 D.t334 4.327
R2206 D.n860 D.t527 4.327
R2207 D.n856 D.t467 4.327
R2208 D.n846 D.t339 4.327
R2209 D.n842 D.t318 4.327
R2210 D.n832 D.t204 4.327
R2211 D.n828 D.t123 4.327
R2212 D.n818 D.t63 4.327
R2213 D.n814 D.t605 4.327
R2214 D.n804 D.t524 4.327
R2215 D.n800 D.t462 4.327
R2216 D.n790 D.t391 4.327
R2217 D.n786 D.t315 4.327
R2218 D.n764 D.t531 4.327
R2219 D.n760 D.t327 4.327
R2220 D.n879 D.t127 4.327
R2221 D.n900 D.t60 4.327
R2222 D.n896 D.t603 4.327
R2223 D.n956 D.t9 4.327
R2224 D.n952 D.t548 4.327
R2225 D.n942 D.t485 4.327
R2226 D.n938 D.t412 4.327
R2227 D.n928 D.t335 4.327
R2228 D.n924 D.t277 4.327
R2229 D.n914 D.t202 4.327
R2230 D.n910 D.t119 4.327
R2231 D.n888 D.t519 4.327
R2232 D.n884 D.t459 4.327
R2233 D.n975 D.t114 4.327
R2234 D.n996 D.t481 4.327
R2235 D.n992 D.t409 4.327
R2236 D.n1024 D.t142 4.327
R2237 D.n1020 D.t78 4.327
R2238 D.n1010 D.t7 4.327
R2239 D.n1006 D.t545 4.327
R2240 D.n984 D.t332 4.327
R2241 D.n980 D.t274 4.327
R2242 D.n1071 D.t289 4.327
R2243 D.n1068 D.t219 4.327
R2244 D.n1052 D.t544 4.327
R2245 D.n1083 D.t352 4.327
R2246 D.n1118 D.t47 4.327
R2247 D.n1115 D.t311 4.327
R2248 D.n1136 D.t368 4.327
R2249 D.n1138 D.t536 4.327
R2250 D.n1155 D.t62 4.091
R2251 D.n1101 D.t46 4.091
R2252 D.n1912 D.t585 4.091
R2253 D.n1733 D.t156 4.091
R2254 D.n1578 D.t349 4.091
R2255 D.n1440 D.t94 4.091
R2256 D.n1325 D.t291 4.091
R2257 D.n1227 D.t484 4.091
R2258 D.n213 D.t331 4.091
R2259 D.n424 D.t137 4.091
R2260 D.n604 D.t561 4.091
R2261 D.n756 D.t373 4.091
R2262 D.n880 D.t186 4.091
R2263 D.n976 D.t534 4.091
R2264 D.n1053 D.t554 4.091
R2265 D.n1084 D.t362 4.091
R2266 D.n194 D.t56 4.084
R2267 D.n1124 D.t341 4.083
R2268 D.n1079 D.t563 4.083
R2269 D.n1104 D.t209 4.083
R2270 D.n1761 D.t512 4.083
R2271 D.n1592 D.t375 4.083
R2272 D.n1468 D.t240 4.083
R2273 D.n1339 D.t145 4.083
R2274 D.n1255 D.t12 4.083
R2275 D.n1166 D.t487 4.083
R2276 D.n9 D.t588 4.083
R2277 D.n412 D.t265 4.083
R2278 D.n595 D.t400 4.083
R2279 D.n747 D.t530 4.083
R2280 D.n871 D.t68 4.083
R2281 D.n967 D.t146 4.083
R2282 D.n1037 D.t292 4.083
R2283 D.n1047 D.t431 4.083
R2284 D.n9 D.t16 4.06
R2285 D.n194 D.t185 4.06
R2286 D.n1156 D.t461 4.057
R2287 D.n1102 D.t254 4.057
R2288 D.n1913 D.t372 4.057
R2289 D.n1734 D.t559 4.057
R2290 D.n1579 D.t169 4.057
R2291 D.n1441 D.t500 4.057
R2292 D.n1326 D.t77 4.057
R2293 D.n1228 D.t276 4.057
R2294 D.n214 D.t543 4.057
R2295 D.n425 D.t351 4.057
R2296 D.n605 D.t157 4.057
R2297 D.n757 D.t586 4.057
R2298 D.n881 D.t356 4.057
R2299 D.n977 D.t131 4.057
R2300 D.n1054 D.t344 4.057
R2301 D.n1085 D.t150 4.057
R2302 D.n1122 D.t281 4.031
R2303 D.n1080 D.t498 4.031
R2304 D.n1105 D.t74 4.031
R2305 D.n1759 D.t447 4.031
R2306 D.n1590 D.t307 4.031
R2307 D.n1466 D.t161 4.031
R2308 D.n1337 D.t79 4.031
R2309 D.n1253 D.t550 4.031
R2310 D.n1164 D.t417 4.031
R2311 D.n413 D.t191 4.031
R2312 D.n596 D.t323 4.031
R2313 D.n748 D.t468 4.031
R2314 D.n872 D.t611 4.031
R2315 D.n968 D.t124 4.031
R2316 D.n1038 D.t222 4.031
R2317 D.n1045 D.t355 4.031
R2318 D.n209 D.n208 0.31
R2319 D.n1107 D.n1106 0.24
R2320 D.n1044 D.n1043 0.225
R2321 D.n418 D.n417 0.225
R2322 D.n598 D.n597 0.225
R2323 D.n750 D.n749 0.225
R2324 D.n874 D.n873 0.225
R2325 D.n970 D.n969 0.225
R2326 D.n1040 D.n1039 0.225
R2327 D.n1050 D.n1049 0.225
R2328 D.n1065 D.n1055 0.203
R2329 D.n177 D.n175 0.174
R2330 D.n1161 D.n1109 0.16
R2331 D.n1922 D.n1921 0.156
R2332 D.n1584 D.n1583 0.156
R2333 D.n1331 D.n1330 0.156
R2334 D.n1158 D.n1157 0.156
R2335 D.n177 D.n176 0.156
R2336 D.n1108 D.n1096 0.143
R2337 D.n1923 D.n1747 0.143
R2338 D.n1744 D.n1743 0.143
R2339 D.n1744 D.n1588 0.143
R2340 D.n1585 D.n1454 0.143
R2341 D.n1451 D.n1450 0.143
R2342 D.n1451 D.n1335 0.143
R2343 D.n1332 D.n1241 0.143
R2344 D.n1238 D.n1237 0.143
R2345 D.n1238 D.n1162 0.143
R2346 D.n1159 D.n1110 0.143
R2347 D.n179 D.n178 0.143
R2348 D.n1088 D.n1087 0.143
R2349 D.n1099 D.n1097 0.133
R2350 D.n1741 D.n1735 0.128
R2351 D.n1448 D.n1442 0.128
R2352 D.n1235 D.n1229 0.128
R2353 D.n1925 D.n1924 0.127
R2354 D.n1746 D.n1745 0.127
R2355 D.n1587 D.n1586 0.127
R2356 D.n1453 D.n1452 0.127
R2357 D.n1334 D.n1333 0.127
R2358 D.n1240 D.n1239 0.127
R2359 D.n1161 D.n1160 0.127
R2360 D.n1088 D.n1076 0.118
R2361 D.n1089 D.n1042 0.117
R2362 D.n1910 D.n1898 0.113
R2363 D.n1731 D.n1720 0.113
R2364 D.n1576 D.n1565 0.113
R2365 D.n1438 D.n1427 0.113
R2366 D.n1323 D.n1312 0.113
R2367 D.n1225 D.n1214 0.113
R2368 D.n1153 D.n1143 0.113
R2369 D.n1094 D.n422 0.112
R2370 D.n1093 D.n602 0.112
R2371 D.n1092 D.n754 0.112
R2372 D.n1091 D.n878 0.112
R2373 D.n1090 D.n974 0.112
R2374 D.n1915 D.n1914 0.096
R2375 D.n416 D.n415 0.092
R2376 D.n191 D.n190 0.092
R2377 D.n209 D.n206 0.091
R2378 D.n1095 D.n211 0.085
R2379 D.n1112 D.n1111 0.083
R2380 D.n1740 D.n1739 0.081
R2381 D.n1447 D.n1446 0.081
R2382 D.n1234 D.n1233 0.081
R2383 D.n1087 D.n1086 0.079
R2384 D.n227 D.n215 0.078
R2385 D.n438 D.n426 0.078
R2386 D.n618 D.n606 0.078
R2387 D.n770 D.n758 0.078
R2388 D.n894 D.n882 0.078
R2389 D.n990 D.n978 0.078
R2390 D.n1742 D.n1741 0.076
R2391 D.n1449 D.n1448 0.076
R2392 D.n1236 D.n1235 0.076
R2393 D.n184 D.n183 0.075
R2394 D.n165 D.n155 0.075
R2395 D.n1750 D.n1749 0.075
R2396 D.n1609 D.n1599 0.075
R2397 D.n1457 D.n1456 0.075
R2398 D.n1356 D.n1346 0.075
R2399 D.n1244 D.n1243 0.075
R2400 D.n1183 D.n1173 0.075
R2401 D.n1906 D.n1905 0.073
R2402 D.n1905 D.n1904 0.073
R2403 D.n1727 D.n1726 0.073
R2404 D.n1726 D.n1725 0.073
R2405 D.n1572 D.n1571 0.073
R2406 D.n1571 D.n1570 0.073
R2407 D.n1434 D.n1433 0.073
R2408 D.n1433 D.n1432 0.073
R2409 D.n1319 D.n1318 0.073
R2410 D.n1318 D.n1317 0.073
R2411 D.n1221 D.n1220 0.073
R2412 D.n1220 D.n1219 0.073
R2413 D.n1149 D.n1148 0.073
R2414 D.n1148 D.n1147 0.073
R2415 D.n1619 D.n1609 0.072
R2416 D.n1366 D.n1356 0.072
R2417 D.n1193 D.n1183 0.072
R2418 D.n1897 D.n1748 0.072
R2419 D.n1629 D.n1619 0.072
R2420 D.n1639 D.n1629 0.072
R2421 D.n1649 D.n1639 0.072
R2422 D.n1659 D.n1649 0.072
R2423 D.n1669 D.n1659 0.072
R2424 D.n1679 D.n1669 0.072
R2425 D.n1689 D.n1679 0.072
R2426 D.n1699 D.n1689 0.072
R2427 D.n1709 D.n1699 0.072
R2428 D.n1719 D.n1709 0.072
R2429 D.n1564 D.n1455 0.072
R2430 D.n1376 D.n1366 0.072
R2431 D.n1386 D.n1376 0.072
R2432 D.n1396 D.n1386 0.072
R2433 D.n1406 D.n1396 0.072
R2434 D.n1416 D.n1406 0.072
R2435 D.n1426 D.n1416 0.072
R2436 D.n1311 D.n1242 0.072
R2437 D.n1203 D.n1193 0.072
R2438 D.n1213 D.n1203 0.072
R2439 D.n1066 D.n1065 0.072
R2440 D.n1142 D.n1112 0.072
R2441 D.n11 D.n10 0.066
R2442 D.n191 D.n184 0.064
R2443 D.n211 D.n210 0.061
R2444 D.n209 D.n193 0.06
R2445 D.n205 D.n204 0.058
R2446 D.n1927 D.n1926 0.058
R2447 D.n1076 D.n1075 0.056
R2448 D.n193 D.n191 0.055
R2449 D.n415 D.n414 0.055
R2450 D.n1027 D.n1026 0.055
R2451 D.n1099 D.n1098 0.053
R2452 D.n1143 D.n1142 0.053
R2453 D.n1029 D.n1028 0.053
R2454 D.n1896 D.n1888 0.053
R2455 D.n1563 D.n1555 0.053
R2456 D.n1310 D.n1302 0.053
R2457 D.n1141 D.n1132 0.053
R2458 D.n143 D.n142 0.053
R2459 D.n1898 D.n1897 0.053
R2460 D.n1720 D.n1719 0.053
R2461 D.n1565 D.n1564 0.053
R2462 D.n1427 D.n1426 0.053
R2463 D.n1312 D.n1311 0.053
R2464 D.n1214 D.n1213 0.053
R2465 D.n1596 D.n1589 0.052
R2466 D.n1343 D.n1336 0.052
R2467 D.n1170 D.n1163 0.052
R2468 D.n1060 D.n1058 0.052
R2469 D.n1063 D.n1062 0.052
R2470 D.n1773 D.n1771 0.052
R2471 D.n1776 D.n1775 0.052
R2472 D.n1793 D.n1791 0.052
R2473 D.n1796 D.n1795 0.052
R2474 D.n1813 D.n1811 0.052
R2475 D.n1816 D.n1815 0.052
R2476 D.n1833 D.n1831 0.052
R2477 D.n1836 D.n1835 0.052
R2478 D.n1853 D.n1851 0.052
R2479 D.n1856 D.n1855 0.052
R2480 D.n1873 D.n1871 0.052
R2481 D.n1876 D.n1875 0.052
R2482 D.n1892 D.n1890 0.052
R2483 D.n1895 D.n1894 0.052
R2484 D.n1885 D.n1884 0.052
R2485 D.n1882 D.n1881 0.052
R2486 D.n1866 D.n1865 0.052
R2487 D.n1863 D.n1862 0.052
R2488 D.n1846 D.n1845 0.052
R2489 D.n1843 D.n1842 0.052
R2490 D.n1826 D.n1825 0.052
R2491 D.n1823 D.n1822 0.052
R2492 D.n1806 D.n1805 0.052
R2493 D.n1803 D.n1802 0.052
R2494 D.n1786 D.n1785 0.052
R2495 D.n1783 D.n1782 0.052
R2496 D.n1756 D.n1755 0.052
R2497 D.n1753 D.n1752 0.052
R2498 D.n1614 D.n1612 0.052
R2499 D.n1617 D.n1616 0.052
R2500 D.n1634 D.n1632 0.052
R2501 D.n1637 D.n1636 0.052
R2502 D.n1654 D.n1652 0.052
R2503 D.n1657 D.n1656 0.052
R2504 D.n1674 D.n1672 0.052
R2505 D.n1677 D.n1676 0.052
R2506 D.n1694 D.n1692 0.052
R2507 D.n1697 D.n1696 0.052
R2508 D.n1714 D.n1712 0.052
R2509 D.n1717 D.n1716 0.052
R2510 D.n1706 D.n1705 0.052
R2511 D.n1703 D.n1702 0.052
R2512 D.n1686 D.n1685 0.052
R2513 D.n1683 D.n1682 0.052
R2514 D.n1666 D.n1665 0.052
R2515 D.n1663 D.n1662 0.052
R2516 D.n1646 D.n1645 0.052
R2517 D.n1643 D.n1642 0.052
R2518 D.n1626 D.n1625 0.052
R2519 D.n1623 D.n1622 0.052
R2520 D.n1606 D.n1605 0.052
R2521 D.n1603 D.n1602 0.052
R2522 D.n1480 D.n1478 0.052
R2523 D.n1483 D.n1482 0.052
R2524 D.n1500 D.n1498 0.052
R2525 D.n1503 D.n1502 0.052
R2526 D.n1520 D.n1518 0.052
R2527 D.n1523 D.n1522 0.052
R2528 D.n1540 D.n1538 0.052
R2529 D.n1543 D.n1542 0.052
R2530 D.n1559 D.n1557 0.052
R2531 D.n1562 D.n1561 0.052
R2532 D.n1552 D.n1551 0.052
R2533 D.n1549 D.n1548 0.052
R2534 D.n1533 D.n1532 0.052
R2535 D.n1530 D.n1529 0.052
R2536 D.n1513 D.n1512 0.052
R2537 D.n1510 D.n1509 0.052
R2538 D.n1493 D.n1492 0.052
R2539 D.n1490 D.n1489 0.052
R2540 D.n1463 D.n1462 0.052
R2541 D.n1460 D.n1459 0.052
R2542 D.n1361 D.n1359 0.052
R2543 D.n1364 D.n1363 0.052
R2544 D.n1381 D.n1379 0.052
R2545 D.n1384 D.n1383 0.052
R2546 D.n1401 D.n1399 0.052
R2547 D.n1404 D.n1403 0.052
R2548 D.n1421 D.n1419 0.052
R2549 D.n1424 D.n1423 0.052
R2550 D.n1413 D.n1412 0.052
R2551 D.n1410 D.n1409 0.052
R2552 D.n1393 D.n1392 0.052
R2553 D.n1390 D.n1389 0.052
R2554 D.n1373 D.n1372 0.052
R2555 D.n1370 D.n1369 0.052
R2556 D.n1353 D.n1352 0.052
R2557 D.n1350 D.n1349 0.052
R2558 D.n1267 D.n1265 0.052
R2559 D.n1270 D.n1269 0.052
R2560 D.n1287 D.n1285 0.052
R2561 D.n1290 D.n1289 0.052
R2562 D.n1306 D.n1304 0.052
R2563 D.n1309 D.n1308 0.052
R2564 D.n1299 D.n1298 0.052
R2565 D.n1296 D.n1295 0.052
R2566 D.n1280 D.n1279 0.052
R2567 D.n1277 D.n1276 0.052
R2568 D.n1250 D.n1249 0.052
R2569 D.n1247 D.n1246 0.052
R2570 D.n1188 D.n1186 0.052
R2571 D.n1191 D.n1190 0.052
R2572 D.n1208 D.n1206 0.052
R2573 D.n1211 D.n1210 0.052
R2574 D.n1200 D.n1199 0.052
R2575 D.n1197 D.n1196 0.052
R2576 D.n1180 D.n1179 0.052
R2577 D.n1177 D.n1176 0.052
R2578 D.n15 D.n13 0.052
R2579 D.n18 D.n17 0.052
R2580 D.n35 D.n33 0.052
R2581 D.n38 D.n37 0.052
R2582 D.n55 D.n53 0.052
R2583 D.n58 D.n57 0.052
R2584 D.n75 D.n73 0.052
R2585 D.n78 D.n77 0.052
R2586 D.n95 D.n93 0.052
R2587 D.n98 D.n97 0.052
R2588 D.n115 D.n113 0.052
R2589 D.n118 D.n117 0.052
R2590 D.n135 D.n133 0.052
R2591 D.n138 D.n137 0.052
R2592 D.n174 D.n173 0.052
R2593 D.n171 D.n170 0.052
R2594 D.n149 D.n148 0.052
R2595 D.n146 D.n145 0.052
R2596 D.n128 D.n127 0.052
R2597 D.n125 D.n124 0.052
R2598 D.n108 D.n107 0.052
R2599 D.n105 D.n104 0.052
R2600 D.n88 D.n87 0.052
R2601 D.n85 D.n84 0.052
R2602 D.n68 D.n67 0.052
R2603 D.n65 D.n64 0.052
R2604 D.n48 D.n47 0.052
R2605 D.n45 D.n44 0.052
R2606 D.n28 D.n27 0.052
R2607 D.n25 D.n24 0.052
R2608 D.n6 D.n5 0.052
R2609 D.n3 D.n2 0.052
R2610 D.n231 D.n229 0.052
R2611 D.n234 D.n233 0.052
R2612 D.n399 D.n397 0.052
R2613 D.n402 D.n401 0.052
R2614 D.n385 D.n383 0.052
R2615 D.n388 D.n387 0.052
R2616 D.n371 D.n369 0.052
R2617 D.n374 D.n373 0.052
R2618 D.n357 D.n355 0.052
R2619 D.n360 D.n359 0.052
R2620 D.n343 D.n341 0.052
R2621 D.n346 D.n345 0.052
R2622 D.n329 D.n327 0.052
R2623 D.n332 D.n331 0.052
R2624 D.n315 D.n313 0.052
R2625 D.n318 D.n317 0.052
R2626 D.n301 D.n299 0.052
R2627 D.n304 D.n303 0.052
R2628 D.n287 D.n285 0.052
R2629 D.n290 D.n289 0.052
R2630 D.n273 D.n271 0.052
R2631 D.n276 D.n275 0.052
R2632 D.n259 D.n257 0.052
R2633 D.n262 D.n261 0.052
R2634 D.n245 D.n243 0.052
R2635 D.n248 D.n247 0.052
R2636 D.n219 D.n217 0.052
R2637 D.n222 D.n221 0.052
R2638 D.n442 D.n440 0.052
R2639 D.n445 D.n444 0.052
R2640 D.n582 D.n580 0.052
R2641 D.n585 D.n584 0.052
R2642 D.n568 D.n566 0.052
R2643 D.n571 D.n570 0.052
R2644 D.n554 D.n552 0.052
R2645 D.n557 D.n556 0.052
R2646 D.n540 D.n538 0.052
R2647 D.n543 D.n542 0.052
R2648 D.n526 D.n524 0.052
R2649 D.n529 D.n528 0.052
R2650 D.n512 D.n510 0.052
R2651 D.n515 D.n514 0.052
R2652 D.n498 D.n496 0.052
R2653 D.n501 D.n500 0.052
R2654 D.n484 D.n482 0.052
R2655 D.n487 D.n486 0.052
R2656 D.n470 D.n468 0.052
R2657 D.n473 D.n472 0.052
R2658 D.n456 D.n454 0.052
R2659 D.n459 D.n458 0.052
R2660 D.n430 D.n428 0.052
R2661 D.n433 D.n432 0.052
R2662 D.n622 D.n620 0.052
R2663 D.n625 D.n624 0.052
R2664 D.n734 D.n732 0.052
R2665 D.n737 D.n736 0.052
R2666 D.n720 D.n718 0.052
R2667 D.n723 D.n722 0.052
R2668 D.n706 D.n704 0.052
R2669 D.n709 D.n708 0.052
R2670 D.n692 D.n690 0.052
R2671 D.n695 D.n694 0.052
R2672 D.n678 D.n676 0.052
R2673 D.n681 D.n680 0.052
R2674 D.n664 D.n662 0.052
R2675 D.n667 D.n666 0.052
R2676 D.n650 D.n648 0.052
R2677 D.n653 D.n652 0.052
R2678 D.n636 D.n634 0.052
R2679 D.n639 D.n638 0.052
R2680 D.n610 D.n608 0.052
R2681 D.n613 D.n612 0.052
R2682 D.n774 D.n772 0.052
R2683 D.n777 D.n776 0.052
R2684 D.n858 D.n856 0.052
R2685 D.n861 D.n860 0.052
R2686 D.n844 D.n842 0.052
R2687 D.n847 D.n846 0.052
R2688 D.n830 D.n828 0.052
R2689 D.n833 D.n832 0.052
R2690 D.n816 D.n814 0.052
R2691 D.n819 D.n818 0.052
R2692 D.n802 D.n800 0.052
R2693 D.n805 D.n804 0.052
R2694 D.n788 D.n786 0.052
R2695 D.n791 D.n790 0.052
R2696 D.n762 D.n760 0.052
R2697 D.n765 D.n764 0.052
R2698 D.n898 D.n896 0.052
R2699 D.n901 D.n900 0.052
R2700 D.n954 D.n952 0.052
R2701 D.n957 D.n956 0.052
R2702 D.n940 D.n938 0.052
R2703 D.n943 D.n942 0.052
R2704 D.n926 D.n924 0.052
R2705 D.n929 D.n928 0.052
R2706 D.n912 D.n910 0.052
R2707 D.n915 D.n914 0.052
R2708 D.n886 D.n884 0.052
R2709 D.n889 D.n888 0.052
R2710 D.n994 D.n992 0.052
R2711 D.n997 D.n996 0.052
R2712 D.n1022 D.n1020 0.052
R2713 D.n1025 D.n1024 0.052
R2714 D.n1008 D.n1006 0.052
R2715 D.n1011 D.n1010 0.052
R2716 D.n982 D.n980 0.052
R2717 D.n985 D.n984 0.052
R2718 D.n1072 D.n1071 0.052
R2719 D.n1069 D.n1068 0.052
R2720 D.n1119 D.n1118 0.052
R2721 D.n1116 D.n1115 0.052
R2722 D.n1137 D.n1136 0.052
R2723 D.n1140 D.n1138 0.052
R2724 D.n206 D.n205 0.052
R2725 D.n1131 D.n1122 0.051
R2726 D.n1082 D.n1080 0.051
R2727 D.n1106 D.n1105 0.051
R2728 D.n1768 D.n1759 0.051
R2729 D.n1593 D.n1590 0.051
R2730 D.n1475 D.n1466 0.051
R2731 D.n1340 D.n1337 0.051
R2732 D.n1262 D.n1253 0.051
R2733 D.n1167 D.n1164 0.051
R2734 D.n421 D.n413 0.051
R2735 D.n601 D.n596 0.051
R2736 D.n753 D.n748 0.051
R2737 D.n877 D.n872 0.051
R2738 D.n973 D.n968 0.051
R2739 D.n1041 D.n1038 0.051
R2740 D.n1051 D.n1045 0.051
R2741 D.n1049 D.n1048 0.051
R2742 D.n186 D.n185 0.051
R2743 D.n187 D.n186 0.051
R2744 D.n188 D.n187 0.051
R2745 D.n189 D.n188 0.051
R2746 D.n190 D.n189 0.051
R2747 D.n417 D.n416 0.051
R2748 D.n193 D.n192 0.049
R2749 D.n21 D.n11 0.049
R2750 D.n1779 D.n1769 0.049
R2751 D.n1888 D.n1879 0.049
R2752 D.n1879 D.n1869 0.049
R2753 D.n1869 D.n1859 0.049
R2754 D.n1859 D.n1849 0.049
R2755 D.n1849 D.n1839 0.049
R2756 D.n1839 D.n1829 0.049
R2757 D.n1829 D.n1819 0.049
R2758 D.n1819 D.n1809 0.049
R2759 D.n1809 D.n1799 0.049
R2760 D.n1799 D.n1789 0.049
R2761 D.n1789 D.n1779 0.049
R2762 D.n1486 D.n1476 0.049
R2763 D.n1555 D.n1546 0.049
R2764 D.n1546 D.n1536 0.049
R2765 D.n1536 D.n1526 0.049
R2766 D.n1526 D.n1516 0.049
R2767 D.n1516 D.n1506 0.049
R2768 D.n1506 D.n1496 0.049
R2769 D.n1496 D.n1486 0.049
R2770 D.n1273 D.n1263 0.049
R2771 D.n1302 D.n1293 0.049
R2772 D.n1293 D.n1283 0.049
R2773 D.n1283 D.n1273 0.049
R2774 D.n180 D.n152 0.049
R2775 D.n152 D.n141 0.049
R2776 D.n141 D.n131 0.049
R2777 D.n131 D.n121 0.049
R2778 D.n121 D.n111 0.049
R2779 D.n111 D.n101 0.049
R2780 D.n101 D.n91 0.049
R2781 D.n91 D.n81 0.049
R2782 D.n81 D.n71 0.049
R2783 D.n71 D.n61 0.049
R2784 D.n61 D.n51 0.049
R2785 D.n51 D.n41 0.049
R2786 D.n41 D.n31 0.049
R2787 D.n31 D.n21 0.049
R2788 D.n409 D.n395 0.049
R2789 D.n395 D.n381 0.049
R2790 D.n381 D.n367 0.049
R2791 D.n367 D.n353 0.049
R2792 D.n353 D.n339 0.049
R2793 D.n339 D.n325 0.049
R2794 D.n325 D.n311 0.049
R2795 D.n311 D.n297 0.049
R2796 D.n297 D.n283 0.049
R2797 D.n283 D.n269 0.049
R2798 D.n269 D.n255 0.049
R2799 D.n255 D.n241 0.049
R2800 D.n241 D.n227 0.049
R2801 D.n592 D.n578 0.049
R2802 D.n578 D.n564 0.049
R2803 D.n564 D.n550 0.049
R2804 D.n550 D.n536 0.049
R2805 D.n536 D.n522 0.049
R2806 D.n522 D.n508 0.049
R2807 D.n508 D.n494 0.049
R2808 D.n494 D.n480 0.049
R2809 D.n480 D.n466 0.049
R2810 D.n466 D.n452 0.049
R2811 D.n452 D.n438 0.049
R2812 D.n744 D.n730 0.049
R2813 D.n730 D.n716 0.049
R2814 D.n716 D.n702 0.049
R2815 D.n702 D.n688 0.049
R2816 D.n688 D.n674 0.049
R2817 D.n674 D.n660 0.049
R2818 D.n660 D.n646 0.049
R2819 D.n646 D.n632 0.049
R2820 D.n632 D.n618 0.049
R2821 D.n868 D.n854 0.049
R2822 D.n854 D.n840 0.049
R2823 D.n840 D.n826 0.049
R2824 D.n826 D.n812 0.049
R2825 D.n812 D.n798 0.049
R2826 D.n798 D.n784 0.049
R2827 D.n784 D.n770 0.049
R2828 D.n964 D.n950 0.049
R2829 D.n950 D.n936 0.049
R2830 D.n936 D.n922 0.049
R2831 D.n922 D.n908 0.049
R2832 D.n908 D.n894 0.049
R2833 D.n1042 D.n1034 0.049
R2834 D.n1034 D.n1018 0.049
R2835 D.n1018 D.n1004 0.049
R2836 D.n1004 D.n990 0.049
R2837 D.n199 D.n198 0.049
R2838 D.n422 D.n409 0.046
R2839 D.n602 D.n592 0.046
R2840 D.n754 D.n744 0.046
R2841 D.n878 D.n868 0.046
R2842 D.n974 D.n964 0.046
R2843 D.n1900 D.n1899 0.045
R2844 D.n1722 D.n1721 0.045
R2845 D.n1567 D.n1566 0.045
R2846 D.n1429 D.n1428 0.045
R2847 D.n1314 D.n1313 0.045
R2848 D.n1216 D.n1215 0.045
R2849 D.n1145 D.n1144 0.045
R2850 D D.n1095 0.044
R2851 D.n210 D.n180 0.044
R2852 D.n1921 D.n1920 0.043
R2853 D.n1583 D.n1582 0.043
R2854 D.n1330 D.n1329 0.043
R2855 D.n205 D.n202 0.043
R2856 D.n240 D.n239 0.042
R2857 D.n254 D.n253 0.042
R2858 D.n268 D.n267 0.042
R2859 D.n282 D.n281 0.042
R2860 D.n296 D.n295 0.042
R2861 D.n310 D.n309 0.042
R2862 D.n324 D.n323 0.042
R2863 D.n338 D.n337 0.042
R2864 D.n352 D.n351 0.042
R2865 D.n366 D.n365 0.042
R2866 D.n380 D.n379 0.042
R2867 D.n394 D.n393 0.042
R2868 D.n408 D.n407 0.042
R2869 D.n451 D.n450 0.042
R2870 D.n465 D.n464 0.042
R2871 D.n479 D.n478 0.042
R2872 D.n493 D.n492 0.042
R2873 D.n507 D.n506 0.042
R2874 D.n521 D.n520 0.042
R2875 D.n535 D.n534 0.042
R2876 D.n549 D.n548 0.042
R2877 D.n563 D.n562 0.042
R2878 D.n577 D.n576 0.042
R2879 D.n591 D.n590 0.042
R2880 D.n631 D.n630 0.042
R2881 D.n645 D.n644 0.042
R2882 D.n659 D.n658 0.042
R2883 D.n673 D.n672 0.042
R2884 D.n687 D.n686 0.042
R2885 D.n701 D.n700 0.042
R2886 D.n715 D.n714 0.042
R2887 D.n729 D.n728 0.042
R2888 D.n743 D.n742 0.042
R2889 D.n783 D.n782 0.042
R2890 D.n797 D.n796 0.042
R2891 D.n811 D.n810 0.042
R2892 D.n825 D.n824 0.042
R2893 D.n839 D.n838 0.042
R2894 D.n853 D.n852 0.042
R2895 D.n867 D.n866 0.042
R2896 D.n907 D.n906 0.042
R2897 D.n921 D.n920 0.042
R2898 D.n935 D.n934 0.042
R2899 D.n949 D.n948 0.042
R2900 D.n963 D.n962 0.042
R2901 D.n1003 D.n1002 0.042
R2902 D.n1017 D.n1016 0.042
R2903 D.n1033 D.n1032 0.042
R2904 D.n1921 D.n1917 0.041
R2905 D.n1904 D.n1903 0.041
R2906 D.n1725 D.n1724 0.041
R2907 D.n1570 D.n1569 0.041
R2908 D.n1432 D.n1431 0.041
R2909 D.n1317 D.n1316 0.041
R2910 D.n1219 D.n1218 0.041
R2911 D.n1132 D.n1131 0.04
R2912 D.n1909 D.n1908 0.039
R2913 D.n1744 D.n1742 0.039
R2914 D.n1730 D.n1729 0.039
R2915 D.n1575 D.n1574 0.039
R2916 D.n1451 D.n1449 0.039
R2917 D.n1437 D.n1436 0.039
R2918 D.n1322 D.n1321 0.039
R2919 D.n1238 D.n1236 0.039
R2920 D.n1224 D.n1223 0.039
R2921 D.n1152 D.n1151 0.039
R2922 D.n179 D.n177 0.039
R2923 D.n179 D.n167 0.039
R2924 D.n1769 D.n1768 0.038
R2925 D.n1476 D.n1475 0.038
R2926 D.n1263 D.n1262 0.038
R2927 D.n1768 D.n1767 0.036
R2928 D.n1594 D.n1593 0.036
R2929 D.n1475 D.n1474 0.036
R2930 D.n1341 D.n1340 0.036
R2931 D.n1262 D.n1261 0.036
R2932 D.n1168 D.n1167 0.036
R2933 D.n1131 D.n1130 0.036
R2934 D.n1923 D.n1922 0.035
R2935 D.n1585 D.n1584 0.035
R2936 D.n1332 D.n1331 0.035
R2937 D.n1159 D.n1158 0.035
R2938 D.n1108 D.n1107 0.035
R2939 D.n1159 D.n1156 0.034
R2940 D.n1108 D.n1102 0.034
R2941 D.n1923 D.n1913 0.034
R2942 D.n1744 D.n1734 0.034
R2943 D.n1739 D.n1738 0.034
R2944 D.n1585 D.n1579 0.034
R2945 D.n1451 D.n1441 0.034
R2946 D.n1446 D.n1445 0.034
R2947 D.n1332 D.n1326 0.034
R2948 D.n1238 D.n1228 0.034
R2949 D.n1233 D.n1232 0.034
R2950 D.n215 D.n214 0.034
R2951 D.n426 D.n425 0.034
R2952 D.n606 D.n605 0.034
R2953 D.n758 D.n757 0.034
R2954 D.n882 D.n881 0.034
R2955 D.n978 D.n977 0.034
R2956 D.n1055 D.n1054 0.034
R2957 D.n1086 D.n1085 0.034
R2958 D.n1925 D.n1746 0.032
R2959 D.n1746 D.n1587 0.032
R2960 D.n1587 D.n1453 0.032
R2961 D.n1453 D.n1334 0.032
R2962 D.n1334 D.n1240 0.032
R2963 D.n1240 D.n1161 0.032
R2964 D D.n1927 0.032
R2965 D.n1927 D.n1925 0.032
R2966 D.n1089 D.n1088 0.031
R2967 D.n1090 D.n1089 0.031
R2968 D.n1091 D.n1090 0.031
R2969 D.n1092 D.n1091 0.031
R2970 D.n1093 D.n1092 0.031
R2971 D.n1094 D.n1093 0.031
R2972 D.n1095 D.n1094 0.031
R2973 D.n166 D.n154 0.029
R2974 D.n1599 D.n1598 0.029
R2975 D.n1346 D.n1345 0.029
R2976 D.n1173 D.n1172 0.029
R2977 D.n164 D.n163 0.028
R2978 D.n1108 D.n1099 0.027
R2979 D.n1766 D.n1765 0.027
R2980 D.n1923 D.n1910 0.027
R2981 D.n1744 D.n1731 0.027
R2982 D.n1473 D.n1472 0.027
R2983 D.n1585 D.n1576 0.027
R2984 D.n1451 D.n1438 0.027
R2985 D.n1260 D.n1259 0.027
R2986 D.n1332 D.n1323 0.027
R2987 D.n1238 D.n1225 0.027
R2988 D.n1159 D.n1153 0.027
R2989 D.n179 D.n168 0.027
R2990 D.n1129 D.n1128 0.027
R2991 D.n164 D.n159 0.027
R2992 D.n199 D.n197 0.026
R2993 D.n184 D.n181 0.026
R2994 D.n1765 D.n1764 0.025
R2995 D.n1598 D.n1597 0.025
R2996 D.n1472 D.n1471 0.025
R2997 D.n1345 D.n1344 0.025
R2998 D.n1259 D.n1258 0.025
R2999 D.n1172 D.n1171 0.025
R3000 D.n1128 D.n1127 0.025
R3001 D.n408 D.n404 0.025
R3002 D.n394 D.n390 0.025
R3003 D.n380 D.n376 0.025
R3004 D.n366 D.n362 0.025
R3005 D.n352 D.n348 0.025
R3006 D.n338 D.n334 0.025
R3007 D.n324 D.n320 0.025
R3008 D.n310 D.n306 0.025
R3009 D.n296 D.n292 0.025
R3010 D.n282 D.n278 0.025
R3011 D.n268 D.n264 0.025
R3012 D.n254 D.n250 0.025
R3013 D.n240 D.n236 0.025
R3014 D.n226 D.n224 0.025
R3015 D.n591 D.n587 0.025
R3016 D.n577 D.n573 0.025
R3017 D.n563 D.n559 0.025
R3018 D.n549 D.n545 0.025
R3019 D.n535 D.n531 0.025
R3020 D.n521 D.n517 0.025
R3021 D.n507 D.n503 0.025
R3022 D.n493 D.n489 0.025
R3023 D.n479 D.n475 0.025
R3024 D.n465 D.n461 0.025
R3025 D.n451 D.n447 0.025
R3026 D.n437 D.n435 0.025
R3027 D.n743 D.n739 0.025
R3028 D.n729 D.n725 0.025
R3029 D.n715 D.n711 0.025
R3030 D.n701 D.n697 0.025
R3031 D.n687 D.n683 0.025
R3032 D.n673 D.n669 0.025
R3033 D.n659 D.n655 0.025
R3034 D.n645 D.n641 0.025
R3035 D.n631 D.n627 0.025
R3036 D.n617 D.n615 0.025
R3037 D.n867 D.n863 0.025
R3038 D.n853 D.n849 0.025
R3039 D.n839 D.n835 0.025
R3040 D.n825 D.n821 0.025
R3041 D.n811 D.n807 0.025
R3042 D.n797 D.n793 0.025
R3043 D.n783 D.n779 0.025
R3044 D.n769 D.n767 0.025
R3045 D.n963 D.n959 0.025
R3046 D.n949 D.n945 0.025
R3047 D.n935 D.n931 0.025
R3048 D.n921 D.n917 0.025
R3049 D.n907 D.n903 0.025
R3050 D.n893 D.n891 0.025
R3051 D.n1033 D.n1029 0.025
R3052 D.n1017 D.n1013 0.025
R3053 D.n1003 D.n999 0.025
R3054 D.n989 D.n987 0.025
R3055 D.n167 D.n166 0.023
R3056 D.n1908 D.n1907 0.023
R3057 D.n1906 D.n1900 0.023
R3058 D.n1740 D.n1736 0.023
R3059 D.n1729 D.n1728 0.023
R3060 D.n1727 D.n1722 0.023
R3061 D.n1574 D.n1573 0.023
R3062 D.n1572 D.n1567 0.023
R3063 D.n1447 D.n1443 0.023
R3064 D.n1436 D.n1435 0.023
R3065 D.n1434 D.n1429 0.023
R3066 D.n1321 D.n1320 0.023
R3067 D.n1319 D.n1314 0.023
R3068 D.n1234 D.n1230 0.023
R3069 D.n1223 D.n1222 0.023
R3070 D.n1221 D.n1216 0.023
R3071 D.n1151 D.n1150 0.023
R3072 D.n1149 D.n1145 0.023
R3073 D.n421 D.n420 0.023
R3074 D.n240 D.n238 0.023
R3075 D.n254 D.n252 0.023
R3076 D.n268 D.n266 0.023
R3077 D.n282 D.n280 0.023
R3078 D.n296 D.n294 0.023
R3079 D.n310 D.n308 0.023
R3080 D.n324 D.n322 0.023
R3081 D.n338 D.n336 0.023
R3082 D.n352 D.n350 0.023
R3083 D.n366 D.n364 0.023
R3084 D.n380 D.n378 0.023
R3085 D.n394 D.n392 0.023
R3086 D.n408 D.n406 0.023
R3087 D.n601 D.n600 0.023
R3088 D.n451 D.n449 0.023
R3089 D.n465 D.n463 0.023
R3090 D.n479 D.n477 0.023
R3091 D.n493 D.n491 0.023
R3092 D.n507 D.n505 0.023
R3093 D.n521 D.n519 0.023
R3094 D.n535 D.n533 0.023
R3095 D.n549 D.n547 0.023
R3096 D.n563 D.n561 0.023
R3097 D.n577 D.n575 0.023
R3098 D.n591 D.n589 0.023
R3099 D.n753 D.n752 0.023
R3100 D.n631 D.n629 0.023
R3101 D.n645 D.n643 0.023
R3102 D.n659 D.n657 0.023
R3103 D.n673 D.n671 0.023
R3104 D.n687 D.n685 0.023
R3105 D.n701 D.n699 0.023
R3106 D.n715 D.n713 0.023
R3107 D.n729 D.n727 0.023
R3108 D.n743 D.n741 0.023
R3109 D.n877 D.n876 0.023
R3110 D.n783 D.n781 0.023
R3111 D.n797 D.n795 0.023
R3112 D.n811 D.n809 0.023
R3113 D.n825 D.n823 0.023
R3114 D.n839 D.n837 0.023
R3115 D.n853 D.n851 0.023
R3116 D.n867 D.n865 0.023
R3117 D.n973 D.n972 0.023
R3118 D.n907 D.n905 0.023
R3119 D.n921 D.n919 0.023
R3120 D.n935 D.n933 0.023
R3121 D.n949 D.n947 0.023
R3122 D.n963 D.n961 0.023
R3123 D.n1003 D.n1001 0.023
R3124 D.n1017 D.n1015 0.023
R3125 D.n1033 D.n1031 0.023
R3126 D.n1599 D.n1596 0.02
R3127 D.n1346 D.n1343 0.02
R3128 D.n1173 D.n1170 0.02
R3129 D.n201 D.n200 0.019
R3130 D.n421 D.n410 0.019
R3131 D.n601 D.n593 0.019
R3132 D.n753 D.n745 0.019
R3133 D.n877 D.n869 0.019
R3134 D.n973 D.n965 0.019
R3135 D.n161 D.n160 0.016
R3136 D.n1082 D.n1081 0.016
R3137 D.n1074 D.n1073 0.016
R3138 D.n408 D.n396 0.016
R3139 D.n394 D.n382 0.016
R3140 D.n380 D.n368 0.016
R3141 D.n366 D.n354 0.016
R3142 D.n352 D.n340 0.016
R3143 D.n338 D.n326 0.016
R3144 D.n324 D.n312 0.016
R3145 D.n310 D.n298 0.016
R3146 D.n296 D.n284 0.016
R3147 D.n282 D.n270 0.016
R3148 D.n268 D.n256 0.016
R3149 D.n254 D.n242 0.016
R3150 D.n591 D.n579 0.016
R3151 D.n577 D.n565 0.016
R3152 D.n563 D.n551 0.016
R3153 D.n549 D.n537 0.016
R3154 D.n535 D.n523 0.016
R3155 D.n521 D.n509 0.016
R3156 D.n507 D.n495 0.016
R3157 D.n493 D.n481 0.016
R3158 D.n479 D.n467 0.016
R3159 D.n465 D.n453 0.016
R3160 D.n743 D.n731 0.016
R3161 D.n729 D.n717 0.016
R3162 D.n715 D.n703 0.016
R3163 D.n701 D.n689 0.016
R3164 D.n687 D.n675 0.016
R3165 D.n673 D.n661 0.016
R3166 D.n659 D.n647 0.016
R3167 D.n645 D.n633 0.016
R3168 D.n867 D.n855 0.016
R3169 D.n853 D.n841 0.016
R3170 D.n839 D.n827 0.016
R3171 D.n825 D.n813 0.016
R3172 D.n811 D.n799 0.016
R3173 D.n797 D.n785 0.016
R3174 D.n963 D.n951 0.016
R3175 D.n949 D.n937 0.016
R3176 D.n935 D.n923 0.016
R3177 D.n921 D.n909 0.016
R3178 D.n1033 D.n1019 0.016
R3179 D.n1017 D.n1005 0.016
R3180 D.n1064 D.n1057 0.016
R3181 D.n1887 D.n1886 0.016
R3182 D.n1868 D.n1867 0.016
R3183 D.n1848 D.n1847 0.016
R3184 D.n1828 D.n1827 0.016
R3185 D.n1808 D.n1807 0.016
R3186 D.n1788 D.n1787 0.016
R3187 D.n1708 D.n1707 0.016
R3188 D.n1688 D.n1687 0.016
R3189 D.n1668 D.n1667 0.016
R3190 D.n1648 D.n1647 0.016
R3191 D.n1628 D.n1627 0.016
R3192 D.n1554 D.n1553 0.016
R3193 D.n1535 D.n1534 0.016
R3194 D.n1515 D.n1514 0.016
R3195 D.n1495 D.n1494 0.016
R3196 D.n1415 D.n1414 0.016
R3197 D.n1395 D.n1394 0.016
R3198 D.n1375 D.n1374 0.016
R3199 D.n1301 D.n1300 0.016
R3200 D.n1282 D.n1281 0.016
R3201 D.n1202 D.n1201 0.016
R3202 D.n151 D.n150 0.016
R3203 D.n130 D.n129 0.016
R3204 D.n110 D.n109 0.016
R3205 D.n90 D.n89 0.016
R3206 D.n70 D.n69 0.016
R3207 D.n50 D.n49 0.016
R3208 D.n30 D.n29 0.016
R3209 D.n226 D.n216 0.016
R3210 D.n437 D.n427 0.016
R3211 D.n617 D.n607 0.016
R3212 D.n769 D.n759 0.016
R3213 D.n893 D.n883 0.016
R3214 D.n989 D.n979 0.016
R3215 D.n421 D.n418 0.016
R3216 D.n601 D.n598 0.016
R3217 D.n753 D.n750 0.016
R3218 D.n877 D.n874 0.016
R3219 D.n973 D.n970 0.016
R3220 D.n1041 D.n1040 0.016
R3221 D.n1051 D.n1044 0.016
R3222 D.n1051 D.n1050 0.016
R3223 D.n1082 D.n1077 0.016
R3224 D.n8 D.n7 0.015
R3225 D.n1121 D.n1120 0.015
R3226 D.n197 D.n196 0.013
R3227 D.n165 D.n164 0.013
R3228 D.n238 D.n237 0.013
R3229 D.n252 D.n251 0.013
R3230 D.n266 D.n265 0.013
R3231 D.n280 D.n279 0.013
R3232 D.n294 D.n293 0.013
R3233 D.n308 D.n307 0.013
R3234 D.n322 D.n321 0.013
R3235 D.n336 D.n335 0.013
R3236 D.n350 D.n349 0.013
R3237 D.n364 D.n363 0.013
R3238 D.n378 D.n377 0.013
R3239 D.n392 D.n391 0.013
R3240 D.n406 D.n405 0.013
R3241 D.n420 D.n419 0.013
R3242 D.n449 D.n448 0.013
R3243 D.n463 D.n462 0.013
R3244 D.n477 D.n476 0.013
R3245 D.n491 D.n490 0.013
R3246 D.n505 D.n504 0.013
R3247 D.n519 D.n518 0.013
R3248 D.n533 D.n532 0.013
R3249 D.n547 D.n546 0.013
R3250 D.n561 D.n560 0.013
R3251 D.n575 D.n574 0.013
R3252 D.n589 D.n588 0.013
R3253 D.n600 D.n599 0.013
R3254 D.n629 D.n628 0.013
R3255 D.n643 D.n642 0.013
R3256 D.n657 D.n656 0.013
R3257 D.n671 D.n670 0.013
R3258 D.n685 D.n684 0.013
R3259 D.n699 D.n698 0.013
R3260 D.n713 D.n712 0.013
R3261 D.n727 D.n726 0.013
R3262 D.n741 D.n740 0.013
R3263 D.n752 D.n751 0.013
R3264 D.n781 D.n780 0.013
R3265 D.n795 D.n794 0.013
R3266 D.n809 D.n808 0.013
R3267 D.n823 D.n822 0.013
R3268 D.n837 D.n836 0.013
R3269 D.n851 D.n850 0.013
R3270 D.n865 D.n864 0.013
R3271 D.n876 D.n875 0.013
R3272 D.n905 D.n904 0.013
R3273 D.n919 D.n918 0.013
R3274 D.n933 D.n932 0.013
R3275 D.n947 D.n946 0.013
R3276 D.n961 D.n960 0.013
R3277 D.n972 D.n971 0.013
R3278 D.n1001 D.n1000 0.013
R3279 D.n1015 D.n1014 0.013
R3280 D.n1031 D.n1030 0.013
R3281 D.n157 D.n156 0.012
R3282 D.n1910 D.n1909 0.012
R3283 D.n1731 D.n1730 0.012
R3284 D.n1576 D.n1575 0.012
R3285 D.n1438 D.n1437 0.012
R3286 D.n1323 D.n1322 0.012
R3287 D.n1225 D.n1224 0.012
R3288 D.n1153 D.n1152 0.012
R3289 D.n8 D.n0 0.011
R3290 D.n1778 D.n1777 0.011
R3291 D.n1788 D.n1780 0.011
R3292 D.n1798 D.n1797 0.011
R3293 D.n1808 D.n1800 0.011
R3294 D.n1818 D.n1817 0.011
R3295 D.n1828 D.n1820 0.011
R3296 D.n1838 D.n1837 0.011
R3297 D.n1848 D.n1840 0.011
R3298 D.n1858 D.n1857 0.011
R3299 D.n1868 D.n1860 0.011
R3300 D.n1878 D.n1877 0.011
R3301 D.n1897 D.n1896 0.011
R3302 D.n1619 D.n1618 0.011
R3303 D.n1629 D.n1628 0.011
R3304 D.n1639 D.n1638 0.011
R3305 D.n1649 D.n1648 0.011
R3306 D.n1659 D.n1658 0.011
R3307 D.n1669 D.n1668 0.011
R3308 D.n1679 D.n1678 0.011
R3309 D.n1689 D.n1688 0.011
R3310 D.n1699 D.n1698 0.011
R3311 D.n1709 D.n1708 0.011
R3312 D.n1719 D.n1718 0.011
R3313 D.n1485 D.n1484 0.011
R3314 D.n1495 D.n1487 0.011
R3315 D.n1505 D.n1504 0.011
R3316 D.n1515 D.n1507 0.011
R3317 D.n1525 D.n1524 0.011
R3318 D.n1535 D.n1527 0.011
R3319 D.n1545 D.n1544 0.011
R3320 D.n1564 D.n1563 0.011
R3321 D.n1366 D.n1365 0.011
R3322 D.n1376 D.n1375 0.011
R3323 D.n1386 D.n1385 0.011
R3324 D.n1396 D.n1395 0.011
R3325 D.n1406 D.n1405 0.011
R3326 D.n1416 D.n1415 0.011
R3327 D.n1426 D.n1425 0.011
R3328 D.n1272 D.n1271 0.011
R3329 D.n1282 D.n1274 0.011
R3330 D.n1292 D.n1291 0.011
R3331 D.n1311 D.n1310 0.011
R3332 D.n1193 D.n1192 0.011
R3333 D.n1203 D.n1202 0.011
R3334 D.n1213 D.n1212 0.011
R3335 D.n20 D.n19 0.011
R3336 D.n30 D.n22 0.011
R3337 D.n40 D.n39 0.011
R3338 D.n50 D.n42 0.011
R3339 D.n60 D.n59 0.011
R3340 D.n70 D.n62 0.011
R3341 D.n80 D.n79 0.011
R3342 D.n90 D.n82 0.011
R3343 D.n100 D.n99 0.011
R3344 D.n110 D.n102 0.011
R3345 D.n120 D.n119 0.011
R3346 D.n130 D.n122 0.011
R3347 D.n140 D.n139 0.011
R3348 D.n151 D.n143 0.011
R3349 D.n1065 D.n1064 0.011
R3350 D.n1041 D.n1035 0.011
R3351 D.n1768 D.n1762 0.011
R3352 D.n1475 D.n1469 0.011
R3353 D.n1262 D.n1256 0.011
R3354 D.n1131 D.n1125 0.011
R3355 D.n183 D.n182 0.01
R3356 D.n1074 D.n1066 0.01
R3357 D.n1142 D.n1141 0.01
R3358 D.n1904 D.n1902 0.01
R3359 D.n226 D.n225 0.01
R3360 D.n437 D.n436 0.01
R3361 D.n617 D.n616 0.01
R3362 D.n769 D.n768 0.01
R3363 D.n893 D.n892 0.01
R3364 D.n989 D.n988 0.01
R3365 D.n1916 D.n1915 0.009
R3366 D.n159 D.n158 0.009
R3367 D.n201 D.n199 0.009
R3368 D.n1758 D.n1757 0.009
R3369 D.n1608 D.n1607 0.009
R3370 D.n1465 D.n1464 0.009
R3371 D.n1355 D.n1354 0.009
R3372 D.n1252 D.n1251 0.009
R3373 D.n1182 D.n1181 0.009
R3374 D.n1919 D.n1918 0.008
R3375 D.n1581 D.n1580 0.008
R3376 D.n1328 D.n1327 0.008
R3377 D.n1758 D.n1750 0.008
R3378 D.n1609 D.n1608 0.008
R3379 D.n1465 D.n1457 0.008
R3380 D.n1356 D.n1355 0.008
R3381 D.n1252 D.n1244 0.008
R3382 D.n1183 D.n1182 0.008
R3383 D.n163 D.n162 0.006
R3384 D.n1741 D.n1740 0.006
R3385 D.n1448 D.n1447 0.006
R3386 D.n1235 D.n1234 0.006
R3387 D.n202 D.n201 0.006
R3388 D.n204 D.n203 0.006
R3389 D.n1896 D.n1889 0.005
R3390 D.n1878 D.n1870 0.005
R3391 D.n1858 D.n1850 0.005
R3392 D.n1838 D.n1830 0.005
R3393 D.n1818 D.n1810 0.005
R3394 D.n1798 D.n1790 0.005
R3395 D.n1778 D.n1770 0.005
R3396 D.n1718 D.n1711 0.005
R3397 D.n1698 D.n1691 0.005
R3398 D.n1678 D.n1671 0.005
R3399 D.n1658 D.n1651 0.005
R3400 D.n1638 D.n1631 0.005
R3401 D.n1618 D.n1611 0.005
R3402 D.n1563 D.n1556 0.005
R3403 D.n1545 D.n1537 0.005
R3404 D.n1525 D.n1517 0.005
R3405 D.n1505 D.n1497 0.005
R3406 D.n1485 D.n1477 0.005
R3407 D.n1425 D.n1418 0.005
R3408 D.n1405 D.n1398 0.005
R3409 D.n1385 D.n1378 0.005
R3410 D.n1365 D.n1358 0.005
R3411 D.n1310 D.n1303 0.005
R3412 D.n1292 D.n1284 0.005
R3413 D.n1272 D.n1264 0.005
R3414 D.n1212 D.n1205 0.005
R3415 D.n1192 D.n1185 0.005
R3416 D.n140 D.n132 0.005
R3417 D.n120 D.n112 0.005
R3418 D.n100 D.n92 0.005
R3419 D.n80 D.n72 0.005
R3420 D.n60 D.n52 0.005
R3421 D.n40 D.n32 0.005
R3422 D.n20 D.n12 0.005
R3423 D.n240 D.n228 0.005
R3424 D.n451 D.n439 0.005
R3425 D.n631 D.n619 0.005
R3426 D.n783 D.n771 0.005
R3427 D.n907 D.n895 0.005
R3428 D.n1003 D.n991 0.005
R3429 D.n1141 D.n1113 0.005
R3430 D.n1905 D.n1901 0.004
R3431 D.n1726 D.n1723 0.004
R3432 D.n1738 D.n1737 0.004
R3433 D.n1571 D.n1568 0.004
R3434 D.n1433 D.n1430 0.004
R3435 D.n1445 D.n1444 0.004
R3436 D.n1318 D.n1315 0.004
R3437 D.n1220 D.n1217 0.004
R3438 D.n1232 D.n1231 0.004
R3439 D.n1148 D.n1146 0.004
R3440 D.n1766 D.n1763 0.004
R3441 D.n1767 D.n1766 0.004
R3442 D.n1596 D.n1595 0.004
R3443 D.n1595 D.n1594 0.004
R3444 D.n1473 D.n1470 0.004
R3445 D.n1474 D.n1473 0.004
R3446 D.n1343 D.n1342 0.004
R3447 D.n1342 D.n1341 0.004
R3448 D.n1260 D.n1257 0.004
R3449 D.n1261 D.n1260 0.004
R3450 D.n1170 D.n1169 0.004
R3451 D.n1169 D.n1168 0.004
R3452 D.n158 D.n157 0.004
R3453 D.n162 D.n161 0.004
R3454 D.n1129 D.n1126 0.004
R3455 D.n1130 D.n1129 0.004
R3456 D.n1155 D.n1154 0.003
R3457 D.n1101 D.n1100 0.003
R3458 D.n1912 D.n1911 0.003
R3459 D.n1733 D.n1732 0.003
R3460 D.n1578 D.n1577 0.003
R3461 D.n1440 D.n1439 0.003
R3462 D.n1325 D.n1324 0.003
R3463 D.n1227 D.n1226 0.003
R3464 D.n213 D.n212 0.003
R3465 D.n424 D.n423 0.003
R3466 D.n604 D.n603 0.003
R3467 D.n756 D.n755 0.003
R3468 D.n880 D.n879 0.003
R3469 D.n976 D.n975 0.003
R3470 D.n1053 D.n1052 0.003
R3471 D.n1084 D.n1083 0.003
R3472 D.n1137 D.n1133 0.003
R3473 D.n1140 D.n1139 0.003
R3474 D.n1124 D.n1123 0.003
R3475 D.n1079 D.n1078 0.003
R3476 D.n1063 D.n1061 0.003
R3477 D.n1060 D.n1059 0.003
R3478 D.n1104 D.n1103 0.003
R3479 D.n1761 D.n1760 0.003
R3480 D.n1776 D.n1774 0.003
R3481 D.n1773 D.n1772 0.003
R3482 D.n1796 D.n1794 0.003
R3483 D.n1793 D.n1792 0.003
R3484 D.n1816 D.n1814 0.003
R3485 D.n1813 D.n1812 0.003
R3486 D.n1836 D.n1834 0.003
R3487 D.n1833 D.n1832 0.003
R3488 D.n1856 D.n1854 0.003
R3489 D.n1853 D.n1852 0.003
R3490 D.n1876 D.n1874 0.003
R3491 D.n1873 D.n1872 0.003
R3492 D.n1895 D.n1893 0.003
R3493 D.n1892 D.n1891 0.003
R3494 D.n1885 D.n1883 0.003
R3495 D.n1882 D.n1880 0.003
R3496 D.n1866 D.n1864 0.003
R3497 D.n1863 D.n1861 0.003
R3498 D.n1846 D.n1844 0.003
R3499 D.n1843 D.n1841 0.003
R3500 D.n1826 D.n1824 0.003
R3501 D.n1823 D.n1821 0.003
R3502 D.n1806 D.n1804 0.003
R3503 D.n1803 D.n1801 0.003
R3504 D.n1786 D.n1784 0.003
R3505 D.n1783 D.n1781 0.003
R3506 D.n1756 D.n1754 0.003
R3507 D.n1753 D.n1751 0.003
R3508 D.n1592 D.n1591 0.003
R3509 D.n1617 D.n1615 0.003
R3510 D.n1614 D.n1613 0.003
R3511 D.n1637 D.n1635 0.003
R3512 D.n1634 D.n1633 0.003
R3513 D.n1657 D.n1655 0.003
R3514 D.n1654 D.n1653 0.003
R3515 D.n1677 D.n1675 0.003
R3516 D.n1674 D.n1673 0.003
R3517 D.n1697 D.n1695 0.003
R3518 D.n1694 D.n1693 0.003
R3519 D.n1717 D.n1715 0.003
R3520 D.n1714 D.n1713 0.003
R3521 D.n1706 D.n1704 0.003
R3522 D.n1703 D.n1701 0.003
R3523 D.n1686 D.n1684 0.003
R3524 D.n1683 D.n1681 0.003
R3525 D.n1666 D.n1664 0.003
R3526 D.n1663 D.n1661 0.003
R3527 D.n1646 D.n1644 0.003
R3528 D.n1643 D.n1641 0.003
R3529 D.n1626 D.n1624 0.003
R3530 D.n1623 D.n1621 0.003
R3531 D.n1606 D.n1604 0.003
R3532 D.n1603 D.n1601 0.003
R3533 D.n1468 D.n1467 0.003
R3534 D.n1483 D.n1481 0.003
R3535 D.n1480 D.n1479 0.003
R3536 D.n1503 D.n1501 0.003
R3537 D.n1500 D.n1499 0.003
R3538 D.n1523 D.n1521 0.003
R3539 D.n1520 D.n1519 0.003
R3540 D.n1543 D.n1541 0.003
R3541 D.n1540 D.n1539 0.003
R3542 D.n1562 D.n1560 0.003
R3543 D.n1559 D.n1558 0.003
R3544 D.n1552 D.n1550 0.003
R3545 D.n1549 D.n1547 0.003
R3546 D.n1533 D.n1531 0.003
R3547 D.n1530 D.n1528 0.003
R3548 D.n1513 D.n1511 0.003
R3549 D.n1510 D.n1508 0.003
R3550 D.n1493 D.n1491 0.003
R3551 D.n1490 D.n1488 0.003
R3552 D.n1463 D.n1461 0.003
R3553 D.n1460 D.n1458 0.003
R3554 D.n1339 D.n1338 0.003
R3555 D.n1364 D.n1362 0.003
R3556 D.n1361 D.n1360 0.003
R3557 D.n1384 D.n1382 0.003
R3558 D.n1381 D.n1380 0.003
R3559 D.n1404 D.n1402 0.003
R3560 D.n1401 D.n1400 0.003
R3561 D.n1424 D.n1422 0.003
R3562 D.n1421 D.n1420 0.003
R3563 D.n1413 D.n1411 0.003
R3564 D.n1410 D.n1408 0.003
R3565 D.n1393 D.n1391 0.003
R3566 D.n1390 D.n1388 0.003
R3567 D.n1373 D.n1371 0.003
R3568 D.n1370 D.n1368 0.003
R3569 D.n1353 D.n1351 0.003
R3570 D.n1350 D.n1348 0.003
R3571 D.n1255 D.n1254 0.003
R3572 D.n1270 D.n1268 0.003
R3573 D.n1267 D.n1266 0.003
R3574 D.n1290 D.n1288 0.003
R3575 D.n1287 D.n1286 0.003
R3576 D.n1309 D.n1307 0.003
R3577 D.n1306 D.n1305 0.003
R3578 D.n1299 D.n1297 0.003
R3579 D.n1296 D.n1294 0.003
R3580 D.n1280 D.n1278 0.003
R3581 D.n1277 D.n1275 0.003
R3582 D.n1250 D.n1248 0.003
R3583 D.n1247 D.n1245 0.003
R3584 D.n1166 D.n1165 0.003
R3585 D.n1191 D.n1189 0.003
R3586 D.n1188 D.n1187 0.003
R3587 D.n1211 D.n1209 0.003
R3588 D.n1208 D.n1207 0.003
R3589 D.n1200 D.n1198 0.003
R3590 D.n1197 D.n1195 0.003
R3591 D.n1180 D.n1178 0.003
R3592 D.n1177 D.n1175 0.003
R3593 D.n18 D.n16 0.003
R3594 D.n15 D.n14 0.003
R3595 D.n38 D.n36 0.003
R3596 D.n35 D.n34 0.003
R3597 D.n58 D.n56 0.003
R3598 D.n55 D.n54 0.003
R3599 D.n78 D.n76 0.003
R3600 D.n75 D.n74 0.003
R3601 D.n98 D.n96 0.003
R3602 D.n95 D.n94 0.003
R3603 D.n118 D.n116 0.003
R3604 D.n115 D.n114 0.003
R3605 D.n138 D.n136 0.003
R3606 D.n135 D.n134 0.003
R3607 D.n174 D.n172 0.003
R3608 D.n171 D.n169 0.003
R3609 D.n149 D.n147 0.003
R3610 D.n146 D.n144 0.003
R3611 D.n128 D.n126 0.003
R3612 D.n125 D.n123 0.003
R3613 D.n108 D.n106 0.003
R3614 D.n105 D.n103 0.003
R3615 D.n88 D.n86 0.003
R3616 D.n85 D.n83 0.003
R3617 D.n68 D.n66 0.003
R3618 D.n65 D.n63 0.003
R3619 D.n48 D.n46 0.003
R3620 D.n45 D.n43 0.003
R3621 D.n28 D.n26 0.003
R3622 D.n25 D.n23 0.003
R3623 D.n6 D.n4 0.003
R3624 D.n3 D.n1 0.003
R3625 D.n234 D.n232 0.003
R3626 D.n231 D.n230 0.003
R3627 D.n412 D.n411 0.003
R3628 D.n402 D.n400 0.003
R3629 D.n399 D.n398 0.003
R3630 D.n388 D.n386 0.003
R3631 D.n385 D.n384 0.003
R3632 D.n374 D.n372 0.003
R3633 D.n371 D.n370 0.003
R3634 D.n360 D.n358 0.003
R3635 D.n357 D.n356 0.003
R3636 D.n346 D.n344 0.003
R3637 D.n343 D.n342 0.003
R3638 D.n332 D.n330 0.003
R3639 D.n329 D.n328 0.003
R3640 D.n318 D.n316 0.003
R3641 D.n315 D.n314 0.003
R3642 D.n304 D.n302 0.003
R3643 D.n301 D.n300 0.003
R3644 D.n290 D.n288 0.003
R3645 D.n287 D.n286 0.003
R3646 D.n276 D.n274 0.003
R3647 D.n273 D.n272 0.003
R3648 D.n262 D.n260 0.003
R3649 D.n259 D.n258 0.003
R3650 D.n248 D.n246 0.003
R3651 D.n245 D.n244 0.003
R3652 D.n222 D.n220 0.003
R3653 D.n219 D.n218 0.003
R3654 D.n445 D.n443 0.003
R3655 D.n442 D.n441 0.003
R3656 D.n595 D.n594 0.003
R3657 D.n585 D.n583 0.003
R3658 D.n582 D.n581 0.003
R3659 D.n571 D.n569 0.003
R3660 D.n568 D.n567 0.003
R3661 D.n557 D.n555 0.003
R3662 D.n554 D.n553 0.003
R3663 D.n543 D.n541 0.003
R3664 D.n540 D.n539 0.003
R3665 D.n529 D.n527 0.003
R3666 D.n526 D.n525 0.003
R3667 D.n515 D.n513 0.003
R3668 D.n512 D.n511 0.003
R3669 D.n501 D.n499 0.003
R3670 D.n498 D.n497 0.003
R3671 D.n487 D.n485 0.003
R3672 D.n484 D.n483 0.003
R3673 D.n473 D.n471 0.003
R3674 D.n470 D.n469 0.003
R3675 D.n459 D.n457 0.003
R3676 D.n456 D.n455 0.003
R3677 D.n433 D.n431 0.003
R3678 D.n430 D.n429 0.003
R3679 D.n625 D.n623 0.003
R3680 D.n622 D.n621 0.003
R3681 D.n747 D.n746 0.003
R3682 D.n737 D.n735 0.003
R3683 D.n734 D.n733 0.003
R3684 D.n723 D.n721 0.003
R3685 D.n720 D.n719 0.003
R3686 D.n709 D.n707 0.003
R3687 D.n706 D.n705 0.003
R3688 D.n695 D.n693 0.003
R3689 D.n692 D.n691 0.003
R3690 D.n681 D.n679 0.003
R3691 D.n678 D.n677 0.003
R3692 D.n667 D.n665 0.003
R3693 D.n664 D.n663 0.003
R3694 D.n653 D.n651 0.003
R3695 D.n650 D.n649 0.003
R3696 D.n639 D.n637 0.003
R3697 D.n636 D.n635 0.003
R3698 D.n613 D.n611 0.003
R3699 D.n610 D.n609 0.003
R3700 D.n777 D.n775 0.003
R3701 D.n774 D.n773 0.003
R3702 D.n871 D.n870 0.003
R3703 D.n861 D.n859 0.003
R3704 D.n858 D.n857 0.003
R3705 D.n847 D.n845 0.003
R3706 D.n844 D.n843 0.003
R3707 D.n833 D.n831 0.003
R3708 D.n830 D.n829 0.003
R3709 D.n819 D.n817 0.003
R3710 D.n816 D.n815 0.003
R3711 D.n805 D.n803 0.003
R3712 D.n802 D.n801 0.003
R3713 D.n791 D.n789 0.003
R3714 D.n788 D.n787 0.003
R3715 D.n765 D.n763 0.003
R3716 D.n762 D.n761 0.003
R3717 D.n901 D.n899 0.003
R3718 D.n898 D.n897 0.003
R3719 D.n967 D.n966 0.003
R3720 D.n957 D.n955 0.003
R3721 D.n954 D.n953 0.003
R3722 D.n943 D.n941 0.003
R3723 D.n940 D.n939 0.003
R3724 D.n929 D.n927 0.003
R3725 D.n926 D.n925 0.003
R3726 D.n915 D.n913 0.003
R3727 D.n912 D.n911 0.003
R3728 D.n889 D.n887 0.003
R3729 D.n886 D.n885 0.003
R3730 D.n997 D.n995 0.003
R3731 D.n994 D.n993 0.003
R3732 D.n1037 D.n1036 0.003
R3733 D.n1025 D.n1023 0.003
R3734 D.n1022 D.n1021 0.003
R3735 D.n1011 D.n1009 0.003
R3736 D.n1008 D.n1007 0.003
R3737 D.n985 D.n983 0.003
R3738 D.n982 D.n981 0.003
R3739 D.n1047 D.n1046 0.003
R3740 D.n1072 D.n1070 0.003
R3741 D.n1069 D.n1067 0.003
R3742 D.n1119 D.n1117 0.003
R3743 D.n1116 D.n1114 0.003
R3744 D.n224 D.n223 0.003
R3745 D.n236 D.n235 0.003
R3746 D.n250 D.n249 0.003
R3747 D.n264 D.n263 0.003
R3748 D.n278 D.n277 0.003
R3749 D.n292 D.n291 0.003
R3750 D.n306 D.n305 0.003
R3751 D.n320 D.n319 0.003
R3752 D.n334 D.n333 0.003
R3753 D.n348 D.n347 0.003
R3754 D.n362 D.n361 0.003
R3755 D.n376 D.n375 0.003
R3756 D.n390 D.n389 0.003
R3757 D.n404 D.n403 0.003
R3758 D.n435 D.n434 0.003
R3759 D.n447 D.n446 0.003
R3760 D.n461 D.n460 0.003
R3761 D.n475 D.n474 0.003
R3762 D.n489 D.n488 0.003
R3763 D.n503 D.n502 0.003
R3764 D.n517 D.n516 0.003
R3765 D.n531 D.n530 0.003
R3766 D.n545 D.n544 0.003
R3767 D.n559 D.n558 0.003
R3768 D.n573 D.n572 0.003
R3769 D.n587 D.n586 0.003
R3770 D.n615 D.n614 0.003
R3771 D.n627 D.n626 0.003
R3772 D.n641 D.n640 0.003
R3773 D.n655 D.n654 0.003
R3774 D.n669 D.n668 0.003
R3775 D.n683 D.n682 0.003
R3776 D.n697 D.n696 0.003
R3777 D.n711 D.n710 0.003
R3778 D.n725 D.n724 0.003
R3779 D.n739 D.n738 0.003
R3780 D.n767 D.n766 0.003
R3781 D.n779 D.n778 0.003
R3782 D.n793 D.n792 0.003
R3783 D.n807 D.n806 0.003
R3784 D.n821 D.n820 0.003
R3785 D.n835 D.n834 0.003
R3786 D.n849 D.n848 0.003
R3787 D.n863 D.n862 0.003
R3788 D.n891 D.n890 0.003
R3789 D.n903 D.n902 0.003
R3790 D.n917 D.n916 0.003
R3791 D.n931 D.n930 0.003
R3792 D.n945 D.n944 0.003
R3793 D.n959 D.n958 0.003
R3794 D.n987 D.n986 0.003
R3795 D.n999 D.n998 0.003
R3796 D.n1013 D.n1012 0.003
R3797 D.n1029 D.n1027 0.003
R3798 D.n1920 D.n1919 0.003
R3799 D.n1582 D.n1581 0.003
R3800 D.n1329 D.n1328 0.003
R3801 D.n1076 D.n1051 0.003
R3802 D.n1718 D.n1710 0.003
R3803 D.n1708 D.n1700 0.003
R3804 D.n1698 D.n1690 0.003
R3805 D.n1688 D.n1680 0.003
R3806 D.n1678 D.n1670 0.003
R3807 D.n1668 D.n1660 0.003
R3808 D.n1658 D.n1650 0.003
R3809 D.n1648 D.n1640 0.003
R3810 D.n1638 D.n1630 0.003
R3811 D.n1628 D.n1620 0.003
R3812 D.n1618 D.n1610 0.003
R3813 D.n1425 D.n1417 0.003
R3814 D.n1415 D.n1407 0.003
R3815 D.n1405 D.n1397 0.003
R3816 D.n1395 D.n1387 0.003
R3817 D.n1385 D.n1377 0.003
R3818 D.n1375 D.n1367 0.003
R3819 D.n1365 D.n1357 0.003
R3820 D.n1212 D.n1204 0.003
R3821 D.n1202 D.n1194 0.003
R3822 D.n1192 D.n1184 0.003
R3823 D.n1608 D.n1600 0.003
R3824 D.n1355 D.n1347 0.003
R3825 D.n1182 D.n1174 0.003
R3826 D.n1064 D.n1056 0.003
R3827 D.n1917 D.n1916 0.002
R3828 D.n1075 D.n1074 0.002
R3829 D.n1924 D.n1923 0.002
R3830 D.n1745 D.n1744 0.002
R3831 D.n1586 D.n1585 0.002
R3832 D.n1452 D.n1451 0.002
R3833 D.n1333 D.n1332 0.002
R3834 D.n1239 D.n1238 0.002
R3835 D.n1160 D.n1159 0.002
R3836 D.n1109 D.n1108 0.002
R3837 D.n1907 D.n1906 0.001
R3838 D.n1728 D.n1727 0.001
R3839 D.n1573 D.n1572 0.001
R3840 D.n1435 D.n1434 0.001
R3841 D.n1320 D.n1319 0.001
R3842 D.n1222 D.n1221 0.001
R3843 D.n1150 D.n1149 0.001
R3844 D.n208 D.n207 0.001
R3845 D.n196 D.n195 0.001
R3846 D.n154 D.n153 0.001
R3847 D.n166 D.n165 0.001
R3848 D.n210 D.n209 0.001
R3849 D.n422 D.n421 0.001
R3850 D.n602 D.n601 0.001
R3851 D.n754 D.n753 0.001
R3852 D.n878 D.n877 0.001
R3853 D.n974 D.n973 0.001
R3854 D.n1087 D.n1082 0.001
R3855 D.n11 D.n8 0.001
R3856 D.n1769 D.n1758 0.001
R3857 D.n1888 D.n1887 0.001
R3858 D.n1879 D.n1878 0.001
R3859 D.n1869 D.n1868 0.001
R3860 D.n1859 D.n1858 0.001
R3861 D.n1849 D.n1848 0.001
R3862 D.n1839 D.n1838 0.001
R3863 D.n1829 D.n1828 0.001
R3864 D.n1819 D.n1818 0.001
R3865 D.n1809 D.n1808 0.001
R3866 D.n1799 D.n1798 0.001
R3867 D.n1789 D.n1788 0.001
R3868 D.n1779 D.n1778 0.001
R3869 D.n1476 D.n1465 0.001
R3870 D.n1555 D.n1554 0.001
R3871 D.n1546 D.n1545 0.001
R3872 D.n1536 D.n1535 0.001
R3873 D.n1526 D.n1525 0.001
R3874 D.n1516 D.n1515 0.001
R3875 D.n1506 D.n1505 0.001
R3876 D.n1496 D.n1495 0.001
R3877 D.n1486 D.n1485 0.001
R3878 D.n1263 D.n1252 0.001
R3879 D.n1302 D.n1301 0.001
R3880 D.n1293 D.n1292 0.001
R3881 D.n1283 D.n1282 0.001
R3882 D.n1273 D.n1272 0.001
R3883 D.n1132 D.n1121 0.001
R3884 D.n180 D.n179 0.001
R3885 D.n152 D.n151 0.001
R3886 D.n141 D.n140 0.001
R3887 D.n131 D.n130 0.001
R3888 D.n121 D.n120 0.001
R3889 D.n111 D.n110 0.001
R3890 D.n101 D.n100 0.001
R3891 D.n91 D.n90 0.001
R3892 D.n81 D.n80 0.001
R3893 D.n71 D.n70 0.001
R3894 D.n61 D.n60 0.001
R3895 D.n51 D.n50 0.001
R3896 D.n41 D.n40 0.001
R3897 D.n31 D.n30 0.001
R3898 D.n21 D.n20 0.001
R3899 D.n409 D.n408 0.001
R3900 D.n395 D.n394 0.001
R3901 D.n381 D.n380 0.001
R3902 D.n367 D.n366 0.001
R3903 D.n353 D.n352 0.001
R3904 D.n339 D.n338 0.001
R3905 D.n325 D.n324 0.001
R3906 D.n311 D.n310 0.001
R3907 D.n297 D.n296 0.001
R3908 D.n283 D.n282 0.001
R3909 D.n269 D.n268 0.001
R3910 D.n255 D.n254 0.001
R3911 D.n241 D.n240 0.001
R3912 D.n227 D.n226 0.001
R3913 D.n592 D.n591 0.001
R3914 D.n578 D.n577 0.001
R3915 D.n564 D.n563 0.001
R3916 D.n550 D.n549 0.001
R3917 D.n536 D.n535 0.001
R3918 D.n522 D.n521 0.001
R3919 D.n508 D.n507 0.001
R3920 D.n494 D.n493 0.001
R3921 D.n480 D.n479 0.001
R3922 D.n466 D.n465 0.001
R3923 D.n452 D.n451 0.001
R3924 D.n438 D.n437 0.001
R3925 D.n744 D.n743 0.001
R3926 D.n730 D.n729 0.001
R3927 D.n716 D.n715 0.001
R3928 D.n702 D.n701 0.001
R3929 D.n688 D.n687 0.001
R3930 D.n674 D.n673 0.001
R3931 D.n660 D.n659 0.001
R3932 D.n646 D.n645 0.001
R3933 D.n632 D.n631 0.001
R3934 D.n618 D.n617 0.001
R3935 D.n868 D.n867 0.001
R3936 D.n854 D.n853 0.001
R3937 D.n840 D.n839 0.001
R3938 D.n826 D.n825 0.001
R3939 D.n812 D.n811 0.001
R3940 D.n798 D.n797 0.001
R3941 D.n784 D.n783 0.001
R3942 D.n770 D.n769 0.001
R3943 D.n964 D.n963 0.001
R3944 D.n950 D.n949 0.001
R3945 D.n936 D.n935 0.001
R3946 D.n922 D.n921 0.001
R3947 D.n908 D.n907 0.001
R3948 D.n894 D.n893 0.001
R3949 D.n1042 D.n1041 0.001
R3950 D.n1034 D.n1033 0.001
R3951 D.n1018 D.n1017 0.001
R3952 D.n1004 D.n1003 0.001
R3953 D.n990 D.n989 0.001
R3954 D.n209 D.n194 0.001
R3955 D.n1131 D.n1124 0.001
R3956 D.n1082 D.n1079 0.001
R3957 D.n1064 D.n1063 0.001
R3958 D.n1064 D.n1060 0.001
R3959 D.n1106 D.n1104 0.001
R3960 D.n1768 D.n1761 0.001
R3961 D.n1778 D.n1776 0.001
R3962 D.n1778 D.n1773 0.001
R3963 D.n1798 D.n1796 0.001
R3964 D.n1798 D.n1793 0.001
R3965 D.n1818 D.n1816 0.001
R3966 D.n1818 D.n1813 0.001
R3967 D.n1838 D.n1836 0.001
R3968 D.n1838 D.n1833 0.001
R3969 D.n1858 D.n1856 0.001
R3970 D.n1858 D.n1853 0.001
R3971 D.n1878 D.n1876 0.001
R3972 D.n1878 D.n1873 0.001
R3973 D.n1896 D.n1895 0.001
R3974 D.n1896 D.n1892 0.001
R3975 D.n1887 D.n1882 0.001
R3976 D.n1887 D.n1885 0.001
R3977 D.n1868 D.n1863 0.001
R3978 D.n1868 D.n1866 0.001
R3979 D.n1848 D.n1843 0.001
R3980 D.n1848 D.n1846 0.001
R3981 D.n1828 D.n1823 0.001
R3982 D.n1828 D.n1826 0.001
R3983 D.n1808 D.n1803 0.001
R3984 D.n1808 D.n1806 0.001
R3985 D.n1788 D.n1783 0.001
R3986 D.n1788 D.n1786 0.001
R3987 D.n1758 D.n1753 0.001
R3988 D.n1758 D.n1756 0.001
R3989 D.n1593 D.n1592 0.001
R3990 D.n1618 D.n1617 0.001
R3991 D.n1618 D.n1614 0.001
R3992 D.n1638 D.n1637 0.001
R3993 D.n1638 D.n1634 0.001
R3994 D.n1658 D.n1657 0.001
R3995 D.n1658 D.n1654 0.001
R3996 D.n1678 D.n1677 0.001
R3997 D.n1678 D.n1674 0.001
R3998 D.n1698 D.n1697 0.001
R3999 D.n1698 D.n1694 0.001
R4000 D.n1718 D.n1717 0.001
R4001 D.n1718 D.n1714 0.001
R4002 D.n1708 D.n1703 0.001
R4003 D.n1708 D.n1706 0.001
R4004 D.n1688 D.n1683 0.001
R4005 D.n1688 D.n1686 0.001
R4006 D.n1668 D.n1663 0.001
R4007 D.n1668 D.n1666 0.001
R4008 D.n1648 D.n1643 0.001
R4009 D.n1648 D.n1646 0.001
R4010 D.n1628 D.n1623 0.001
R4011 D.n1628 D.n1626 0.001
R4012 D.n1608 D.n1603 0.001
R4013 D.n1608 D.n1606 0.001
R4014 D.n1475 D.n1468 0.001
R4015 D.n1485 D.n1483 0.001
R4016 D.n1485 D.n1480 0.001
R4017 D.n1505 D.n1503 0.001
R4018 D.n1505 D.n1500 0.001
R4019 D.n1525 D.n1523 0.001
R4020 D.n1525 D.n1520 0.001
R4021 D.n1545 D.n1543 0.001
R4022 D.n1545 D.n1540 0.001
R4023 D.n1563 D.n1562 0.001
R4024 D.n1563 D.n1559 0.001
R4025 D.n1554 D.n1549 0.001
R4026 D.n1554 D.n1552 0.001
R4027 D.n1535 D.n1530 0.001
R4028 D.n1535 D.n1533 0.001
R4029 D.n1515 D.n1510 0.001
R4030 D.n1515 D.n1513 0.001
R4031 D.n1495 D.n1490 0.001
R4032 D.n1495 D.n1493 0.001
R4033 D.n1465 D.n1460 0.001
R4034 D.n1465 D.n1463 0.001
R4035 D.n1340 D.n1339 0.001
R4036 D.n1365 D.n1364 0.001
R4037 D.n1365 D.n1361 0.001
R4038 D.n1385 D.n1384 0.001
R4039 D.n1385 D.n1381 0.001
R4040 D.n1405 D.n1404 0.001
R4041 D.n1405 D.n1401 0.001
R4042 D.n1425 D.n1424 0.001
R4043 D.n1425 D.n1421 0.001
R4044 D.n1415 D.n1410 0.001
R4045 D.n1415 D.n1413 0.001
R4046 D.n1395 D.n1390 0.001
R4047 D.n1395 D.n1393 0.001
R4048 D.n1375 D.n1370 0.001
R4049 D.n1375 D.n1373 0.001
R4050 D.n1355 D.n1350 0.001
R4051 D.n1355 D.n1353 0.001
R4052 D.n1262 D.n1255 0.001
R4053 D.n1272 D.n1270 0.001
R4054 D.n1272 D.n1267 0.001
R4055 D.n1292 D.n1290 0.001
R4056 D.n1292 D.n1287 0.001
R4057 D.n1310 D.n1309 0.001
R4058 D.n1310 D.n1306 0.001
R4059 D.n1301 D.n1296 0.001
R4060 D.n1301 D.n1299 0.001
R4061 D.n1282 D.n1277 0.001
R4062 D.n1282 D.n1280 0.001
R4063 D.n1252 D.n1247 0.001
R4064 D.n1252 D.n1250 0.001
R4065 D.n1167 D.n1166 0.001
R4066 D.n1192 D.n1191 0.001
R4067 D.n1192 D.n1188 0.001
R4068 D.n1212 D.n1211 0.001
R4069 D.n1212 D.n1208 0.001
R4070 D.n1202 D.n1197 0.001
R4071 D.n1202 D.n1200 0.001
R4072 D.n1182 D.n1177 0.001
R4073 D.n1182 D.n1180 0.001
R4074 D.n10 D.n9 0.001
R4075 D.n20 D.n18 0.001
R4076 D.n20 D.n15 0.001
R4077 D.n40 D.n38 0.001
R4078 D.n40 D.n35 0.001
R4079 D.n60 D.n58 0.001
R4080 D.n60 D.n55 0.001
R4081 D.n80 D.n78 0.001
R4082 D.n80 D.n75 0.001
R4083 D.n100 D.n98 0.001
R4084 D.n100 D.n95 0.001
R4085 D.n120 D.n118 0.001
R4086 D.n120 D.n115 0.001
R4087 D.n140 D.n138 0.001
R4088 D.n140 D.n135 0.001
R4089 D.n179 D.n171 0.001
R4090 D.n179 D.n174 0.001
R4091 D.n151 D.n146 0.001
R4092 D.n151 D.n149 0.001
R4093 D.n130 D.n125 0.001
R4094 D.n130 D.n128 0.001
R4095 D.n110 D.n105 0.001
R4096 D.n110 D.n108 0.001
R4097 D.n90 D.n85 0.001
R4098 D.n90 D.n88 0.001
R4099 D.n70 D.n65 0.001
R4100 D.n70 D.n68 0.001
R4101 D.n50 D.n45 0.001
R4102 D.n50 D.n48 0.001
R4103 D.n30 D.n25 0.001
R4104 D.n30 D.n28 0.001
R4105 D.n8 D.n3 0.001
R4106 D.n8 D.n6 0.001
R4107 D.n240 D.n234 0.001
R4108 D.n240 D.n231 0.001
R4109 D.n421 D.n412 0.001
R4110 D.n408 D.n402 0.001
R4111 D.n408 D.n399 0.001
R4112 D.n394 D.n388 0.001
R4113 D.n394 D.n385 0.001
R4114 D.n380 D.n374 0.001
R4115 D.n380 D.n371 0.001
R4116 D.n366 D.n360 0.001
R4117 D.n366 D.n357 0.001
R4118 D.n352 D.n346 0.001
R4119 D.n352 D.n343 0.001
R4120 D.n338 D.n332 0.001
R4121 D.n338 D.n329 0.001
R4122 D.n324 D.n318 0.001
R4123 D.n324 D.n315 0.001
R4124 D.n310 D.n304 0.001
R4125 D.n310 D.n301 0.001
R4126 D.n296 D.n290 0.001
R4127 D.n296 D.n287 0.001
R4128 D.n282 D.n276 0.001
R4129 D.n282 D.n273 0.001
R4130 D.n268 D.n262 0.001
R4131 D.n268 D.n259 0.001
R4132 D.n254 D.n248 0.001
R4133 D.n254 D.n245 0.001
R4134 D.n226 D.n222 0.001
R4135 D.n226 D.n219 0.001
R4136 D.n451 D.n445 0.001
R4137 D.n451 D.n442 0.001
R4138 D.n601 D.n595 0.001
R4139 D.n591 D.n585 0.001
R4140 D.n591 D.n582 0.001
R4141 D.n577 D.n571 0.001
R4142 D.n577 D.n568 0.001
R4143 D.n563 D.n557 0.001
R4144 D.n563 D.n554 0.001
R4145 D.n549 D.n543 0.001
R4146 D.n549 D.n540 0.001
R4147 D.n535 D.n529 0.001
R4148 D.n535 D.n526 0.001
R4149 D.n521 D.n515 0.001
R4150 D.n521 D.n512 0.001
R4151 D.n507 D.n501 0.001
R4152 D.n507 D.n498 0.001
R4153 D.n493 D.n487 0.001
R4154 D.n493 D.n484 0.001
R4155 D.n479 D.n473 0.001
R4156 D.n479 D.n470 0.001
R4157 D.n465 D.n459 0.001
R4158 D.n465 D.n456 0.001
R4159 D.n437 D.n433 0.001
R4160 D.n437 D.n430 0.001
R4161 D.n631 D.n625 0.001
R4162 D.n631 D.n622 0.001
R4163 D.n753 D.n747 0.001
R4164 D.n743 D.n737 0.001
R4165 D.n743 D.n734 0.001
R4166 D.n729 D.n723 0.001
R4167 D.n729 D.n720 0.001
R4168 D.n715 D.n709 0.001
R4169 D.n715 D.n706 0.001
R4170 D.n701 D.n695 0.001
R4171 D.n701 D.n692 0.001
R4172 D.n687 D.n681 0.001
R4173 D.n687 D.n678 0.001
R4174 D.n673 D.n667 0.001
R4175 D.n673 D.n664 0.001
R4176 D.n659 D.n653 0.001
R4177 D.n659 D.n650 0.001
R4178 D.n645 D.n639 0.001
R4179 D.n645 D.n636 0.001
R4180 D.n617 D.n613 0.001
R4181 D.n617 D.n610 0.001
R4182 D.n783 D.n777 0.001
R4183 D.n783 D.n774 0.001
R4184 D.n877 D.n871 0.001
R4185 D.n867 D.n861 0.001
R4186 D.n867 D.n858 0.001
R4187 D.n853 D.n847 0.001
R4188 D.n853 D.n844 0.001
R4189 D.n839 D.n833 0.001
R4190 D.n839 D.n830 0.001
R4191 D.n825 D.n819 0.001
R4192 D.n825 D.n816 0.001
R4193 D.n811 D.n805 0.001
R4194 D.n811 D.n802 0.001
R4195 D.n797 D.n791 0.001
R4196 D.n797 D.n788 0.001
R4197 D.n769 D.n765 0.001
R4198 D.n769 D.n762 0.001
R4199 D.n907 D.n901 0.001
R4200 D.n907 D.n898 0.001
R4201 D.n973 D.n967 0.001
R4202 D.n963 D.n957 0.001
R4203 D.n963 D.n954 0.001
R4204 D.n949 D.n943 0.001
R4205 D.n949 D.n940 0.001
R4206 D.n935 D.n929 0.001
R4207 D.n935 D.n926 0.001
R4208 D.n921 D.n915 0.001
R4209 D.n921 D.n912 0.001
R4210 D.n893 D.n889 0.001
R4211 D.n893 D.n886 0.001
R4212 D.n1003 D.n997 0.001
R4213 D.n1003 D.n994 0.001
R4214 D.n1041 D.n1037 0.001
R4215 D.n1033 D.n1025 0.001
R4216 D.n1033 D.n1022 0.001
R4217 D.n1017 D.n1011 0.001
R4218 D.n1017 D.n1008 0.001
R4219 D.n989 D.n985 0.001
R4220 D.n989 D.n982 0.001
R4221 D.n1051 D.n1047 0.001
R4222 D.n1074 D.n1069 0.001
R4223 D.n1074 D.n1072 0.001
R4224 D.n1121 D.n1116 0.001
R4225 D.n1121 D.n1119 0.001
R4226 D.n1141 D.n1137 0.001
R4227 D.n1141 D.n1140 0.001
R4228 D.n1159 D.n1155 0.001
R4229 D.n1108 D.n1101 0.001
R4230 D.n1923 D.n1912 0.001
R4231 D.n1744 D.n1733 0.001
R4232 D.n1585 D.n1578 0.001
R4233 D.n1451 D.n1440 0.001
R4234 D.n1332 D.n1325 0.001
R4235 D.n1238 D.n1227 0.001
R4236 D.n215 D.n213 0.001
R4237 D.n426 D.n424 0.001
R4238 D.n606 D.n604 0.001
R4239 D.n758 D.n756 0.001
R4240 D.n882 D.n880 0.001
R4241 D.n978 D.n976 0.001
R4242 D.n1055 D.n1053 0.001
R4243 D.n1086 D.n1084 0.001
C0 DNW S 1825.11fF
C1 DNW G 4.69fF
C2 DNW D 274.03fF
C3 S G 826.28fF
C4 S D 1281.65fF
C5 G D 582.15fF
C6 D VSUBS -23.80fF $ **FLOATING
C7 G VSUBS -70.07fF
C8 S VSUBS 171.22fF $ **FLOATING
C9 DNW VSUBS 5160.69fF $ **FLOATING
C10 D.n0 VSUBS 2.16fF $ **FLOATING
C11 D.t122 VSUBS -0.02fF
C12 D.n1 VSUBS 0.20fF $ **FLOATING
C13 D.t571 VSUBS -0.06fF
C14 D.n2 VSUBS 0.61fF $ **FLOATING
C15 D.t296 VSUBS -0.02fF
C16 D.n4 VSUBS 0.20fF $ **FLOATING
C17 D.t304 VSUBS -0.06fF
C18 D.n5 VSUBS 0.61fF $ **FLOATING
C19 D.n7 VSUBS 1.37fF $ **FLOATING
C20 D.n8 VSUBS 1.67fF $ **FLOATING
C21 D.t588 VSUBS -0.01fF
C22 D.t16 VSUBS 0.00fF
C23 D.n9 VSUBS 0.73fF $ **FLOATING
C24 D.n10 VSUBS 8.52fF $ **FLOATING
C25 D.n11 VSUBS 2.25fF $ **FLOATING
C26 D.n12 VSUBS 2.95fF $ **FLOATING
C27 D.t490 VSUBS -0.06fF
C28 D.n13 VSUBS 0.61fF $ **FLOATING
C29 D.t130 VSUBS -0.02fF
C30 D.n14 VSUBS 0.20fF $ **FLOATING
C31 D.t533 VSUBS -0.02fF
C32 D.n16 VSUBS 0.20fF $ **FLOATING
C33 D.t82 VSUBS -0.06fF
C34 D.n17 VSUBS 0.61fF $ **FLOATING
C35 D.n19 VSUBS 2.27fF $ **FLOATING
C36 D.n20 VSUBS 2.07fF $ **FLOATING
C37 D.n21 VSUBS 1.75fF $ **FLOATING
C38 D.n22 VSUBS 2.27fF $ **FLOATING
C39 D.t135 VSUBS -0.02fF
C40 D.n23 VSUBS 0.20fF $ **FLOATING
C41 D.t495 VSUBS -0.06fF
C42 D.n24 VSUBS 0.61fF $ **FLOATING
C43 D.t541 VSUBS -0.02fF
C44 D.n26 VSUBS 0.20fF $ **FLOATING
C45 D.t84 VSUBS -0.06fF
C46 D.n27 VSUBS 0.61fF $ **FLOATING
C47 D.n29 VSUBS 1.44fF $ **FLOATING
C48 D.n30 VSUBS 1.67fF $ **FLOATING
C49 D.n31 VSUBS 1.75fF $ **FLOATING
C50 D.n32 VSUBS 2.90fF $ **FLOATING
C51 D.t501 VSUBS -0.06fF
C52 D.n33 VSUBS 0.61fF $ **FLOATING
C53 D.t143 VSUBS -0.02fF
C54 D.n34 VSUBS 0.20fF $ **FLOATING
C55 D.t547 VSUBS -0.02fF
C56 D.n36 VSUBS 0.20fF $ **FLOATING
C57 D.t90 VSUBS -0.06fF
C58 D.n37 VSUBS 0.61fF $ **FLOATING
C59 D.n39 VSUBS 2.27fF $ **FLOATING
C60 D.n40 VSUBS 2.07fF $ **FLOATING
C61 D.n41 VSUBS 1.75fF $ **FLOATING
C62 D.n42 VSUBS 2.27fF $ **FLOATING
C63 D.t148 VSUBS -0.02fF
C64 D.n43 VSUBS 0.20fF $ **FLOATING
C65 D.t503 VSUBS -0.06fF
C66 D.n44 VSUBS 0.61fF $ **FLOATING
C67 D.t552 VSUBS -0.02fF
C68 D.n46 VSUBS 0.20fF $ **FLOATING
C69 D.t95 VSUBS -0.06fF
C70 D.n47 VSUBS 0.61fF $ **FLOATING
C71 D.n49 VSUBS 1.44fF $ **FLOATING
C72 D.n50 VSUBS 1.67fF $ **FLOATING
C73 D.n51 VSUBS 1.75fF $ **FLOATING
C74 D.n52 VSUBS 2.90fF $ **FLOATING
C75 D.t509 VSUBS -0.06fF
C76 D.n53 VSUBS 0.61fF $ **FLOATING
C77 D.t153 VSUBS -0.02fF
C78 D.n54 VSUBS 0.20fF $ **FLOATING
C79 D.t557 VSUBS -0.02fF
C80 D.n56 VSUBS 0.20fF $ **FLOATING
C81 D.t98 VSUBS -0.06fF
C82 D.n57 VSUBS 0.61fF $ **FLOATING
C83 D.n59 VSUBS 2.27fF $ **FLOATING
C84 D.n60 VSUBS 2.07fF $ **FLOATING
C85 D.n61 VSUBS 1.75fF $ **FLOATING
C86 D.n62 VSUBS 2.27fF $ **FLOATING
C87 D.t160 VSUBS -0.02fF
C88 D.n63 VSUBS 0.20fF $ **FLOATING
C89 D.t3 VSUBS -0.06fF
C90 D.n64 VSUBS 0.61fF $ **FLOATING
C91 D.t565 VSUBS -0.02fF
C92 D.n66 VSUBS 0.20fF $ **FLOATING
C93 D.t105 VSUBS -0.06fF
C94 D.n67 VSUBS 0.61fF $ **FLOATING
C95 D.n69 VSUBS 1.44fF $ **FLOATING
C96 D.n70 VSUBS 1.67fF $ **FLOATING
C97 D.n71 VSUBS 1.75fF $ **FLOATING
C98 D.n72 VSUBS 2.90fF $ **FLOATING
C99 D.t8 VSUBS -0.06fF
C100 D.n73 VSUBS 0.61fF $ **FLOATING
C101 D.t273 VSUBS -0.02fF
C102 D.n74 VSUBS 0.20fF $ **FLOATING
C103 D.t58 VSUBS -0.02fF
C104 D.n76 VSUBS 0.20fF $ **FLOATING
C105 D.t213 VSUBS -0.06fF
C106 D.n77 VSUBS 0.61fF $ **FLOATING
C107 D.n79 VSUBS 2.27fF $ **FLOATING
C108 D.n80 VSUBS 2.07fF $ **FLOATING
C109 D.n81 VSUBS 1.75fF $ **FLOATING
C110 D.n82 VSUBS 2.27fF $ **FLOATING
C111 D.t280 VSUBS -0.02fF
C112 D.n83 VSUBS 0.20fF $ **FLOATING
C113 D.t14 VSUBS -0.06fF
C114 D.n84 VSUBS 0.61fF $ **FLOATING
C115 D.t67 VSUBS -0.02fF
C116 D.n86 VSUBS 0.20fF $ **FLOATING
C117 D.t217 VSUBS -0.06fF
C118 D.n87 VSUBS 0.61fF $ **FLOATING
C119 D.n89 VSUBS 1.44fF $ **FLOATING
C120 D.n90 VSUBS 1.67fF $ **FLOATING
C121 D.n91 VSUBS 1.75fF $ **FLOATING
C122 D.n92 VSUBS 2.90fF $ **FLOATING
C123 D.t22 VSUBS -0.06fF
C124 D.n93 VSUBS 0.61fF $ **FLOATING
C125 D.t324 VSUBS -0.02fF
C126 D.n94 VSUBS 0.20fF $ **FLOATING
C127 D.t71 VSUBS -0.02fF
C128 D.n96 VSUBS 0.20fF $ **FLOATING
C129 D.t226 VSUBS -0.06fF
C130 D.n97 VSUBS 0.61fF $ **FLOATING
C131 D.n99 VSUBS 2.27fF $ **FLOATING
C132 D.n100 VSUBS 2.07fF $ **FLOATING
C133 D.n101 VSUBS 1.75fF $ **FLOATING
C134 D.n102 VSUBS 2.27fF $ **FLOATING
C135 D.t440 VSUBS -0.02fF
C136 D.n103 VSUBS 0.20fF $ **FLOATING
C137 D.t429 VSUBS -0.06fF
C138 D.n104 VSUBS 0.61fF $ **FLOATING
C139 D.t266 VSUBS -0.02fF
C140 D.n106 VSUBS 0.20fF $ **FLOATING
C141 D.t496 VSUBS -0.06fF
C142 D.n107 VSUBS 0.61fF $ **FLOATING
C143 D.n109 VSUBS 1.44fF $ **FLOATING
C144 D.n110 VSUBS 1.67fF $ **FLOATING
C145 D.n111 VSUBS 1.75fF $ **FLOATING
C146 D.n112 VSUBS 2.90fF $ **FLOATING
C147 D.t564 VSUBS -0.06fF
C148 D.n113 VSUBS 0.61fF $ **FLOATING
C149 D.t578 VSUBS -0.02fF
C150 D.n114 VSUBS 0.20fF $ **FLOATING
C151 D.t364 VSUBS -0.02fF
C152 D.n116 VSUBS 0.20fF $ **FLOATING
C153 D.t30 VSUBS -0.06fF
C154 D.n117 VSUBS 0.61fF $ **FLOATING
C155 D.n119 VSUBS 2.27fF $ **FLOATING
C156 D.n120 VSUBS 2.07fF $ **FLOATING
C157 D.n121 VSUBS 1.75fF $ **FLOATING
C158 D.n122 VSUBS 2.27fF $ **FLOATING
C159 D.t102 VSUBS -0.02fF
C160 D.n123 VSUBS 0.20fF $ **FLOATING
C161 D.t93 VSUBS -0.06fF
C162 D.n124 VSUBS 0.61fF $ **FLOATING
C163 D.t507 VSUBS -0.02fF
C164 D.n126 VSUBS 0.20fF $ **FLOATING
C165 D.t159 VSUBS -0.06fF
C166 D.n127 VSUBS 0.61fF $ **FLOATING
C167 D.n129 VSUBS 1.44fF $ **FLOATING
C168 D.n130 VSUBS 1.67fF $ **FLOATING
C169 D.n131 VSUBS 1.75fF $ **FLOATING
C170 D.n132 VSUBS 2.90fF $ **FLOATING
C171 D.t242 VSUBS -0.06fF
C172 D.n133 VSUBS 0.61fF $ **FLOATING
C173 D.t259 VSUBS -0.02fF
C174 D.n134 VSUBS 0.20fF $ **FLOATING
C175 D.t43 VSUBS -0.02fF
C176 D.n136 VSUBS 0.20fF $ **FLOATING
C177 D.t308 VSUBS -0.06fF
C178 D.n137 VSUBS 0.61fF $ **FLOATING
C179 D.n139 VSUBS 2.27fF $ **FLOATING
C180 D.n140 VSUBS 2.07fF $ **FLOATING
C181 D.n141 VSUBS 1.75fF $ **FLOATING
C182 D.n142 VSUBS 1.23fF $ **FLOATING
C183 D.n143 VSUBS 1.95fF $ **FLOATING
C184 D.t396 VSUBS -0.02fF
C185 D.n144 VSUBS 0.20fF $ **FLOATING
C186 D.t378 VSUBS -0.06fF
C187 D.n145 VSUBS 0.61fF $ **FLOATING
C188 D.t182 VSUBS -0.02fF
C189 D.n147 VSUBS 0.20fF $ **FLOATING
C190 D.t450 VSUBS -0.06fF
C191 D.n148 VSUBS 0.61fF $ **FLOATING
C192 D.n150 VSUBS 1.88fF $ **FLOATING
C193 D.n151 VSUBS 1.67fF $ **FLOATING
C194 D.n152 VSUBS 1.75fF $ **FLOATING
C195 D.n153 VSUBS 0.09fF $ **FLOATING
C196 D.n154 VSUBS 0.09fF $ **FLOATING
C197 D.n155 VSUBS 0.07fF $ **FLOATING
C198 D.n156 VSUBS 0.06fF $ **FLOATING
C199 D.n157 VSUBS 0.04fF $ **FLOATING
C200 D.n158 VSUBS 0.03fF $ **FLOATING
C201 D.n159 VSUBS 0.06fF $ **FLOATING
C202 D.n160 VSUBS 0.20fF $ **FLOATING
C203 D.n161 VSUBS 0.06fF $ **FLOATING
C204 D.n162 VSUBS 0.08fF $ **FLOATING
C205 D.n163 VSUBS 0.40fF $ **FLOATING
C206 D.n164 VSUBS 0.14fF $ **FLOATING
C207 D.n165 VSUBS 0.24fF $ **FLOATING
C208 D.n166 VSUBS 0.32fF $ **FLOATING
C209 D.n167 VSUBS 0.19fF $ **FLOATING
C210 D.n168 VSUBS 0.13fF $ **FLOATING
C211 D.t488 VSUBS -0.02fF
C212 D.n169 VSUBS 0.20fF $ **FLOATING
C213 D.t456 VSUBS -0.06fF
C214 D.n170 VSUBS 0.61fF $ **FLOATING
C215 D.t282 VSUBS -0.02fF
C216 D.n172 VSUBS 0.20fF $ **FLOATING
C217 D.t594 VSUBS -0.06fF
C218 D.n173 VSUBS 0.61fF $ **FLOATING
C219 D.n175 VSUBS 0.11fF $ **FLOATING
C220 D.n176 VSUBS 0.10fF $ **FLOATING
C221 D.n177 VSUBS 0.10fF $ **FLOATING
C222 D.n178 VSUBS 1.16fF $ **FLOATING
C223 D.n179 VSUBS 1.48fF $ **FLOATING
C224 D.n180 VSUBS 1.64fF $ **FLOATING
C225 D.n181 VSUBS 0.33fF $ **FLOATING
C226 D.n182 VSUBS 3.26fF $ **FLOATING
C227 D.n183 VSUBS 11.54fF $ **FLOATING
C228 D.n184 VSUBS 1.32fF $ **FLOATING
C229 D.n185 VSUBS 9.63fF $ **FLOATING
C230 D.n186 VSUBS 9.63fF $ **FLOATING
C231 D.n187 VSUBS 9.63fF $ **FLOATING
C232 D.n188 VSUBS 9.63fF $ **FLOATING
C233 D.n189 VSUBS 9.63fF $ **FLOATING
C234 D.n190 VSUBS 14.39fF $ **FLOATING
C235 D.n191 VSUBS 2.02fF $ **FLOATING
C236 D.n192 VSUBS 0.08fF $ **FLOATING
C237 D.n193 VSUBS 0.24fF $ **FLOATING
C238 D.t185 VSUBS 0.00fF
C239 D.t56 VSUBS -0.01fF
C240 D.n194 VSUBS 0.73fF $ **FLOATING
C241 D.n195 VSUBS 0.30fF $ **FLOATING
C242 D.n196 VSUBS 0.24fF $ **FLOATING
C243 D.n197 VSUBS 0.14fF $ **FLOATING
C244 D.n198 VSUBS 0.07fF $ **FLOATING
C245 D.n199 VSUBS 0.06fF $ **FLOATING
C246 D.n200 VSUBS 0.41fF $ **FLOATING
C247 D.n201 VSUBS 0.03fF $ **FLOATING
C248 D.n202 VSUBS 0.08fF $ **FLOATING
C249 D.n203 VSUBS 0.08fF $ **FLOATING
C250 D.n204 VSUBS 0.28fF $ **FLOATING
C251 D.n205 VSUBS 0.05fF $ **FLOATING
C252 D.n206 VSUBS 0.09fF $ **FLOATING
C253 D.n207 VSUBS 0.20fF $ **FLOATING
C254 D.n208 VSUBS 0.31fF $ **FLOATING
C255 D.n209 VSUBS 2.26fF $ **FLOATING
C256 D.n210 VSUBS 0.95fF $ **FLOATING
C257 D.n211 VSUBS 1.64fF $ **FLOATING
C258 D.t331 VSUBS 0.00fF
C259 D.t288 VSUBS -0.06fF
C260 D.n212 VSUBS 0.25fF $ **FLOATING
C261 D.n213 VSUBS 0.33fF $ **FLOATING
C262 D.t543 VSUBS 0.00fF
C263 D.n214 VSUBS 0.33fF $ **FLOATING
C264 D.n215 VSUBS 10.45fF $ **FLOATING
C265 D.n216 VSUBS 1.87fF $ **FLOATING
C266 D.t295 VSUBS -0.06fF
C267 D.n217 VSUBS 0.61fF $ **FLOATING
C268 D.t549 VSUBS -0.02fF
C269 D.n218 VSUBS 0.20fF $ **FLOATING
C270 D.t340 VSUBS -0.02fF
C271 D.n220 VSUBS 0.20fF $ **FLOATING
C272 D.t497 VSUBS -0.06fF
C273 D.n221 VSUBS 0.61fF $ **FLOATING
C274 D.n223 VSUBS 0.41fF $ **FLOATING
C275 D.n224 VSUBS 0.31fF $ **FLOATING
C276 D.n225 VSUBS 1.33fF $ **FLOATING
C277 D.n226 VSUBS 2.21fF $ **FLOATING
C278 D.n227 VSUBS 2.03fF $ **FLOATING
C279 D.n228 VSUBS 2.90fF $ **FLOATING
C280 D.t298 VSUBS -0.06fF
C281 D.n229 VSUBS 0.61fF $ **FLOATING
C282 D.t553 VSUBS -0.02fF
C283 D.n230 VSUBS 0.20fF $ **FLOATING
C284 D.t343 VSUBS -0.02fF
C285 D.n232 VSUBS 0.20fF $ **FLOATING
C286 D.t502 VSUBS -0.06fF
C287 D.n233 VSUBS 0.61fF $ **FLOATING
C288 D.n235 VSUBS 0.26fF $ **FLOATING
C289 D.n236 VSUBS 0.31fF $ **FLOATING
C290 D.n237 VSUBS 0.75fF $ **FLOATING
C291 D.n238 VSUBS 0.44fF $ **FLOATING
C292 D.n239 VSUBS 0.25fF $ **FLOATING
C293 D.n240 VSUBS 2.49fF $ **FLOATING
C294 D.n241 VSUBS 1.75fF $ **FLOATING
C295 D.n242 VSUBS 2.08fF $ **FLOATING
C296 D.t303 VSUBS -0.06fF
C297 D.n243 VSUBS 0.61fF $ **FLOATING
C298 D.t558 VSUBS -0.02fF
C299 D.n244 VSUBS 0.20fF $ **FLOATING
C300 D.t348 VSUBS -0.02fF
C301 D.n246 VSUBS 0.20fF $ **FLOATING
C302 D.t505 VSUBS -0.06fF
C303 D.n247 VSUBS 0.61fF $ **FLOATING
C304 D.n249 VSUBS 0.26fF $ **FLOATING
C305 D.n250 VSUBS 0.31fF $ **FLOATING
C306 D.n251 VSUBS 0.75fF $ **FLOATING
C307 D.n252 VSUBS 0.44fF $ **FLOATING
C308 D.n253 VSUBS 0.25fF $ **FLOATING
C309 D.n254 VSUBS 2.09fF $ **FLOATING
C310 D.n255 VSUBS 1.75fF $ **FLOATING
C311 D.n256 VSUBS 2.36fF $ **FLOATING
C312 D.t309 VSUBS -0.06fF
C313 D.n257 VSUBS 0.61fF $ **FLOATING
C314 D.t566 VSUBS -0.02fF
C315 D.n258 VSUBS 0.20fF $ **FLOATING
C316 D.t357 VSUBS -0.02fF
C317 D.n260 VSUBS 0.20fF $ **FLOATING
C318 D.t511 VSUBS -0.06fF
C319 D.n261 VSUBS 0.61fF $ **FLOATING
C320 D.n263 VSUBS 0.26fF $ **FLOATING
C321 D.n264 VSUBS 0.31fF $ **FLOATING
C322 D.n265 VSUBS 0.75fF $ **FLOATING
C323 D.n266 VSUBS 0.44fF $ **FLOATING
C324 D.n267 VSUBS 0.25fF $ **FLOATING
C325 D.n268 VSUBS 2.09fF $ **FLOATING
C326 D.n269 VSUBS 1.75fF $ **FLOATING
C327 D.n270 VSUBS 2.36fF $ **FLOATING
C328 D.t312 VSUBS -0.06fF
C329 D.n271 VSUBS 0.61fF $ **FLOATING
C330 D.t570 VSUBS -0.02fF
C331 D.n272 VSUBS 0.20fF $ **FLOATING
C332 D.t360 VSUBS -0.02fF
C333 D.n274 VSUBS 0.20fF $ **FLOATING
C334 D.t517 VSUBS -0.06fF
C335 D.n275 VSUBS 0.61fF $ **FLOATING
C336 D.n277 VSUBS 0.26fF $ **FLOATING
C337 D.n278 VSUBS 0.31fF $ **FLOATING
C338 D.n279 VSUBS 0.75fF $ **FLOATING
C339 D.n280 VSUBS 0.44fF $ **FLOATING
C340 D.n281 VSUBS 0.25fF $ **FLOATING
C341 D.n282 VSUBS 2.09fF $ **FLOATING
C342 D.n283 VSUBS 1.75fF $ **FLOATING
C343 D.n284 VSUBS 2.36fF $ **FLOATING
C344 D.t319 VSUBS -0.06fF
C345 D.n285 VSUBS 0.61fF $ **FLOATING
C346 D.t579 VSUBS -0.02fF
C347 D.n286 VSUBS 0.20fF $ **FLOATING
C348 D.t366 VSUBS -0.02fF
C349 D.n288 VSUBS 0.20fF $ **FLOATING
C350 D.t520 VSUBS -0.06fF
C351 D.n289 VSUBS 0.61fF $ **FLOATING
C352 D.n291 VSUBS 0.26fF $ **FLOATING
C353 D.n292 VSUBS 0.31fF $ **FLOATING
C354 D.n293 VSUBS 0.75fF $ **FLOATING
C355 D.n294 VSUBS 0.44fF $ **FLOATING
C356 D.n295 VSUBS 0.25fF $ **FLOATING
C357 D.n296 VSUBS 2.09fF $ **FLOATING
C358 D.n297 VSUBS 1.75fF $ **FLOATING
C359 D.n298 VSUBS 2.36fF $ **FLOATING
C360 D.t422 VSUBS -0.06fF
C361 D.n299 VSUBS 0.61fF $ **FLOATING
C362 D.t591 VSUBS -0.02fF
C363 D.n300 VSUBS 0.20fF $ **FLOATING
C364 D.t377 VSUBS -0.02fF
C365 D.n302 VSUBS 0.20fF $ **FLOATING
C366 D.t528 VSUBS -0.06fF
C367 D.n303 VSUBS 0.61fF $ **FLOATING
C368 D.n305 VSUBS 0.26fF $ **FLOATING
C369 D.n306 VSUBS 0.31fF $ **FLOATING
C370 D.n307 VSUBS 0.75fF $ **FLOATING
C371 D.n308 VSUBS 0.44fF $ **FLOATING
C372 D.n309 VSUBS 0.25fF $ **FLOATING
C373 D.n310 VSUBS 2.09fF $ **FLOATING
C374 D.n311 VSUBS 1.75fF $ **FLOATING
C375 D.n312 VSUBS 2.36fF $ **FLOATING
C376 D.t430 VSUBS -0.06fF
C377 D.n313 VSUBS 0.61fF $ **FLOATING
C378 D.t469 VSUBS -0.02fF
C379 D.n314 VSUBS 0.20fF $ **FLOATING
C380 D.t479 VSUBS -0.02fF
C381 D.n316 VSUBS 0.20fF $ **FLOATING
C382 D.t24 VSUBS -0.06fF
C383 D.n317 VSUBS 0.61fF $ **FLOATING
C384 D.n319 VSUBS 0.26fF $ **FLOATING
C385 D.n320 VSUBS 0.31fF $ **FLOATING
C386 D.n321 VSUBS 0.75fF $ **FLOATING
C387 D.n322 VSUBS 0.44fF $ **FLOATING
C388 D.n323 VSUBS 0.25fF $ **FLOATING
C389 D.n324 VSUBS 2.09fF $ **FLOATING
C390 D.n325 VSUBS 1.75fF $ **FLOATING
C391 D.n326 VSUBS 2.36fF $ **FLOATING
C392 D.t562 VSUBS -0.06fF
C393 D.n327 VSUBS 0.61fF $ **FLOATING
C394 D.t575 VSUBS -0.02fF
C395 D.n328 VSUBS 0.20fF $ **FLOATING
C396 D.t401 VSUBS -0.02fF
C397 D.n330 VSUBS 0.20fF $ **FLOATING
C398 D.t29 VSUBS -0.06fF
C399 D.n331 VSUBS 0.61fF $ **FLOATING
C400 D.n333 VSUBS 0.26fF $ **FLOATING
C401 D.n334 VSUBS 0.31fF $ **FLOATING
C402 D.n335 VSUBS 0.75fF $ **FLOATING
C403 D.n336 VSUBS 0.44fF $ **FLOATING
C404 D.n337 VSUBS 0.25fF $ **FLOATING
C405 D.n338 VSUBS 2.09fF $ **FLOATING
C406 D.n339 VSUBS 1.75fF $ **FLOATING
C407 D.n340 VSUBS 2.36fF $ **FLOATING
C408 D.t91 VSUBS -0.06fF
C409 D.n341 VSUBS 0.61fF $ **FLOATING
C410 D.t99 VSUBS -0.02fF
C411 D.n342 VSUBS 0.20fF $ **FLOATING
C412 D.t504 VSUBS -0.02fF
C413 D.n344 VSUBS 0.20fF $ **FLOATING
C414 D.t158 VSUBS -0.06fF
C415 D.n345 VSUBS 0.61fF $ **FLOATING
C416 D.n347 VSUBS 0.26fF $ **FLOATING
C417 D.n348 VSUBS 0.31fF $ **FLOATING
C418 D.n349 VSUBS 0.75fF $ **FLOATING
C419 D.n350 VSUBS 0.44fF $ **FLOATING
C420 D.n351 VSUBS 0.25fF $ **FLOATING
C421 D.n352 VSUBS 2.09fF $ **FLOATING
C422 D.n353 VSUBS 1.75fF $ **FLOATING
C423 D.n354 VSUBS 2.36fF $ **FLOATING
C424 D.t238 VSUBS -0.06fF
C425 D.n355 VSUBS 0.61fF $ **FLOATING
C426 D.t255 VSUBS -0.02fF
C427 D.n356 VSUBS 0.20fF $ **FLOATING
C428 D.t40 VSUBS -0.02fF
C429 D.n358 VSUBS 0.20fF $ **FLOATING
C430 D.t305 VSUBS -0.06fF
C431 D.n359 VSUBS 0.61fF $ **FLOATING
C432 D.n361 VSUBS 0.26fF $ **FLOATING
C433 D.n362 VSUBS 0.31fF $ **FLOATING
C434 D.n363 VSUBS 0.75fF $ **FLOATING
C435 D.n364 VSUBS 0.44fF $ **FLOATING
C436 D.n365 VSUBS 0.25fF $ **FLOATING
C437 D.n366 VSUBS 2.09fF $ **FLOATING
C438 D.n367 VSUBS 1.75fF $ **FLOATING
C439 D.n368 VSUBS 2.36fF $ **FLOATING
C440 D.t376 VSUBS -0.06fF
C441 D.n369 VSUBS 0.61fF $ **FLOATING
C442 D.t393 VSUBS -0.02fF
C443 D.n370 VSUBS 0.20fF $ **FLOATING
C444 D.t179 VSUBS -0.02fF
C445 D.n372 VSUBS 0.20fF $ **FLOATING
C446 D.t448 VSUBS -0.06fF
C447 D.n373 VSUBS 0.61fF $ **FLOATING
C448 D.n375 VSUBS 0.26fF $ **FLOATING
C449 D.n376 VSUBS 0.31fF $ **FLOATING
C450 D.n377 VSUBS 0.75fF $ **FLOATING
C451 D.n378 VSUBS 0.44fF $ **FLOATING
C452 D.n379 VSUBS 0.25fF $ **FLOATING
C453 D.n380 VSUBS 2.09fF $ **FLOATING
C454 D.n381 VSUBS 1.75fF $ **FLOATING
C455 D.n382 VSUBS 2.36fF $ **FLOATING
C456 D.t514 VSUBS -0.06fF
C457 D.n383 VSUBS 0.61fF $ **FLOATING
C458 D.t525 VSUBS -0.02fF
C459 D.n384 VSUBS 0.20fF $ **FLOATING
C460 D.t316 VSUBS -0.02fF
C461 D.n386 VSUBS 0.20fF $ **FLOATING
C462 D.t590 VSUBS -0.06fF
C463 D.n387 VSUBS 0.61fF $ **FLOATING
C464 D.n389 VSUBS 0.26fF $ **FLOATING
C465 D.n390 VSUBS 0.31fF $ **FLOATING
C466 D.n391 VSUBS 0.75fF $ **FLOATING
C467 D.n392 VSUBS 0.44fF $ **FLOATING
C468 D.n393 VSUBS 0.25fF $ **FLOATING
C469 D.n394 VSUBS 2.09fF $ **FLOATING
C470 D.n395 VSUBS 1.75fF $ **FLOATING
C471 D.n396 VSUBS 2.36fF $ **FLOATING
C472 D.t52 VSUBS -0.06fF
C473 D.n397 VSUBS 0.61fF $ **FLOATING
C474 D.t65 VSUBS -0.02fF
C475 D.n398 VSUBS 0.20fF $ **FLOATING
C476 D.t464 VSUBS -0.02fF
C477 D.n400 VSUBS 0.20fF $ **FLOATING
C478 D.t109 VSUBS -0.06fF
C479 D.n401 VSUBS 0.61fF $ **FLOATING
C480 D.n403 VSUBS 0.26fF $ **FLOATING
C481 D.n404 VSUBS 0.31fF $ **FLOATING
C482 D.n405 VSUBS 0.75fF $ **FLOATING
C483 D.n406 VSUBS 0.44fF $ **FLOATING
C484 D.n407 VSUBS 0.25fF $ **FLOATING
C485 D.n408 VSUBS 2.09fF $ **FLOATING
C486 D.n409 VSUBS 1.69fF $ **FLOATING
C487 D.n410 VSUBS 0.80fF $ **FLOATING
C488 D.t606 VSUBS -0.02fF
C489 D.n411 VSUBS 0.20fF $ **FLOATING
C490 D.t265 VSUBS -0.01fF
C491 D.n412 VSUBS 0.55fF $ **FLOATING
C492 D.t191 VSUBS -0.02fF
C493 D.n413 VSUBS 0.56fF $ **FLOATING
C494 D.n414 VSUBS 0.19fF $ **FLOATING
C495 D.n415 VSUBS 2.02fF $ **FLOATING
C496 D.n416 VSUBS 14.23fF $ **FLOATING
C497 D.n417 VSUBS 9.31fF $ **FLOATING
C498 D.n418 VSUBS 2.16fF $ **FLOATING
C499 D.n419 VSUBS 0.83fF $ **FLOATING
C500 D.n420 VSUBS 0.44fF $ **FLOATING
C501 D.n421 VSUBS 2.31fF $ **FLOATING
C502 D.n422 VSUBS 2.40fF $ **FLOATING
C503 D.t137 VSUBS 0.00fF
C504 D.t92 VSUBS -0.06fF
C505 D.n423 VSUBS 0.25fF $ **FLOATING
C506 D.n424 VSUBS 0.33fF $ **FLOATING
C507 D.t351 VSUBS 0.00fF
C508 D.n425 VSUBS 0.33fF $ **FLOATING
C509 D.n426 VSUBS 10.45fF $ **FLOATING
C510 D.n427 VSUBS 1.87fF $ **FLOATING
C511 D.t96 VSUBS -0.06fF
C512 D.n428 VSUBS 0.61fF $ **FLOATING
C513 D.t359 VSUBS -0.02fF
C514 D.n429 VSUBS 0.20fF $ **FLOATING
C515 D.t144 VSUBS -0.02fF
C516 D.n431 VSUBS 0.20fF $ **FLOATING
C517 D.t306 VSUBS -0.06fF
C518 D.n432 VSUBS 0.61fF $ **FLOATING
C519 D.n434 VSUBS 0.41fF $ **FLOATING
C520 D.n435 VSUBS 0.31fF $ **FLOATING
C521 D.n436 VSUBS 1.33fF $ **FLOATING
C522 D.n437 VSUBS 2.21fF $ **FLOATING
C523 D.n438 VSUBS 2.03fF $ **FLOATING
C524 D.n439 VSUBS 2.90fF $ **FLOATING
C525 D.t100 VSUBS -0.06fF
C526 D.n440 VSUBS 0.61fF $ **FLOATING
C527 D.t361 VSUBS -0.02fF
C528 D.n441 VSUBS 0.20fF $ **FLOATING
C529 D.t149 VSUBS -0.02fF
C530 D.n443 VSUBS 0.20fF $ **FLOATING
C531 D.t310 VSUBS -0.06fF
C532 D.n444 VSUBS 0.61fF $ **FLOATING
C533 D.n446 VSUBS 0.26fF $ **FLOATING
C534 D.n447 VSUBS 0.31fF $ **FLOATING
C535 D.n448 VSUBS 0.75fF $ **FLOATING
C536 D.n449 VSUBS 0.44fF $ **FLOATING
C537 D.n450 VSUBS 0.25fF $ **FLOATING
C538 D.n451 VSUBS 2.49fF $ **FLOATING
C539 D.n452 VSUBS 1.75fF $ **FLOATING
C540 D.n453 VSUBS 2.08fF $ **FLOATING
C541 D.t106 VSUBS -0.06fF
C542 D.n454 VSUBS 0.61fF $ **FLOATING
C543 D.t369 VSUBS -0.02fF
C544 D.n455 VSUBS 0.20fF $ **FLOATING
C545 D.t155 VSUBS -0.02fF
C546 D.n457 VSUBS 0.20fF $ **FLOATING
C547 D.t314 VSUBS -0.06fF
C548 D.n458 VSUBS 0.61fF $ **FLOATING
C549 D.n460 VSUBS 0.26fF $ **FLOATING
C550 D.n461 VSUBS 0.31fF $ **FLOATING
C551 D.n462 VSUBS 0.75fF $ **FLOATING
C552 D.n463 VSUBS 0.44fF $ **FLOATING
C553 D.n464 VSUBS 0.25fF $ **FLOATING
C554 D.n465 VSUBS 2.09fF $ **FLOATING
C555 D.n466 VSUBS 1.75fF $ **FLOATING
C556 D.n467 VSUBS 2.36fF $ **FLOATING
C557 D.t111 VSUBS -0.06fF
C558 D.n468 VSUBS 0.61fF $ **FLOATING
C559 D.t379 VSUBS -0.02fF
C560 D.n469 VSUBS 0.20fF $ **FLOATING
C561 D.t163 VSUBS -0.02fF
C562 D.n471 VSUBS 0.20fF $ **FLOATING
C563 D.t320 VSUBS -0.06fF
C564 D.n472 VSUBS 0.61fF $ **FLOATING
C565 D.n474 VSUBS 0.26fF $ **FLOATING
C566 D.n475 VSUBS 0.31fF $ **FLOATING
C567 D.n476 VSUBS 0.75fF $ **FLOATING
C568 D.n477 VSUBS 0.44fF $ **FLOATING
C569 D.n478 VSUBS 0.25fF $ **FLOATING
C570 D.n479 VSUBS 2.09fF $ **FLOATING
C571 D.n480 VSUBS 1.75fF $ **FLOATING
C572 D.n481 VSUBS 2.36fF $ **FLOATING
C573 D.t115 VSUBS -0.06fF
C574 D.n482 VSUBS 0.61fF $ **FLOATING
C575 D.t385 VSUBS -0.02fF
C576 D.n483 VSUBS 0.20fF $ **FLOATING
C577 D.t170 VSUBS -0.02fF
C578 D.n485 VSUBS 0.20fF $ **FLOATING
C579 D.t325 VSUBS -0.06fF
C580 D.n486 VSUBS 0.61fF $ **FLOATING
C581 D.n488 VSUBS 0.26fF $ **FLOATING
C582 D.n489 VSUBS 0.31fF $ **FLOATING
C583 D.n490 VSUBS 0.75fF $ **FLOATING
C584 D.n491 VSUBS 0.44fF $ **FLOATING
C585 D.n492 VSUBS 0.25fF $ **FLOATING
C586 D.n493 VSUBS 2.09fF $ **FLOATING
C587 D.n494 VSUBS 1.75fF $ **FLOATING
C588 D.n495 VSUBS 2.36fF $ **FLOATING
C589 D.t125 VSUBS -0.06fF
C590 D.n496 VSUBS 0.61fF $ **FLOATING
C591 D.t551 VSUBS -0.02fF
C592 D.n497 VSUBS 0.20fF $ **FLOATING
C593 D.t180 VSUBS -0.02fF
C594 D.n499 VSUBS 0.20fF $ **FLOATING
C595 D.t333 VSUBS -0.06fF
C596 D.n500 VSUBS 0.61fF $ **FLOATING
C597 D.n502 VSUBS 0.26fF $ **FLOATING
C598 D.n503 VSUBS 0.31fF $ **FLOATING
C599 D.n504 VSUBS 0.75fF $ **FLOATING
C600 D.n505 VSUBS 0.44fF $ **FLOATING
C601 D.n506 VSUBS 0.25fF $ **FLOATING
C602 D.n507 VSUBS 2.09fF $ **FLOATING
C603 D.n508 VSUBS 1.75fF $ **FLOATING
C604 D.n509 VSUBS 2.36fF $ **FLOATING
C605 D.t87 VSUBS -0.06fF
C606 D.n510 VSUBS 0.61fF $ **FLOATING
C607 D.t55 VSUBS -0.02fF
C608 D.n511 VSUBS 0.20fF $ **FLOATING
C609 D.t486 VSUBS -0.02fF
C610 D.n513 VSUBS 0.20fF $ **FLOATING
C611 D.t101 VSUBS -0.06fF
C612 D.n514 VSUBS 0.61fF $ **FLOATING
C613 D.n516 VSUBS 0.26fF $ **FLOATING
C614 D.n517 VSUBS 0.31fF $ **FLOATING
C615 D.n518 VSUBS 0.75fF $ **FLOATING
C616 D.n519 VSUBS 0.44fF $ **FLOATING
C617 D.n520 VSUBS 0.25fF $ **FLOATING
C618 D.n521 VSUBS 2.09fF $ **FLOATING
C619 D.n522 VSUBS 1.75fF $ **FLOATING
C620 D.n523 VSUBS 2.36fF $ **FLOATING
C621 D.t237 VSUBS -0.06fF
C622 D.n524 VSUBS 0.61fF $ **FLOATING
C623 D.t251 VSUBS -0.02fF
C624 D.n525 VSUBS 0.20fF $ **FLOATING
C625 D.t39 VSUBS -0.02fF
C626 D.n527 VSUBS 0.20fF $ **FLOATING
C627 D.t301 VSUBS -0.06fF
C628 D.n528 VSUBS 0.61fF $ **FLOATING
C629 D.n530 VSUBS 0.26fF $ **FLOATING
C630 D.n531 VSUBS 0.31fF $ **FLOATING
C631 D.n532 VSUBS 0.75fF $ **FLOATING
C632 D.n533 VSUBS 0.44fF $ **FLOATING
C633 D.n534 VSUBS 0.25fF $ **FLOATING
C634 D.n535 VSUBS 2.09fF $ **FLOATING
C635 D.n536 VSUBS 1.75fF $ **FLOATING
C636 D.n537 VSUBS 2.36fF $ **FLOATING
C637 D.t371 VSUBS -0.06fF
C638 D.n538 VSUBS 0.61fF $ **FLOATING
C639 D.t389 VSUBS -0.02fF
C640 D.n539 VSUBS 0.20fF $ **FLOATING
C641 D.t174 VSUBS -0.02fF
C642 D.n541 VSUBS 0.20fF $ **FLOATING
C643 D.t446 VSUBS -0.06fF
C644 D.n542 VSUBS 0.61fF $ **FLOATING
C645 D.n544 VSUBS 0.26fF $ **FLOATING
C646 D.n545 VSUBS 0.31fF $ **FLOATING
C647 D.n546 VSUBS 0.75fF $ **FLOATING
C648 D.n547 VSUBS 0.44fF $ **FLOATING
C649 D.n548 VSUBS 0.25fF $ **FLOATING
C650 D.n549 VSUBS 2.09fF $ **FLOATING
C651 D.n550 VSUBS 1.75fF $ **FLOATING
C652 D.n551 VSUBS 2.36fF $ **FLOATING
C653 D.t510 VSUBS -0.06fF
C654 D.n552 VSUBS 0.61fF $ **FLOATING
C655 D.t522 VSUBS -0.02fF
C656 D.n553 VSUBS 0.20fF $ **FLOATING
C657 D.t313 VSUBS -0.02fF
C658 D.n555 VSUBS 0.20fF $ **FLOATING
C659 D.t584 VSUBS -0.06fF
C660 D.n556 VSUBS 0.61fF $ **FLOATING
C661 D.n558 VSUBS 0.26fF $ **FLOATING
C662 D.n559 VSUBS 0.31fF $ **FLOATING
C663 D.n560 VSUBS 0.75fF $ **FLOATING
C664 D.n561 VSUBS 0.44fF $ **FLOATING
C665 D.n562 VSUBS 0.25fF $ **FLOATING
C666 D.n563 VSUBS 2.09fF $ **FLOATING
C667 D.n564 VSUBS 1.75fF $ **FLOATING
C668 D.n565 VSUBS 2.36fF $ **FLOATING
C669 D.t49 VSUBS -0.06fF
C670 D.n566 VSUBS 0.61fF $ **FLOATING
C671 D.t61 VSUBS -0.02fF
C672 D.n567 VSUBS 0.20fF $ **FLOATING
C673 D.t460 VSUBS -0.02fF
C674 D.n569 VSUBS 0.20fF $ **FLOATING
C675 D.t107 VSUBS -0.06fF
C676 D.n570 VSUBS 0.61fF $ **FLOATING
C677 D.n572 VSUBS 0.26fF $ **FLOATING
C678 D.n573 VSUBS 0.31fF $ **FLOATING
C679 D.n574 VSUBS 0.75fF $ **FLOATING
C680 D.n575 VSUBS 0.44fF $ **FLOATING
C681 D.n576 VSUBS 0.25fF $ **FLOATING
C682 D.n577 VSUBS 2.09fF $ **FLOATING
C683 D.n578 VSUBS 1.75fF $ **FLOATING
C684 D.n579 VSUBS 2.36fF $ **FLOATING
C685 D.t189 VSUBS -0.06fF
C686 D.n580 VSUBS 0.61fF $ **FLOATING
C687 D.t203 VSUBS -0.02fF
C688 D.n581 VSUBS 0.20fF $ **FLOATING
C689 D.t604 VSUBS -0.02fF
C690 D.n583 VSUBS 0.20fF $ **FLOATING
C691 D.t263 VSUBS -0.06fF
C692 D.n584 VSUBS 0.61fF $ **FLOATING
C693 D.n586 VSUBS 0.26fF $ **FLOATING
C694 D.n587 VSUBS 0.31fF $ **FLOATING
C695 D.n588 VSUBS 0.75fF $ **FLOATING
C696 D.n589 VSUBS 0.44fF $ **FLOATING
C697 D.n590 VSUBS 0.25fF $ **FLOATING
C698 D.n591 VSUBS 2.09fF $ **FLOATING
C699 D.n592 VSUBS 1.69fF $ **FLOATING
C700 D.n593 VSUBS 0.80fF $ **FLOATING
C701 D.t121 VSUBS -0.02fF
C702 D.n594 VSUBS 0.20fF $ **FLOATING
C703 D.t400 VSUBS -0.01fF
C704 D.n595 VSUBS 0.55fF $ **FLOATING
C705 D.t323 VSUBS -0.02fF
C706 D.n596 VSUBS 0.56fF $ **FLOATING
C707 D.n597 VSUBS 9.31fF $ **FLOATING
C708 D.n598 VSUBS 2.16fF $ **FLOATING
C709 D.n599 VSUBS 0.83fF $ **FLOATING
C710 D.n600 VSUBS 0.44fF $ **FLOATING
C711 D.n601 VSUBS 2.31fF $ **FLOATING
C712 D.n602 VSUBS 2.40fF $ **FLOATING
C713 D.t561 VSUBS 0.00fF
C714 D.t513 VSUBS -0.06fF
C715 D.n603 VSUBS 0.25fF $ **FLOATING
C716 D.n604 VSUBS 0.33fF $ **FLOATING
C717 D.t157 VSUBS 0.00fF
C718 D.n605 VSUBS 0.33fF $ **FLOATING
C719 D.n606 VSUBS 10.45fF $ **FLOATING
C720 D.n607 VSUBS 1.87fF $ **FLOATING
C721 D.t518 VSUBS -0.06fF
C722 D.n608 VSUBS 0.61fF $ **FLOATING
C723 D.t166 VSUBS -0.02fF
C724 D.n609 VSUBS 0.20fF $ **FLOATING
C725 D.t568 VSUBS -0.02fF
C726 D.n611 VSUBS 0.20fF $ **FLOATING
C727 D.t108 VSUBS -0.06fF
C728 D.n612 VSUBS 0.61fF $ **FLOATING
C729 D.n614 VSUBS 0.41fF $ **FLOATING
C730 D.n615 VSUBS 0.31fF $ **FLOATING
C731 D.n616 VSUBS 1.33fF $ **FLOATING
C732 D.n617 VSUBS 2.21fF $ **FLOATING
C733 D.n618 VSUBS 2.03fF $ **FLOATING
C734 D.n619 VSUBS 2.90fF $ **FLOATING
C735 D.t523 VSUBS -0.06fF
C736 D.n620 VSUBS 0.61fF $ **FLOATING
C737 D.t172 VSUBS -0.02fF
C738 D.n621 VSUBS 0.20fF $ **FLOATING
C739 D.t573 VSUBS -0.02fF
C740 D.n623 VSUBS 0.20fF $ **FLOATING
C741 D.t112 VSUBS -0.06fF
C742 D.n624 VSUBS 0.61fF $ **FLOATING
C743 D.n626 VSUBS 0.26fF $ **FLOATING
C744 D.n627 VSUBS 0.31fF $ **FLOATING
C745 D.n628 VSUBS 0.75fF $ **FLOATING
C746 D.n629 VSUBS 0.44fF $ **FLOATING
C747 D.n630 VSUBS 0.25fF $ **FLOATING
C748 D.n631 VSUBS 2.49fF $ **FLOATING
C749 D.n632 VSUBS 1.75fF $ **FLOATING
C750 D.n633 VSUBS 2.08fF $ **FLOATING
C751 D.t529 VSUBS -0.06fF
C752 D.n634 VSUBS 0.61fF $ **FLOATING
C753 D.t183 VSUBS -0.02fF
C754 D.n635 VSUBS 0.20fF $ **FLOATING
C755 D.t582 VSUBS -0.02fF
C756 D.n637 VSUBS 0.20fF $ **FLOATING
C757 D.t117 VSUBS -0.06fF
C758 D.n638 VSUBS 0.61fF $ **FLOATING
C759 D.n640 VSUBS 0.26fF $ **FLOATING
C760 D.n641 VSUBS 0.31fF $ **FLOATING
C761 D.n642 VSUBS 0.75fF $ **FLOATING
C762 D.n643 VSUBS 0.44fF $ **FLOATING
C763 D.n644 VSUBS 0.25fF $ **FLOATING
C764 D.n645 VSUBS 2.09fF $ **FLOATING
C765 D.n646 VSUBS 1.75fF $ **FLOATING
C766 D.n647 VSUBS 2.36fF $ **FLOATING
C767 D.t537 VSUBS -0.06fF
C768 D.n648 VSUBS 0.61fF $ **FLOATING
C769 D.t81 VSUBS -0.02fF
C770 D.n649 VSUBS 0.20fF $ **FLOATING
C771 D.t592 VSUBS -0.02fF
C772 D.n651 VSUBS 0.20fF $ **FLOATING
C773 D.t126 VSUBS -0.06fF
C774 D.n652 VSUBS 0.61fF $ **FLOATING
C775 D.n654 VSUBS 0.26fF $ **FLOATING
C776 D.n655 VSUBS 0.31fF $ **FLOATING
C777 D.n656 VSUBS 0.75fF $ **FLOATING
C778 D.n657 VSUBS 0.44fF $ **FLOATING
C779 D.n658 VSUBS 0.25fF $ **FLOATING
C780 D.n659 VSUBS 2.09fF $ **FLOATING
C781 D.n660 VSUBS 1.75fF $ **FLOATING
C782 D.n661 VSUBS 2.36fF $ **FLOATING
C783 D.t178 VSUBS -0.06fF
C784 D.n662 VSUBS 0.61fF $ **FLOATING
C785 D.t196 VSUBS -0.02fF
C786 D.n663 VSUBS 0.20fF $ **FLOATING
C787 D.t13 VSUBS -0.02fF
C788 D.n665 VSUBS 0.20fF $ **FLOATING
C789 D.t257 VSUBS -0.06fF
C790 D.n666 VSUBS 0.61fF $ **FLOATING
C791 D.n668 VSUBS 0.26fF $ **FLOATING
C792 D.n669 VSUBS 0.31fF $ **FLOATING
C793 D.n670 VSUBS 0.75fF $ **FLOATING
C794 D.n671 VSUBS 0.44fF $ **FLOATING
C795 D.n672 VSUBS 0.25fF $ **FLOATING
C796 D.n673 VSUBS 2.09fF $ **FLOATING
C797 D.n674 VSUBS 1.75fF $ **FLOATING
C798 D.n675 VSUBS 2.36fF $ **FLOATING
C799 D.t317 VSUBS -0.06fF
C800 D.n676 VSUBS 0.61fF $ **FLOATING
C801 D.t330 VSUBS -0.02fF
C802 D.n677 VSUBS 0.20fF $ **FLOATING
C803 D.t113 VSUBS -0.02fF
C804 D.n679 VSUBS 0.20fF $ **FLOATING
C805 D.t394 VSUBS -0.06fF
C806 D.n680 VSUBS 0.61fF $ **FLOATING
C807 D.n682 VSUBS 0.26fF $ **FLOATING
C808 D.n683 VSUBS 0.31fF $ **FLOATING
C809 D.n684 VSUBS 0.75fF $ **FLOATING
C810 D.n685 VSUBS 0.44fF $ **FLOATING
C811 D.n686 VSUBS 0.25fF $ **FLOATING
C812 D.n687 VSUBS 2.09fF $ **FLOATING
C813 D.n688 VSUBS 1.75fF $ **FLOATING
C814 D.n689 VSUBS 2.36fF $ **FLOATING
C815 D.t508 VSUBS -0.06fF
C816 D.n690 VSUBS 0.61fF $ **FLOATING
C817 D.t478 VSUBS -0.02fF
C818 D.n691 VSUBS 0.20fF $ **FLOATING
C819 D.t270 VSUBS -0.02fF
C820 D.n693 VSUBS 0.20fF $ **FLOATING
C821 D.t526 VSUBS -0.06fF
C822 D.n694 VSUBS 0.61fF $ **FLOATING
C823 D.n696 VSUBS 0.26fF $ **FLOATING
C824 D.n697 VSUBS 0.31fF $ **FLOATING
C825 D.n698 VSUBS 0.75fF $ **FLOATING
C826 D.n699 VSUBS 0.44fF $ **FLOATING
C827 D.n700 VSUBS 0.25fF $ **FLOATING
C828 D.n701 VSUBS 2.09fF $ **FLOATING
C829 D.n702 VSUBS 1.75fF $ **FLOATING
C830 D.n703 VSUBS 2.36fF $ **FLOATING
C831 D.t45 VSUBS -0.06fF
C832 D.n704 VSUBS 0.61fF $ **FLOATING
C833 D.t59 VSUBS -0.02fF
C834 D.n705 VSUBS 0.20fF $ **FLOATING
C835 D.t458 VSUBS -0.02fF
C836 D.n707 VSUBS 0.20fF $ **FLOATING
C837 D.t104 VSUBS -0.06fF
C838 D.n708 VSUBS 0.61fF $ **FLOATING
C839 D.n710 VSUBS 0.26fF $ **FLOATING
C840 D.n711 VSUBS 0.31fF $ **FLOATING
C841 D.n712 VSUBS 0.75fF $ **FLOATING
C842 D.n713 VSUBS 0.44fF $ **FLOATING
C843 D.n714 VSUBS 0.25fF $ **FLOATING
C844 D.n715 VSUBS 2.09fF $ **FLOATING
C845 D.n716 VSUBS 1.75fF $ **FLOATING
C846 D.n717 VSUBS 2.36fF $ **FLOATING
C847 D.t188 VSUBS -0.06fF
C848 D.n718 VSUBS 0.61fF $ **FLOATING
C849 D.t200 VSUBS -0.02fF
C850 D.n719 VSUBS 0.20fF $ **FLOATING
C851 D.t601 VSUBS -0.02fF
C852 D.n721 VSUBS 0.20fF $ **FLOATING
C853 D.t261 VSUBS -0.06fF
C854 D.n722 VSUBS 0.61fF $ **FLOATING
C855 D.n724 VSUBS 0.26fF $ **FLOATING
C856 D.n725 VSUBS 0.31fF $ **FLOATING
C857 D.n726 VSUBS 0.75fF $ **FLOATING
C858 D.n727 VSUBS 0.44fF $ **FLOATING
C859 D.n728 VSUBS 0.25fF $ **FLOATING
C860 D.n729 VSUBS 2.09fF $ **FLOATING
C861 D.n730 VSUBS 1.75fF $ **FLOATING
C862 D.n731 VSUBS 2.36fF $ **FLOATING
C863 D.t321 VSUBS -0.06fF
C864 D.n732 VSUBS 0.61fF $ **FLOATING
C865 D.t336 VSUBS -0.02fF
C866 D.n733 VSUBS 0.20fF $ **FLOATING
C867 D.t116 VSUBS -0.02fF
C868 D.n735 VSUBS 0.20fF $ **FLOATING
C869 D.t399 VSUBS -0.06fF
C870 D.n736 VSUBS 0.61fF $ **FLOATING
C871 D.n738 VSUBS 0.26fF $ **FLOATING
C872 D.n739 VSUBS 0.31fF $ **FLOATING
C873 D.n740 VSUBS 0.75fF $ **FLOATING
C874 D.n741 VSUBS 0.44fF $ **FLOATING
C875 D.n742 VSUBS 0.25fF $ **FLOATING
C876 D.n743 VSUBS 2.09fF $ **FLOATING
C877 D.n744 VSUBS 1.69fF $ **FLOATING
C878 D.n745 VSUBS 0.80fF $ **FLOATING
C879 D.t275 VSUBS -0.02fF
C880 D.n746 VSUBS 0.20fF $ **FLOATING
C881 D.t530 VSUBS -0.01fF
C882 D.n747 VSUBS 0.55fF $ **FLOATING
C883 D.t468 VSUBS -0.02fF
C884 D.n748 VSUBS 0.56fF $ **FLOATING
C885 D.n749 VSUBS 9.31fF $ **FLOATING
C886 D.n750 VSUBS 2.16fF $ **FLOATING
C887 D.n751 VSUBS 0.83fF $ **FLOATING
C888 D.n752 VSUBS 0.44fF $ **FLOATING
C889 D.n753 VSUBS 2.31fF $ **FLOATING
C890 D.n754 VSUBS 2.40fF $ **FLOATING
C891 D.t373 VSUBS 0.00fF
C892 D.t322 VSUBS -0.06fF
C893 D.n755 VSUBS 0.25fF $ **FLOATING
C894 D.n756 VSUBS 0.33fF $ **FLOATING
C895 D.t586 VSUBS 0.00fF
C896 D.n757 VSUBS 0.33fF $ **FLOATING
C897 D.n758 VSUBS 10.45fF $ **FLOATING
C898 D.n759 VSUBS 1.87fF $ **FLOATING
C899 D.t327 VSUBS -0.06fF
C900 D.n760 VSUBS 0.61fF $ **FLOATING
C901 D.t595 VSUBS -0.02fF
C902 D.n761 VSUBS 0.20fF $ **FLOATING
C903 D.t381 VSUBS -0.02fF
C904 D.n763 VSUBS 0.20fF $ **FLOATING
C905 D.t531 VSUBS -0.06fF
C906 D.n764 VSUBS 0.61fF $ **FLOATING
C907 D.n766 VSUBS 0.41fF $ **FLOATING
C908 D.n767 VSUBS 0.31fF $ **FLOATING
C909 D.n768 VSUBS 1.33fF $ **FLOATING
C910 D.n769 VSUBS 2.21fF $ **FLOATING
C911 D.n770 VSUBS 2.03fF $ **FLOATING
C912 D.n771 VSUBS 2.90fF $ **FLOATING
C913 D.t334 VSUBS -0.06fF
C914 D.n772 VSUBS 0.61fF $ **FLOATING
C915 D.t223 VSUBS -0.02fF
C916 D.n773 VSUBS 0.20fF $ **FLOATING
C917 D.t387 VSUBS -0.02fF
C918 D.n775 VSUBS 0.20fF $ **FLOATING
C919 D.t538 VSUBS -0.06fF
C920 D.n776 VSUBS 0.61fF $ **FLOATING
C921 D.n778 VSUBS 0.26fF $ **FLOATING
C922 D.n779 VSUBS 0.31fF $ **FLOATING
C923 D.n780 VSUBS 0.75fF $ **FLOATING
C924 D.n781 VSUBS 0.44fF $ **FLOATING
C925 D.n782 VSUBS 0.25fF $ **FLOATING
C926 D.n783 VSUBS 2.49fF $ **FLOATING
C927 D.n784 VSUBS 1.75fF $ **FLOATING
C928 D.n785 VSUBS 2.08fF $ **FLOATING
C929 D.t315 VSUBS -0.06fF
C930 D.n786 VSUBS 0.61fF $ **FLOATING
C931 D.t326 VSUBS -0.02fF
C932 D.n787 VSUBS 0.20fF $ **FLOATING
C933 D.t147 VSUBS -0.02fF
C934 D.n789 VSUBS 0.20fF $ **FLOATING
C935 D.t391 VSUBS -0.06fF
C936 D.n790 VSUBS 0.61fF $ **FLOATING
C937 D.n792 VSUBS 0.26fF $ **FLOATING
C938 D.n793 VSUBS 0.31fF $ **FLOATING
C939 D.n794 VSUBS 0.75fF $ **FLOATING
C940 D.n795 VSUBS 0.44fF $ **FLOATING
C941 D.n796 VSUBS 0.25fF $ **FLOATING
C942 D.n797 VSUBS 2.09fF $ **FLOATING
C943 D.n798 VSUBS 1.75fF $ **FLOATING
C944 D.n799 VSUBS 2.36fF $ **FLOATING
C945 D.t462 VSUBS -0.06fF
C946 D.n800 VSUBS 0.61fF $ **FLOATING
C947 D.t475 VSUBS -0.02fF
C948 D.n801 VSUBS 0.20fF $ **FLOATING
C949 D.t268 VSUBS -0.02fF
C950 D.n803 VSUBS 0.20fF $ **FLOATING
C951 D.t524 VSUBS -0.06fF
C952 D.n804 VSUBS 0.61fF $ **FLOATING
C953 D.n806 VSUBS 0.26fF $ **FLOATING
C954 D.n807 VSUBS 0.31fF $ **FLOATING
C955 D.n808 VSUBS 0.75fF $ **FLOATING
C956 D.n809 VSUBS 0.44fF $ **FLOATING
C957 D.n810 VSUBS 0.25fF $ **FLOATING
C958 D.n811 VSUBS 2.09fF $ **FLOATING
C959 D.n812 VSUBS 1.75fF $ **FLOATING
C960 D.n813 VSUBS 2.36fF $ **FLOATING
C961 D.t605 VSUBS -0.06fF
C962 D.n814 VSUBS 0.61fF $ **FLOATING
C963 D.t4 VSUBS -0.02fF
C964 D.n815 VSUBS 0.20fF $ **FLOATING
C965 D.t406 VSUBS -0.02fF
C966 D.n817 VSUBS 0.20fF $ **FLOATING
C967 D.t63 VSUBS -0.06fF
C968 D.n818 VSUBS 0.61fF $ **FLOATING
C969 D.n820 VSUBS 0.26fF $ **FLOATING
C970 D.n821 VSUBS 0.31fF $ **FLOATING
C971 D.n822 VSUBS 0.75fF $ **FLOATING
C972 D.n823 VSUBS 0.44fF $ **FLOATING
C973 D.n824 VSUBS 0.25fF $ **FLOATING
C974 D.n825 VSUBS 2.09fF $ **FLOATING
C975 D.n826 VSUBS 1.75fF $ **FLOATING
C976 D.n827 VSUBS 2.36fF $ **FLOATING
C977 D.t123 VSUBS -0.06fF
C978 D.n828 VSUBS 0.61fF $ **FLOATING
C979 D.t136 VSUBS -0.02fF
C980 D.n829 VSUBS 0.20fF $ **FLOATING
C981 D.t542 VSUBS -0.02fF
C982 D.n831 VSUBS 0.20fF $ **FLOATING
C983 D.t204 VSUBS -0.06fF
C984 D.n832 VSUBS 0.61fF $ **FLOATING
C985 D.n834 VSUBS 0.26fF $ **FLOATING
C986 D.n835 VSUBS 0.31fF $ **FLOATING
C987 D.n836 VSUBS 0.75fF $ **FLOATING
C988 D.n837 VSUBS 0.44fF $ **FLOATING
C989 D.n838 VSUBS 0.25fF $ **FLOATING
C990 D.n839 VSUBS 2.09fF $ **FLOATING
C991 D.n840 VSUBS 1.75fF $ **FLOATING
C992 D.n841 VSUBS 2.36fF $ **FLOATING
C993 D.t318 VSUBS -0.06fF
C994 D.n842 VSUBS 0.61fF $ **FLOATING
C995 D.t286 VSUBS -0.02fF
C996 D.n843 VSUBS 0.20fF $ **FLOATING
C997 D.t75 VSUBS -0.02fF
C998 D.n845 VSUBS 0.20fF $ **FLOATING
C999 D.t339 VSUBS -0.06fF
C1000 D.n846 VSUBS 0.61fF $ **FLOATING
C1001 D.n848 VSUBS 0.26fF $ **FLOATING
C1002 D.n849 VSUBS 0.31fF $ **FLOATING
C1003 D.n850 VSUBS 0.75fF $ **FLOATING
C1004 D.n851 VSUBS 0.44fF $ **FLOATING
C1005 D.n852 VSUBS 0.25fF $ **FLOATING
C1006 D.n853 VSUBS 2.09fF $ **FLOATING
C1007 D.n854 VSUBS 1.75fF $ **FLOATING
C1008 D.n855 VSUBS 2.36fF $ **FLOATING
C1009 D.t467 VSUBS -0.06fF
C1010 D.n856 VSUBS 0.61fF $ **FLOATING
C1011 D.t482 VSUBS -0.02fF
C1012 D.n857 VSUBS 0.20fF $ **FLOATING
C1013 D.t272 VSUBS -0.02fF
C1014 D.n859 VSUBS 0.20fF $ **FLOATING
C1015 D.t527 VSUBS -0.06fF
C1016 D.n860 VSUBS 0.61fF $ **FLOATING
C1017 D.n862 VSUBS 0.26fF $ **FLOATING
C1018 D.n863 VSUBS 0.31fF $ **FLOATING
C1019 D.n864 VSUBS 0.75fF $ **FLOATING
C1020 D.n865 VSUBS 0.44fF $ **FLOATING
C1021 D.n866 VSUBS 0.25fF $ **FLOATING
C1022 D.n867 VSUBS 2.09fF $ **FLOATING
C1023 D.n868 VSUBS 1.69fF $ **FLOATING
C1024 D.n869 VSUBS 0.80fF $ **FLOATING
C1025 D.t410 VSUBS -0.02fF
C1026 D.n870 VSUBS 0.20fF $ **FLOATING
C1027 D.t68 VSUBS -0.01fF
C1028 D.n871 VSUBS 0.55fF $ **FLOATING
C1029 D.t611 VSUBS -0.02fF
C1030 D.n872 VSUBS 0.56fF $ **FLOATING
C1031 D.n873 VSUBS 9.31fF $ **FLOATING
C1032 D.n874 VSUBS 2.16fF $ **FLOATING
C1033 D.n875 VSUBS 0.83fF $ **FLOATING
C1034 D.n876 VSUBS 0.44fF $ **FLOATING
C1035 D.n877 VSUBS 2.31fF $ **FLOATING
C1036 D.n878 VSUBS 2.40fF $ **FLOATING
C1037 D.t186 VSUBS 0.00fF
C1038 D.t127 VSUBS -0.06fF
C1039 D.n879 VSUBS 0.25fF $ **FLOATING
C1040 D.n880 VSUBS 0.33fF $ **FLOATING
C1041 D.t356 VSUBS 0.00fF
C1042 D.n881 VSUBS 0.33fF $ **FLOATING
C1043 D.n882 VSUBS 10.45fF $ **FLOATING
C1044 D.n883 VSUBS 1.87fF $ **FLOATING
C1045 D.t459 VSUBS -0.06fF
C1046 D.n884 VSUBS 0.61fF $ **FLOATING
C1047 D.t474 VSUBS -0.02fF
C1048 D.n885 VSUBS 0.20fF $ **FLOATING
C1049 D.t293 VSUBS -0.02fF
C1050 D.n887 VSUBS 0.20fF $ **FLOATING
C1051 D.t519 VSUBS -0.06fF
C1052 D.n888 VSUBS 0.61fF $ **FLOATING
C1053 D.n890 VSUBS 0.41fF $ **FLOATING
C1054 D.n891 VSUBS 0.31fF $ **FLOATING
C1055 D.n892 VSUBS 1.33fF $ **FLOATING
C1056 D.n893 VSUBS 2.21fF $ **FLOATING
C1057 D.n894 VSUBS 2.03fF $ **FLOATING
C1058 D.n895 VSUBS 2.90fF $ **FLOATING
C1059 D.t603 VSUBS -0.06fF
C1060 D.n896 VSUBS 0.61fF $ **FLOATING
C1061 D.t2 VSUBS -0.02fF
C1062 D.n897 VSUBS 0.20fF $ **FLOATING
C1063 D.t404 VSUBS -0.02fF
C1064 D.n899 VSUBS 0.20fF $ **FLOATING
C1065 D.t60 VSUBS -0.06fF
C1066 D.n900 VSUBS 0.61fF $ **FLOATING
C1067 D.n902 VSUBS 0.26fF $ **FLOATING
C1068 D.n903 VSUBS 0.31fF $ **FLOATING
C1069 D.n904 VSUBS 0.75fF $ **FLOATING
C1070 D.n905 VSUBS 0.44fF $ **FLOATING
C1071 D.n906 VSUBS 0.25fF $ **FLOATING
C1072 D.n907 VSUBS 2.49fF $ **FLOATING
C1073 D.n908 VSUBS 1.75fF $ **FLOATING
C1074 D.n909 VSUBS 2.08fF $ **FLOATING
C1075 D.t119 VSUBS -0.06fF
C1076 D.n910 VSUBS 0.61fF $ **FLOATING
C1077 D.t133 VSUBS -0.02fF
C1078 D.n911 VSUBS 0.20fF $ **FLOATING
C1079 D.t539 VSUBS -0.02fF
C1080 D.n913 VSUBS 0.20fF $ **FLOATING
C1081 D.t202 VSUBS -0.06fF
C1082 D.n914 VSUBS 0.61fF $ **FLOATING
C1083 D.n916 VSUBS 0.26fF $ **FLOATING
C1084 D.n917 VSUBS 0.31fF $ **FLOATING
C1085 D.n918 VSUBS 0.75fF $ **FLOATING
C1086 D.n919 VSUBS 0.44fF $ **FLOATING
C1087 D.n920 VSUBS 0.25fF $ **FLOATING
C1088 D.n921 VSUBS 2.09fF $ **FLOATING
C1089 D.n922 VSUBS 1.75fF $ **FLOATING
C1090 D.n923 VSUBS 2.36fF $ **FLOATING
C1091 D.t277 VSUBS -0.06fF
C1092 D.n924 VSUBS 0.61fF $ **FLOATING
C1093 D.t284 VSUBS -0.02fF
C1094 D.n925 VSUBS 0.20fF $ **FLOATING
C1095 D.t73 VSUBS -0.02fF
C1096 D.n927 VSUBS 0.20fF $ **FLOATING
C1097 D.t335 VSUBS -0.06fF
C1098 D.n928 VSUBS 0.61fF $ **FLOATING
C1099 D.n930 VSUBS 0.26fF $ **FLOATING
C1100 D.n931 VSUBS 0.31fF $ **FLOATING
C1101 D.n932 VSUBS 0.75fF $ **FLOATING
C1102 D.n933 VSUBS 0.44fF $ **FLOATING
C1103 D.n934 VSUBS 0.25fF $ **FLOATING
C1104 D.n935 VSUBS 2.09fF $ **FLOATING
C1105 D.n936 VSUBS 1.75fF $ **FLOATING
C1106 D.n937 VSUBS 2.36fF $ **FLOATING
C1107 D.t412 VSUBS -0.06fF
C1108 D.n938 VSUBS 0.61fF $ **FLOATING
C1109 D.t425 VSUBS -0.02fF
C1110 D.n939 VSUBS 0.20fF $ **FLOATING
C1111 D.t214 VSUBS -0.02fF
C1112 D.n941 VSUBS 0.20fF $ **FLOATING
C1113 D.t485 VSUBS -0.06fF
C1114 D.n942 VSUBS 0.61fF $ **FLOATING
C1115 D.n944 VSUBS 0.26fF $ **FLOATING
C1116 D.n945 VSUBS 0.31fF $ **FLOATING
C1117 D.n946 VSUBS 0.75fF $ **FLOATING
C1118 D.n947 VSUBS 0.44fF $ **FLOATING
C1119 D.n948 VSUBS 0.25fF $ **FLOATING
C1120 D.n949 VSUBS 2.09fF $ **FLOATING
C1121 D.n950 VSUBS 1.75fF $ **FLOATING
C1122 D.n951 VSUBS 2.36fF $ **FLOATING
C1123 D.t548 VSUBS -0.06fF
C1124 D.n952 VSUBS 0.61fF $ **FLOATING
C1125 D.t560 VSUBS -0.02fF
C1126 D.n953 VSUBS 0.20fF $ **FLOATING
C1127 D.t350 VSUBS -0.02fF
C1128 D.n955 VSUBS 0.20fF $ **FLOATING
C1129 D.t9 VSUBS -0.06fF
C1130 D.n956 VSUBS 0.61fF $ **FLOATING
C1131 D.n958 VSUBS 0.26fF $ **FLOATING
C1132 D.n959 VSUBS 0.31fF $ **FLOATING
C1133 D.n960 VSUBS 0.75fF $ **FLOATING
C1134 D.n961 VSUBS 0.44fF $ **FLOATING
C1135 D.n962 VSUBS 0.25fF $ **FLOATING
C1136 D.n963 VSUBS 2.09fF $ **FLOATING
C1137 D.n964 VSUBS 1.69fF $ **FLOATING
C1138 D.n965 VSUBS 0.80fF $ **FLOATING
C1139 D.t494 VSUBS -0.02fF
C1140 D.n966 VSUBS 0.20fF $ **FLOATING
C1141 D.t146 VSUBS -0.01fF
C1142 D.n967 VSUBS 0.55fF $ **FLOATING
C1143 D.t124 VSUBS -0.02fF
C1144 D.n968 VSUBS 0.56fF $ **FLOATING
C1145 D.n969 VSUBS 9.31fF $ **FLOATING
C1146 D.n970 VSUBS 2.16fF $ **FLOATING
C1147 D.n971 VSUBS 0.83fF $ **FLOATING
C1148 D.n972 VSUBS 0.44fF $ **FLOATING
C1149 D.n973 VSUBS 2.31fF $ **FLOATING
C1150 D.n974 VSUBS 2.40fF $ **FLOATING
C1151 D.t534 VSUBS 0.00fF
C1152 D.t114 VSUBS -0.06fF
C1153 D.n975 VSUBS 0.25fF $ **FLOATING
C1154 D.n976 VSUBS 0.33fF $ **FLOATING
C1155 D.t131 VSUBS 0.00fF
C1156 D.n977 VSUBS 0.33fF $ **FLOATING
C1157 D.n978 VSUBS 10.45fF $ **FLOATING
C1158 D.n979 VSUBS 1.87fF $ **FLOATING
C1159 D.t274 VSUBS -0.06fF
C1160 D.n980 VSUBS 0.61fF $ **FLOATING
C1161 D.t283 VSUBS -0.02fF
C1162 D.n981 VSUBS 0.20fF $ **FLOATING
C1163 D.t72 VSUBS -0.02fF
C1164 D.n983 VSUBS 0.20fF $ **FLOATING
C1165 D.t332 VSUBS -0.06fF
C1166 D.n984 VSUBS 0.61fF $ **FLOATING
C1167 D.n986 VSUBS 0.41fF $ **FLOATING
C1168 D.n987 VSUBS 0.31fF $ **FLOATING
C1169 D.n988 VSUBS 1.33fF $ **FLOATING
C1170 D.n989 VSUBS 2.21fF $ **FLOATING
C1171 D.n990 VSUBS 2.03fF $ **FLOATING
C1172 D.n991 VSUBS 2.90fF $ **FLOATING
C1173 D.t409 VSUBS -0.06fF
C1174 D.n992 VSUBS 0.61fF $ **FLOATING
C1175 D.t421 VSUBS -0.02fF
C1176 D.n993 VSUBS 0.20fF $ **FLOATING
C1177 D.t212 VSUBS -0.02fF
C1178 D.n995 VSUBS 0.20fF $ **FLOATING
C1179 D.t481 VSUBS -0.06fF
C1180 D.n996 VSUBS 0.61fF $ **FLOATING
C1181 D.n998 VSUBS 0.26fF $ **FLOATING
C1182 D.n999 VSUBS 0.31fF $ **FLOATING
C1183 D.n1000 VSUBS 0.75fF $ **FLOATING
C1184 D.n1001 VSUBS 0.44fF $ **FLOATING
C1185 D.n1002 VSUBS 0.25fF $ **FLOATING
C1186 D.n1003 VSUBS 2.49fF $ **FLOATING
C1187 D.n1004 VSUBS 1.75fF $ **FLOATING
C1188 D.n1005 VSUBS 2.08fF $ **FLOATING
C1189 D.t545 VSUBS -0.06fF
C1190 D.n1006 VSUBS 0.61fF $ **FLOATING
C1191 D.t556 VSUBS -0.02fF
C1192 D.n1007 VSUBS 0.20fF $ **FLOATING
C1193 D.t346 VSUBS -0.02fF
C1194 D.n1009 VSUBS 0.20fF $ **FLOATING
C1195 D.t7 VSUBS -0.06fF
C1196 D.n1010 VSUBS 0.61fF $ **FLOATING
C1197 D.n1012 VSUBS 0.26fF $ **FLOATING
C1198 D.n1013 VSUBS 0.31fF $ **FLOATING
C1199 D.n1014 VSUBS 0.75fF $ **FLOATING
C1200 D.n1015 VSUBS 0.44fF $ **FLOATING
C1201 D.n1016 VSUBS 0.25fF $ **FLOATING
C1202 D.n1017 VSUBS 2.09fF $ **FLOATING
C1203 D.n1018 VSUBS 1.75fF $ **FLOATING
C1204 D.n1019 VSUBS 2.36fF $ **FLOATING
C1205 D.t78 VSUBS -0.06fF
C1206 D.n1020 VSUBS 0.61fF $ **FLOATING
C1207 D.t86 VSUBS -0.02fF
C1208 D.n1021 VSUBS 0.20fF $ **FLOATING
C1209 D.t492 VSUBS -0.02fF
C1210 D.n1023 VSUBS 0.20fF $ **FLOATING
C1211 D.t142 VSUBS -0.06fF
C1212 D.n1024 VSUBS 0.61fF $ **FLOATING
C1213 D.n1026 VSUBS 0.98fF $ **FLOATING
C1214 D.n1027 VSUBS 0.26fF $ **FLOATING
C1215 D.n1028 VSUBS 0.14fF $ **FLOATING
C1216 D.n1029 VSUBS 0.34fF $ **FLOATING
C1217 D.n1030 VSUBS 0.75fF $ **FLOATING
C1218 D.n1031 VSUBS 0.44fF $ **FLOATING
C1219 D.n1032 VSUBS 0.25fF $ **FLOATING
C1220 D.n1033 VSUBS 2.09fF $ **FLOATING
C1221 D.n1034 VSUBS 1.75fF $ **FLOATING
C1222 D.n1035 VSUBS 0.67fF $ **FLOATING
C1223 D.t28 VSUBS -0.02fF
C1224 D.n1036 VSUBS 0.20fF $ **FLOATING
C1225 D.t292 VSUBS -0.01fF
C1226 D.n1037 VSUBS 0.55fF $ **FLOATING
C1227 D.t222 VSUBS -0.02fF
C1228 D.n1038 VSUBS 0.56fF $ **FLOATING
C1229 D.n1039 VSUBS 9.31fF $ **FLOATING
C1230 D.n1040 VSUBS 2.16fF $ **FLOATING
C1231 D.n1041 VSUBS 2.40fF $ **FLOATING
C1232 D.n1042 VSUBS 2.37fF $ **FLOATING
C1233 D.n1043 VSUBS 19.11fF $ **FLOATING
C1234 D.n1044 VSUBS 2.16fF $ **FLOATING
C1235 D.t355 VSUBS -0.02fF
C1236 D.n1045 VSUBS 0.56fF $ **FLOATING
C1237 D.t152 VSUBS -0.02fF
C1238 D.n1046 VSUBS 0.20fF $ **FLOATING
C1239 D.t431 VSUBS -0.01fF
C1240 D.n1047 VSUBS 0.55fF $ **FLOATING
C1241 D.n1048 VSUBS 9.71fF $ **FLOATING
C1242 D.n1049 VSUBS 19.12fF $ **FLOATING
C1243 D.n1050 VSUBS 1.87fF $ **FLOATING
C1244 D.n1051 VSUBS 1.57fF $ **FLOATING
C1245 D.t544 VSUBS -0.06fF
C1246 D.n1052 VSUBS 0.25fF $ **FLOATING
C1247 D.t554 VSUBS 0.00fF
C1248 D.n1053 VSUBS 0.33fF $ **FLOATING
C1249 D.t344 VSUBS 0.00fF
C1250 D.n1054 VSUBS 0.33fF $ **FLOATING
C1251 D.n1055 VSUBS 11.55fF $ **FLOATING
C1252 D.n1056 VSUBS 1.71fF $ **FLOATING
C1253 D.n1057 VSUBS 2.50fF $ **FLOATING
C1254 D.t76 VSUBS -0.06fF
C1255 D.n1058 VSUBS 0.61fF $ **FLOATING
C1256 D.t85 VSUBS -0.02fF
C1257 D.n1059 VSUBS 0.20fF $ **FLOATING
C1258 D.t491 VSUBS -0.02fF
C1259 D.n1061 VSUBS 0.20fF $ **FLOATING
C1260 D.t139 VSUBS -0.06fF
C1261 D.n1062 VSUBS 0.61fF $ **FLOATING
C1262 D.n1064 VSUBS 1.85fF $ **FLOATING
C1263 D.n1065 VSUBS 2.74fF $ **FLOATING
C1264 D.n1066 VSUBS 2.67fF $ **FLOATING
C1265 D.t232 VSUBS -0.02fF
C1266 D.n1067 VSUBS 0.20fF $ **FLOATING
C1267 D.t219 VSUBS -0.06fF
C1268 D.n1068 VSUBS 0.61fF $ **FLOATING
C1269 D.t23 VSUBS -0.02fF
C1270 D.n1070 VSUBS 0.20fF $ **FLOATING
C1271 D.t289 VSUBS -0.06fF
C1272 D.n1071 VSUBS 0.61fF $ **FLOATING
C1273 D.n1073 VSUBS 2.36fF $ **FLOATING
C1274 D.n1074 VSUBS 1.69fF $ **FLOATING
C1275 D.n1075 VSUBS 1.37fF $ **FLOATING
C1276 D.n1076 VSUBS 2.20fF $ **FLOATING
C1277 D.n1077 VSUBS 4.41fF $ **FLOATING
C1278 D.t299 VSUBS -0.02fF
C1279 D.n1078 VSUBS 0.20fF $ **FLOATING
C1280 D.t563 VSUBS -0.01fF
C1281 D.n1079 VSUBS 0.55fF $ **FLOATING
C1282 D.t498 VSUBS -0.02fF
C1283 D.n1080 VSUBS 0.56fF $ **FLOATING
C1284 D.n1081 VSUBS 4.95fF $ **FLOATING
C1285 D.n1082 VSUBS 1.62fF $ **FLOATING
C1286 D.t352 VSUBS -0.06fF
C1287 D.n1083 VSUBS 0.25fF $ **FLOATING
C1288 D.t362 VSUBS 0.00fF
C1289 D.n1084 VSUBS 0.33fF $ **FLOATING
C1290 D.t150 VSUBS 0.00fF
C1291 D.n1085 VSUBS 0.33fF $ **FLOATING
C1292 D.n1086 VSUBS 10.85fF $ **FLOATING
C1293 D.n1087 VSUBS 5.06fF $ **FLOATING
C1294 D.n1088 VSUBS 16.73fF $ **FLOATING
C1295 D.n1089 VSUBS 8.10fF $ **FLOATING
C1296 D.n1090 VSUBS 8.06fF $ **FLOATING
C1297 D.n1091 VSUBS 8.06fF $ **FLOATING
C1298 D.n1092 VSUBS 8.06fF $ **FLOATING
C1299 D.n1093 VSUBS 8.06fF $ **FLOATING
C1300 D.n1094 VSUBS 8.06fF $ **FLOATING
C1301 D.n1095 VSUBS 9.06fF $ **FLOATING
C1302 D.n1096 VSUBS 0.13fF $ **FLOATING
C1303 D.n1097 VSUBS 0.70fF $ **FLOATING
C1304 D.n1098 VSUBS 4.84fF $ **FLOATING
C1305 D.n1099 VSUBS 0.24fF $ **FLOATING
C1306 D.t46 VSUBS 0.00fF
C1307 D.t535 VSUBS -0.06fF
C1308 D.n1100 VSUBS 0.25fF $ **FLOATING
C1309 D.n1101 VSUBS 0.33fF $ **FLOATING
C1310 D.t254 VSUBS 0.00fF
C1311 D.n1102 VSUBS 0.33fF $ **FLOATING
C1312 D.t253 VSUBS -0.02fF
C1313 D.n1103 VSUBS 0.20fF $ **FLOATING
C1314 D.t209 VSUBS -0.01fF
C1315 D.n1104 VSUBS 0.55fF $ **FLOATING
C1316 D.t74 VSUBS -0.02fF
C1317 D.n1105 VSUBS 0.56fF $ **FLOATING
C1318 D.n1106 VSUBS 11.93fF $ **FLOATING
C1319 D.n1107 VSUBS 4.77fF $ **FLOATING
C1320 D.n1108 VSUBS 2.16fF $ **FLOATING
C1321 D.n1109 VSUBS 3.87fF $ **FLOATING
C1322 D.n1110 VSUBS 0.09fF $ **FLOATING
C1323 D.n1111 VSUBS 0.90fF $ **FLOATING
C1324 D.n1112 VSUBS 1.78fF $ **FLOATING
C1325 D.n1113 VSUBS 3.16fF $ **FLOATING
C1326 D.t420 VSUBS -0.02fF
C1327 D.n1114 VSUBS 0.20fF $ **FLOATING
C1328 D.t311 VSUBS -0.06fF
C1329 D.n1115 VSUBS 0.61fF $ **FLOATING
C1330 D.t367 VSUBS -0.02fF
C1331 D.n1117 VSUBS 0.20fF $ **FLOATING
C1332 D.t47 VSUBS -0.06fF
C1333 D.n1118 VSUBS 0.61fF $ **FLOATING
C1334 D.n1120 VSUBS 1.42fF $ **FLOATING
C1335 D.n1121 VSUBS 1.67fF $ **FLOATING
C1336 D.t281 VSUBS -0.02fF
C1337 D.n1122 VSUBS 0.56fF $ **FLOATING
C1338 D.t89 VSUBS -0.02fF
C1339 D.n1123 VSUBS 0.20fF $ **FLOATING
C1340 D.t341 VSUBS -0.01fF
C1341 D.n1124 VSUBS 0.55fF $ **FLOATING
C1342 D.n1125 VSUBS 1.77fF $ **FLOATING
C1343 D.n1126 VSUBS 0.86fF $ **FLOATING
C1344 D.n1127 VSUBS 0.26fF $ **FLOATING
C1345 D.n1128 VSUBS 0.14fF $ **FLOATING
C1346 D.n1129 VSUBS 0.05fF $ **FLOATING
C1347 D.n1130 VSUBS 0.07fF $ **FLOATING
C1348 D.n1131 VSUBS 7.97fF $ **FLOATING
C1349 D.n1132 VSUBS 1.82fF $ **FLOATING
C1350 D.t207 VSUBS -0.02fF
C1351 D.n1133 VSUBS 0.20fF $ **FLOATING
C1352 D.n1134 VSUBS 0.01fF $ **FLOATING
C1353 D.t368 VSUBS -0.06fF
C1354 D.n1136 VSUBS 0.60fF $ **FLOATING
C1355 D.t536 VSUBS -0.06fF
C1356 D.n1138 VSUBS 0.61fF $ **FLOATING
C1357 D.t610 VSUBS -0.02fF
C1358 D.n1139 VSUBS 0.20fF $ **FLOATING
C1359 D.n1141 VSUBS 4.39fF $ **FLOATING
C1360 D.n1142 VSUBS 1.93fF $ **FLOATING
C1361 D.n1143 VSUBS 1.20fF $ **FLOATING
C1362 D.n1144 VSUBS 0.03fF $ **FLOATING
C1363 D.n1145 VSUBS 0.04fF $ **FLOATING
C1364 D.n1146 VSUBS 0.24fF $ **FLOATING
C1365 D.n1147 VSUBS 13.51fF $ **FLOATING
C1366 D.n1148 VSUBS 1.39fF $ **FLOATING
C1367 D.n1149 VSUBS 0.67fF $ **FLOATING
C1368 D.n1150 VSUBS 0.25fF $ **FLOATING
C1369 D.n1151 VSUBS 0.08fF $ **FLOATING
C1370 D.n1152 VSUBS 0.10fF $ **FLOATING
C1371 D.n1153 VSUBS 0.11fF $ **FLOATING
C1372 D.t132 VSUBS -0.06fF
C1373 D.n1154 VSUBS 0.25fF $ **FLOATING
C1374 D.t62 VSUBS 0.00fF
C1375 D.n1155 VSUBS 0.33fF $ **FLOATING
C1376 D.t461 VSUBS 0.00fF
C1377 D.n1156 VSUBS 0.33fF $ **FLOATING
C1378 D.n1157 VSUBS 16.87fF $ **FLOATING
C1379 D.n1158 VSUBS 1.91fF $ **FLOATING
C1380 D.n1159 VSUBS 2.16fF $ **FLOATING
C1381 D.n1160 VSUBS 1.36fF $ **FLOATING
C1382 D.n1161 VSUBS 17.07fF $ **FLOATING
C1383 D.n1162 VSUBS 0.09fF $ **FLOATING
C1384 D.n1163 VSUBS 1.77fF $ **FLOATING
C1385 D.t417 VSUBS -0.02fF
C1386 D.n1164 VSUBS 0.56fF $ **FLOATING
C1387 D.t138 VSUBS -0.02fF
C1388 D.n1165 VSUBS 0.20fF $ **FLOATING
C1389 D.t487 VSUBS -0.01fF
C1390 D.n1166 VSUBS 0.55fF $ **FLOATING
C1391 D.n1167 VSUBS 8.51fF $ **FLOATING
C1392 D.n1168 VSUBS 0.07fF $ **FLOATING
C1393 D.n1169 VSUBS 0.05fF $ **FLOATING
C1394 D.n1170 VSUBS 0.81fF $ **FLOATING
C1395 D.n1171 VSUBS 0.26fF $ **FLOATING
C1396 D.n1172 VSUBS 0.14fF $ **FLOATING
C1397 D.n1173 VSUBS 0.91fF $ **FLOATING
C1398 D.n1174 VSUBS 1.61fF $ **FLOATING
C1399 D.t218 VSUBS -0.02fF
C1400 D.n1175 VSUBS 0.20fF $ **FLOATING
C1401 D.t384 VSUBS -0.06fF
C1402 D.n1176 VSUBS 0.61fF $ **FLOATING
C1403 D.t426 VSUBS -0.02fF
C1404 D.n1178 VSUBS 0.20fF $ **FLOATING
C1405 D.t103 VSUBS -0.06fF
C1406 D.n1179 VSUBS 0.61fF $ **FLOATING
C1407 D.n1181 VSUBS 1.41fF $ **FLOATING
C1408 D.n1182 VSUBS 1.96fF $ **FLOATING
C1409 D.n1183 VSUBS 1.76fF $ **FLOATING
C1410 D.n1184 VSUBS 1.59fF $ **FLOATING
C1411 D.n1185 VSUBS 3.09fF $ **FLOATING
C1412 D.t572 VSUBS -0.06fF
C1413 D.n1186 VSUBS 0.61fF $ **FLOATING
C1414 D.t228 VSUBS -0.02fF
C1415 D.n1187 VSUBS 0.20fF $ **FLOATING
C1416 D.t17 VSUBS -0.02fF
C1417 D.n1189 VSUBS 0.20fF $ **FLOATING
C1418 D.t165 VSUBS -0.06fF
C1419 D.n1190 VSUBS 0.61fF $ **FLOATING
C1420 D.n1192 VSUBS 2.24fF $ **FLOATING
C1421 D.n1193 VSUBS 2.27fF $ **FLOATING
C1422 D.n1194 VSUBS 1.59fF $ **FLOATING
C1423 D.t233 VSUBS -0.02fF
C1424 D.n1195 VSUBS 0.20fF $ **FLOATING
C1425 D.t580 VSUBS -0.06fF
C1426 D.n1196 VSUBS 0.61fF $ **FLOATING
C1427 D.t25 VSUBS -0.02fF
C1428 D.n1198 VSUBS 0.20fF $ **FLOATING
C1429 D.t171 VSUBS -0.06fF
C1430 D.n1199 VSUBS 0.61fF $ **FLOATING
C1431 D.n1201 VSUBS 1.44fF $ **FLOATING
C1432 D.n1202 VSUBS 1.85fF $ **FLOATING
C1433 D.n1203 VSUBS 2.27fF $ **FLOATING
C1434 D.n1204 VSUBS 1.59fF $ **FLOATING
C1435 D.n1205 VSUBS 2.99fF $ **FLOATING
C1436 D.t345 VSUBS -0.06fF
C1437 D.n1206 VSUBS 0.61fF $ **FLOATING
C1438 D.t15 VSUBS -0.02fF
C1439 D.n1207 VSUBS 0.20fF $ **FLOATING
C1440 D.t415 VSUBS -0.02fF
C1441 D.n1209 VSUBS 0.20fF $ **FLOATING
C1442 D.t181 VSUBS -0.06fF
C1443 D.n1210 VSUBS 0.61fF $ **FLOATING
C1444 D.n1212 VSUBS 2.24fF $ **FLOATING
C1445 D.n1213 VSUBS 1.95fF $ **FLOATING
C1446 D.n1214 VSUBS 1.19fF $ **FLOATING
C1447 D.n1215 VSUBS 0.03fF $ **FLOATING
C1448 D.n1216 VSUBS 0.04fF $ **FLOATING
C1449 D.n1217 VSUBS 0.24fF $ **FLOATING
C1450 D.n1218 VSUBS 3.48fF $ **FLOATING
C1451 D.n1219 VSUBS 4.16fF $ **FLOATING
C1452 D.n1220 VSUBS 1.39fF $ **FLOATING
C1453 D.n1221 VSUBS 0.67fF $ **FLOATING
C1454 D.n1222 VSUBS 0.25fF $ **FLOATING
C1455 D.n1223 VSUBS 0.08fF $ **FLOATING
C1456 D.n1224 VSUBS 0.10fF $ **FLOATING
C1457 D.n1225 VSUBS 0.11fF $ **FLOATING
C1458 D.t555 VSUBS -0.06fF
C1459 D.n1226 VSUBS 0.25fF $ **FLOATING
C1460 D.t484 VSUBS 0.00fF
C1461 D.n1227 VSUBS 0.33fF $ **FLOATING
C1462 D.t276 VSUBS 0.00fF
C1463 D.n1228 VSUBS 0.33fF $ **FLOATING
C1464 D.n1229 VSUBS 0.24fF $ **FLOATING
C1465 D.n1230 VSUBS 0.04fF $ **FLOATING
C1466 D.n1231 VSUBS 0.22fF $ **FLOATING
C1467 D.n1232 VSUBS 0.18fF $ **FLOATING
C1468 D.n1233 VSUBS 1.24fF $ **FLOATING
C1469 D.n1234 VSUBS 0.65fF $ **FLOATING
C1470 D.n1235 VSUBS 0.10fF $ **FLOATING
C1471 D.n1236 VSUBS 0.10fF $ **FLOATING
C1472 D.n1237 VSUBS 0.57fF $ **FLOATING
C1473 D.n1238 VSUBS 2.09fF $ **FLOATING
C1474 D.n1239 VSUBS 1.34fF $ **FLOATING
C1475 D.n1240 VSUBS 8.16fF $ **FLOATING
C1476 D.n1241 VSUBS 0.09fF $ **FLOATING
C1477 D.n1242 VSUBS 2.27fF $ **FLOATING
C1478 D.n1243 VSUBS 0.91fF $ **FLOATING
C1479 D.n1244 VSUBS 1.76fF $ **FLOATING
C1480 D.t18 VSUBS -0.02fF
C1481 D.n1245 VSUBS 0.20fF $ **FLOATING
C1482 D.t452 VSUBS -0.06fF
C1483 D.n1246 VSUBS 0.61fF $ **FLOATING
C1484 D.t480 VSUBS -0.02fF
C1485 D.n1248 VSUBS 0.20fF $ **FLOATING
C1486 D.t176 VSUBS -0.06fF
C1487 D.n1249 VSUBS 0.61fF $ **FLOATING
C1488 D.n1251 VSUBS 1.41fF $ **FLOATING
C1489 D.n1252 VSUBS 1.78fF $ **FLOATING
C1490 D.t550 VSUBS -0.02fF
C1491 D.n1253 VSUBS 0.56fF $ **FLOATING
C1492 D.t199 VSUBS -0.02fF
C1493 D.n1254 VSUBS 0.20fF $ **FLOATING
C1494 D.t12 VSUBS -0.01fF
C1495 D.n1255 VSUBS 0.55fF $ **FLOATING
C1496 D.n1256 VSUBS 1.77fF $ **FLOATING
C1497 D.n1257 VSUBS 0.81fF $ **FLOATING
C1498 D.n1258 VSUBS 0.26fF $ **FLOATING
C1499 D.n1259 VSUBS 0.14fF $ **FLOATING
C1500 D.n1260 VSUBS 0.05fF $ **FLOATING
C1501 D.n1261 VSUBS 0.07fF $ **FLOATING
C1502 D.n1262 VSUBS 7.81fF $ **FLOATING
C1503 D.n1263 VSUBS 1.86fF $ **FLOATING
C1504 D.n1264 VSUBS 3.09fF $ **FLOATING
C1505 D.t370 VSUBS -0.06fF
C1506 D.n1265 VSUBS 0.61fF $ **FLOATING
C1507 D.t26 VSUBS -0.02fF
C1508 D.n1266 VSUBS 0.20fF $ **FLOATING
C1509 D.t423 VSUBS -0.02fF
C1510 D.n1268 VSUBS 0.20fF $ **FLOATING
C1511 D.t574 VSUBS -0.06fF
C1512 D.n1269 VSUBS 0.61fF $ **FLOATING
C1513 D.n1271 VSUBS 2.27fF $ **FLOATING
C1514 D.n1272 VSUBS 2.07fF $ **FLOATING
C1515 D.n1273 VSUBS 1.75fF $ **FLOATING
C1516 D.n1274 VSUBS 2.27fF $ **FLOATING
C1517 D.t31 VSUBS -0.02fF
C1518 D.n1275 VSUBS 0.20fF $ **FLOATING
C1519 D.t380 VSUBS -0.06fF
C1520 D.n1276 VSUBS 0.61fF $ **FLOATING
C1521 D.t432 VSUBS -0.02fF
C1522 D.n1278 VSUBS 0.20fF $ **FLOATING
C1523 D.t583 VSUBS -0.06fF
C1524 D.n1279 VSUBS 0.61fF $ **FLOATING
C1525 D.n1281 VSUBS 1.44fF $ **FLOATING
C1526 D.n1282 VSUBS 1.67fF $ **FLOATING
C1527 D.n1283 VSUBS 1.75fF $ **FLOATING
C1528 D.n1284 VSUBS 2.90fF $ **FLOATING
C1529 D.t386 VSUBS -0.06fF
C1530 D.n1285 VSUBS 0.61fF $ **FLOATING
C1531 D.t35 VSUBS -0.02fF
C1532 D.n1286 VSUBS 0.20fF $ **FLOATING
C1533 D.t436 VSUBS -0.02fF
C1534 D.n1288 VSUBS 0.20fF $ **FLOATING
C1535 D.t593 VSUBS -0.06fF
C1536 D.n1289 VSUBS 0.61fF $ **FLOATING
C1537 D.n1291 VSUBS 2.27fF $ **FLOATING
C1538 D.n1292 VSUBS 2.07fF $ **FLOATING
C1539 D.n1293 VSUBS 1.75fF $ **FLOATING
C1540 D.t41 VSUBS -0.02fF
C1541 D.n1294 VSUBS 0.20fF $ **FLOATING
C1542 D.t395 VSUBS -0.06fF
C1543 D.n1295 VSUBS 0.61fF $ **FLOATING
C1544 D.t441 VSUBS -0.02fF
C1545 D.n1297 VSUBS 0.20fF $ **FLOATING
C1546 D.t599 VSUBS -0.06fF
C1547 D.n1298 VSUBS 0.61fF $ **FLOATING
C1548 D.n1300 VSUBS 1.44fF $ **FLOATING
C1549 D.n1301 VSUBS 1.67fF $ **FLOATING
C1550 D.n1302 VSUBS 1.76fF $ **FLOATING
C1551 D.n1303 VSUBS 3.11fF $ **FLOATING
C1552 D.t151 VSUBS -0.06fF
C1553 D.n1304 VSUBS 0.61fF $ **FLOATING
C1554 D.t435 VSUBS -0.02fF
C1555 D.n1305 VSUBS 0.20fF $ **FLOATING
C1556 D.t227 VSUBS -0.02fF
C1557 D.n1307 VSUBS 0.20fF $ **FLOATING
C1558 D.t607 VSUBS -0.06fF
C1559 D.n1308 VSUBS 0.61fF $ **FLOATING
C1560 D.n1310 VSUBS 4.38fF $ **FLOATING
C1561 D.n1311 VSUBS 1.95fF $ **FLOATING
C1562 D.n1312 VSUBS 1.19fF $ **FLOATING
C1563 D.n1313 VSUBS 0.03fF $ **FLOATING
C1564 D.n1314 VSUBS 0.04fF $ **FLOATING
C1565 D.n1315 VSUBS 0.24fF $ **FLOATING
C1566 D.n1316 VSUBS 3.48fF $ **FLOATING
C1567 D.n1317 VSUBS 4.16fF $ **FLOATING
C1568 D.n1318 VSUBS 1.39fF $ **FLOATING
C1569 D.n1319 VSUBS 0.67fF $ **FLOATING
C1570 D.n1320 VSUBS 0.25fF $ **FLOATING
C1571 D.n1321 VSUBS 0.08fF $ **FLOATING
C1572 D.n1322 VSUBS 0.10fF $ **FLOATING
C1573 D.n1323 VSUBS 0.11fF $ **FLOATING
C1574 D.t363 VSUBS -0.06fF
C1575 D.n1324 VSUBS 0.25fF $ **FLOATING
C1576 D.t291 VSUBS 0.00fF
C1577 D.n1325 VSUBS 0.33fF $ **FLOATING
C1578 D.t77 VSUBS 0.00fF
C1579 D.n1326 VSUBS 0.33fF $ **FLOATING
C1580 D.n1327 VSUBS 4.43fF $ **FLOATING
C1581 D.n1328 VSUBS 0.93fF $ **FLOATING
C1582 D.n1329 VSUBS 3.17fF $ **FLOATING
C1583 D.n1330 VSUBS 8.07fF $ **FLOATING
C1584 D.n1331 VSUBS 1.91fF $ **FLOATING
C1585 D.n1332 VSUBS 2.16fF $ **FLOATING
C1586 D.n1333 VSUBS 1.36fF $ **FLOATING
C1587 D.n1334 VSUBS 8.16fF $ **FLOATING
C1588 D.n1335 VSUBS 0.09fF $ **FLOATING
C1589 D.n1336 VSUBS 1.77fF $ **FLOATING
C1590 D.t79 VSUBS -0.02fF
C1591 D.n1337 VSUBS 0.56fF $ **FLOATING
C1592 D.t252 VSUBS -0.02fF
C1593 D.n1338 VSUBS 0.20fF $ **FLOATING
C1594 D.t145 VSUBS -0.01fF
C1595 D.n1339 VSUBS 0.55fF $ **FLOATING
C1596 D.n1340 VSUBS 8.51fF $ **FLOATING
C1597 D.n1341 VSUBS 0.07fF $ **FLOATING
C1598 D.n1342 VSUBS 0.05fF $ **FLOATING
C1599 D.n1343 VSUBS 0.81fF $ **FLOATING
C1600 D.n1344 VSUBS 0.26fF $ **FLOATING
C1601 D.n1345 VSUBS 0.14fF $ **FLOATING
C1602 D.n1346 VSUBS 0.91fF $ **FLOATING
C1603 D.n1347 VSUBS 1.61fF $ **FLOATING
C1604 D.t424 VSUBS -0.02fF
C1605 D.n1348 VSUBS 0.20fF $ **FLOATING
C1606 D.t515 VSUBS -0.06fF
C1607 D.n1349 VSUBS 0.61fF $ **FLOATING
C1608 D.t521 VSUBS -0.02fF
C1609 D.n1351 VSUBS 0.20fF $ **FLOATING
C1610 D.t250 VSUBS -0.06fF
C1611 D.n1352 VSUBS 0.61fF $ **FLOATING
C1612 D.n1354 VSUBS 1.41fF $ **FLOATING
C1613 D.n1355 VSUBS 1.96fF $ **FLOATING
C1614 D.n1356 VSUBS 1.76fF $ **FLOATING
C1615 D.n1357 VSUBS 1.59fF $ **FLOATING
C1616 D.n1358 VSUBS 3.09fF $ **FLOATING
C1617 D.t167 VSUBS -0.06fF
C1618 D.n1359 VSUBS 0.61fF $ **FLOATING
C1619 D.t433 VSUBS -0.02fF
C1620 D.n1360 VSUBS 0.20fF $ **FLOATING
C1621 D.t220 VSUBS -0.02fF
C1622 D.n1362 VSUBS 0.20fF $ **FLOATING
C1623 D.t374 VSUBS -0.06fF
C1624 D.n1363 VSUBS 0.61fF $ **FLOATING
C1625 D.n1365 VSUBS 2.24fF $ **FLOATING
C1626 D.n1366 VSUBS 2.27fF $ **FLOATING
C1627 D.n1367 VSUBS 1.59fF $ **FLOATING
C1628 D.t437 VSUBS -0.02fF
C1629 D.n1368 VSUBS 0.20fF $ **FLOATING
C1630 D.t173 VSUBS -0.06fF
C1631 D.n1369 VSUBS 0.61fF $ **FLOATING
C1632 D.t230 VSUBS -0.02fF
C1633 D.n1371 VSUBS 0.20fF $ **FLOATING
C1634 D.t382 VSUBS -0.06fF
C1635 D.n1372 VSUBS 0.61fF $ **FLOATING
C1636 D.n1374 VSUBS 1.44fF $ **FLOATING
C1637 D.n1375 VSUBS 1.85fF $ **FLOATING
C1638 D.n1376 VSUBS 2.27fF $ **FLOATING
C1639 D.n1377 VSUBS 1.59fF $ **FLOATING
C1640 D.n1378 VSUBS 2.90fF $ **FLOATING
C1641 D.t184 VSUBS -0.06fF
C1642 D.n1379 VSUBS 0.61fF $ **FLOATING
C1643 D.t443 VSUBS -0.02fF
C1644 D.n1380 VSUBS 0.20fF $ **FLOATING
C1645 D.t235 VSUBS -0.02fF
C1646 D.n1382 VSUBS 0.20fF $ **FLOATING
C1647 D.t388 VSUBS -0.06fF
C1648 D.n1383 VSUBS 0.61fF $ **FLOATING
C1649 D.n1385 VSUBS 2.24fF $ **FLOATING
C1650 D.n1386 VSUBS 2.27fF $ **FLOATING
C1651 D.n1387 VSUBS 1.59fF $ **FLOATING
C1652 D.t449 VSUBS -0.02fF
C1653 D.n1388 VSUBS 0.20fF $ **FLOATING
C1654 D.t190 VSUBS -0.06fF
C1655 D.n1389 VSUBS 0.61fF $ **FLOATING
C1656 D.t239 VSUBS -0.02fF
C1657 D.n1391 VSUBS 0.20fF $ **FLOATING
C1658 D.t397 VSUBS -0.06fF
C1659 D.n1392 VSUBS 0.61fF $ **FLOATING
C1660 D.n1394 VSUBS 1.44fF $ **FLOATING
C1661 D.n1395 VSUBS 1.85fF $ **FLOATING
C1662 D.n1396 VSUBS 2.27fF $ **FLOATING
C1663 D.n1397 VSUBS 1.59fF $ **FLOATING
C1664 D.n1398 VSUBS 2.90fF $ **FLOATING
C1665 D.t197 VSUBS -0.06fF
C1666 D.n1399 VSUBS 0.61fF $ **FLOATING
C1667 D.t454 VSUBS -0.02fF
C1668 D.n1400 VSUBS 0.20fF $ **FLOATING
C1669 D.t246 VSUBS -0.02fF
C1670 D.n1402 VSUBS 0.20fF $ **FLOATING
C1671 D.t402 VSUBS -0.06fF
C1672 D.n1403 VSUBS 0.61fF $ **FLOATING
C1673 D.n1405 VSUBS 2.24fF $ **FLOATING
C1674 D.n1406 VSUBS 2.27fF $ **FLOATING
C1675 D.n1407 VSUBS 1.59fF $ **FLOATING
C1676 D.t463 VSUBS -0.02fF
C1677 D.n1408 VSUBS 0.20fF $ **FLOATING
C1678 D.t205 VSUBS -0.06fF
C1679 D.n1409 VSUBS 0.61fF $ **FLOATING
C1680 D.t256 VSUBS -0.02fF
C1681 D.n1411 VSUBS 0.20fF $ **FLOATING
C1682 D.t407 VSUBS -0.06fF
C1683 D.n1412 VSUBS 0.61fF $ **FLOATING
C1684 D.n1414 VSUBS 1.44fF $ **FLOATING
C1685 D.n1415 VSUBS 1.85fF $ **FLOATING
C1686 D.n1416 VSUBS 2.27fF $ **FLOATING
C1687 D.n1417 VSUBS 1.59fF $ **FLOATING
C1688 D.n1418 VSUBS 2.99fF $ **FLOATING
C1689 D.t577 VSUBS -0.06fF
C1690 D.n1419 VSUBS 0.61fF $ **FLOATING
C1691 D.t245 VSUBS -0.02fF
C1692 D.n1420 VSUBS 0.20fF $ **FLOATING
C1693 D.t34 VSUBS -0.02fF
C1694 D.n1422 VSUBS 0.20fF $ **FLOATING
C1695 D.t413 VSUBS -0.06fF
C1696 D.n1423 VSUBS 0.61fF $ **FLOATING
C1697 D.n1425 VSUBS 2.24fF $ **FLOATING
C1698 D.n1426 VSUBS 1.95fF $ **FLOATING
C1699 D.n1427 VSUBS 1.19fF $ **FLOATING
C1700 D.n1428 VSUBS 0.03fF $ **FLOATING
C1701 D.n1429 VSUBS 0.04fF $ **FLOATING
C1702 D.n1430 VSUBS 0.24fF $ **FLOATING
C1703 D.n1431 VSUBS 3.48fF $ **FLOATING
C1704 D.n1432 VSUBS 4.16fF $ **FLOATING
C1705 D.n1433 VSUBS 1.39fF $ **FLOATING
C1706 D.n1434 VSUBS 0.67fF $ **FLOATING
C1707 D.n1435 VSUBS 0.25fF $ **FLOATING
C1708 D.n1436 VSUBS 0.08fF $ **FLOATING
C1709 D.n1437 VSUBS 0.10fF $ **FLOATING
C1710 D.n1438 VSUBS 0.11fF $ **FLOATING
C1711 D.t177 VSUBS -0.06fF
C1712 D.n1439 VSUBS 0.25fF $ **FLOATING
C1713 D.t94 VSUBS 0.00fF
C1714 D.n1440 VSUBS 0.33fF $ **FLOATING
C1715 D.t500 VSUBS 0.00fF
C1716 D.n1441 VSUBS 0.33fF $ **FLOATING
C1717 D.n1442 VSUBS 0.24fF $ **FLOATING
C1718 D.n1443 VSUBS 0.04fF $ **FLOATING
C1719 D.n1444 VSUBS 0.22fF $ **FLOATING
C1720 D.n1445 VSUBS 0.18fF $ **FLOATING
C1721 D.n1446 VSUBS 1.24fF $ **FLOATING
C1722 D.n1447 VSUBS 0.65fF $ **FLOATING
C1723 D.n1448 VSUBS 0.10fF $ **FLOATING
C1724 D.n1449 VSUBS 0.10fF $ **FLOATING
C1725 D.n1450 VSUBS 0.57fF $ **FLOATING
C1726 D.n1451 VSUBS 2.09fF $ **FLOATING
C1727 D.n1452 VSUBS 1.34fF $ **FLOATING
C1728 D.n1453 VSUBS 8.16fF $ **FLOATING
C1729 D.n1454 VSUBS 0.09fF $ **FLOATING
C1730 D.n1455 VSUBS 2.27fF $ **FLOATING
C1731 D.n1456 VSUBS 0.91fF $ **FLOATING
C1732 D.n1457 VSUBS 1.76fF $ **FLOATING
C1733 D.t118 VSUBS -0.02fF
C1734 D.n1458 VSUBS 0.20fF $ **FLOATING
C1735 D.t589 VSUBS -0.06fF
C1736 D.n1459 VSUBS 0.61fF $ **FLOATING
C1737 D.t129 VSUBS -0.02fF
C1738 D.n1461 VSUBS 0.20fF $ **FLOATING
C1739 D.t97 VSUBS -0.06fF
C1740 D.n1462 VSUBS 0.61fF $ **FLOATING
C1741 D.n1464 VSUBS 1.41fF $ **FLOATING
C1742 D.n1465 VSUBS 1.78fF $ **FLOATING
C1743 D.t161 VSUBS -0.02fF
C1744 D.n1466 VSUBS 0.56fF $ **FLOATING
C1745 D.t473 VSUBS -0.02fF
C1746 D.n1467 VSUBS 0.20fF $ **FLOATING
C1747 D.t240 VSUBS -0.01fF
C1748 D.n1468 VSUBS 0.55fF $ **FLOATING
C1749 D.n1469 VSUBS 1.77fF $ **FLOATING
C1750 D.n1470 VSUBS 0.81fF $ **FLOATING
C1751 D.n1471 VSUBS 0.26fF $ **FLOATING
C1752 D.n1472 VSUBS 0.14fF $ **FLOATING
C1753 D.n1473 VSUBS 0.05fF $ **FLOATING
C1754 D.n1474 VSUBS 0.07fF $ **FLOATING
C1755 D.n1475 VSUBS 7.81fF $ **FLOATING
C1756 D.n1476 VSUBS 1.86fF $ **FLOATING
C1757 D.n1477 VSUBS 3.09fF $ **FLOATING
C1758 D.t576 VSUBS -0.06fF
C1759 D.n1478 VSUBS 0.61fF $ **FLOATING
C1760 D.t231 VSUBS -0.02fF
C1761 D.n1479 VSUBS 0.20fF $ **FLOATING
C1762 D.t20 VSUBS -0.02fF
C1763 D.n1481 VSUBS 0.20fF $ **FLOATING
C1764 D.t168 VSUBS -0.06fF
C1765 D.n1482 VSUBS 0.61fF $ **FLOATING
C1766 D.n1484 VSUBS 2.27fF $ **FLOATING
C1767 D.n1485 VSUBS 2.07fF $ **FLOATING
C1768 D.n1486 VSUBS 1.75fF $ **FLOATING
C1769 D.n1487 VSUBS 2.27fF $ **FLOATING
C1770 D.t236 VSUBS -0.02fF
C1771 D.n1488 VSUBS 0.20fF $ **FLOATING
C1772 D.t587 VSUBS -0.06fF
C1773 D.n1489 VSUBS 0.61fF $ **FLOATING
C1774 D.t27 VSUBS -0.02fF
C1775 D.n1491 VSUBS 0.20fF $ **FLOATING
C1776 D.t175 VSUBS -0.06fF
C1777 D.n1492 VSUBS 0.61fF $ **FLOATING
C1778 D.n1494 VSUBS 1.44fF $ **FLOATING
C1779 D.n1495 VSUBS 1.67fF $ **FLOATING
C1780 D.n1496 VSUBS 1.75fF $ **FLOATING
C1781 D.n1497 VSUBS 2.90fF $ **FLOATING
C1782 D.t596 VSUBS -0.06fF
C1783 D.n1498 VSUBS 0.61fF $ **FLOATING
C1784 D.t243 VSUBS -0.02fF
C1785 D.n1499 VSUBS 0.20fF $ **FLOATING
C1786 D.t33 VSUBS -0.02fF
C1787 D.n1501 VSUBS 0.20fF $ **FLOATING
C1788 D.t187 VSUBS -0.06fF
C1789 D.n1502 VSUBS 0.61fF $ **FLOATING
C1790 D.n1504 VSUBS 2.27fF $ **FLOATING
C1791 D.n1505 VSUBS 2.07fF $ **FLOATING
C1792 D.n1506 VSUBS 1.75fF $ **FLOATING
C1793 D.n1507 VSUBS 2.27fF $ **FLOATING
C1794 D.t247 VSUBS -0.02fF
C1795 D.n1508 VSUBS 0.20fF $ **FLOATING
C1796 D.t600 VSUBS -0.06fF
C1797 D.n1509 VSUBS 0.61fF $ **FLOATING
C1798 D.t36 VSUBS -0.02fF
C1799 D.n1511 VSUBS 0.20fF $ **FLOATING
C1800 D.t193 VSUBS -0.06fF
C1801 D.n1512 VSUBS 0.61fF $ **FLOATING
C1802 D.n1514 VSUBS 1.44fF $ **FLOATING
C1803 D.n1515 VSUBS 1.67fF $ **FLOATING
C1804 D.n1516 VSUBS 1.75fF $ **FLOATING
C1805 D.n1517 VSUBS 2.90fF $ **FLOATING
C1806 D.t608 VSUBS -0.06fF
C1807 D.n1518 VSUBS 0.61fF $ **FLOATING
C1808 D.t258 VSUBS -0.02fF
C1809 D.n1519 VSUBS 0.20fF $ **FLOATING
C1810 D.t42 VSUBS -0.02fF
C1811 D.n1521 VSUBS 0.20fF $ **FLOATING
C1812 D.t198 VSUBS -0.06fF
C1813 D.n1522 VSUBS 0.61fF $ **FLOATING
C1814 D.n1524 VSUBS 2.27fF $ **FLOATING
C1815 D.n1525 VSUBS 2.07fF $ **FLOATING
C1816 D.n1526 VSUBS 1.75fF $ **FLOATING
C1817 D.n1527 VSUBS 2.27fF $ **FLOATING
C1818 D.t264 VSUBS -0.02fF
C1819 D.n1528 VSUBS 0.20fF $ **FLOATING
C1820 D.t0 VSUBS -0.06fF
C1821 D.n1529 VSUBS 0.61fF $ **FLOATING
C1822 D.t50 VSUBS -0.02fF
C1823 D.n1531 VSUBS 0.20fF $ **FLOATING
C1824 D.t206 VSUBS -0.06fF
C1825 D.n1532 VSUBS 0.61fF $ **FLOATING
C1826 D.n1534 VSUBS 1.44fF $ **FLOATING
C1827 D.n1535 VSUBS 1.67fF $ **FLOATING
C1828 D.n1536 VSUBS 1.75fF $ **FLOATING
C1829 D.n1537 VSUBS 2.90fF $ **FLOATING
C1830 D.t5 VSUBS -0.06fF
C1831 D.n1538 VSUBS 0.61fF $ **FLOATING
C1832 D.t269 VSUBS -0.02fF
C1833 D.n1539 VSUBS 0.20fF $ **FLOATING
C1834 D.t54 VSUBS -0.02fF
C1835 D.n1541 VSUBS 0.20fF $ **FLOATING
C1836 D.t210 VSUBS -0.06fF
C1837 D.n1542 VSUBS 0.61fF $ **FLOATING
C1838 D.n1544 VSUBS 2.27fF $ **FLOATING
C1839 D.n1545 VSUBS 2.07fF $ **FLOATING
C1840 D.n1546 VSUBS 1.75fF $ **FLOATING
C1841 D.t278 VSUBS -0.02fF
C1842 D.n1547 VSUBS 0.20fF $ **FLOATING
C1843 D.t10 VSUBS -0.06fF
C1844 D.n1548 VSUBS 0.61fF $ **FLOATING
C1845 D.t64 VSUBS -0.02fF
C1846 D.n1550 VSUBS 0.20fF $ **FLOATING
C1847 D.t215 VSUBS -0.06fF
C1848 D.n1551 VSUBS 0.61fF $ **FLOATING
C1849 D.n1553 VSUBS 1.44fF $ **FLOATING
C1850 D.n1554 VSUBS 1.67fF $ **FLOATING
C1851 D.n1555 VSUBS 1.76fF $ **FLOATING
C1852 D.n1556 VSUBS 3.11fF $ **FLOATING
C1853 D.t392 VSUBS -0.06fF
C1854 D.n1557 VSUBS 0.61fF $ **FLOATING
C1855 D.t483 VSUBS -0.02fF
C1856 D.n1558 VSUBS 0.20fF $ **FLOATING
C1857 D.t453 VSUBS -0.02fF
C1858 D.n1560 VSUBS 0.20fF $ **FLOATING
C1859 D.t224 VSUBS -0.06fF
C1860 D.n1561 VSUBS 0.61fF $ **FLOATING
C1861 D.n1563 VSUBS 4.38fF $ **FLOATING
C1862 D.n1564 VSUBS 1.95fF $ **FLOATING
C1863 D.n1565 VSUBS 1.19fF $ **FLOATING
C1864 D.n1566 VSUBS 0.03fF $ **FLOATING
C1865 D.n1567 VSUBS 0.04fF $ **FLOATING
C1866 D.n1568 VSUBS 0.24fF $ **FLOATING
C1867 D.n1569 VSUBS 3.48fF $ **FLOATING
C1868 D.n1570 VSUBS 4.16fF $ **FLOATING
C1869 D.n1571 VSUBS 1.39fF $ **FLOATING
C1870 D.n1572 VSUBS 0.67fF $ **FLOATING
C1871 D.n1573 VSUBS 0.25fF $ **FLOATING
C1872 D.n1574 VSUBS 0.08fF $ **FLOATING
C1873 D.n1575 VSUBS 0.10fF $ **FLOATING
C1874 D.n1576 VSUBS 0.11fF $ **FLOATING
C1875 D.t19 VSUBS -0.06fF
C1876 D.n1577 VSUBS 0.25fF $ **FLOATING
C1877 D.t349 VSUBS 0.00fF
C1878 D.n1578 VSUBS 0.33fF $ **FLOATING
C1879 D.t169 VSUBS 0.00fF
C1880 D.n1579 VSUBS 0.33fF $ **FLOATING
C1881 D.n1580 VSUBS 4.43fF $ **FLOATING
C1882 D.n1581 VSUBS 0.93fF $ **FLOATING
C1883 D.n1582 VSUBS 3.17fF $ **FLOATING
C1884 D.n1583 VSUBS 8.07fF $ **FLOATING
C1885 D.n1584 VSUBS 1.91fF $ **FLOATING
C1886 D.n1585 VSUBS 2.16fF $ **FLOATING
C1887 D.n1586 VSUBS 1.36fF $ **FLOATING
C1888 D.n1587 VSUBS 8.16fF $ **FLOATING
C1889 D.n1588 VSUBS 0.09fF $ **FLOATING
C1890 D.n1589 VSUBS 1.77fF $ **FLOATING
C1891 D.t307 VSUBS -0.02fF
C1892 D.n1590 VSUBS 0.56fF $ **FLOATING
C1893 D.t516 VSUBS -0.02fF
C1894 D.n1591 VSUBS 0.20fF $ **FLOATING
C1895 D.t375 VSUBS -0.01fF
C1896 D.n1592 VSUBS 0.55fF $ **FLOATING
C1897 D.n1593 VSUBS 8.51fF $ **FLOATING
C1898 D.n1594 VSUBS 0.07fF $ **FLOATING
C1899 D.n1595 VSUBS 0.05fF $ **FLOATING
C1900 D.n1596 VSUBS 0.81fF $ **FLOATING
C1901 D.n1597 VSUBS 0.26fF $ **FLOATING
C1902 D.n1598 VSUBS 0.14fF $ **FLOATING
C1903 D.n1599 VSUBS 0.91fF $ **FLOATING
C1904 D.n1600 VSUBS 1.61fF $ **FLOATING
C1905 D.t532 VSUBS -0.02fF
C1906 D.n1601 VSUBS 0.20fF $ **FLOATING
C1907 D.t444 VSUBS -0.06fF
C1908 D.n1602 VSUBS 0.61fF $ **FLOATING
C1909 D.t194 VSUBS -0.02fF
C1910 D.n1604 VSUBS 0.20fF $ **FLOATING
C1911 D.t164 VSUBS -0.06fF
C1912 D.n1605 VSUBS 0.61fF $ **FLOATING
C1913 D.n1607 VSUBS 1.41fF $ **FLOATING
C1914 D.n1608 VSUBS 1.96fF $ **FLOATING
C1915 D.n1609 VSUBS 1.76fF $ **FLOATING
C1916 D.n1610 VSUBS 1.59fF $ **FLOATING
C1917 D.n1611 VSUBS 3.09fF $ **FLOATING
C1918 D.t285 VSUBS -0.06fF
C1919 D.n1612 VSUBS 0.61fF $ **FLOATING
C1920 D.t540 VSUBS -0.02fF
C1921 D.n1613 VSUBS 0.20fF $ **FLOATING
C1922 D.t328 VSUBS -0.02fF
C1923 D.n1615 VSUBS 0.20fF $ **FLOATING
C1924 D.t489 VSUBS -0.06fF
C1925 D.n1616 VSUBS 0.61fF $ **FLOATING
C1926 D.n1618 VSUBS 2.24fF $ **FLOATING
C1927 D.n1619 VSUBS 2.27fF $ **FLOATING
C1928 D.n1620 VSUBS 1.59fF $ **FLOATING
C1929 D.t546 VSUBS -0.02fF
C1930 D.n1621 VSUBS 0.20fF $ **FLOATING
C1931 D.t383 VSUBS -0.06fF
C1932 D.n1622 VSUBS 0.61fF $ **FLOATING
C1933 D.t337 VSUBS -0.02fF
C1934 D.n1624 VSUBS 0.20fF $ **FLOATING
C1935 D.t493 VSUBS -0.06fF
C1936 D.n1625 VSUBS 0.61fF $ **FLOATING
C1937 D.n1627 VSUBS 1.44fF $ **FLOATING
C1938 D.n1628 VSUBS 1.85fF $ **FLOATING
C1939 D.n1629 VSUBS 2.27fF $ **FLOATING
C1940 D.n1630 VSUBS 1.59fF $ **FLOATING
C1941 D.n1631 VSUBS 2.90fF $ **FLOATING
C1942 D.t390 VSUBS -0.06fF
C1943 D.n1632 VSUBS 0.61fF $ **FLOATING
C1944 D.t38 VSUBS -0.02fF
C1945 D.n1633 VSUBS 0.20fF $ **FLOATING
C1946 D.t439 VSUBS -0.02fF
C1947 D.n1635 VSUBS 0.20fF $ **FLOATING
C1948 D.t597 VSUBS -0.06fF
C1949 D.n1636 VSUBS 0.61fF $ **FLOATING
C1950 D.n1638 VSUBS 2.24fF $ **FLOATING
C1951 D.n1639 VSUBS 2.27fF $ **FLOATING
C1952 D.n1640 VSUBS 1.59fF $ **FLOATING
C1953 D.t44 VSUBS -0.02fF
C1954 D.n1641 VSUBS 0.20fF $ **FLOATING
C1955 D.t398 VSUBS -0.06fF
C1956 D.n1642 VSUBS 0.61fF $ **FLOATING
C1957 D.t445 VSUBS -0.02fF
C1958 D.n1644 VSUBS 0.20fF $ **FLOATING
C1959 D.t602 VSUBS -0.06fF
C1960 D.n1645 VSUBS 0.61fF $ **FLOATING
C1961 D.n1647 VSUBS 1.44fF $ **FLOATING
C1962 D.n1648 VSUBS 1.85fF $ **FLOATING
C1963 D.n1649 VSUBS 2.27fF $ **FLOATING
C1964 D.n1650 VSUBS 1.59fF $ **FLOATING
C1965 D.n1651 VSUBS 2.90fF $ **FLOATING
C1966 D.t403 VSUBS -0.06fF
C1967 D.n1652 VSUBS 0.61fF $ **FLOATING
C1968 D.t51 VSUBS -0.02fF
C1969 D.n1653 VSUBS 0.20fF $ **FLOATING
C1970 D.t451 VSUBS -0.02fF
C1971 D.n1655 VSUBS 0.20fF $ **FLOATING
C1972 D.t609 VSUBS -0.06fF
C1973 D.n1656 VSUBS 0.61fF $ **FLOATING
C1974 D.n1658 VSUBS 2.24fF $ **FLOATING
C1975 D.n1659 VSUBS 2.27fF $ **FLOATING
C1976 D.n1660 VSUBS 1.59fF $ **FLOATING
C1977 D.t57 VSUBS -0.02fF
C1978 D.n1661 VSUBS 0.20fF $ **FLOATING
C1979 D.t408 VSUBS -0.06fF
C1980 D.n1662 VSUBS 0.61fF $ **FLOATING
C1981 D.t455 VSUBS -0.02fF
C1982 D.n1664 VSUBS 0.20fF $ **FLOATING
C1983 D.t1 VSUBS -0.06fF
C1984 D.n1665 VSUBS 0.61fF $ **FLOATING
C1985 D.n1667 VSUBS 1.44fF $ **FLOATING
C1986 D.n1668 VSUBS 1.85fF $ **FLOATING
C1987 D.n1669 VSUBS 2.27fF $ **FLOATING
C1988 D.n1670 VSUBS 1.59fF $ **FLOATING
C1989 D.n1671 VSUBS 2.90fF $ **FLOATING
C1990 D.t414 VSUBS -0.06fF
C1991 D.n1672 VSUBS 0.61fF $ **FLOATING
C1992 D.t66 VSUBS -0.02fF
C1993 D.n1673 VSUBS 0.20fF $ **FLOATING
C1994 D.t465 VSUBS -0.02fF
C1995 D.n1675 VSUBS 0.20fF $ **FLOATING
C1996 D.t6 VSUBS -0.06fF
C1997 D.n1676 VSUBS 0.61fF $ **FLOATING
C1998 D.n1678 VSUBS 2.24fF $ **FLOATING
C1999 D.n1679 VSUBS 2.27fF $ **FLOATING
C2000 D.n1680 VSUBS 1.59fF $ **FLOATING
C2001 D.t70 VSUBS -0.02fF
C2002 D.n1681 VSUBS 0.20fF $ **FLOATING
C2003 D.t418 VSUBS -0.06fF
C2004 D.n1682 VSUBS 0.61fF $ **FLOATING
C2005 D.t471 VSUBS -0.02fF
C2006 D.n1684 VSUBS 0.20fF $ **FLOATING
C2007 D.t11 VSUBS -0.06fF
C2008 D.n1685 VSUBS 0.61fF $ **FLOATING
C2009 D.n1687 VSUBS 1.44fF $ **FLOATING
C2010 D.n1688 VSUBS 1.85fF $ **FLOATING
C2011 D.n1689 VSUBS 2.27fF $ **FLOATING
C2012 D.n1690 VSUBS 1.59fF $ **FLOATING
C2013 D.n1691 VSUBS 2.90fF $ **FLOATING
C2014 D.t427 VSUBS -0.06fF
C2015 D.n1692 VSUBS 0.61fF $ **FLOATING
C2016 D.t53 VSUBS -0.02fF
C2017 D.n1693 VSUBS 0.20fF $ **FLOATING
C2018 D.t476 VSUBS -0.02fF
C2019 D.n1695 VSUBS 0.20fF $ **FLOATING
C2020 D.t21 VSUBS -0.06fF
C2021 D.n1696 VSUBS 0.61fF $ **FLOATING
C2022 D.n1698 VSUBS 2.24fF $ **FLOATING
C2023 D.n1699 VSUBS 2.27fF $ **FLOATING
C2024 D.n1700 VSUBS 1.59fF $ **FLOATING
C2025 D.t154 VSUBS -0.02fF
C2026 D.n1701 VSUBS 0.20fF $ **FLOATING
C2027 D.t141 VSUBS -0.06fF
C2028 D.n1702 VSUBS 0.61fF $ **FLOATING
C2029 D.t598 VSUBS -0.02fF
C2030 D.n1704 VSUBS 0.20fF $ **FLOATING
C2031 D.t221 VSUBS -0.06fF
C2032 D.n1705 VSUBS 0.61fF $ **FLOATING
C2033 D.n1707 VSUBS 1.44fF $ **FLOATING
C2034 D.n1708 VSUBS 1.85fF $ **FLOATING
C2035 D.n1709 VSUBS 2.27fF $ **FLOATING
C2036 D.n1710 VSUBS 1.59fF $ **FLOATING
C2037 D.n1711 VSUBS 2.99fF $ **FLOATING
C2038 D.t229 VSUBS -0.06fF
C2039 D.n1712 VSUBS 0.61fF $ **FLOATING
C2040 D.t262 VSUBS -0.02fF
C2041 D.n1713 VSUBS 0.20fF $ **FLOATING
C2042 D.t48 VSUBS -0.02fF
C2043 D.n1715 VSUBS 0.20fF $ **FLOATING
C2044 D.t358 VSUBS -0.06fF
C2045 D.n1716 VSUBS 0.61fF $ **FLOATING
C2046 D.n1718 VSUBS 2.24fF $ **FLOATING
C2047 D.n1719 VSUBS 1.95fF $ **FLOATING
C2048 D.n1720 VSUBS 1.19fF $ **FLOATING
C2049 D.n1721 VSUBS 0.03fF $ **FLOATING
C2050 D.n1722 VSUBS 0.04fF $ **FLOATING
C2051 D.n1723 VSUBS 0.24fF $ **FLOATING
C2052 D.n1724 VSUBS 3.48fF $ **FLOATING
C2053 D.n1725 VSUBS 4.16fF $ **FLOATING
C2054 D.n1726 VSUBS 1.39fF $ **FLOATING
C2055 D.n1727 VSUBS 0.67fF $ **FLOATING
C2056 D.n1728 VSUBS 0.25fF $ **FLOATING
C2057 D.n1729 VSUBS 0.08fF $ **FLOATING
C2058 D.n1730 VSUBS 0.10fF $ **FLOATING
C2059 D.n1731 VSUBS 0.11fF $ **FLOATING
C2060 D.t438 VSUBS -0.06fF
C2061 D.n1732 VSUBS 0.25fF $ **FLOATING
C2062 D.t156 VSUBS 0.00fF
C2063 D.n1733 VSUBS 0.33fF $ **FLOATING
C2064 D.t559 VSUBS 0.00fF
C2065 D.n1734 VSUBS 0.33fF $ **FLOATING
C2066 D.n1735 VSUBS 0.24fF $ **FLOATING
C2067 D.n1736 VSUBS 0.04fF $ **FLOATING
C2068 D.n1737 VSUBS 0.22fF $ **FLOATING
C2069 D.n1738 VSUBS 0.18fF $ **FLOATING
C2070 D.n1739 VSUBS 1.24fF $ **FLOATING
C2071 D.n1740 VSUBS 0.65fF $ **FLOATING
C2072 D.n1741 VSUBS 0.10fF $ **FLOATING
C2073 D.n1742 VSUBS 0.10fF $ **FLOATING
C2074 D.n1743 VSUBS 0.57fF $ **FLOATING
C2075 D.n1744 VSUBS 2.09fF $ **FLOATING
C2076 D.n1745 VSUBS 1.34fF $ **FLOATING
C2077 D.n1746 VSUBS 8.16fF $ **FLOATING
C2078 D.n1747 VSUBS 0.09fF $ **FLOATING
C2079 D.n1748 VSUBS 2.27fF $ **FLOATING
C2080 D.n1749 VSUBS 0.91fF $ **FLOATING
C2081 D.n1750 VSUBS 1.76fF $ **FLOATING
C2082 D.t329 VSUBS -0.02fF
C2083 D.n1751 VSUBS 0.20fF $ **FLOATING
C2084 D.t506 VSUBS -0.06fF
C2085 D.n1752 VSUBS 0.61fF $ **FLOATING
C2086 D.t244 VSUBS -0.02fF
C2087 D.n1754 VSUBS 0.20fF $ **FLOATING
C2088 D.t241 VSUBS -0.06fF
C2089 D.n1755 VSUBS 0.61fF $ **FLOATING
C2090 D.n1757 VSUBS 1.41fF $ **FLOATING
C2091 D.n1758 VSUBS 1.78fF $ **FLOATING
C2092 D.t447 VSUBS -0.02fF
C2093 D.n1759 VSUBS 0.56fF $ **FLOATING
C2094 D.t569 VSUBS -0.02fF
C2095 D.n1760 VSUBS 0.20fF $ **FLOATING
C2096 D.t512 VSUBS -0.01fF
C2097 D.n1761 VSUBS 0.55fF $ **FLOATING
C2098 D.n1762 VSUBS 1.77fF $ **FLOATING
C2099 D.n1763 VSUBS 0.81fF $ **FLOATING
C2100 D.n1764 VSUBS 0.26fF $ **FLOATING
C2101 D.n1765 VSUBS 0.14fF $ **FLOATING
C2102 D.n1766 VSUBS 0.05fF $ **FLOATING
C2103 D.n1767 VSUBS 0.07fF $ **FLOATING
C2104 D.n1768 VSUBS 7.81fF $ **FLOATING
C2105 D.n1769 VSUBS 1.86fF $ **FLOATING
C2106 D.n1770 VSUBS 3.09fF $ **FLOATING
C2107 D.t80 VSUBS -0.06fF
C2108 D.n1771 VSUBS 0.61fF $ **FLOATING
C2109 D.t338 VSUBS -0.02fF
C2110 D.n1772 VSUBS 0.20fF $ **FLOATING
C2111 D.t120 VSUBS -0.02fF
C2112 D.n1774 VSUBS 0.20fF $ **FLOATING
C2113 D.t287 VSUBS -0.06fF
C2114 D.n1775 VSUBS 0.61fF $ **FLOATING
C2115 D.n1777 VSUBS 2.27fF $ **FLOATING
C2116 D.n1778 VSUBS 2.07fF $ **FLOATING
C2117 D.n1779 VSUBS 1.75fF $ **FLOATING
C2118 D.n1780 VSUBS 2.27fF $ **FLOATING
C2119 D.t342 VSUBS -0.02fF
C2120 D.n1781 VSUBS 0.20fF $ **FLOATING
C2121 D.t83 VSUBS -0.06fF
C2122 D.n1782 VSUBS 0.61fF $ **FLOATING
C2123 D.t128 VSUBS -0.02fF
C2124 D.n1784 VSUBS 0.20fF $ **FLOATING
C2125 D.t294 VSUBS -0.06fF
C2126 D.n1785 VSUBS 0.61fF $ **FLOATING
C2127 D.n1787 VSUBS 1.44fF $ **FLOATING
C2128 D.n1788 VSUBS 1.67fF $ **FLOATING
C2129 D.n1789 VSUBS 1.75fF $ **FLOATING
C2130 D.n1790 VSUBS 2.90fF $ **FLOATING
C2131 D.t88 VSUBS -0.06fF
C2132 D.n1791 VSUBS 0.61fF $ **FLOATING
C2133 D.t347 VSUBS -0.02fF
C2134 D.n1792 VSUBS 0.20fF $ **FLOATING
C2135 D.t134 VSUBS -0.02fF
C2136 D.n1794 VSUBS 0.20fF $ **FLOATING
C2137 D.t297 VSUBS -0.06fF
C2138 D.n1795 VSUBS 0.61fF $ **FLOATING
C2139 D.n1797 VSUBS 2.27fF $ **FLOATING
C2140 D.n1798 VSUBS 2.07fF $ **FLOATING
C2141 D.n1799 VSUBS 1.75fF $ **FLOATING
C2142 D.n1800 VSUBS 2.27fF $ **FLOATING
C2143 D.t354 VSUBS -0.02fF
C2144 D.n1801 VSUBS 0.20fF $ **FLOATING
C2145 D.t195 VSUBS -0.06fF
C2146 D.n1802 VSUBS 0.61fF $ **FLOATING
C2147 D.t140 VSUBS -0.02fF
C2148 D.n1804 VSUBS 0.20fF $ **FLOATING
C2149 D.t302 VSUBS -0.06fF
C2150 D.n1805 VSUBS 0.61fF $ **FLOATING
C2151 D.n1807 VSUBS 1.44fF $ **FLOATING
C2152 D.n1808 VSUBS 1.67fF $ **FLOATING
C2153 D.n1809 VSUBS 1.75fF $ **FLOATING
C2154 D.n1810 VSUBS 2.90fF $ **FLOATING
C2155 D.t201 VSUBS -0.06fF
C2156 D.n1811 VSUBS 0.61fF $ **FLOATING
C2157 D.t457 VSUBS -0.02fF
C2158 D.n1812 VSUBS 0.20fF $ **FLOATING
C2159 D.t249 VSUBS -0.02fF
C2160 D.n1814 VSUBS 0.20fF $ **FLOATING
C2161 D.t405 VSUBS -0.06fF
C2162 D.n1815 VSUBS 0.61fF $ **FLOATING
C2163 D.n1817 VSUBS 2.27fF $ **FLOATING
C2164 D.n1818 VSUBS 2.07fF $ **FLOATING
C2165 D.n1819 VSUBS 1.75fF $ **FLOATING
C2166 D.n1820 VSUBS 2.27fF $ **FLOATING
C2167 D.t466 VSUBS -0.02fF
C2168 D.n1821 VSUBS 0.20fF $ **FLOATING
C2169 D.t208 VSUBS -0.06fF
C2170 D.n1822 VSUBS 0.61fF $ **FLOATING
C2171 D.t260 VSUBS -0.02fF
C2172 D.n1824 VSUBS 0.20fF $ **FLOATING
C2173 D.t411 VSUBS -0.06fF
C2174 D.n1825 VSUBS 0.61fF $ **FLOATING
C2175 D.n1827 VSUBS 1.44fF $ **FLOATING
C2176 D.n1828 VSUBS 1.67fF $ **FLOATING
C2177 D.n1829 VSUBS 1.75fF $ **FLOATING
C2178 D.n1830 VSUBS 2.90fF $ **FLOATING
C2179 D.t211 VSUBS -0.06fF
C2180 D.n1831 VSUBS 0.61fF $ **FLOATING
C2181 D.t472 VSUBS -0.02fF
C2182 D.n1832 VSUBS 0.20fF $ **FLOATING
C2183 D.t267 VSUBS -0.02fF
C2184 D.n1834 VSUBS 0.20fF $ **FLOATING
C2185 D.t416 VSUBS -0.06fF
C2186 D.n1835 VSUBS 0.61fF $ **FLOATING
C2187 D.n1837 VSUBS 2.27fF $ **FLOATING
C2188 D.n1838 VSUBS 2.07fF $ **FLOATING
C2189 D.n1839 VSUBS 1.75fF $ **FLOATING
C2190 D.n1840 VSUBS 2.27fF $ **FLOATING
C2191 D.t477 VSUBS -0.02fF
C2192 D.n1841 VSUBS 0.20fF $ **FLOATING
C2193 D.t216 VSUBS -0.06fF
C2194 D.n1842 VSUBS 0.61fF $ **FLOATING
C2195 D.t271 VSUBS -0.02fF
C2196 D.n1844 VSUBS 0.20fF $ **FLOATING
C2197 D.t419 VSUBS -0.06fF
C2198 D.n1845 VSUBS 0.61fF $ **FLOATING
C2199 D.n1847 VSUBS 1.44fF $ **FLOATING
C2200 D.n1848 VSUBS 1.67fF $ **FLOATING
C2201 D.n1849 VSUBS 1.75fF $ **FLOATING
C2202 D.n1850 VSUBS 2.90fF $ **FLOATING
C2203 D.t225 VSUBS -0.06fF
C2204 D.n1851 VSUBS 0.61fF $ **FLOATING
C2205 D.t192 VSUBS -0.02fF
C2206 D.n1852 VSUBS 0.20fF $ **FLOATING
C2207 D.t279 VSUBS -0.02fF
C2208 D.n1854 VSUBS 0.20fF $ **FLOATING
C2209 D.t428 VSUBS -0.06fF
C2210 D.n1855 VSUBS 0.61fF $ **FLOATING
C2211 D.n1857 VSUBS 2.27fF $ **FLOATING
C2212 D.n1858 VSUBS 2.07fF $ **FLOATING
C2213 D.n1859 VSUBS 1.75fF $ **FLOATING
C2214 D.n1860 VSUBS 2.27fF $ **FLOATING
C2215 D.t300 VSUBS -0.02fF
C2216 D.n1861 VSUBS 0.20fF $ **FLOATING
C2217 D.t290 VSUBS -0.06fF
C2218 D.n1862 VSUBS 0.61fF $ **FLOATING
C2219 D.t110 VSUBS -0.02fF
C2220 D.n1864 VSUBS 0.20fF $ **FLOATING
C2221 D.t353 VSUBS -0.06fF
C2222 D.n1865 VSUBS 0.61fF $ **FLOATING
C2223 D.n1867 VSUBS 1.44fF $ **FLOATING
C2224 D.n1868 VSUBS 1.67fF $ **FLOATING
C2225 D.n1869 VSUBS 1.75fF $ **FLOATING
C2226 D.n1870 VSUBS 2.90fF $ **FLOATING
C2227 D.t434 VSUBS -0.06fF
C2228 D.n1871 VSUBS 0.61fF $ **FLOATING
C2229 D.t442 VSUBS -0.02fF
C2230 D.n1872 VSUBS 0.20fF $ **FLOATING
C2231 D.t234 VSUBS -0.02fF
C2232 D.n1874 VSUBS 0.20fF $ **FLOATING
C2233 D.t499 VSUBS -0.06fF
C2234 D.n1875 VSUBS 0.61fF $ **FLOATING
C2235 D.n1877 VSUBS 2.27fF $ **FLOATING
C2236 D.n1878 VSUBS 2.07fF $ **FLOATING
C2237 D.n1879 VSUBS 1.75fF $ **FLOATING
C2238 D.t581 VSUBS -0.02fF
C2239 D.n1880 VSUBS 0.20fF $ **FLOATING
C2240 D.t567 VSUBS -0.06fF
C2241 D.n1881 VSUBS 0.61fF $ **FLOATING
C2242 D.t365 VSUBS -0.02fF
C2243 D.n1883 VSUBS 0.20fF $ **FLOATING
C2244 D.t32 VSUBS -0.06fF
C2245 D.n1884 VSUBS 0.61fF $ **FLOATING
C2246 D.n1886 VSUBS 1.44fF $ **FLOATING
C2247 D.n1887 VSUBS 1.67fF $ **FLOATING
C2248 D.n1888 VSUBS 1.76fF $ **FLOATING
C2249 D.n1889 VSUBS 3.11fF $ **FLOATING
C2250 D.t37 VSUBS -0.06fF
C2251 D.n1890 VSUBS 0.61fF $ **FLOATING
C2252 D.t69 VSUBS -0.02fF
C2253 D.n1891 VSUBS 0.20fF $ **FLOATING
C2254 D.t470 VSUBS -0.02fF
C2255 D.n1893 VSUBS 0.20fF $ **FLOATING
C2256 D.t162 VSUBS -0.06fF
C2257 D.n1894 VSUBS 0.61fF $ **FLOATING
C2258 D.n1896 VSUBS 4.38fF $ **FLOATING
C2259 D.n1897 VSUBS 1.95fF $ **FLOATING
C2260 D.n1898 VSUBS 1.19fF $ **FLOATING
C2261 D.n1899 VSUBS 0.03fF $ **FLOATING
C2262 D.n1900 VSUBS 0.04fF $ **FLOATING
C2263 D.n1901 VSUBS 0.24fF $ **FLOATING
C2264 D.n1902 VSUBS 2.98fF $ **FLOATING
C2265 D.n1903 VSUBS 3.48fF $ **FLOATING
C2266 D.n1904 VSUBS 4.16fF $ **FLOATING
C2267 D.n1905 VSUBS 1.39fF $ **FLOATING
C2268 D.n1906 VSUBS 0.67fF $ **FLOATING
C2269 D.n1907 VSUBS 0.25fF $ **FLOATING
C2270 D.n1908 VSUBS 0.08fF $ **FLOATING
C2271 D.n1909 VSUBS 0.10fF $ **FLOATING
C2272 D.n1910 VSUBS 0.11fF $ **FLOATING
C2273 D.t248 VSUBS -0.06fF
C2274 D.n1911 VSUBS 0.25fF $ **FLOATING
C2275 D.t585 VSUBS 0.00fF
C2276 D.n1912 VSUBS 0.33fF $ **FLOATING
C2277 D.t372 VSUBS 0.00fF
C2278 D.n1913 VSUBS 0.33fF $ **FLOATING
C2279 D.n1914 VSUBS 1.13fF $ **FLOATING
C2280 D.n1915 VSUBS 11.41fF $ **FLOATING
C2281 D.n1916 VSUBS 1.03fF $ **FLOATING
C2282 D.n1917 VSUBS 3.12fF $ **FLOATING
C2283 D.n1918 VSUBS 4.43fF $ **FLOATING
C2284 D.n1919 VSUBS 0.93fF $ **FLOATING
C2285 D.n1920 VSUBS 3.17fF $ **FLOATING
C2286 D.n1921 VSUBS 7.61fF $ **FLOATING
C2287 D.n1922 VSUBS 1.91fF $ **FLOATING
C2288 D.n1923 VSUBS 2.16fF $ **FLOATING
C2289 D.n1924 VSUBS 1.36fF $ **FLOATING
C2290 D.n1925 VSUBS 8.10fF $ **FLOATING
C2291 D.n1926 VSUBS 1.05fF $ **FLOATING
C2292 D.n1927 VSUBS 7.59fF $ **FLOATING
C2293 S.n0 VSUBS 0.24fF $ **FLOATING
C2294 S.n1 VSUBS 0.20fF $ **FLOATING
C2295 S.t94 VSUBS 108.06fF
C2296 S.t99 VSUBS 108.64fF
C2297 S.n2 VSUBS 0.09fF $ **FLOATING
C2298 S.t144 VSUBS 98.77fF
C2299 S.t32 VSUBS 98.52fF
C2300 S.n3 VSUBS 15.21fF $ **FLOATING
C2301 S.n4 VSUBS 15.21fF $ **FLOATING
C2302 S.n5 VSUBS 15.21fF $ **FLOATING
C2303 S.n6 VSUBS 15.21fF $ **FLOATING
C2304 S.n7 VSUBS 17.10fF $ **FLOATING
C2305 S.n8 VSUBS 0.86fF $ **FLOATING
C2306 S.n9 VSUBS 16.56fF $ **FLOATING
C2307 S.n10 VSUBS 0.87fF $ **FLOATING
C2308 S.n11 VSUBS 0.87fF $ **FLOATING
C2309 S.n12 VSUBS 0.87fF $ **FLOATING
C2310 S.n13 VSUBS 0.87fF $ **FLOATING
C2311 S.n14 VSUBS 0.87fF $ **FLOATING
C2312 S.n15 VSUBS 0.87fF $ **FLOATING
C2313 S.n16 VSUBS 0.87fF $ **FLOATING
C2314 S.n17 VSUBS 0.87fF $ **FLOATING
C2315 S.n18 VSUBS 0.87fF $ **FLOATING
C2316 S.n19 VSUBS 0.87fF $ **FLOATING
C2317 S.n20 VSUBS 0.87fF $ **FLOATING
C2318 S.n21 VSUBS 0.87fF $ **FLOATING
C2319 S.n22 VSUBS 0.87fF $ **FLOATING
C2320 S.n23 VSUBS 0.87fF $ **FLOATING
C2321 S.n24 VSUBS 0.87fF $ **FLOATING
C2322 S.n25 VSUBS 0.87fF $ **FLOATING
C2323 S.t0 VSUBS 783.05fF
C2324 S.n26 VSUBS 0.87fF $ **FLOATING
C2325 S.n27 VSUBS 0.87fF $ **FLOATING
C2326 S.n28 VSUBS 0.87fF $ **FLOATING
C2327 S.n29 VSUBS 0.87fF $ **FLOATING
C2328 S.n30 VSUBS 0.87fF $ **FLOATING
C2329 S.n31 VSUBS 0.87fF $ **FLOATING
C2330 S.n32 VSUBS 0.87fF $ **FLOATING
C2331 S.n33 VSUBS 0.87fF $ **FLOATING
C2332 S.n34 VSUBS 0.87fF $ **FLOATING
C2333 S.n35 VSUBS 0.87fF $ **FLOATING
C2334 S.n36 VSUBS 0.87fF $ **FLOATING
C2335 S.n37 VSUBS 0.38fF $ **FLOATING
C2336 S.n38 VSUBS 0.87fF $ **FLOATING
C2337 S.n39 VSUBS 0.87fF $ **FLOATING
C2338 S.n40 VSUBS 0.38fF $ **FLOATING
C2339 S.n41 VSUBS 0.87fF $ **FLOATING
C2340 S.n42 VSUBS 0.87fF $ **FLOATING
C2341 S.n43 VSUBS 1.03fF $ **FLOATING
C2342 S.t2 VSUBS 196.12fF
C2343 S.t47 VSUBS 98.16fF
C2344 S.n44 VSUBS 1.54fF $ **FLOATING
C2345 S.n45 VSUBS 1.32fF $ **FLOATING
C2346 S.n46 VSUBS 0.09fF $ **FLOATING
C2347 S.t34 VSUBS 113.11fF
C2348 S.n47 VSUBS 0.09fF $ **FLOATING
C2349 S.n48 VSUBS 2.87fF $ **FLOATING
C2350 S.n49 VSUBS 2.87fF $ **FLOATING
C2351 S.t41 VSUBS 104.79fF
C2352 S.t78 VSUBS 106.32fF
C2353 S.n50 VSUBS 2.87fF $ **FLOATING
C2354 S.n51 VSUBS 0.26fF $ **FLOATING
C2355 S.t52 VSUBS 109.80fF
C2356 S.n52 VSUBS 1.85fF $ **FLOATING
C2357 S.n53 VSUBS 1.56fF $ **FLOATING
C2358 S.t139 VSUBS 96.42fF
C2359 S.n54 VSUBS 2.63fF $ **FLOATING
C2360 S.n55 VSUBS 12.69fF $ **FLOATING
C2361 S.n56 VSUBS 1.06fF $ **FLOATING
C2362 S.n57 VSUBS 0.14fF $ **FLOATING
C2363 S.n58 VSUBS 0.90fF $ **FLOATING
C2364 S.n59 VSUBS 16.29fF $ **FLOATING
C2365 S.n60 VSUBS 1.73fF $ **FLOATING
C2366 S.n61 VSUBS 16.15fF $ **FLOATING
C2367 S.n62 VSUBS 1.73fF $ **FLOATING
C2368 S.n63 VSUBS 16.22fF $ **FLOATING
C2369 S.n64 VSUBS 1.73fF $ **FLOATING
C2370 S.n65 VSUBS 16.29fF $ **FLOATING
C2371 S.n66 VSUBS 1.73fF $ **FLOATING
C2372 S.n67 VSUBS 0.14fF $ **FLOATING
C2373 S.t45 VSUBS 106.90fF
C2374 S.n68 VSUBS 0.14fF $ **FLOATING
C2375 S.n69 VSUBS 0.19fF $ **FLOATING
C2376 S.n70 VSUBS 2.87fF $ **FLOATING
C2377 S.n71 VSUBS 0.26fF $ **FLOATING
C2378 S.n72 VSUBS 0.96fF $ **FLOATING
C2379 S.n73 VSUBS 2.87fF $ **FLOATING
C2380 S.n74 VSUBS 0.14fF $ **FLOATING
C2381 S.n75 VSUBS 0.20fF $ **FLOATING
C2382 S.n76 VSUBS 0.20fF $ **FLOATING
C2383 S.t55 VSUBS 100.32fF
C2384 S.t49 VSUBS 110.48fF
C2385 S.n77 VSUBS 0.14fF $ **FLOATING
C2386 S.n78 VSUBS 8.54fF $ **FLOATING
C2387 S.n79 VSUBS 0.96fF $ **FLOATING
C2388 S.n80 VSUBS 0.20fF $ **FLOATING
C2389 S.n81 VSUBS 0.20fF $ **FLOATING
C2390 S.n82 VSUBS 0.24fF $ **FLOATING
C2391 S.t18 VSUBS 106.17fF
C2392 S.n83 VSUBS 0.14fF $ **FLOATING
C2393 S.n84 VSUBS 1.32fF $ **FLOATING
C2394 S.n85 VSUBS 0.89fF $ **FLOATING
C2395 S.n86 VSUBS 0.90fF $ **FLOATING
C2396 S.n87 VSUBS 0.32fF $ **FLOATING
C2397 S.n88 VSUBS 0.14fF $ **FLOATING
C2398 S.n89 VSUBS 0.14fF $ **FLOATING
C2399 S.t14 VSUBS 104.20fF
C2400 S.n90 VSUBS 9.85fF $ **FLOATING
C2401 S.n91 VSUBS 0.60fF $ **FLOATING
C2402 S.n92 VSUBS 0.60fF $ **FLOATING
C2403 S.n93 VSUBS 0.60fF $ **FLOATING
C2404 S.n94 VSUBS 0.60fF $ **FLOATING
C2405 S.n95 VSUBS 0.60fF $ **FLOATING
C2406 S.n96 VSUBS 1.64fF $ **FLOATING
C2407 S.n97 VSUBS 0.16fF $ **FLOATING
C2408 S.n98 VSUBS 0.16fF $ **FLOATING
C2409 S.n99 VSUBS 0.16fF $ **FLOATING
C2410 S.n100 VSUBS 0.16fF $ **FLOATING
C2411 S.n101 VSUBS 0.16fF $ **FLOATING
C2412 S.n102 VSUBS 1.64fF $ **FLOATING
C2413 S.n103 VSUBS 1.31fF $ **FLOATING
C2414 S.n104 VSUBS 1.33fF $ **FLOATING
C2415 S.n105 VSUBS 1.77fF $ **FLOATING
C2416 S.n106 VSUBS 8.77fF $ **FLOATING
C2417 S.n107 VSUBS 8.77fF $ **FLOATING
C2418 S.n108 VSUBS 94.27fF $ **FLOATING
C2419 S.n109 VSUBS 8.77fF $ **FLOATING
C2420 S.n110 VSUBS 8.77fF $ **FLOATING
C2421 S.n111 VSUBS 5.32fF $ **FLOATING
C2422 S.n112 VSUBS 13.30fF $ **FLOATING
C2423 S.n113 VSUBS 13.30fF $ **FLOATING
C2424 S.n114 VSUBS 5.26fF $ **FLOATING
C2425 S.t395 VSUBS 0.02fF
C2426 S.n115 VSUBS 8.77fF $ **FLOATING
C2427 S.n116 VSUBS 8.77fF $ **FLOATING
C2428 S.n117 VSUBS 5.35fF $ **FLOATING
C2429 S.t160 VSUBS 0.02fF
C2430 S.t377 VSUBS 0.02fF
C2431 S.n118 VSUBS 0.02fF $ **FLOATING
C2432 S.t368 VSUBS 0.02fF
C2433 S.n119 VSUBS 8.77fF $ **FLOATING
C2434 S.n120 VSUBS 8.77fF $ **FLOATING
C2435 S.n121 VSUBS 5.35fF $ **FLOATING
C2436 S.t616 VSUBS 0.02fF
C2437 S.t221 VSUBS 0.02fF
C2438 S.n122 VSUBS 5.78fF $ **FLOATING
C2439 S.n123 VSUBS 0.02fF $ **FLOATING
C2440 S.t563 VSUBS 0.02fF
C2441 S.n124 VSUBS 8.77fF $ **FLOATING
C2442 S.n125 VSUBS 8.77fF $ **FLOATING
C2443 S.t385 VSUBS 0.02fF
C2444 S.t592 VSUBS 0.02fF
C2445 S.n126 VSUBS 0.02fF $ **FLOATING
C2446 S.t333 VSUBS 0.02fF
C2447 S.n127 VSUBS 8.77fF $ **FLOATING
C2448 S.n128 VSUBS 8.77fF $ **FLOATING
C2449 S.n129 VSUBS 5.38fF $ **FLOATING
C2450 S.t574 VSUBS 0.02fF
C2451 S.t164 VSUBS 0.02fF
C2452 S.n130 VSUBS 0.02fF $ **FLOATING
C2453 S.t533 VSUBS 0.02fF
C2454 S.n131 VSUBS 20.33fF $ **FLOATING
C2455 S.n132 VSUBS 20.33fF $ **FLOATING
C2456 S.n133 VSUBS 5.68fF $ **FLOATING
C2457 S.t30 VSUBS 0.02fF
C2458 S.t367 VSUBS 0.02fF
C2459 S.n134 VSUBS 0.02fF $ **FLOATING
C2460 S.t329 VSUBS 0.02fF
C2461 S.t177 VSUBS 0.02fF
C2462 S.n135 VSUBS 0.02fF $ **FLOATING
C2463 S.t166 VSUBS 0.02fF
C2464 S.t494 VSUBS 0.02fF
C2465 S.t570 VSUBS 0.02fF
C2466 S.n136 VSUBS 0.02fF $ **FLOATING
C2467 S.t557 VSUBS 0.02fF
C2468 S.t389 VSUBS 0.02fF
C2469 S.t397 VSUBS 0.02fF
C2470 S.n137 VSUBS 0.02fF $ **FLOATING
C2471 S.t134 VSUBS 0.02fF
C2472 S.t184 VSUBS 0.02fF
C2473 S.t595 VSUBS 0.02fF
C2474 S.n138 VSUBS 1.28fF $ **FLOATING
C2475 S.n139 VSUBS 19.67fF $ **FLOATING
C2476 S.n140 VSUBS 5.75fF $ **FLOATING
C2477 S.n141 VSUBS 0.12fF $ **FLOATING
C2478 S.t313 VSUBS 0.02fF
C2479 S.n142 VSUBS 0.89fF $ **FLOATING
C2480 S.t521 VSUBS 0.02fF
C2481 S.n143 VSUBS 0.23fF $ **FLOATING
C2482 S.t578 VSUBS 0.02fF
C2483 S.n144 VSUBS 0.23fF $ **FLOATING
C2484 S.n145 VSUBS 0.89fF $ **FLOATING
C2485 S.t527 VSUBS 0.02fF
C2486 S.n146 VSUBS 0.12fF $ **FLOATING
C2487 S.n147 VSUBS 0.09fF $ **FLOATING
C2488 S.n148 VSUBS 0.18fF $ **FLOATING
C2489 S.n149 VSUBS 0.12fF $ **FLOATING
C2490 S.t510 VSUBS 0.02fF
C2491 S.n150 VSUBS 0.89fF $ **FLOATING
C2492 S.t86 VSUBS 0.02fF
C2493 S.n151 VSUBS 0.23fF $ **FLOATING
C2494 S.t3 VSUBS 0.02fF
C2495 S.n152 VSUBS 0.23fF $ **FLOATING
C2496 S.n153 VSUBS 0.89fF $ **FLOATING
C2497 S.t95 VSUBS 0.02fF
C2498 S.n154 VSUBS 0.12fF $ **FLOATING
C2499 S.n155 VSUBS 0.12fF $ **FLOATING
C2500 S.t622 VSUBS 0.02fF
C2501 S.n156 VSUBS 0.89fF $ **FLOATING
C2502 S.t493 VSUBS 0.02fF
C2503 S.n157 VSUBS 0.23fF $ **FLOATING
C2504 S.t157 VSUBS 0.02fF
C2505 S.n158 VSUBS 0.23fF $ **FLOATING
C2506 S.n159 VSUBS 0.89fF $ **FLOATING
C2507 S.t320 VSUBS 0.02fF
C2508 S.n160 VSUBS 0.12fF $ **FLOATING
C2509 S.n161 VSUBS 0.09fF $ **FLOATING
C2510 S.n162 VSUBS 0.18fF $ **FLOATING
C2511 S.n163 VSUBS 0.12fF $ **FLOATING
C2512 S.t200 VSUBS 0.02fF
C2513 S.n164 VSUBS 0.89fF $ **FLOATING
C2514 S.t138 VSUBS 0.02fF
C2515 S.n165 VSUBS 0.23fF $ **FLOATING
C2516 S.t355 VSUBS 0.02fF
C2517 S.n166 VSUBS 0.23fF $ **FLOATING
C2518 S.n167 VSUBS 0.89fF $ **FLOATING
C2519 S.t414 VSUBS 0.02fF
C2520 S.n168 VSUBS 0.12fF $ **FLOATING
C2521 S.n169 VSUBS 0.12fF $ **FLOATING
C2522 S.t392 VSUBS 0.02fF
C2523 S.t461 VSUBS 0.02fF
C2524 S.n170 VSUBS 1.19fF $ **FLOATING
C2525 S.n171 VSUBS 0.58fF $ **FLOATING
C2526 S.n172 VSUBS 0.58fF $ **FLOATING
C2527 S.t23 VSUBS 11.07fF
C2528 S.n173 VSUBS 0.01fF $ **FLOATING
C2529 S.t264 VSUBS 0.02fF
C2530 S.t536 VSUBS 0.04fF
C2531 S.n174 VSUBS 0.12fF $ **FLOATING
C2532 S.t419 VSUBS 0.02fF
C2533 S.n175 VSUBS 0.89fF $ **FLOATING
C2534 S.t24 VSUBS 0.02fF
C2535 S.n176 VSUBS 0.23fF $ **FLOATING
C2536 S.t8 VSUBS 0.02fF
C2537 S.n177 VSUBS 0.23fF $ **FLOATING
C2538 S.n178 VSUBS 0.89fF $ **FLOATING
C2539 S.t40 VSUBS 0.02fF
C2540 S.n179 VSUBS 0.12fF $ **FLOATING
C2541 S.n180 VSUBS 0.12fF $ **FLOATING
C2542 S.t15 VSUBS 0.02fF
C2543 S.n181 VSUBS 0.89fF $ **FLOATING
C2544 S.t238 VSUBS 0.02fF
C2545 S.n182 VSUBS 0.23fF $ **FLOATING
C2546 S.t303 VSUBS 0.02fF
C2547 S.n183 VSUBS 0.23fF $ **FLOATING
C2548 S.n184 VSUBS 0.89fF $ **FLOATING
C2549 S.t251 VSUBS 0.02fF
C2550 S.n185 VSUBS 0.12fF $ **FLOATING
C2551 S.n186 VSUBS 0.12fF $ **FLOATING
C2552 S.t259 VSUBS 0.02fF
C2553 S.n187 VSUBS 0.89fF $ **FLOATING
C2554 S.t426 VSUBS 0.02fF
C2555 S.n188 VSUBS 0.23fF $ **FLOATING
C2556 S.t486 VSUBS 0.02fF
C2557 S.n189 VSUBS 0.23fF $ **FLOATING
C2558 S.n190 VSUBS 0.89fF $ **FLOATING
C2559 S.t436 VSUBS 0.02fF
C2560 S.n191 VSUBS 0.12fF $ **FLOATING
C2561 S.n192 VSUBS 0.12fF $ **FLOATING
C2562 S.t206 VSUBS 0.02fF
C2563 S.n193 VSUBS 0.89fF $ **FLOATING
C2564 S.t146 VSUBS 0.02fF
C2565 S.n194 VSUBS 0.23fF $ **FLOATING
C2566 S.n195 VSUBS 0.13fF $ **FLOATING
C2567 S.t364 VSUBS 0.02fF
C2568 S.n196 VSUBS 0.23fF $ **FLOATING
C2569 S.n197 VSUBS 0.89fF $ **FLOATING
C2570 S.t422 VSUBS 0.02fF
C2571 S.n198 VSUBS 0.12fF $ **FLOATING
C2572 S.n199 VSUBS 0.12fF $ **FLOATING
C2573 S.t587 VSUBS 0.02fF
C2574 S.n200 VSUBS 0.89fF $ **FLOATING
C2575 S.t542 VSUBS 0.02fF
C2576 S.n201 VSUBS 0.23fF $ **FLOATING
C2577 S.t105 VSUBS 0.02fF
C2578 S.n202 VSUBS 0.23fF $ **FLOATING
C2579 S.n203 VSUBS 0.89fF $ **FLOATING
C2580 S.t176 VSUBS 0.02fF
C2581 S.n204 VSUBS 0.12fF $ **FLOATING
C2582 S.n205 VSUBS 0.12fF $ **FLOATING
C2583 S.t159 VSUBS 0.02fF
C2584 S.n206 VSUBS 0.89fF $ **FLOATING
C2585 S.t110 VSUBS 0.02fF
C2586 S.n207 VSUBS 0.23fF $ **FLOATING
C2587 S.t322 VSUBS 0.02fF
C2588 S.n208 VSUBS 0.23fF $ **FLOATING
C2589 S.n209 VSUBS 0.89fF $ **FLOATING
C2590 S.t376 VSUBS 0.02fF
C2591 S.n210 VSUBS 0.12fF $ **FLOATING
C2592 S.n211 VSUBS 10.74fF $ **FLOATING
C2593 S.n212 VSUBS 0.12fF $ **FLOATING
C2594 S.t597 VSUBS 0.02fF
C2595 S.n213 VSUBS 0.89fF $ **FLOATING
C2596 S.t274 VSUBS 0.02fF
C2597 S.n214 VSUBS 0.23fF $ **FLOATING
C2598 S.t569 VSUBS 0.02fF
C2599 S.n215 VSUBS 0.12fF $ **FLOATING
C2600 S.t603 VSUBS 0.02fF
C2601 S.n216 VSUBS 0.23fF $ **FLOATING
C2602 S.n217 VSUBS 0.89fF $ **FLOATING
C2603 S.t577 VSUBS 0.02fF
C2604 S.n218 VSUBS 0.12fF $ **FLOATING
C2605 S.t556 VSUBS 0.02fF
C2606 S.n219 VSUBS 0.23fF $ **FLOATING
C2607 S.n220 VSUBS 0.89fF $ **FLOATING
C2608 S.n221 VSUBS 0.89fF $ **FLOATING
C2609 S.t351 VSUBS 0.02fF
C2610 S.n222 VSUBS 0.23fF $ **FLOATING
C2611 S.n223 VSUBS 0.12fF $ **FLOATING
C2612 S.t394 VSUBS 0.02fF
C2613 S.n224 VSUBS 0.89fF $ **FLOATING
C2614 S.t344 VSUBS 0.02fF
C2615 S.n225 VSUBS 0.23fF $ **FLOATING
C2616 S.n226 VSUBS 1.73fF $ **FLOATING
C2617 S.t549 VSUBS 0.02fF
C2618 S.n227 VSUBS 0.23fF $ **FLOATING
C2619 S.n228 VSUBS 0.89fF $ **FLOATING
C2620 S.t598 VSUBS 0.02fF
C2621 S.n229 VSUBS 0.12fF $ **FLOATING
C2622 S.n230 VSUBS 1.01fF $ **FLOATING
C2623 S.n231 VSUBS 0.12fF $ **FLOATING
C2624 S.t580 VSUBS 0.02fF
C2625 S.n232 VSUBS 0.89fF $ **FLOATING
C2626 S.t539 VSUBS 0.02fF
C2627 S.n233 VSUBS 0.23fF $ **FLOATING
C2628 S.n234 VSUBS 0.09fF $ **FLOATING
C2629 S.n235 VSUBS 0.42fF $ **FLOATING
C2630 S.n236 VSUBS 1.08fF $ **FLOATING
C2631 S.t121 VSUBS 0.02fF
C2632 S.n237 VSUBS 0.23fF $ **FLOATING
C2633 S.n238 VSUBS 0.89fF $ **FLOATING
C2634 S.t172 VSUBS 0.02fF
C2635 S.n239 VSUBS 0.12fF $ **FLOATING
C2636 S.n240 VSUBS 0.09fF $ **FLOATING
C2637 S.n241 VSUBS 0.18fF $ **FLOATING
C2638 S.n242 VSUBS 0.75fF $ **FLOATING
C2639 S.n243 VSUBS 0.75fF $ **FLOATING
C2640 S.n244 VSUBS 0.12fF $ **FLOATING
C2641 S.t151 VSUBS 0.02fF
C2642 S.n245 VSUBS 0.89fF $ **FLOATING
C2643 S.t109 VSUBS 0.02fF
C2644 S.n246 VSUBS 0.23fF $ **FLOATING
C2645 S.t182 VSUBS 0.02fF
C2646 S.n247 VSUBS 0.23fF $ **FLOATING
C2647 S.n248 VSUBS 0.89fF $ **FLOATING
C2648 S.t375 VSUBS 0.02fF
C2649 S.n249 VSUBS 0.12fF $ **FLOATING
C2650 S.t326 VSUBS 0.02fF
C2651 S.n250 VSUBS 0.12fF $ **FLOATING
C2652 S.n251 VSUBS 0.12fF $ **FLOATING
C2653 S.t113 VSUBS 0.02fF
C2654 S.n252 VSUBS 0.89fF $ **FLOATING
C2655 S.t316 VSUBS 0.02fF
C2656 S.n253 VSUBS 0.23fF $ **FLOATING
C2657 S.n254 VSUBS 1.16fF $ **FLOATING
C2658 S.t386 VSUBS 0.02fF
C2659 S.n255 VSUBS 0.23fF $ **FLOATING
C2660 S.n256 VSUBS 0.89fF $ **FLOATING
C2661 S.t323 VSUBS 0.02fF
C2662 S.n257 VSUBS 0.01fF $ **FLOATING
C2663 S.t617 VSUBS 0.02fF
C2664 S.n258 VSUBS 1.17fF $ **FLOATING
C2665 S.n259 VSUBS 1.17fF $ **FLOATING
C2666 S.t550 VSUBS 0.02fF
C2667 S.n260 VSUBS 19.91fF $ **FLOATING
C2668 S.n261 VSUBS 19.91fF $ **FLOATING
C2669 S.n262 VSUBS 0.20fF $ **FLOATING
C2670 S.t7 VSUBS 11.07fF
C2671 S.n263 VSUBS 0.86fF $ **FLOATING
C2672 S.n264 VSUBS 0.08fF $ **FLOATING
C2673 S.n265 VSUBS 0.86fF $ **FLOATING
C2674 S.n266 VSUBS 0.48fF $ **FLOATING
C2675 S.n267 VSUBS 0.09fF $ **FLOATING
C2676 S.n268 VSUBS 0.24fF $ **FLOATING
C2677 S.n269 VSUBS 0.67fF $ **FLOATING
C2678 S.n270 VSUBS 0.12fF $ **FLOATING
C2679 S.t145 VSUBS 0.02fF
C2680 S.n271 VSUBS 0.89fF $ **FLOATING
C2681 S.t359 VSUBS 0.02fF
C2682 S.n272 VSUBS 0.23fF $ **FLOATING
C2683 S.n273 VSUBS 0.43fF $ **FLOATING
C2684 S.n274 VSUBS 0.02fF $ **FLOATING
C2685 S.t441 VSUBS 0.02fF
C2686 S.n275 VSUBS 0.23fF $ **FLOATING
C2687 S.n276 VSUBS 0.89fF $ **FLOATING
C2688 S.t382 VSUBS 0.02fF
C2689 S.n277 VSUBS 0.12fF $ **FLOATING
C2690 S.n278 VSUBS 0.09fF $ **FLOATING
C2691 S.n279 VSUBS 0.25fF $ **FLOATING
C2692 S.n280 VSUBS 0.12fF $ **FLOATING
C2693 S.t361 VSUBS 0.02fF
C2694 S.n281 VSUBS 0.89fF $ **FLOATING
C2695 S.t561 VSUBS 0.02fF
C2696 S.n282 VSUBS 0.23fF $ **FLOATING
C2697 S.n283 VSUBS 0.43fF $ **FLOATING
C2698 S.n284 VSUBS 0.02fF $ **FLOATING
C2699 S.t631 VSUBS 0.02fF
C2700 S.n285 VSUBS 0.23fF $ **FLOATING
C2701 S.n286 VSUBS 0.89fF $ **FLOATING
C2702 S.t571 VSUBS 0.02fF
C2703 S.n287 VSUBS 0.12fF $ **FLOATING
C2704 S.n288 VSUBS 0.09fF $ **FLOATING
C2705 S.n289 VSUBS 0.24fF $ **FLOATING
C2706 S.n290 VSUBS 0.67fF $ **FLOATING
C2707 S.n291 VSUBS 0.12fF $ **FLOATING
C2708 S.t217 VSUBS 0.02fF
C2709 S.n292 VSUBS 0.89fF $ **FLOATING
C2710 S.t156 VSUBS 0.02fF
C2711 S.n293 VSUBS 0.23fF $ **FLOATING
C2712 S.n294 VSUBS 0.46fF $ **FLOATING
C2713 S.n295 VSUBS 0.02fF $ **FLOATING
C2714 S.t362 VSUBS 0.02fF
C2715 S.n296 VSUBS 0.23fF $ **FLOATING
C2716 S.n297 VSUBS 0.89fF $ **FLOATING
C2717 S.t174 VSUBS 0.02fF
C2718 S.n298 VSUBS 0.12fF $ **FLOATING
C2719 S.n299 VSUBS 0.89fF $ **FLOATING
C2720 S.t353 VSUBS 0.02fF
C2721 S.n300 VSUBS 0.23fF $ **FLOATING
C2722 S.n301 VSUBS 0.12fF $ **FLOATING
C2723 S.t405 VSUBS 0.02fF
C2724 S.n302 VSUBS 1.12fF $ **FLOATING
C2725 S.t560 VSUBS 0.02fF
C2726 S.n303 VSUBS 0.23fF $ **FLOATING
C2727 S.n304 VSUBS 0.89fF $ **FLOATING
C2728 S.t611 VSUBS 0.02fF
C2729 S.n305 VSUBS 0.12fF $ **FLOATING
C2730 S.n306 VSUBS 0.12fF $ **FLOATING
C2731 S.t590 VSUBS 0.02fF
C2732 S.n307 VSUBS 0.89fF $ **FLOATING
C2733 S.t547 VSUBS 0.02fF
C2734 S.n308 VSUBS 0.23fF $ **FLOATING
C2735 S.n309 VSUBS 0.41fF $ **FLOATING
C2736 S.n310 VSUBS 0.50fF $ **FLOATING
C2737 S.t126 VSUBS 0.02fF
C2738 S.n311 VSUBS 0.23fF $ **FLOATING
C2739 S.n312 VSUBS 0.89fF $ **FLOATING
C2740 S.t193 VSUBS 0.02fF
C2741 S.n313 VSUBS 0.12fF $ **FLOATING
C2742 S.n314 VSUBS 0.09fF $ **FLOATING
C2743 S.n315 VSUBS 0.24fF $ **FLOATING
C2744 S.n316 VSUBS 0.67fF $ **FLOATING
C2745 S.n317 VSUBS 0.12fF $ **FLOATING
C2746 S.t162 VSUBS 0.02fF
C2747 S.n318 VSUBS 0.89fF $ **FLOATING
C2748 S.t120 VSUBS 0.02fF
C2749 S.n319 VSUBS 0.23fF $ **FLOATING
C2750 S.t324 VSUBS 0.02fF
C2751 S.n320 VSUBS 0.23fF $ **FLOATING
C2752 S.n321 VSUBS 0.89fF $ **FLOATING
C2753 S.t380 VSUBS 0.02fF
C2754 S.n322 VSUBS 0.12fF $ **FLOATING
C2755 S.n323 VSUBS 10.74fF $ **FLOATING
C2756 S.n324 VSUBS 0.09fF $ **FLOATING
C2757 S.n325 VSUBS 0.20fF $ **FLOATING
C2758 S.n326 VSUBS 0.06fF $ **FLOATING
C2759 S.n327 VSUBS 0.20fF $ **FLOATING
C2760 S.n328 VSUBS 0.12fF $ **FLOATING
C2761 S.t488 VSUBS 0.02fF
C2762 S.n329 VSUBS 0.89fF $ **FLOATING
C2763 S.t169 VSUBS 0.02fF
C2764 S.n330 VSUBS 0.23fF $ **FLOATING
C2765 S.n331 VSUBS 0.89fF $ **FLOATING
C2766 S.n332 VSUBS 0.41fF $ **FLOATING
C2767 S.t179 VSUBS 0.02fF
C2768 S.n333 VSUBS 0.12fF $ **FLOATING
C2769 S.t247 VSUBS 0.02fF
C2770 S.n334 VSUBS 0.23fF $ **FLOATING
C2771 S.n335 VSUBS 0.89fF $ **FLOATING
C2772 S.n336 VSUBS 0.12fF $ **FLOATING
C2773 S.t371 VSUBS 0.02fF
C2774 S.t321 VSUBS 0.02fF
C2775 S.n337 VSUBS 1.19fF $ **FLOATING
C2776 S.n338 VSUBS 0.58fF $ **FLOATING
C2777 S.n339 VSUBS 0.58fF $ **FLOATING
C2778 S.t88 VSUBS 11.07fF
C2779 S.n340 VSUBS 0.01fF $ **FLOATING
C2780 S.t114 VSUBS 0.02fF
C2781 S.t388 VSUBS 0.04fF
C2782 S.n341 VSUBS 0.12fF $ **FLOATING
C2783 S.t314 VSUBS 0.02fF
C2784 S.n342 VSUBS 0.89fF $ **FLOATING
C2785 S.t523 VSUBS 0.02fF
C2786 S.n343 VSUBS 0.23fF $ **FLOATING
C2787 S.t579 VSUBS 0.02fF
C2788 S.n344 VSUBS 0.23fF $ **FLOATING
C2789 S.n345 VSUBS 0.89fF $ **FLOATING
C2790 S.t528 VSUBS 0.02fF
C2791 S.n346 VSUBS 0.12fF $ **FLOATING
C2792 S.n347 VSUBS 0.89fF $ **FLOATING
C2793 S.t89 VSUBS 0.02fF
C2794 S.n348 VSUBS 0.23fF $ **FLOATING
C2795 S.n349 VSUBS 0.12fF $ **FLOATING
C2796 S.t511 VSUBS 0.02fF
C2797 S.n350 VSUBS 0.09fF $ **FLOATING
C2798 S.n351 VSUBS 0.25fF $ **FLOATING
C2799 S.t148 VSUBS 0.02fF
C2800 S.n352 VSUBS 0.23fF $ **FLOATING
C2801 S.n353 VSUBS 0.89fF $ **FLOATING
C2802 S.t100 VSUBS 0.02fF
C2803 S.n354 VSUBS 0.12fF $ **FLOATING
C2804 S.n355 VSUBS 0.12fF $ **FLOATING
C2805 S.t108 VSUBS 0.02fF
C2806 S.n356 VSUBS 0.89fF $ **FLOATING
C2807 S.t288 VSUBS 0.02fF
C2808 S.n357 VSUBS 0.23fF $ **FLOATING
C2809 S.t345 VSUBS 0.02fF
C2810 S.n358 VSUBS 0.23fF $ **FLOATING
C2811 S.n359 VSUBS 0.89fF $ **FLOATING
C2812 S.t298 VSUBS 0.02fF
C2813 S.n360 VSUBS 0.12fF $ **FLOATING
C2814 S.n361 VSUBS 0.89fF $ **FLOATING
C2815 S.t358 VSUBS 0.02fF
C2816 S.n362 VSUBS 0.23fF $ **FLOATING
C2817 S.n363 VSUBS 0.12fF $ **FLOATING
C2818 S.t412 VSUBS 0.02fF
C2819 S.n364 VSUBS 0.09fF $ **FLOATING
C2820 S.n365 VSUBS 0.25fF $ **FLOATING
C2821 S.t567 VSUBS 0.02fF
C2822 S.n366 VSUBS 0.23fF $ **FLOATING
C2823 S.n367 VSUBS 0.89fF $ **FLOATING
C2824 S.t572 VSUBS 0.02fF
C2825 S.n368 VSUBS 0.12fF $ **FLOATING
C2826 S.n369 VSUBS 0.89fF $ **FLOATING
C2827 S.t555 VSUBS 0.02fF
C2828 S.n370 VSUBS 0.23fF $ **FLOATING
C2829 S.n371 VSUBS 0.12fF $ **FLOATING
C2830 S.t600 VSUBS 0.02fF
C2831 S.t132 VSUBS 0.02fF
C2832 S.n372 VSUBS 0.23fF $ **FLOATING
C2833 S.n373 VSUBS 0.89fF $ **FLOATING
C2834 S.t188 VSUBS 0.02fF
C2835 S.n374 VSUBS 0.12fF $ **FLOATING
C2836 S.n375 VSUBS 0.12fF $ **FLOATING
C2837 S.t170 VSUBS 0.02fF
C2838 S.n376 VSUBS 0.89fF $ **FLOATING
C2839 S.t111 VSUBS 0.02fF
C2840 S.n377 VSUBS 0.23fF $ **FLOATING
C2841 S.t330 VSUBS 0.02fF
C2842 S.n378 VSUBS 0.23fF $ **FLOATING
C2843 S.n379 VSUBS 0.89fF $ **FLOATING
C2844 S.t390 VSUBS 0.02fF
C2845 S.n380 VSUBS 0.12fF $ **FLOATING
C2846 S.n381 VSUBS 10.74fF $ **FLOATING
C2847 S.n382 VSUBS 0.12fF $ **FLOATING
C2848 S.t552 VSUBS 0.02fF
C2849 S.n383 VSUBS 0.89fF $ **FLOATING
C2850 S.t183 VSUBS 0.02fF
C2851 S.n384 VSUBS 0.23fF $ **FLOATING
C2852 S.t150 VSUBS 0.02fF
C2853 S.n385 VSUBS 0.12fF $ **FLOATING
C2854 S.t535 VSUBS 0.02fF
C2855 S.n386 VSUBS 0.23fF $ **FLOATING
C2856 S.n387 VSUBS 0.89fF $ **FLOATING
C2857 S.t582 VSUBS 0.02fF
C2858 S.n388 VSUBS 0.12fF $ **FLOATING
C2859 S.t530 VSUBS 0.02fF
C2860 S.n389 VSUBS 0.23fF $ **FLOATING
C2861 S.n390 VSUBS 0.89fF $ **FLOATING
C2862 S.n391 VSUBS 0.89fF $ **FLOATING
C2863 S.t319 VSUBS 0.02fF
C2864 S.n392 VSUBS 0.23fF $ **FLOATING
C2865 S.n393 VSUBS 0.12fF $ **FLOATING
C2866 S.t366 VSUBS 0.02fF
C2867 S.n394 VSUBS 0.89fF $ **FLOATING
C2868 S.t185 VSUBS 0.02fF
C2869 S.n395 VSUBS 0.23fF $ **FLOATING
C2870 S.t575 VSUBS 0.02fF
C2871 S.n396 VSUBS 0.12fF $ **FLOATING
C2872 S.t515 VSUBS 0.02fF
C2873 S.n397 VSUBS 0.23fF $ **FLOATING
C2874 S.n398 VSUBS 0.89fF $ **FLOATING
C2875 S.t276 VSUBS 0.02fF
C2876 S.n399 VSUBS 0.01fF $ **FLOATING
C2877 S.t474 VSUBS 0.02fF
C2878 S.n400 VSUBS 1.17fF $ **FLOATING
C2879 S.n401 VSUBS 1.17fF $ **FLOATING
C2880 S.t409 VSUBS 0.02fF
C2881 S.n402 VSUBS 8.77fF $ **FLOATING
C2882 S.t119 VSUBS 11.07fF
C2883 S.n403 VSUBS 0.58fF $ **FLOATING
C2884 S.n404 VSUBS 0.08fF $ **FLOATING
C2885 S.n405 VSUBS 0.48fF $ **FLOATING
C2886 S.n406 VSUBS 5.02fF $ **FLOATING
C2887 S.n407 VSUBS 8.77fF $ **FLOATING
C2888 S.n408 VSUBS 0.43fF $ **FLOATING
C2889 S.n409 VSUBS 0.02fF $ **FLOATING
C2890 S.n410 VSUBS 0.89fF $ **FLOATING
C2891 S.t239 VSUBS 0.02fF
C2892 S.n411 VSUBS 0.23fF $ **FLOATING
C2893 S.n412 VSUBS 1.50fF $ **FLOATING
C2894 S.n413 VSUBS 0.12fF $ **FLOATING
C2895 S.t19 VSUBS 0.02fF
C2896 S.n414 VSUBS 0.09fF $ **FLOATING
C2897 S.n415 VSUBS 0.25fF $ **FLOATING
C2898 S.t307 VSUBS 0.02fF
C2899 S.n416 VSUBS 0.23fF $ **FLOATING
C2900 S.n417 VSUBS 0.89fF $ **FLOATING
C2901 S.t249 VSUBS 0.02fF
C2902 S.n418 VSUBS 0.12fF $ **FLOATING
C2903 S.n419 VSUBS 0.09fF $ **FLOATING
C2904 S.n420 VSUBS 0.24fF $ **FLOATING
C2905 S.n421 VSUBS 0.12fF $ **FLOATING
C2906 S.t232 VSUBS 0.02fF
C2907 S.n422 VSUBS 0.89fF $ **FLOATING
C2908 S.t431 VSUBS 0.02fF
C2909 S.n423 VSUBS 0.23fF $ **FLOATING
C2910 S.t500 VSUBS 0.02fF
C2911 S.n424 VSUBS 0.23fF $ **FLOATING
C2912 S.n425 VSUBS 0.89fF $ **FLOATING
C2913 S.t438 VSUBS 0.02fF
C2914 S.n426 VSUBS 0.12fF $ **FLOATING
C2915 S.n427 VSUBS 0.89fF $ **FLOATING
C2916 S.t369 VSUBS 0.02fF
C2917 S.n428 VSUBS 0.23fF $ **FLOATING
C2918 S.n429 VSUBS 1.50fF $ **FLOATING
C2919 S.n430 VSUBS 0.12fF $ **FLOATING
C2920 S.t415 VSUBS 0.02fF
C2921 S.n431 VSUBS 0.09fF $ **FLOATING
C2922 S.n432 VSUBS 0.25fF $ **FLOATING
C2923 S.t495 VSUBS 0.02fF
C2924 S.n433 VSUBS 0.23fF $ **FLOATING
C2925 S.n434 VSUBS 0.89fF $ **FLOATING
C2926 S.t28 VSUBS 0.02fF
C2927 S.n435 VSUBS 0.12fF $ **FLOATING
C2928 S.n436 VSUBS 0.60fF $ **FLOATING
C2929 S.n437 VSUBS 0.41fF $ **FLOATING
C2930 S.n438 VSUBS 0.89fF $ **FLOATING
C2931 S.t558 VSUBS 0.02fF
C2932 S.n439 VSUBS 0.23fF $ **FLOATING
C2933 S.n440 VSUBS 0.12fF $ **FLOATING
C2934 S.t602 VSUBS 0.02fF
C2935 S.t137 VSUBS 0.02fF
C2936 S.n441 VSUBS 0.23fF $ **FLOATING
C2937 S.n442 VSUBS 0.89fF $ **FLOATING
C2938 S.t202 VSUBS 0.02fF
C2939 S.n443 VSUBS 0.12fF $ **FLOATING
C2940 S.n444 VSUBS 0.09fF $ **FLOATING
C2941 S.n445 VSUBS 0.24fF $ **FLOATING
C2942 S.n446 VSUBS 0.12fF $ **FLOATING
C2943 S.t175 VSUBS 0.02fF
C2944 S.n447 VSUBS 0.89fF $ **FLOATING
C2945 S.t124 VSUBS 0.02fF
C2946 S.n448 VSUBS 0.23fF $ **FLOATING
C2947 S.t347 VSUBS 0.02fF
C2948 S.n449 VSUBS 0.23fF $ **FLOATING
C2949 S.n450 VSUBS 0.89fF $ **FLOATING
C2950 S.t393 VSUBS 0.02fF
C2951 S.n451 VSUBS 0.12fF $ **FLOATING
C2952 S.n452 VSUBS 10.74fF $ **FLOATING
C2953 S.n453 VSUBS 0.24fF $ **FLOATING
C2954 S.n454 VSUBS 0.20fF $ **FLOATING
C2955 S.n455 VSUBS 0.12fF $ **FLOATING
C2956 S.t454 VSUBS 0.02fF
C2957 S.n456 VSUBS 0.89fF $ **FLOATING
C2958 S.t21 VSUBS 0.02fF
C2959 S.n457 VSUBS 0.23fF $ **FLOATING
C2960 S.t38 VSUBS 0.02fF
C2961 S.n458 VSUBS 0.12fF $ **FLOATING
C2962 S.t104 VSUBS 0.02fF
C2963 S.n459 VSUBS 0.23fF $ **FLOATING
C2964 S.n460 VSUBS 0.89fF $ **FLOATING
C2965 S.n461 VSUBS 0.12fF $ **FLOATING
C2966 S.t383 VSUBS 0.02fF
C2967 S.t589 VSUBS 0.02fF
C2968 S.n462 VSUBS 0.12fF $ **FLOATING
C2969 S.t540 VSUBS 0.02fF
C2970 S.n463 VSUBS 0.23fF $ **FLOATING
C2971 S.n464 VSUBS 0.89fF $ **FLOATING
C2972 S.n465 VSUBS 0.89fF $ **FLOATING
C2973 S.t331 VSUBS 0.02fF
C2974 S.n466 VSUBS 0.23fF $ **FLOATING
C2975 S.n467 VSUBS 0.12fF $ **FLOATING
C2976 S.t373 VSUBS 0.02fF
C2977 S.n468 VSUBS 0.89fF $ **FLOATING
C2978 S.t325 VSUBS 0.02fF
C2979 S.n469 VSUBS 0.23fF $ **FLOATING
C2980 S.t586 VSUBS 0.02fF
C2981 S.n470 VSUBS 0.12fF $ **FLOATING
C2982 S.t534 VSUBS 0.02fF
C2983 S.n471 VSUBS 0.23fF $ **FLOATING
C2984 S.n472 VSUBS 0.89fF $ **FLOATING
C2985 S.n473 VSUBS 0.12fF $ **FLOATING
C2986 S.t573 VSUBS 0.02fF
C2987 S.t171 VSUBS 0.02fF
C2988 S.n474 VSUBS 1.19fF $ **FLOATING
C2989 S.n475 VSUBS 0.58fF $ **FLOATING
C2990 S.n476 VSUBS 0.58fF $ **FLOATING
C2991 S.t5 VSUBS 11.07fF
C2992 S.n477 VSUBS 0.01fF $ **FLOATING
C2993 S.t593 VSUBS 0.02fF
C2994 S.t258 VSUBS 0.04fF
C2995 S.n478 VSUBS 0.89fF $ **FLOATING
C2996 S.t372 VSUBS 0.02fF
C2997 S.n479 VSUBS 0.23fF $ **FLOATING
C2998 S.n480 VSUBS 0.12fF $ **FLOATING
C2999 S.t163 VSUBS 0.02fF
C3000 S.n481 VSUBS 0.09fF $ **FLOATING
C3001 S.n482 VSUBS 0.25fF $ **FLOATING
C3002 S.t444 VSUBS 0.02fF
C3003 S.n483 VSUBS 0.23fF $ **FLOATING
C3004 S.n484 VSUBS 0.89fF $ **FLOATING
C3005 S.t384 VSUBS 0.02fF
C3006 S.n485 VSUBS 0.12fF $ **FLOATING
C3007 S.n486 VSUBS 0.12fF $ **FLOATING
C3008 S.t363 VSUBS 0.02fF
C3009 S.n487 VSUBS 0.89fF $ **FLOATING
C3010 S.t562 VSUBS 0.02fF
C3011 S.n488 VSUBS 0.23fF $ **FLOATING
C3012 S.t632 VSUBS 0.02fF
C3013 S.n489 VSUBS 0.23fF $ **FLOATING
C3014 S.n490 VSUBS 0.89fF $ **FLOATING
C3015 S.t576 VSUBS 0.02fF
C3016 S.n491 VSUBS 0.12fF $ **FLOATING
C3017 S.n492 VSUBS 0.89fF $ **FLOATING
C3018 S.t128 VSUBS 0.02fF
C3019 S.n493 VSUBS 0.23fF $ **FLOATING
C3020 S.n494 VSUBS 0.12fF $ **FLOATING
C3021 S.t585 VSUBS 0.02fF
C3022 S.n495 VSUBS 0.09fF $ **FLOATING
C3023 S.n496 VSUBS 0.25fF $ **FLOATING
C3024 S.t213 VSUBS 0.02fF
C3025 S.n497 VSUBS 0.23fF $ **FLOATING
C3026 S.n498 VSUBS 0.89fF $ **FLOATING
C3027 S.t140 VSUBS 0.02fF
C3028 S.n499 VSUBS 0.12fF $ **FLOATING
C3029 S.n500 VSUBS 0.89fF $ **FLOATING
C3030 S.t566 VSUBS 0.02fF
C3031 S.n501 VSUBS 0.23fF $ **FLOATING
C3032 S.n502 VSUBS 0.12fF $ **FLOATING
C3033 S.t609 VSUBS 0.02fF
C3034 S.t141 VSUBS 0.02fF
C3035 S.n503 VSUBS 0.23fF $ **FLOATING
C3036 S.n504 VSUBS 0.89fF $ **FLOATING
C3037 S.t215 VSUBS 0.02fF
C3038 S.n505 VSUBS 0.12fF $ **FLOATING
C3039 S.n506 VSUBS 0.12fF $ **FLOATING
C3040 S.t180 VSUBS 0.02fF
C3041 S.n507 VSUBS 0.89fF $ **FLOATING
C3042 S.t131 VSUBS 0.02fF
C3043 S.n508 VSUBS 0.23fF $ **FLOATING
C3044 S.t349 VSUBS 0.02fF
C3045 S.n509 VSUBS 0.23fF $ **FLOATING
C3046 S.n510 VSUBS 0.89fF $ **FLOATING
C3047 S.t404 VSUBS 0.02fF
C3048 S.n511 VSUBS 0.12fF $ **FLOATING
C3049 S.n512 VSUBS 10.74fF $ **FLOATING
C3050 S.n513 VSUBS 0.12fF $ **FLOATING
C3051 S.t509 VSUBS 0.02fF
C3052 S.n514 VSUBS 0.37fF $ **FLOATING
C3053 S.n515 VSUBS 0.89fF $ **FLOATING
C3054 S.t6 VSUBS 0.02fF
C3055 S.n516 VSUBS 0.23fF $ **FLOATING
C3056 S.t365 VSUBS 0.02fF
C3057 S.n517 VSUBS 0.12fF $ **FLOATING
C3058 S.t471 VSUBS 0.02fF
C3059 S.n518 VSUBS 0.23fF $ **FLOATING
C3060 S.n519 VSUBS 0.89fF $ **FLOATING
C3061 S.t142 VSUBS 0.02fF
C3062 S.n520 VSUBS 0.12fF $ **FLOATING
C3063 S.t112 VSUBS 0.02fF
C3064 S.n521 VSUBS 0.23fF $ **FLOATING
C3065 S.n522 VSUBS 0.89fF $ **FLOATING
C3066 S.n523 VSUBS 0.89fF $ **FLOATING
C3067 S.t529 VSUBS 0.02fF
C3068 S.n524 VSUBS 0.23fF $ **FLOATING
C3069 S.n525 VSUBS 0.12fF $ **FLOATING
C3070 S.t568 VSUBS 0.02fF
C3071 S.n526 VSUBS 0.89fF $ **FLOATING
C3072 S.t526 VSUBS 0.02fF
C3073 S.n527 VSUBS 0.23fF $ **FLOATING
C3074 S.t154 VSUBS 0.02fF
C3075 S.n528 VSUBS 0.12fF $ **FLOATING
C3076 S.t107 VSUBS 0.02fF
C3077 S.n529 VSUBS 0.23fF $ **FLOATING
C3078 S.n530 VSUBS 0.89fF $ **FLOATING
C3079 S.t231 VSUBS 0.02fF
C3080 S.n531 VSUBS 0.01fF $ **FLOATING
C3081 S.t342 VSUBS 0.02fF
C3082 S.n532 VSUBS 1.17fF $ **FLOATING
C3083 S.n533 VSUBS 1.17fF $ **FLOATING
C3084 S.t273 VSUBS 0.02fF
C3085 S.n534 VSUBS 5.08fF $ **FLOATING
C3086 S.n535 VSUBS 8.77fF $ **FLOATING
C3087 S.n536 VSUBS 8.77fF $ **FLOATING
C3088 S.t20 VSUBS 11.07fF
C3089 S.n537 VSUBS 0.58fF $ **FLOATING
C3090 S.n538 VSUBS 0.08fF $ **FLOATING
C3091 S.n539 VSUBS 0.48fF $ **FLOATING
C3092 S.n540 VSUBS 0.01fF $ **FLOATING
C3093 S.n541 VSUBS 0.07fF $ **FLOATING
C3094 S.n542 VSUBS 0.23fF $ **FLOATING
C3095 S.n543 VSUBS 0.01fF $ **FLOATING
C3096 S.n544 VSUBS 0.09fF $ **FLOATING
C3097 S.n545 VSUBS 0.24fF $ **FLOATING
C3098 S.n546 VSUBS 0.12fF $ **FLOATING
C3099 S.t514 VSUBS 0.02fF
C3100 S.n547 VSUBS 0.89fF $ **FLOATING
C3101 S.t130 VSUBS 0.02fF
C3102 S.n548 VSUBS 0.23fF $ **FLOATING
C3103 S.t152 VSUBS 0.02fF
C3104 S.n549 VSUBS 0.23fF $ **FLOATING
C3105 S.n550 VSUBS 0.89fF $ **FLOATING
C3106 S.t102 VSUBS 0.02fF
C3107 S.n551 VSUBS 0.12fF $ **FLOATING
C3108 S.n552 VSUBS 0.89fF $ **FLOATING
C3109 S.t328 VSUBS 0.02fF
C3110 S.n553 VSUBS 0.23fF $ **FLOATING
C3111 S.n554 VSUBS 1.50fF $ **FLOATING
C3112 S.n555 VSUBS 0.12fF $ **FLOATING
C3113 S.t79 VSUBS 0.02fF
C3114 S.n556 VSUBS 0.09fF $ **FLOATING
C3115 S.n557 VSUBS 0.25fF $ **FLOATING
C3116 S.t341 VSUBS 0.02fF
C3117 S.n558 VSUBS 0.23fF $ **FLOATING
C3118 S.n559 VSUBS 0.89fF $ **FLOATING
C3119 S.t187 VSUBS 0.02fF
C3120 S.n560 VSUBS 0.12fF $ **FLOATING
C3121 S.n561 VSUBS 0.60fF $ **FLOATING
C3122 S.n562 VSUBS 0.41fF $ **FLOATING
C3123 S.n563 VSUBS 0.89fF $ **FLOATING
C3124 S.t39 VSUBS 0.02fF
C3125 S.n564 VSUBS 0.23fF $ **FLOATING
C3126 S.n565 VSUBS 0.12fF $ **FLOATING
C3127 S.t620 VSUBS 0.02fF
C3128 S.t155 VSUBS 0.02fF
C3129 S.n566 VSUBS 0.23fF $ **FLOATING
C3130 S.n567 VSUBS 0.89fF $ **FLOATING
C3131 S.t524 VSUBS 0.02fF
C3132 S.n568 VSUBS 0.12fF $ **FLOATING
C3133 S.n569 VSUBS 0.09fF $ **FLOATING
C3134 S.n570 VSUBS 0.24fF $ **FLOATING
C3135 S.n571 VSUBS 0.12fF $ **FLOATING
C3136 S.t197 VSUBS 0.02fF
C3137 S.n572 VSUBS 0.89fF $ **FLOATING
C3138 S.t252 VSUBS 0.02fF
C3139 S.n573 VSUBS 0.23fF $ **FLOATING
C3140 S.t352 VSUBS 0.02fF
C3141 S.n574 VSUBS 0.23fF $ **FLOATING
C3142 S.n575 VSUBS 0.89fF $ **FLOATING
C3143 S.t410 VSUBS 0.02fF
C3144 S.n576 VSUBS 0.12fF $ **FLOATING
C3145 S.n577 VSUBS 10.74fF $ **FLOATING
C3146 S.n578 VSUBS 0.89fF $ **FLOATING
C3147 S.t564 VSUBS 0.02fF
C3148 S.n579 VSUBS 0.23fF $ **FLOATING
C3149 S.n580 VSUBS 1.21fF $ **FLOATING
C3150 S.n581 VSUBS 0.12fF $ **FLOATING
C3151 S.t304 VSUBS 0.02fF
C3152 S.n582 VSUBS 0.20fF $ **FLOATING
C3153 S.n583 VSUBS 0.09fF $ **FLOATING
C3154 S.n584 VSUBS 0.20fF $ **FLOATING
C3155 S.n585 VSUBS 0.06fF $ **FLOATING
C3156 S.t531 VSUBS 0.02fF
C3157 S.n586 VSUBS 0.12fF $ **FLOATING
C3158 S.t583 VSUBS 0.02fF
C3159 S.n587 VSUBS 0.23fF $ **FLOATING
C3160 S.n588 VSUBS 0.89fF $ **FLOATING
C3161 S.n589 VSUBS 0.12fF $ **FLOATING
C3162 S.t387 VSUBS 0.02fF
C3163 S.n590 VSUBS 0.89fF $ **FLOATING
C3164 S.t437 VSUBS 0.02fF
C3165 S.n591 VSUBS 0.23fF $ **FLOATING
C3166 S.t599 VSUBS 0.02fF
C3167 S.n592 VSUBS 0.12fF $ **FLOATING
C3168 S.t545 VSUBS 0.02fF
C3169 S.n593 VSUBS 0.23fF $ **FLOATING
C3170 S.n594 VSUBS 0.89fF $ **FLOATING
C3171 S.n595 VSUBS 0.12fF $ **FLOATING
C3172 S.t581 VSUBS 0.02fF
C3173 S.n596 VSUBS 0.89fF $ **FLOATING
C3174 S.t624 VSUBS 0.02fF
C3175 S.n597 VSUBS 0.23fF $ **FLOATING
C3176 S.t168 VSUBS 0.02fF
C3177 S.n598 VSUBS 0.12fF $ **FLOATING
C3178 S.t117 VSUBS 0.02fF
C3179 S.n599 VSUBS 0.23fF $ **FLOATING
C3180 S.n600 VSUBS 0.89fF $ **FLOATING
C3181 S.n601 VSUBS 0.12fF $ **FLOATING
C3182 S.t189 VSUBS 0.02fF
C3183 S.t93 VSUBS 0.02fF
C3184 S.n602 VSUBS 1.19fF $ **FLOATING
C3185 S.n603 VSUBS 0.58fF $ **FLOATING
C3186 S.n604 VSUBS 0.58fF $ **FLOATING
C3187 S.t25 VSUBS 11.07fF
C3188 S.n605 VSUBS 0.01fF $ **FLOATING
C3189 S.t518 VSUBS 0.02fF
C3190 S.t153 VSUBS 0.04fF
C3191 S.n606 VSUBS 0.12fF $ **FLOATING
C3192 S.t85 VSUBS 0.02fF
C3193 S.n607 VSUBS 0.89fF $ **FLOATING
C3194 S.t293 VSUBS 0.02fF
C3195 S.n608 VSUBS 0.23fF $ **FLOATING
C3196 S.t335 VSUBS 0.02fF
C3197 S.n609 VSUBS 0.23fF $ **FLOATING
C3198 S.n610 VSUBS 0.89fF $ **FLOATING
C3199 S.t301 VSUBS 0.02fF
C3200 S.n611 VSUBS 0.12fF $ **FLOATING
C3201 S.n612 VSUBS 0.89fF $ **FLOATING
C3202 S.t472 VSUBS 0.02fF
C3203 S.n613 VSUBS 0.23fF $ **FLOATING
C3204 S.n614 VSUBS 0.12fF $ **FLOATING
C3205 S.t282 VSUBS 0.02fF
C3206 S.n615 VSUBS 0.09fF $ **FLOATING
C3207 S.n616 VSUBS 0.25fF $ **FLOATING
C3208 S.t544 VSUBS 0.02fF
C3209 S.n617 VSUBS 0.23fF $ **FLOATING
C3210 S.n618 VSUBS 0.89fF $ **FLOATING
C3211 S.t485 VSUBS 0.02fF
C3212 S.n619 VSUBS 0.12fF $ **FLOATING
C3213 S.n620 VSUBS 0.89fF $ **FLOATING
C3214 S.t37 VSUBS 0.02fF
C3215 S.n621 VSUBS 0.23fF $ **FLOATING
C3216 S.n622 VSUBS 0.12fF $ **FLOATING
C3217 S.t505 VSUBS 0.02fF
C3218 S.t116 VSUBS 0.02fF
C3219 S.n623 VSUBS 0.23fF $ **FLOATING
C3220 S.n624 VSUBS 0.89fF $ **FLOATING
C3221 S.t64 VSUBS 0.02fF
C3222 S.n625 VSUBS 0.12fF $ **FLOATING
C3223 S.n626 VSUBS 0.12fF $ **FLOATING
C3224 S.t305 VSUBS 0.02fF
C3225 S.n627 VSUBS 0.89fF $ **FLOATING
C3226 S.t254 VSUBS 0.02fF
C3227 S.n628 VSUBS 0.23fF $ **FLOATING
C3228 S.t418 VSUBS 0.02fF
C3229 S.n629 VSUBS 0.23fF $ **FLOATING
C3230 S.n630 VSUBS 0.89fF $ **FLOATING
C3231 S.t519 VSUBS 0.02fF
C3232 S.n631 VSUBS 0.12fF $ **FLOATING
C3233 S.n632 VSUBS 10.74fF $ **FLOATING
C3234 S.n633 VSUBS 0.12fF $ **FLOATING
C3235 S.t482 VSUBS 0.02fF
C3236 S.n634 VSUBS 0.89fF $ **FLOATING
C3237 S.t443 VSUBS 0.02fF
C3238 S.n635 VSUBS 0.23fF $ **FLOATING
C3239 S.t84 VSUBS 0.02fF
C3240 S.n636 VSUBS 0.12fF $ **FLOATING
C3241 S.t17 VSUBS 0.02fF
C3242 S.n637 VSUBS 0.23fF $ **FLOATING
C3243 S.n638 VSUBS 0.89fF $ **FLOATING
C3244 S.n639 VSUBS 0.12fF $ **FLOATING
C3245 S.t61 VSUBS 0.02fF
C3246 S.n640 VSUBS 0.89fF $ **FLOATING
C3247 S.t629 VSUBS 0.02fF
C3248 S.n641 VSUBS 0.23fF $ **FLOATING
C3249 S.t280 VSUBS 0.02fF
C3250 S.n642 VSUBS 0.12fF $ **FLOATING
C3251 S.t228 VSUBS 0.02fF
C3252 S.n643 VSUBS 0.23fF $ **FLOATING
C3253 S.n644 VSUBS 0.89fF $ **FLOATING
C3254 S.n645 VSUBS 0.12fF $ **FLOATING
C3255 S.t283 VSUBS 0.02fF
C3256 S.n646 VSUBS 0.37fF $ **FLOATING
C3257 S.n647 VSUBS 0.89fF $ **FLOATING
C3258 S.t281 VSUBS 0.02fF
C3259 S.n648 VSUBS 0.23fF $ **FLOATING
C3260 S.t42 VSUBS 0.02fF
C3261 S.n649 VSUBS 0.12fF $ **FLOATING
C3262 S.t618 VSUBS 0.02fF
C3263 S.n650 VSUBS 0.23fF $ **FLOATING
C3264 S.n651 VSUBS 0.89fF $ **FLOATING
C3265 S.t340 VSUBS 0.02fF
C3266 S.n652 VSUBS 0.12fF $ **FLOATING
C3267 S.t334 VSUBS 0.02fF
C3268 S.n653 VSUBS 0.23fF $ **FLOATING
C3269 S.n654 VSUBS 0.89fF $ **FLOATING
C3270 S.n655 VSUBS 0.89fF $ **FLOATING
C3271 S.t210 VSUBS 0.02fF
C3272 S.n656 VSUBS 0.23fF $ **FLOATING
C3273 S.n657 VSUBS 0.12fF $ **FLOATING
C3274 S.t147 VSUBS 0.02fF
C3275 S.n658 VSUBS 0.89fF $ **FLOATING
C3276 S.t204 VSUBS 0.02fF
C3277 S.n659 VSUBS 0.23fF $ **FLOATING
C3278 S.t360 VSUBS 0.02fF
C3279 S.n660 VSUBS 0.12fF $ **FLOATING
C3280 S.t315 VSUBS 0.02fF
C3281 S.n661 VSUBS 0.23fF $ **FLOATING
C3282 S.n662 VSUBS 0.89fF $ **FLOATING
C3283 S.t158 VSUBS 0.02fF
C3284 S.n663 VSUBS 0.01fF $ **FLOATING
C3285 S.t198 VSUBS 0.02fF
C3286 S.n664 VSUBS 1.17fF $ **FLOATING
C3287 S.n665 VSUBS 1.17fF $ **FLOATING
C3288 S.t173 VSUBS 0.02fF
C3289 S.n666 VSUBS 5.08fF $ **FLOATING
C3290 S.n667 VSUBS 8.77fF $ **FLOATING
C3291 S.n668 VSUBS 8.77fF $ **FLOATING
C3292 S.t16 VSUBS 11.07fF
C3293 S.n669 VSUBS 0.58fF $ **FLOATING
C3294 S.n670 VSUBS 0.08fF $ **FLOATING
C3295 S.n671 VSUBS 0.48fF $ **FLOATING
C3296 S.n672 VSUBS 0.07fF $ **FLOATING
C3297 S.n673 VSUBS 0.23fF $ **FLOATING
C3298 S.n674 VSUBS 0.01fF $ **FLOATING
C3299 S.n675 VSUBS 0.01fF $ **FLOATING
C3300 S.n676 VSUBS 0.05fF $ **FLOATING
C3301 S.n677 VSUBS 0.08fF $ **FLOATING
C3302 S.n678 VSUBS 0.05fF $ **FLOATING
C3303 S.n679 VSUBS 0.22fF $ **FLOATING
C3304 S.n680 VSUBS 0.95fF $ **FLOATING
C3305 S.t10 VSUBS 11.07fF
C3306 S.n681 VSUBS 0.58fF $ **FLOATING
C3307 S.n682 VSUBS 0.08fF $ **FLOATING
C3308 S.n683 VSUBS 0.48fF $ **FLOATING
C3309 S.n684 VSUBS 0.89fF $ **FLOATING
C3310 S.t613 VSUBS 0.02fF
C3311 S.n685 VSUBS 0.23fF $ **FLOATING
C3312 S.n686 VSUBS 1.50fF $ **FLOATING
C3313 S.n687 VSUBS 0.12fF $ **FLOATING
C3314 S.t424 VSUBS 0.02fF
C3315 S.n688 VSUBS 0.09fF $ **FLOATING
C3316 S.n689 VSUBS 0.25fF $ **FLOATING
C3317 S.t71 VSUBS 0.02fF
C3318 S.n690 VSUBS 0.23fF $ **FLOATING
C3319 S.n691 VSUBS 0.89fF $ **FLOATING
C3320 S.t628 VSUBS 0.02fF
C3321 S.n692 VSUBS 0.12fF $ **FLOATING
C3322 S.n693 VSUBS 0.60fF $ **FLOATING
C3323 S.n694 VSUBS 0.41fF $ **FLOATING
C3324 S.n695 VSUBS 0.89fF $ **FLOATING
C3325 S.t195 VSUBS 0.02fF
C3326 S.n696 VSUBS 0.23fF $ **FLOATING
C3327 S.n697 VSUBS 0.12fF $ **FLOATING
C3328 S.t491 VSUBS 0.02fF
C3329 S.t267 VSUBS 0.02fF
C3330 S.n698 VSUBS 0.23fF $ **FLOATING
C3331 S.n699 VSUBS 0.89fF $ **FLOATING
C3332 S.t209 VSUBS 0.02fF
C3333 S.n700 VSUBS 0.12fF $ **FLOATING
C3334 S.n701 VSUBS 0.09fF $ **FLOATING
C3335 S.n702 VSUBS 0.24fF $ **FLOATING
C3336 S.n703 VSUBS 0.12fF $ **FLOATING
C3337 S.t312 VSUBS 0.02fF
C3338 S.n704 VSUBS 0.89fF $ **FLOATING
C3339 S.t261 VSUBS 0.02fF
C3340 S.n705 VSUBS 0.23fF $ **FLOATING
C3341 S.t459 VSUBS 0.02fF
C3342 S.n706 VSUBS 0.23fF $ **FLOATING
C3343 S.n707 VSUBS 0.89fF $ **FLOATING
C3344 S.t421 VSUBS 0.02fF
C3345 S.n708 VSUBS 0.12fF $ **FLOATING
C3346 S.n709 VSUBS 10.74fF $ **FLOATING
C3347 S.n710 VSUBS 0.24fF $ **FLOATING
C3348 S.n711 VSUBS 0.20fF $ **FLOATING
C3349 S.n712 VSUBS 0.12fF $ **FLOATING
C3350 S.t227 VSUBS 0.02fF
C3351 S.n713 VSUBS 0.89fF $ **FLOATING
C3352 S.t434 VSUBS 0.02fF
C3353 S.n714 VSUBS 0.23fF $ **FLOATING
C3354 S.t442 VSUBS 0.02fF
C3355 S.n715 VSUBS 0.12fF $ **FLOATING
C3356 S.t504 VSUBS 0.02fF
C3357 S.n716 VSUBS 0.23fF $ **FLOATING
C3358 S.n717 VSUBS 0.89fF $ **FLOATING
C3359 S.n718 VSUBS 0.12fF $ **FLOATING
C3360 S.t503 VSUBS 0.02fF
C3361 S.n719 VSUBS 0.89fF $ **FLOATING
C3362 S.t446 VSUBS 0.02fF
C3363 S.n720 VSUBS 0.23fF $ **FLOATING
C3364 S.t92 VSUBS 0.02fF
C3365 S.n721 VSUBS 0.12fF $ **FLOATING
C3366 S.t26 VSUBS 0.02fF
C3367 S.n722 VSUBS 0.23fF $ **FLOATING
C3368 S.n723 VSUBS 0.89fF $ **FLOATING
C3369 S.n724 VSUBS 0.12fF $ **FLOATING
C3370 S.t70 VSUBS 0.02fF
C3371 S.n725 VSUBS 0.89fF $ **FLOATING
C3372 S.t636 VSUBS 0.02fF
C3373 S.n726 VSUBS 0.23fF $ **FLOATING
C3374 S.t292 VSUBS 0.02fF
C3375 S.n727 VSUBS 0.12fF $ **FLOATING
C3376 S.t236 VSUBS 0.02fF
C3377 S.n728 VSUBS 0.23fF $ **FLOATING
C3378 S.n729 VSUBS 0.89fF $ **FLOATING
C3379 S.n730 VSUBS 0.12fF $ **FLOATING
C3380 S.t269 VSUBS 0.02fF
C3381 S.n731 VSUBS 0.89fF $ **FLOATING
C3382 S.t222 VSUBS 0.02fF
C3383 S.n732 VSUBS 0.23fF $ **FLOATING
C3384 S.t473 VSUBS 0.02fF
C3385 S.n733 VSUBS 0.12fF $ **FLOATING
C3386 S.t425 VSUBS 0.02fF
C3387 S.n734 VSUBS 0.23fF $ **FLOATING
C3388 S.n735 VSUBS 0.89fF $ **FLOATING
C3389 S.n736 VSUBS 0.12fF $ **FLOATING
C3390 S.t463 VSUBS 0.02fF
C3391 S.t243 VSUBS 0.02fF
C3392 S.n737 VSUBS 0.23fF $ **FLOATING
C3393 S.t191 VSUBS 0.02fF
C3394 S.n738 VSUBS 0.12fF $ **FLOATING
C3395 S.n739 VSUBS 0.12fF $ **FLOATING
C3396 S.t74 VSUBS 0.02fF
C3397 S.t565 VSUBS 0.02fF
C3398 S.n740 VSUBS 1.19fF $ **FLOATING
C3399 S.n741 VSUBS 0.58fF $ **FLOATING
C3400 S.t12 VSUBS 11.07fF
C3401 S.n742 VSUBS 0.01fF $ **FLOATING
C3402 S.t370 VSUBS 0.02fF
C3403 S.t638 VSUBS 0.04fF
C3404 S.n743 VSUBS 0.89fF $ **FLOATING
C3405 S.t133 VSUBS 0.02fF
C3406 S.n744 VSUBS 0.23fF $ **FLOATING
C3407 S.n745 VSUBS 0.12fF $ **FLOATING
C3408 S.t559 VSUBS 0.02fF
C3409 S.n746 VSUBS 0.09fF $ **FLOATING
C3410 S.n747 VSUBS 0.25fF $ **FLOATING
C3411 S.t223 VSUBS 0.02fF
C3412 S.n748 VSUBS 0.23fF $ **FLOATING
C3413 S.n749 VSUBS 0.89fF $ **FLOATING
C3414 S.t143 VSUBS 0.02fF
C3415 S.n750 VSUBS 0.12fF $ **FLOATING
C3416 S.n751 VSUBS 0.89fF $ **FLOATING
C3417 S.t332 VSUBS 0.02fF
C3418 S.n752 VSUBS 0.23fF $ **FLOATING
C3419 S.n753 VSUBS 0.12fF $ **FLOATING
C3420 S.t125 VSUBS 0.02fF
C3421 S.t407 VSUBS 0.02fF
C3422 S.n754 VSUBS 0.23fF $ **FLOATING
C3423 S.n755 VSUBS 0.89fF $ **FLOATING
C3424 S.t350 VSUBS 0.02fF
C3425 S.n756 VSUBS 0.12fF $ **FLOATING
C3426 S.n757 VSUBS 0.12fF $ **FLOATING
C3427 S.t357 VSUBS 0.02fF
C3428 S.n758 VSUBS 0.89fF $ **FLOATING
C3429 S.t532 VSUBS 0.02fF
C3430 S.n759 VSUBS 0.23fF $ **FLOATING
C3431 S.t594 VSUBS 0.02fF
C3432 S.n760 VSUBS 0.23fF $ **FLOATING
C3433 S.n761 VSUBS 0.89fF $ **FLOATING
C3434 S.t541 VSUBS 0.02fF
C3435 S.n762 VSUBS 0.12fF $ **FLOATING
C3436 S.n763 VSUBS 10.74fF $ **FLOATING
C3437 S.n764 VSUBS 0.12fF $ **FLOATING
C3438 S.t508 VSUBS 0.02fF
C3439 S.n765 VSUBS 0.89fF $ **FLOATING
C3440 S.t451 VSUBS 0.02fF
C3441 S.n766 VSUBS 0.23fF $ **FLOATING
C3442 S.t98 VSUBS 0.02fF
C3443 S.n767 VSUBS 0.12fF $ **FLOATING
C3444 S.t29 VSUBS 0.02fF
C3445 S.n768 VSUBS 0.23fF $ **FLOATING
C3446 S.n769 VSUBS 0.89fF $ **FLOATING
C3447 S.n770 VSUBS 0.12fF $ **FLOATING
C3448 S.t272 VSUBS 0.02fF
C3449 S.n771 VSUBS 0.89fF $ **FLOATING
C3450 S.t230 VSUBS 0.02fF
C3451 S.n772 VSUBS 0.23fF $ **FLOATING
C3452 S.t478 VSUBS 0.02fF
C3453 S.n773 VSUBS 0.12fF $ **FLOATING
C3454 S.t433 VSUBS 0.02fF
C3455 S.n774 VSUBS 0.23fF $ **FLOATING
C3456 S.n775 VSUBS 0.89fF $ **FLOATING
C3457 S.n776 VSUBS 0.09fF $ **FLOATING
C3458 S.n777 VSUBS 0.25fF $ **FLOATING
C3459 S.n778 VSUBS 0.12fF $ **FLOATING
C3460 S.t235 VSUBS 0.02fF
C3461 S.n779 VSUBS 0.89fF $ **FLOATING
C3462 S.t211 VSUBS 0.02fF
C3463 S.n780 VSUBS 0.23fF $ **FLOATING
C3464 S.n781 VSUBS 0.60fF $ **FLOATING
C3465 S.t256 VSUBS 0.02fF
C3466 S.n782 VSUBS 0.12fF $ **FLOATING
C3467 S.t551 VSUBS 0.02fF
C3468 S.n783 VSUBS 0.23fF $ **FLOATING
C3469 S.n784 VSUBS 0.89fF $ **FLOATING
C3470 S.n785 VSUBS 0.23fF $ **FLOATING
C3471 S.t13 VSUBS 0.02fF
C3472 S.t56 VSUBS 0.02fF
C3473 S.n786 VSUBS 0.12fF $ **FLOATING
C3474 S.t614 VSUBS 0.02fF
C3475 S.n787 VSUBS 0.23fF $ **FLOATING
C3476 S.n788 VSUBS 0.89fF $ **FLOATING
C3477 S.n789 VSUBS 0.89fF $ **FLOATING
C3478 S.t343 VSUBS 0.02fF
C3479 S.n790 VSUBS 0.23fF $ **FLOATING
C3480 S.n791 VSUBS 0.12fF $ **FLOATING
C3481 S.t453 VSUBS 0.02fF
C3482 S.n792 VSUBS 0.89fF $ **FLOATING
C3483 S.t408 VSUBS 0.02fF
C3484 S.n793 VSUBS 0.23fF $ **FLOATING
C3485 S.t50 VSUBS 0.02fF
C3486 S.n794 VSUBS 0.12fF $ **FLOATING
C3487 S.t487 VSUBS 0.02fF
C3488 S.n795 VSUBS 0.23fF $ **FLOATING
C3489 S.n796 VSUBS 0.89fF $ **FLOATING
C3490 S.t553 VSUBS 0.02fF
C3491 S.n797 VSUBS 0.01fF $ **FLOATING
C3492 S.t106 VSUBS 0.02fF
C3493 S.n798 VSUBS 1.17fF $ **FLOATING
C3494 S.n799 VSUBS 1.17fF $ **FLOATING
C3495 S.t11 VSUBS 0.02fF
C3496 S.n800 VSUBS 0.05fF $ **FLOATING
C3497 S.n801 VSUBS 0.08fF $ **FLOATING
C3498 S.n802 VSUBS 0.05fF $ **FLOATING
C3499 S.n803 VSUBS 0.09fF $ **FLOATING
C3500 S.n804 VSUBS 0.24fF $ **FLOATING
C3501 S.n805 VSUBS 0.12fF $ **FLOATING
C3502 S.t127 VSUBS 0.02fF
C3503 S.n806 VSUBS 0.89fF $ **FLOATING
C3504 S.t346 VSUBS 0.02fF
C3505 S.n807 VSUBS 0.23fF $ **FLOATING
C3506 S.t411 VSUBS 0.02fF
C3507 S.n808 VSUBS 0.23fF $ **FLOATING
C3508 S.n809 VSUBS 0.89fF $ **FLOATING
C3509 S.t337 VSUBS 0.02fF
C3510 S.n810 VSUBS 0.12fF $ **FLOATING
C3511 S.n811 VSUBS 0.89fF $ **FLOATING
C3512 S.t205 VSUBS 0.02fF
C3513 S.n812 VSUBS 0.23fF $ **FLOATING
C3514 S.t296 VSUBS 0.02fF
C3515 S.n813 VSUBS 0.01fF $ **FLOATING
C3516 S.t91 VSUBS 0.02fF
C3517 S.t356 VSUBS 0.04fF
C3518 S.n814 VSUBS 0.12fF $ **FLOATING
C3519 S.t291 VSUBS 0.02fF
C3520 S.n815 VSUBS 0.89fF $ **FLOATING
C3521 S.t477 VSUBS 0.02fF
C3522 S.n816 VSUBS 0.23fF $ **FLOATING
C3523 S.t548 VSUBS 0.02fF
C3524 S.n817 VSUBS 0.23fF $ **FLOATING
C3525 S.n818 VSUBS 0.89fF $ **FLOATING
C3526 S.t501 VSUBS 0.02fF
C3527 S.n819 VSUBS 0.12fF $ **FLOATING
C3528 S.n820 VSUBS 0.37fF $ **FLOATING
C3529 S.n821 VSUBS 0.89fF $ **FLOATING
C3530 S.t73 VSUBS 0.02fF
C3531 S.n822 VSUBS 0.23fF $ **FLOATING
C3532 S.n823 VSUBS 0.12fF $ **FLOATING
C3533 S.t118 VSUBS 0.02fF
C3534 S.t338 VSUBS 0.02fF
C3535 S.n824 VSUBS 0.23fF $ **FLOATING
C3536 S.n825 VSUBS 0.89fF $ **FLOATING
C3537 S.t33 VSUBS 0.02fF
C3538 S.n826 VSUBS 0.12fF $ **FLOATING
C3539 S.n827 VSUBS 0.12fF $ **FLOATING
C3540 S.t469 VSUBS 0.02fF
C3541 S.n828 VSUBS 0.89fF $ **FLOATING
C3542 S.t54 VSUBS 0.02fF
C3543 S.n829 VSUBS 0.23fF $ **FLOATING
C3544 S.t62 VSUBS 0.02fF
C3545 S.n830 VSUBS 0.12fF $ **FLOATING
C3546 S.t122 VSUBS 0.02fF
C3547 S.n831 VSUBS 0.23fF $ **FLOATING
C3548 S.n832 VSUBS 0.89fF $ **FLOATING
C3549 S.n833 VSUBS 0.89fF $ **FLOATING
C3550 S.t257 VSUBS 0.02fF
C3551 S.n834 VSUBS 0.23fF $ **FLOATING
C3552 S.n835 VSUBS 0.12fF $ **FLOATING
C3553 S.t76 VSUBS 0.02fF
C3554 S.t266 VSUBS 0.02fF
C3555 S.n836 VSUBS 0.12fF $ **FLOATING
C3556 S.t317 VSUBS 0.02fF
C3557 S.n837 VSUBS 0.23fF $ **FLOATING
C3558 S.n838 VSUBS 0.89fF $ **FLOATING
C3559 S.n839 VSUBS 0.12fF $ **FLOATING
C3560 S.t299 VSUBS 0.02fF
C3561 S.n840 VSUBS 0.89fF $ **FLOATING
C3562 S.t248 VSUBS 0.02fF
C3563 S.n841 VSUBS 0.23fF $ **FLOATING
C3564 S.t512 VSUBS 0.02fF
C3565 S.n842 VSUBS 0.12fF $ **FLOATING
C3566 S.t450 VSUBS 0.02fF
C3567 S.n843 VSUBS 0.23fF $ **FLOATING
C3568 S.n844 VSUBS 0.89fF $ **FLOATING
C3569 S.n845 VSUBS 0.12fF $ **FLOATING
C3570 S.t481 VSUBS 0.02fF
C3571 S.n846 VSUBS 0.89fF $ **FLOATING
C3572 S.t439 VSUBS 0.02fF
C3573 S.n847 VSUBS 0.23fF $ **FLOATING
C3574 S.t77 VSUBS 0.02fF
C3575 S.n848 VSUBS 0.12fF $ **FLOATING
C3576 S.t1 VSUBS 0.02fF
C3577 S.n849 VSUBS 0.23fF $ **FLOATING
C3578 S.n850 VSUBS 0.89fF $ **FLOATING
C3579 S.n851 VSUBS 0.12fF $ **FLOATING
C3580 S.t57 VSUBS 0.02fF
C3581 S.n852 VSUBS 0.89fF $ **FLOATING
C3582 S.t625 VSUBS 0.02fF
C3583 S.n853 VSUBS 0.23fF $ **FLOATING
C3584 S.t278 VSUBS 0.02fF
C3585 S.n854 VSUBS 0.12fF $ **FLOATING
C3586 S.t225 VSUBS 0.02fF
C3587 S.n855 VSUBS 0.23fF $ **FLOATING
C3588 S.n856 VSUBS 0.89fF $ **FLOATING
C3589 S.t413 VSUBS 0.02fF
C3590 S.n857 VSUBS 0.23fF $ **FLOATING
C3591 S.n858 VSUBS 0.89fF $ **FLOATING
C3592 S.t465 VSUBS 0.02fF
C3593 S.n859 VSUBS 0.12fF $ **FLOATING
C3594 S.n860 VSUBS 0.12fF $ **FLOATING
C3595 S.t263 VSUBS 0.02fF
C3596 S.n861 VSUBS 0.12fF $ **FLOATING
C3597 S.t255 VSUBS 0.02fF
C3598 S.n862 VSUBS 0.89fF $ **FLOATING
C3599 S.t199 VSUBS 0.02fF
C3600 S.n863 VSUBS 0.23fF $ **FLOATING
C3601 S.t406 VSUBS 0.02fF
C3602 S.n864 VSUBS 0.23fF $ **FLOATING
C3603 S.n865 VSUBS 0.89fF $ **FLOATING
C3604 S.t462 VSUBS 0.02fF
C3605 S.n866 VSUBS 0.12fF $ **FLOATING
C3606 S.n867 VSUBS 0.89fF $ **FLOATING
C3607 S.t135 VSUBS 0.02fF
C3608 S.n868 VSUBS 0.23fF $ **FLOATING
C3609 S.n869 VSUBS 0.12fF $ **FLOATING
C3610 S.t554 VSUBS 0.02fF
C3611 S.n870 VSUBS 1.40fF $ **FLOATING
C3612 S.t149 VSUBS 0.02fF
C3613 S.n871 VSUBS 0.12fF $ **FLOATING
C3614 S.t224 VSUBS 0.02fF
C3615 S.n872 VSUBS 0.23fF $ **FLOATING
C3616 S.n873 VSUBS 0.89fF $ **FLOATING
C3617 S.n874 VSUBS 0.12fF $ **FLOATING
C3618 S.t327 VSUBS 0.02fF
C3619 S.n875 VSUBS 0.89fF $ **FLOATING
C3620 S.t537 VSUBS 0.02fF
C3621 S.n876 VSUBS 0.23fF $ **FLOATING
C3622 S.t543 VSUBS 0.02fF
C3623 S.n877 VSUBS 0.12fF $ **FLOATING
C3624 S.t596 VSUBS 0.02fF
C3625 S.n878 VSUBS 0.23fF $ **FLOATING
C3626 S.n879 VSUBS 0.89fF $ **FLOATING
C3627 S.n880 VSUBS 0.89fF $ **FLOATING
C3628 S.t43 VSUBS 0.02fF
C3629 S.n881 VSUBS 0.23fF $ **FLOATING
C3630 S.n882 VSUBS 0.12fF $ **FLOATING
C3631 S.t97 VSUBS 0.02fF
C3632 S.t136 VSUBS 0.02fF
C3633 S.n883 VSUBS 0.12fF $ **FLOATING
C3634 S.t260 VSUBS 0.02fF
C3635 S.n884 VSUBS 0.23fF $ **FLOATING
C3636 S.n885 VSUBS 0.89fF $ **FLOATING
C3637 S.n886 VSUBS 0.12fF $ **FLOATING
C3638 S.t295 VSUBS 0.02fF
C3639 S.n887 VSUBS 0.89fF $ **FLOATING
C3640 S.t245 VSUBS 0.02fF
C3641 S.n888 VSUBS 0.23fF $ **FLOATING
C3642 S.t507 VSUBS 0.02fF
C3643 S.n889 VSUBS 0.12fF $ **FLOATING
C3644 S.t448 VSUBS 0.02fF
C3645 S.n890 VSUBS 0.23fF $ **FLOATING
C3646 S.n891 VSUBS 0.89fF $ **FLOATING
C3647 S.n892 VSUBS 0.12fF $ **FLOATING
C3648 S.t476 VSUBS 0.02fF
C3649 S.n893 VSUBS 0.89fF $ **FLOATING
C3650 S.t417 VSUBS 0.02fF
C3651 S.n894 VSUBS 0.23fF $ **FLOATING
C3652 S.t63 VSUBS 0.02fF
C3653 S.n895 VSUBS 0.12fF $ **FLOATING
C3654 S.t635 VSUBS 0.02fF
C3655 S.n896 VSUBS 0.23fF $ **FLOATING
C3656 S.n897 VSUBS 0.89fF $ **FLOATING
C3657 S.n898 VSUBS 0.09fF $ **FLOATING
C3658 S.n899 VSUBS 0.25fF $ **FLOATING
C3659 S.n900 VSUBS 0.12fF $ **FLOATING
C3660 S.t53 VSUBS 0.02fF
C3661 S.n901 VSUBS 0.89fF $ **FLOATING
C3662 S.t621 VSUBS 0.02fF
C3663 S.n902 VSUBS 0.23fF $ **FLOATING
C3664 S.t271 VSUBS 0.02fF
C3665 S.n903 VSUBS 0.12fF $ **FLOATING
C3666 S.t218 VSUBS 0.02fF
C3667 S.n904 VSUBS 0.23fF $ **FLOATING
C3668 S.n905 VSUBS 0.89fF $ **FLOATING
C3669 S.t456 VSUBS 0.02fF
C3670 S.n906 VSUBS 0.01fF $ **FLOATING
C3671 S.t449 VSUBS 0.02fF
C3672 S.n907 VSUBS 1.17fF $ **FLOATING
C3673 S.n908 VSUBS 1.17fF $ **FLOATING
C3674 S.n909 VSUBS 0.16fF $ **FLOATING
C3675 S.t374 VSUBS 0.02fF
C3676 S.t244 VSUBS 0.02fF
C3677 S.n910 VSUBS 1.19fF $ **FLOATING
C3678 S.n911 VSUBS 0.89fF $ **FLOATING
C3679 S.t400 VSUBS 0.02fF
C3680 S.n912 VSUBS 0.23fF $ **FLOATING
C3681 S.n913 VSUBS 1.32fF $ **FLOATING
C3682 S.n914 VSUBS 0.12fF $ **FLOATING
C3683 S.t420 VSUBS 0.02fF
C3684 S.t604 VSUBS 0.02fF
C3685 S.n915 VSUBS 0.23fF $ **FLOATING
C3686 S.n916 VSUBS 0.89fF $ **FLOATING
C3687 S.t46 VSUBS 0.02fF
C3688 S.n917 VSUBS 0.12fF $ **FLOATING
C3689 S.n918 VSUBS 0.89fF $ **FLOATING
C3690 S.t207 VSUBS 0.02fF
C3691 S.n919 VSUBS 0.23fF $ **FLOATING
C3692 S.n920 VSUBS 0.12fF $ **FLOATING
C3693 S.t265 VSUBS 0.02fF
C3694 S.t416 VSUBS 0.02fF
C3695 S.n921 VSUBS 0.23fF $ **FLOATING
C3696 S.n922 VSUBS 0.89fF $ **FLOATING
C3697 S.t339 VSUBS 0.02fF
C3698 S.n923 VSUBS 0.12fF $ **FLOATING
C3699 S.n924 VSUBS 0.12fF $ **FLOATING
C3700 S.t430 VSUBS 0.02fF
C3701 S.n925 VSUBS 0.89fF $ **FLOATING
C3702 S.t492 VSUBS 0.02fF
C3703 S.n926 VSUBS 0.23fF $ **FLOATING
C3704 S.t633 VSUBS 0.02fF
C3705 S.n927 VSUBS 0.12fF $ **FLOATING
C3706 S.t75 VSUBS 0.02fF
C3707 S.n928 VSUBS 0.23fF $ **FLOATING
C3708 S.n929 VSUBS 0.89fF $ **FLOATING
C3709 S.n930 VSUBS 0.12fF $ **FLOATING
C3710 S.t610 VSUBS 0.02fF
C3711 S.n931 VSUBS 0.89fF $ **FLOATING
C3712 S.t190 VSUBS 0.02fF
C3713 S.n932 VSUBS 0.23fF $ **FLOATING
C3714 S.n933 VSUBS 0.85fF $ **FLOATING
C3715 S.t216 VSUBS 0.02fF
C3716 S.n934 VSUBS 0.12fF $ **FLOATING
C3717 S.t275 VSUBS 0.02fF
C3718 S.n935 VSUBS 0.23fF $ **FLOATING
C3719 S.n936 VSUBS 0.89fF $ **FLOATING
C3720 S.n937 VSUBS 0.89fF $ **FLOATING
C3721 S.t391 VSUBS 0.02fF
C3722 S.n938 VSUBS 0.23fF $ **FLOATING
C3723 S.n939 VSUBS 0.12fF $ **FLOATING
C3724 S.t192 VSUBS 0.02fF
C3725 S.t403 VSUBS 0.02fF
C3726 S.n940 VSUBS 0.12fF $ **FLOATING
C3727 S.t460 VSUBS 0.02fF
C3728 S.n941 VSUBS 0.23fF $ **FLOATING
C3729 S.n942 VSUBS 0.89fF $ **FLOATING
C3730 S.n943 VSUBS 0.12fF $ **FLOATING
C3731 S.t308 VSUBS 0.02fF
C3732 S.n944 VSUBS 0.89fF $ **FLOATING
C3733 S.t246 VSUBS 0.02fF
C3734 S.n945 VSUBS 0.23fF $ **FLOATING
C3735 S.t626 VSUBS 0.02fF
C3736 S.n946 VSUBS 0.12fF $ **FLOATING
C3737 S.t457 VSUBS 0.02fF
C3738 S.n947 VSUBS 0.23fF $ **FLOATING
C3739 S.n948 VSUBS 0.89fF $ **FLOATING
C3740 S.n949 VSUBS 0.12fF $ **FLOATING
C3741 S.t489 VSUBS 0.02fF
C3742 S.n950 VSUBS 0.89fF $ **FLOATING
C3743 S.t445 VSUBS 0.02fF
C3744 S.n951 VSUBS 0.23fF $ **FLOATING
C3745 S.t90 VSUBS 0.02fF
C3746 S.n952 VSUBS 0.12fF $ **FLOATING
C3747 S.t4 VSUBS 0.02fF
C3748 S.n953 VSUBS 0.23fF $ **FLOATING
C3749 S.n954 VSUBS 0.89fF $ **FLOATING
C3750 S.n955 VSUBS 0.12fF $ **FLOATING
C3751 S.t66 VSUBS 0.02fF
C3752 S.n956 VSUBS 0.89fF $ **FLOATING
C3753 S.t634 VSUBS 0.02fF
C3754 S.n957 VSUBS 0.23fF $ **FLOATING
C3755 S.t287 VSUBS 0.02fF
C3756 S.n958 VSUBS 0.12fF $ **FLOATING
C3757 S.t233 VSUBS 0.02fF
C3758 S.n959 VSUBS 0.23fF $ **FLOATING
C3759 S.n960 VSUBS 0.89fF $ **FLOATING
C3760 S.t311 VSUBS 0.04fF
C3761 S.t401 VSUBS 0.02fF
C3762 S.n961 VSUBS 0.01fF $ **FLOATING
C3763 S.t101 VSUBS 0.02fF
C3764 S.n962 VSUBS 1.25fF $ **FLOATING
C3765 S.t83 VSUBS 0.02fF
C3766 S.t306 VSUBS 0.02fF
C3767 S.t381 VSUBS 0.02fF
C3768 S.n963 VSUBS 0.02fF $ **FLOATING
C3769 S.t522 VSUBS 0.02fF
C3770 S.t103 VSUBS 0.02fF
C3771 S.t178 VSUBS 0.02fF
C3772 S.n964 VSUBS 0.02fF $ **FLOATING
C3773 S.t220 VSUBS 0.02fF
C3774 S.t483 VSUBS 0.02fF
C3775 S.n965 VSUBS 0.02fF $ **FLOATING
C3776 S.t615 VSUBS 0.02fF
C3777 S.t399 VSUBS 0.02fF
C3778 S.t60 VSUBS 0.02fF
C3779 S.n966 VSUBS 0.02fF $ **FLOATING
C3780 S.t194 VSUBS 0.02fF
C3781 S.t591 VSUBS 0.02fF
C3782 S.t219 VSUBS 0.02fF
C3783 S.n967 VSUBS 0.02fF $ **FLOATING
C3784 S.t379 VSUBS 0.02fF
C3785 S.t203 VSUBS 0.02fF
C3786 S.t427 VSUBS 0.02fF
C3787 S.n968 VSUBS 0.02fF $ **FLOATING
C3788 S.t123 VSUBS 0.02fF
C3789 S.t538 VSUBS 0.02fF
C3790 S.t606 VSUBS 0.02fF
C3791 S.n969 VSUBS 0.02fF $ **FLOATING
C3792 S.t318 VSUBS 0.02fF
C3793 S.t72 VSUBS 0.02fF
C3794 S.t496 VSUBS 0.02fF
C3795 S.n970 VSUBS 0.02fF $ **FLOATING
C3796 S.t286 VSUBS 0.02fF
C3797 S.t499 VSUBS 0.02fF
C3798 S.n971 VSUBS 15.72fF $ **FLOATING
C3799 S.n972 VSUBS 9.26fF $ **FLOATING
C3800 S.n973 VSUBS 0.03fF $ **FLOATING
C3801 S.n974 VSUBS 1.06fF $ **FLOATING
C3802 S.n975 VSUBS 0.03fF $ **FLOATING
C3803 S.n976 VSUBS 0.60fF $ **FLOATING
C3804 S.n977 VSUBS 0.41fF $ **FLOATING
C3805 S.n978 VSUBS 0.89fF $ **FLOATING
C3806 S.t475 VSUBS 0.02fF
C3807 S.n979 VSUBS 0.23fF $ **FLOATING
C3808 S.n980 VSUBS 0.12fF $ **FLOATING
C3809 S.t285 VSUBS 0.02fF
C3810 S.t546 VSUBS 0.02fF
C3811 S.n981 VSUBS 0.23fF $ **FLOATING
C3812 S.n982 VSUBS 0.89fF $ **FLOATING
C3813 S.t498 VSUBS 0.02fF
C3814 S.n983 VSUBS 0.12fF $ **FLOATING
C3815 S.n984 VSUBS 0.09fF $ **FLOATING
C3816 S.n985 VSUBS 0.24fF $ **FLOATING
C3817 S.n986 VSUBS 0.12fF $ **FLOATING
C3818 S.t468 VSUBS 0.02fF
C3819 S.n987 VSUBS 0.89fF $ **FLOATING
C3820 S.t51 VSUBS 0.02fF
C3821 S.n988 VSUBS 0.23fF $ **FLOATING
C3822 S.t115 VSUBS 0.02fF
C3823 S.n989 VSUBS 0.23fF $ **FLOATING
C3824 S.n990 VSUBS 0.89fF $ **FLOATING
C3825 S.t65 VSUBS 0.02fF
C3826 S.n991 VSUBS 0.12fF $ **FLOATING
C3827 S.n992 VSUBS 10.74fF $ **FLOATING
C3828 S.n993 VSUBS 0.89fF $ **FLOATING
C3829 S.t290 VSUBS 0.02fF
C3830 S.n994 VSUBS 0.23fF $ **FLOATING
C3831 S.n995 VSUBS 1.21fF $ **FLOATING
C3832 S.n996 VSUBS 0.12fF $ **FLOATING
C3833 S.t87 VSUBS 0.02fF
C3834 S.n997 VSUBS 0.20fF $ **FLOATING
C3835 S.n998 VSUBS 0.09fF $ **FLOATING
C3836 S.n999 VSUBS 0.20fF $ **FLOATING
C3837 S.n1000 VSUBS 0.06fF $ **FLOATING
C3838 S.t302 VSUBS 0.02fF
C3839 S.n1001 VSUBS 0.12fF $ **FLOATING
C3840 S.t354 VSUBS 0.02fF
C3841 S.n1002 VSUBS 0.23fF $ **FLOATING
C3842 S.n1003 VSUBS 0.89fF $ **FLOATING
C3843 S.n1004 VSUBS 0.12fF $ **FLOATING
C3844 S.t229 VSUBS 0.02fF
C3845 S.t435 VSUBS 0.02fF
C3846 S.n1005 VSUBS 1.19fF $ **FLOATING
C3847 S.n1006 VSUBS 0.01fF $ **FLOATING
C3848 S.t237 VSUBS 0.02fF
C3849 S.t490 VSUBS 0.04fF
C3850 S.n1007 VSUBS 0.89fF $ **FLOATING
C3851 S.t619 VSUBS 0.02fF
C3852 S.n1008 VSUBS 0.23fF $ **FLOATING
C3853 S.n1009 VSUBS 0.12fF $ **FLOATING
C3854 S.t428 VSUBS 0.02fF
C3855 S.t68 VSUBS 0.02fF
C3856 S.n1010 VSUBS 0.23fF $ **FLOATING
C3857 S.n1011 VSUBS 0.89fF $ **FLOATING
C3858 S.t630 VSUBS 0.02fF
C3859 S.n1012 VSUBS 0.12fF $ **FLOATING
C3860 S.n1013 VSUBS 0.12fF $ **FLOATING
C3861 S.t607 VSUBS 0.02fF
C3862 S.n1014 VSUBS 0.89fF $ **FLOATING
C3863 S.t196 VSUBS 0.02fF
C3864 S.n1015 VSUBS 0.23fF $ **FLOATING
C3865 S.t270 VSUBS 0.02fF
C3866 S.n1016 VSUBS 0.23fF $ **FLOATING
C3867 S.n1017 VSUBS 0.89fF $ **FLOATING
C3868 S.t214 VSUBS 0.02fF
C3869 S.n1018 VSUBS 0.12fF $ **FLOATING
C3870 S.n1019 VSUBS 0.12fF $ **FLOATING
C3871 S.t165 VSUBS 0.02fF
C3872 S.n1020 VSUBS 0.89fF $ **FLOATING
C3873 S.t129 VSUBS 0.02fF
C3874 S.n1021 VSUBS 0.23fF $ **FLOATING
C3875 S.n1022 VSUBS 0.01fF $ **FLOATING
C3876 S.n1023 VSUBS 0.05fF $ **FLOATING
C3877 S.n1024 VSUBS 0.02fF $ **FLOATING
C3878 S.t479 VSUBS 0.02fF
C3879 S.n1025 VSUBS 0.23fF $ **FLOATING
C3880 S.n1026 VSUBS 0.89fF $ **FLOATING
C3881 S.t452 VSUBS 0.02fF
C3882 S.n1027 VSUBS 0.12fF $ **FLOATING
C3883 S.n1028 VSUBS 0.12fF $ **FLOATING
C3884 S.t289 VSUBS 0.02fF
C3885 S.n1029 VSUBS 0.89fF $ **FLOATING
C3886 S.t241 VSUBS 0.02fF
C3887 S.n1030 VSUBS 0.23fF $ **FLOATING
C3888 S.t502 VSUBS 0.02fF
C3889 S.n1031 VSUBS 0.12fF $ **FLOATING
C3890 S.t440 VSUBS 0.02fF
C3891 S.n1032 VSUBS 0.23fF $ **FLOATING
C3892 S.n1033 VSUBS 0.89fF $ **FLOATING
C3893 S.n1034 VSUBS 0.12fF $ **FLOATING
C3894 S.t470 VSUBS 0.02fF
C3895 S.n1035 VSUBS 0.89fF $ **FLOATING
C3896 S.t429 VSUBS 0.02fF
C3897 S.n1036 VSUBS 0.23fF $ **FLOATING
C3898 S.t67 VSUBS 0.02fF
C3899 S.n1037 VSUBS 0.12fF $ **FLOATING
C3900 S.t627 VSUBS 0.02fF
C3901 S.n1038 VSUBS 0.23fF $ **FLOATING
C3902 S.n1039 VSUBS 0.89fF $ **FLOATING
C3903 S.n1040 VSUBS 0.09fF $ **FLOATING
C3904 S.n1041 VSUBS 0.25fF $ **FLOATING
C3905 S.n1042 VSUBS 0.12fF $ **FLOATING
C3906 S.t48 VSUBS 0.02fF
C3907 S.n1043 VSUBS 0.89fF $ **FLOATING
C3908 S.t612 VSUBS 0.02fF
C3909 S.n1044 VSUBS 0.23fF $ **FLOATING
C3910 S.t268 VSUBS 0.02fF
C3911 S.n1045 VSUBS 0.12fF $ **FLOATING
C3912 S.t208 VSUBS 0.02fF
C3913 S.n1046 VSUBS 0.23fF $ **FLOATING
C3914 S.n1047 VSUBS 0.89fF $ **FLOATING
C3915 S.t402 VSUBS 0.02fF
C3916 S.n1048 VSUBS 0.12fF $ **FLOATING
C3917 S.t458 VSUBS 0.02fF
C3918 S.n1049 VSUBS 0.23fF $ **FLOATING
C3919 S.n1050 VSUBS 0.89fF $ **FLOATING
C3920 S.n1051 VSUBS 0.89fF $ **FLOATING
C3921 S.t378 VSUBS 0.02fF
C3922 S.n1052 VSUBS 0.23fF $ **FLOATING
C3923 S.n1053 VSUBS 0.12fF $ **FLOATING
C3924 S.t513 VSUBS 0.02fF
C3925 S.n1054 VSUBS 0.89fF $ **FLOATING
C3926 S.t455 VSUBS 0.02fF
C3927 S.n1055 VSUBS 0.23fF $ **FLOATING
C3928 S.t297 VSUBS 0.02fF
C3929 S.n1056 VSUBS 0.12fF $ **FLOATING
C3930 S.t44 VSUBS 0.02fF
C3931 S.n1057 VSUBS 0.23fF $ **FLOATING
C3932 S.n1058 VSUBS 0.89fF $ **FLOATING
C3933 S.n1059 VSUBS 0.89fF $ **FLOATING
C3934 S.t22 VSUBS 0.02fF
C3935 S.n1060 VSUBS 0.23fF $ **FLOATING
C3936 S.n1061 VSUBS 0.12fF $ **FLOATING
C3937 S.t81 VSUBS 0.02fF
C3938 S.n1062 VSUBS 0.89fF $ **FLOATING
C3939 S.t27 VSUBS 0.02fF
C3940 S.n1063 VSUBS 0.23fF $ **FLOATING
C3941 S.t253 VSUBS 0.02fF
C3942 S.n1064 VSUBS 0.23fF $ **FLOATING
C3943 S.n1065 VSUBS 0.89fF $ **FLOATING
C3944 S.t309 VSUBS 0.02fF
C3945 S.n1066 VSUBS 0.12fF $ **FLOATING
C3946 S.n1067 VSUBS 0.12fF $ **FLOATING
C3947 S.t82 VSUBS 0.02fF
C3948 S.t300 VSUBS 0.02fF
C3949 S.n1068 VSUBS 0.12fF $ **FLOATING
C3950 S.t250 VSUBS 0.02fF
C3951 S.n1069 VSUBS 0.23fF $ **FLOATING
C3952 S.n1070 VSUBS 0.89fF $ **FLOATING
C3953 S.n1071 VSUBS 0.12fF $ **FLOATING
C3954 S.t279 VSUBS 0.02fF
C3955 S.n1072 VSUBS 0.89fF $ **FLOATING
C3956 S.t234 VSUBS 0.02fF
C3957 S.n1073 VSUBS 0.23fF $ **FLOATING
C3958 S.t484 VSUBS 0.02fF
C3959 S.n1074 VSUBS 0.12fF $ **FLOATING
C3960 S.t336 VSUBS 0.02fF
C3961 S.n1075 VSUBS 0.23fF $ **FLOATING
C3962 S.n1076 VSUBS 0.89fF $ **FLOATING
C3963 S.n1077 VSUBS 0.12fF $ **FLOATING
C3964 S.t466 VSUBS 0.02fF
C3965 S.n1078 VSUBS 0.89fF $ **FLOATING
C3966 S.t423 VSUBS 0.02fF
C3967 S.n1079 VSUBS 0.23fF $ **FLOATING
C3968 S.t59 VSUBS 0.02fF
C3969 S.n1080 VSUBS 0.12fF $ **FLOATING
C3970 S.t623 VSUBS 0.02fF
C3971 S.n1081 VSUBS 0.23fF $ **FLOATING
C3972 S.n1082 VSUBS 0.89fF $ **FLOATING
C3973 S.n1083 VSUBS 0.09fF $ **FLOATING
C3974 S.n1084 VSUBS 0.25fF $ **FLOATING
C3975 S.n1085 VSUBS 0.12fF $ **FLOATING
C3976 S.t35 VSUBS 0.02fF
C3977 S.n1086 VSUBS 0.89fF $ **FLOATING
C3978 S.t605 VSUBS 0.02fF
C3979 S.n1087 VSUBS 0.23fF $ **FLOATING
C3980 S.t186 VSUBS 0.02fF
C3981 S.n1088 VSUBS 0.12fF $ **FLOATING
C3982 S.t201 VSUBS 0.02fF
C3983 S.n1089 VSUBS 0.23fF $ **FLOATING
C3984 S.n1090 VSUBS 0.89fF $ **FLOATING
C3985 S.t520 VSUBS 0.02fF
C3986 S.n1091 VSUBS 0.01fF $ **FLOATING
C3987 S.n1092 VSUBS 1.17fF $ **FLOATING
C3988 S.t516 VSUBS 0.02fF
C3989 S.t584 VSUBS 0.02fF
C3990 S.n1093 VSUBS 1.17fF $ **FLOATING
C3991 S.n1094 VSUBS 9.08fF $ **FLOATING
C3992 S.n1095 VSUBS 9.08fF $ **FLOATING
C3993 S.n1096 VSUBS 9.08fF $ **FLOATING
C3994 S.n1097 VSUBS 9.08fF $ **FLOATING
C3995 S.n1098 VSUBS 9.13fF $ **FLOATING
C3996 S.n1099 VSUBS 11.71fF $ **FLOATING
.ends

