* NGSPICE file created from nmos_36x36_flat.ext - technology: sky130A

.subckt nmos_36x36_flat
X0 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=3.50005e+15p pd=2.37328e+10u as=0p ps=0u w=4.38e+06u l=500000u
X1 D G S.t2581 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 D G S.t2580 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 D G S.t2578 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 S.t2577 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 D G S.t2576 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 S.t2575 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 S.t2574 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 S.t2573 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 D G S.t2572 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 D G S.t2571 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 D G S.t2570 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D G S.t2569 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 S.t2568 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 S.t2567 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 S.t2566 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 S.t2565 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 S.t2564 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 S.t2563 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 S.t2562 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 S.t2561 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 D G S.t2560 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D G S.t2559 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 D G S.t2558 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D G S.t2556 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 S.t2555 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D G S.t2554 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 S.t2553 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 S.t2552 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 S.t2551 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 S.t2550 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 S.t2549 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 D G S.t2548 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 D G S.t2547 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 D G S.t2546 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t2545 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 S.t2544 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 D G S.t2543 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D G S.t2542 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 D G S.t2541 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 S.t2540 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 D G S.t2539 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 S.t2538 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 D G S.t2537 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 S.t2536 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 S.t2535 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 S.t2534 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 S.t2533 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 D G S.t2532 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D G S.t2531 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 D G S.t2530 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 D G S.t2529 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 D G S.t2528 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 D G S.t2527 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 S.t2526 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 D G S.t2525 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 S.t2524 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 S.t2523 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 S.t2522 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 D G S.t2521 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 D G S.t2520 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 D G S.t2519 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 S.t2518 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 D G S.t2517 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 D G S.t2516 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 D G S.t2515 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 D G S.t2514 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 D G S.t2513 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 S.t2512 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D G S.t2511 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 D G S.t2510 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 D G S.t2509 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 S.t2508 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 S.t2507 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 D G S.t2506 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 S.t2505 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 S.t2504 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 D G S.t2503 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 D G S.t2502 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 S.t2501 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 D G S.t2500 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 S.t2498 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 S.t2497 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 S.t2496 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 S.t2495 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 S.t2494 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 D G S.t2493 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D G S.t2492 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 S.t2491 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 S.t2490 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 S.t2489 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 S.t2488 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 S.t2487 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D G S.t2486 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 D G S.t2484 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 D G S.t2483 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 D G S.t2482 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 S.t2481 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 D G S.t2480 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 D G S.t2479 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 S.t2478 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 S.t2477 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 S.t2476 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 S.t2475 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 S.t2474 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 D G S.t2473 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 S.t2472 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 D G S.t2471 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t2470 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 S.t2468 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 S.t2467 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 S.t2466 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 S.t2465 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 S.t2464 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 S.t2463 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 D G S.t2462 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 S.t2461 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 S.t2460 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 D G S.t2459 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 S.t2458 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 D G S.t2457 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 S.t2456 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 D G S.t2455 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 D G S.t2454 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 S.t2453 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 D G S.t2452 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 D G S.t2451 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t2449 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 S.t2448 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t2447 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 D G S.t2446 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 S.t2445 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 S.t2444 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 S.t2443 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 S.t2442 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 D G S.t2441 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 D G S.t2440 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 D G S.t2439 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 D G S.t2438 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 D G S.t2437 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 S.t2436 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 S.t2435 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 S.t2434 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 S.t2433 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 S.t2432 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 D G S.t2431 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 D G S.t2430 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 S.t2429 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 S.t2428 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 S.t2427 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 S.t2426 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 S.t2425 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 S.t2424 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 D G S.t2423 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 D G S.t2422 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 D G S.t2421 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 D G S.t2420 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 D G S.t2419 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 D G S.t2418 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 S.t2417 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 S.t2416 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 S.t2415 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 D G S.t2413 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 D G S.t2412 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 D G S.t2410 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 D G S.t2409 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 S.t2408 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 S.t2407 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 D G S.t2406 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 D G S.t2405 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 D G S.t2404 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 D G S.t2403 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 D G S.t2402 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 D G S.t2401 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 S.t2400 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 S.t2399 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 D G S.t2398 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 D G S.t2397 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 D G S.t2396 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 D G S.t2395 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 D G S.t2394 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 D G S.t2393 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 D G S.t2392 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 S.t2391 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 S.t2390 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 D G S.t2389 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 S.t2388 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 S.t2387 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 D G S.t2386 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 S.t2385 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 D G S.t2384 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 D G S.t2383 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 D G S.t2382 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 D G S.t2381 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 S.t2380 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 S.t2379 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 S.t2378 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 D G S.t2377 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 D G S.t2376 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 S.t2375 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 D G S.t2373 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 D G S.t2372 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 S.t2371 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 S.t2370 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 D G S.t2369 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 D G S.t2368 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 D G S.t2367 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 S.t2366 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 D G S.t2365 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 S.t2364 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 S.t2363 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 D G S.t2362 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 D G S.t2361 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 D G S.t2360 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 D G S.t2359 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 S.t2358 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 S.t2357 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 S.t2356 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 S.t2355 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 S.t2354 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 D G S.t2353 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 S.t2352 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 S.t2351 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 S.t2350 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 D G S.t2349 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 D G S.t2348 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 D G S.t2347 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 D G S.t2346 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 D G S.t2345 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 S.t2344 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 S.t2343 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 S.t2342 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 S.t2341 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 S.t2340 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 S.t2339 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 D G S.t2338 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 D G S.t2337 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 D G S.t2336 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 D G S.t2335 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 D G S.t2334 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 D G S.t2333 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 S.t2332 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 S.t2331 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 S.t2330 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 S.t2329 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 D G S.t2328 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 D G S.t2327 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 D G S.t2326 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 D G S.t2325 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 S.t2324 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 S.t2323 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 S.t2322 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 S.t2321 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 S.t2320 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 S.t2319 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 D G S.t2318 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 D G S.t2317 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 D G S.t2316 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 S.t2315 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 S.t2314 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 S.t2313 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 D G S.t2312 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 D G S.t2311 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 S.t2310 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 D G S.t2309 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 D G S.t2308 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 D G S.t2307 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 S.t2306 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 S.t2305 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 D G S.t2304 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 S.t2303 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 S.t2302 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 D G S.t2301 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 D G S.t2300 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D G S.t2299 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 D G S.t2298 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 D G S.t2297 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 D G S.t2296 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 D G S.t2295 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 S.t2294 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 S.t2293 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 S.t2291 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 S.t2290 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 D G S.t2289 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 D G S.t2288 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 D G S.t2286 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 D G S.t2285 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 S.t2284 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 S.t2283 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 S.t2282 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 D G S.t2281 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 S.t2280 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 D G S.t2279 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 S.t2278 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 D G S.t2277 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 D G S.t2276 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 D G S.t2275 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 D G S.t2274 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 S.t2273 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 S.t2272 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 D G S.t2271 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 D G S.t2270 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 S.t2269 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 D G S.t2268 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 D G S.t2267 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 D G S.t2266 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 S.t2265 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 S.t2264 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 S.t2263 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 S.t2262 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 D G S.t2261 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 S.t2260 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 D G S.t2259 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 S.t2258 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 S.t2257 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 S.t2256 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 S.t2255 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 S.t2254 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 S.t2253 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 D G S.t2252 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 D G S.t2251 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 D G S.t2250 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 S.t2249 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 D G S.t2248 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 D G S.t2247 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 S.t2246 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 S.t2245 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 S.t2244 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 D G S.t2243 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 D G S.t2242 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 S.t2241 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 S.t2240 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 S.t2239 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 D G S.t2238 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 S.t2237 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 D G S.t2236 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 S.t2235 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 S.t2234 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t2233 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 S.t2232 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 S.t2231 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 S.t2230 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 S.t2229 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 S.t2228 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 D G S.t2227 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 S.t2226 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 D G S.t2225 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 D G S.t2224 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 S.t2223 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 S.t2222 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 S.t2221 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 S.t2220 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 S.t2219 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 D G S.t2218 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 D G S.t2217 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 D G S.t2216 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 D G S.t2215 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 D G S.t2214 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 S.t2213 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 S.t2212 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 S.t2211 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 D G S.t2210 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 D G S.t2209 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 D G S.t2208 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 D G S.t2207 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 D G S.t2206 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 D G S.t2205 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 D G S.t2204 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 S.t2203 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 S.t2202 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 S.t2201 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 S.t2200 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 D G S.t2199 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 D G S.t2198 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 D G S.t2197 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 D G S.t2196 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 S.t2195 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 S.t2194 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 D G S.t2193 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 D G S.t2192 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 D G S.t2191 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 D G S.t2190 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 D G S.t2189 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 D G S.t2188 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 D G S.t2187 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 D G S.t2186 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 S.t2185 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 S.t2184 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 D G S.t2183 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 D G S.t2182 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 D G S.t2181 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 D G S.t2180 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 D G S.t2179 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 D G S.t2178 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 D G S.t2177 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 D G S.t2176 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 S.t2175 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 S.t2174 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 S.t2173 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 S.t2172 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 D G S.t2171 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 S.t2170 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 D G S.t2169 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 D G S.t2168 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 D G S.t2167 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 D G S.t2166 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 S.t2165 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 S.t2164 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 S.t2163 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 D G S.t2162 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 D G S.t2161 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 S.t2160 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 D G S.t2159 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 D G S.t2158 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 D G S.t2157 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 D G S.t2156 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 S.t2155 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 S.t2154 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 D G S.t2153 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 D G S.t2152 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 D G S.t2151 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 D G S.t2150 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 D G S.t2149 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 S.t2148 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 S.t2147 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 S.t2145 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 S.t2144 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 S.t2143 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 D G S.t2142 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 D G S.t2141 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 S.t2140 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 D G S.t2139 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 S.t2138 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 S.t2137 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 S.t2136 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 S.t2135 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 D G S.t2134 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 D G S.t2133 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 D G S.t2132 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 S.t2131 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 S.t2130 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 S.t2129 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 S.t2128 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 S.t2127 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 S.t2126 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 S.t2125 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 D G S.t2124 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 D G S.t2123 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 S.t2122 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 D G S.t2121 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 S.t2120 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t2119 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 S.t2118 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 S.t2117 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 S.t2116 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 S.t2115 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 D G S.t2114 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 D G S.t2113 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 D G S.t2112 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 S.t2110 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 S.t2109 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 S.t2108 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 S.t2107 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 S.t2106 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 D G S.t2105 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 D G S.t2104 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 S.t2103 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 D G S.t2102 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 D G S.t2101 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 S.t2100 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 S.t2099 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 S.t2098 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 S.t2097 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 S.t2096 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 S.t2095 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 D G S.t2094 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 D G S.t2093 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 D G S.t2092 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 D G S.t2091 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 S.t2090 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 S.t2089 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t2088 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 S.t2087 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 D G S.t2086 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 S.t2085 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 D G S.t2084 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 D G S.t2083 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 D G S.t2081 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 S.t2080 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 S.t2079 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 D G S.t2078 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 D G S.t2077 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 D G S.t2076 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 S.t2075 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 S.t2074 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 D G S.t2073 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t2072 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 S.t2071 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 S.t2070 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 D G S.t2069 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 D G S.t2066 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 D G S.t2065 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 D G S.t2064 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 S.t2063 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 S.t2062 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 S.t2061 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 S.t2060 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 D G S.t2059 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 D G S.t2058 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 S.t2057 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 D G S.t2056 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 S.t2055 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 S.t2054 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 S.t2053 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 S.t2052 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D G S.t2051 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 D G S.t2050 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 D G S.t2049 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 D G S.t2047 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 D G S.t2046 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 D G S.t2045 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 S.t2044 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 S.t2043 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 D G S.t2042 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 D G S.t2041 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 D G S.t2040 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 S.t2039 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 S.t2038 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t2037 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 D G S.t2035 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 D G S.t2034 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 S.t2033 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 D G S.t2032 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 S.t2031 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 S.t2030 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 D G S.t2029 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 D G S.t2028 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 D G S.t2027 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 D G S.t2026 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 S.t2025 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 D G S.t2024 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 S.t2023 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 S.t2022 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 S.t2021 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 S.t2020 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 S.t2019 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 S.t2018 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 D G S.t2017 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 D G S.t2016 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 D G S.t2015 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 S.t2014 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 S.t2013 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 S.t2012 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 S.t2011 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 S.t2010 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 S.t2009 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 D G S.t2008 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 D G S.t2007 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 D G S.t2006 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 D G S.t2005 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 S.t2004 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 S.t2003 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 S.t2002 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 S.t2001 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 D G S.t1999 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 D G S.t1998 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 S.t1997 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 S.t1996 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 S.t1995 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 S.t1994 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 S.t1993 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 S.t1992 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 D G S.t1991 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 D G S.t1990 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 S.t1989 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 D G S.t1988 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 D G S.t1987 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 S.t1986 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 D G S.t1985 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 S.t1984 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 S.t1983 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 D G S.t1982 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D G S.t1981 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 D G S.t1980 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 D G S.t1979 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 D G S.t1978 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 S.t1977 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 S.t1976 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 S.t1975 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 S.t1974 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 D G S.t1973 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 D G S.t1972 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 D G S.t1971 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 D G S.t1970 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 S.t1969 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 S.t1968 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 S.t1967 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 D G S.t1966 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 D G S.t1965 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 S.t1964 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 D G S.t1963 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 D G S.t1962 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 D G S.t1961 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 D G S.t1960 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 D G S.t1959 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 D G S.t1958 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 S.t1957 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 S.t1956 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 D G S.t1955 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 D G S.t1954 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 D G S.t1953 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 S.t1952 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 D G S.t1951 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 D G S.t1950 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 D G S.t1949 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 S.t1947 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 S.t1946 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 D G S.t1945 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 D G S.t1944 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 D G S.t1943 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 D G S.t1941 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 S.t1940 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 S.t1939 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 S.t1938 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 S.t1937 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 D G S.t1936 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 D G S.t1935 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 D G S.t1934 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 D G S.t1933 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 D G S.t1932 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 S.t1931 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 D G S.t1930 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 S.t1929 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 S.t1928 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 S.t1927 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 S.t1926 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 S.t1925 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 D G S.t1924 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 D G S.t1923 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 D G S.t1922 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 S.t1921 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 S.t1920 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 D G S.t1919 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 S.t1918 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 D G S.t1917 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 D G S.t1916 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 D G S.t1915 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 S.t1914 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 S.t1913 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 D G S.t1912 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 S.t1911 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 D G S.t1910 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 S.t1909 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 S.t1908 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 S.t1907 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 S.t1906 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 D G S.t1905 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 S.t1904 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 S.t1903 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 D G S.t1902 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 S.t1901 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 D G S.t1900 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 S.t1899 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 D G S.t1898 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 S.t1897 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 S.t1896 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 S.t1895 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 S.t1894 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 D G S.t1893 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 D G S.t1892 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 D G S.t1891 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 D G S.t1890 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 D G S.t1889 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 S.t1888 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 S.t1887 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 S.t1886 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 D G S.t1885 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 D G S.t1884 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 D G S.t1883 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 D G S.t1882 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 D G S.t1881 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 S.t1880 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 D G S.t1879 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 S.t1878 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 S.t1877 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 S.t1876 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 S.t1875 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 S.t1874 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 S.t1873 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 S.t1872 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 S.t1871 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 D G S.t1870 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 D G S.t1868 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 D G S.t1867 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 D G S.t1866 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 S.t1865 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 S.t1864 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 S.t1863 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 S.t1862 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 D G S.t1860 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 D G S.t1859 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 D G S.t1858 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 S.t1857 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 D G S.t1856 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 D G S.t1855 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 D G S.t1854 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 D G S.t1853 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 S.t1852 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 S.t1851 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 S.t1850 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 S.t1849 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 D G S.t1848 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 S.t1847 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 S.t1846 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 D G S.t1845 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 D G S.t1844 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 D G S.t1843 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 D G S.t1842 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 D G S.t1841 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 S.t1840 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 D G S.t1839 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 D G S.t1838 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 S.t1837 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 S.t1836 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 D G S.t1835 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 D G S.t1834 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 D G S.t1833 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 D G S.t1832 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 S.t1831 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 D G S.t1830 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 D G S.t1829 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 D G S.t1828 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 D G S.t1827 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 S.t1826 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 D G S.t1825 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 S.t1824 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 S.t1823 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 D G S.t1822 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 D G S.t1821 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 D G S.t1820 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 D G S.t1819 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 S.t1818 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 D G S.t1817 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 S.t1816 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 D G S.t1815 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 D G S.t1814 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 S.t1813 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 S.t1812 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 D G S.t1811 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 S.t1810 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 D G S.t1809 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 D G S.t1808 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 D G S.t1807 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 S.t1806 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 S.t1805 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 S.t1804 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 S.t1803 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 S.t1802 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 S.t1801 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 S.t1800 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 D G S.t1799 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 D G S.t1798 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 D G S.t1797 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 D G S.t1796 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 S.t1795 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 D G S.t1794 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 S.t1793 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 S.t1792 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 S.t1791 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 D G S.t1790 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 D G S.t1789 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 D G S.t1788 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 D G S.t1787 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 S.t1786 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 S.t1785 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 S.t1784 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 S.t1783 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 D G S.t1782 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 S.t1781 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 D G S.t1780 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 D G S.t1778 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 S.t1777 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 D G S.t1776 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 S.t1775 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 S.t1774 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 S.t1773 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 S.t1772 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 D G S.t1771 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 S.t1770 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 D G S.t1769 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 D G S.t1768 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 S.t1767 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 S.t1766 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 D G S.t1765 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 S.t1764 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 D G S.t1763 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 S.t1762 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 D G S.t1761 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 D G S.t1760 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 S.t1759 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 D G S.t1758 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 S.t1757 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 D G S.t1756 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 S.t1755 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 S.t1754 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 D G S.t1753 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 S.t1752 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 S.t1751 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 S.t1750 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 D G S.t1749 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 D G S.t1748 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 D G S.t1747 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 D G S.t1746 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 D G S.t1745 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 D G S.t1744 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 S.t1743 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 S.t1742 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 S.t1741 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 S.t1740 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 S.t1739 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 S.t1738 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 D G S.t1737 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 D G S.t1736 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 S.t1735 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 D G S.t1734 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 S.t1733 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 S.t1732 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 S.t1731 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 D G S.t1730 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 D G S.t1729 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 D G S.t1728 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 D G S.t1727 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 D G S.t1726 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 D G S.t1725 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 S.t1724 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 D G S.t1723 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 D G S.t1722 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 S.t1721 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 D G S.t1720 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 S.t1719 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 D G S.t1718 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 D G S.t1717 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 D G S.t1716 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 S.t1715 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 D G S.t1714 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 S.t1713 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 S.t1711 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 S.t1710 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 S.t1709 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 D G S.t1708 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 S.t1707 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 D G S.t1706 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 D G S.t1705 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 D G S.t1704 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 D G S.t1703 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 S.t1702 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 S.t1701 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 S.t1700 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 S.t1699 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 D G S.t1698 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 D G S.t1697 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 D G S.t1696 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 D G S.t1695 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 D G S.t1693 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 D G S.t1692 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 S.t1691 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 S.t1690 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 S.t1689 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 D G S.t1688 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 S.t1687 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 S.t1686 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 D G S.t1685 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 D G S.t1684 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 D G S.t1683 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 S.t1681 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 S.t1680 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 S.t1679 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 S.t1678 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 D G S.t1677 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 D G S.t1676 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 S.t1675 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 D G S.t1673 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 S.t1672 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 S.t1671 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 S.t1670 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 D G S.t1669 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 D G S.t1668 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 S.t1667 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 D G S.t1666 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 D G S.t1665 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 S.t1664 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 S.t1663 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 S.t1662 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 S.t1661 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 S.t1660 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 S.t1659 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 D G S.t1658 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 D G S.t1657 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 S.t1656 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 D G S.t1655 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 S.t1654 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 D G S.t1653 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 D G S.t1652 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 S.t1651 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 S.t1650 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 S.t1649 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 S.t1648 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 D G S.t1647 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 D G S.t1646 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 S.t1645 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 S.t1644 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 D G S.t1643 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 S.t1642 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 S.t1641 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 S.t1640 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 D G S.t1639 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 D G S.t1638 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 D G S.t1637 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 D G S.t1636 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 S.t1635 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 D G S.t1634 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 D G S.t1633 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 S.t1632 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 S.t1631 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 D G S.t1630 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 S.t1629 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 S.t1628 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 D G S.t1626 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 D G S.t1625 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 D G S.t1623 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 D G S.t1622 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 S.t1621 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 S.t1620 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 D G S.t1619 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 D G S.t1618 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 D G S.t1617 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 D G S.t1616 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 D G S.t1615 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 S.t1614 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 S.t1613 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 S.t1612 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 D G S.t1611 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 S.t1610 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 D G S.t1609 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 D G S.t1608 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 D G S.t1607 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 D G S.t1606 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 D G S.t1605 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 D G S.t1604 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 D G S.t1603 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 S.t1602 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 D G S.t1601 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 S.t1600 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 S.t1599 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 D G S.t1598 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 D G S.t1597 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 S.t1596 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 D G S.t1595 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 D G S.t1594 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 D G S.t1593 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 D G S.t1592 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 S.t1591 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 D G S.t1590 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 S.t1589 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 S.t1588 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 D G S.t1587 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 D G S.t1586 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 S.t1585 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 D G S.t1583 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 S.t1582 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 D G S.t1581 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 S.t1580 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 D G S.t1579 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 S.t1578 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 S.t1577 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 D G S.t1576 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 D G S.t1575 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 D G S.t1574 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 D G S.t1573 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 S.t1572 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 S.t1571 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 D G S.t1570 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 D G S.t1569 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 S.t1568 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 S.t1567 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 D G S.t1566 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 D G S.t1565 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 D G S.t1564 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 D G S.t1563 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 S.t1562 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 D G S.t1561 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 S.t1560 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 D G S.t1559 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 D G S.t1558 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 D G S.t1557 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 S.t1556 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 S.t1555 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 S.t1554 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 S.t1553 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 S.t1552 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 S.t1551 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 D G S.t1550 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 D G S.t1549 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 D G S.t1548 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 S.t1547 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 S.t1546 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 S.t1545 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 S.t1544 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 D G S.t1543 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 S.t1542 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 S.t1541 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 D G S.t1540 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 S.t1539 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 S.t1538 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 S.t1537 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 S.t1536 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 S.t1535 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 S.t1534 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 S.t1533 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 D G S.t1532 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 D G S.t1531 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 S.t1530 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 S.t1529 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 S.t1528 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 S.t1527 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 S.t1526 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 S.t1525 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 D G S.t1524 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 S.t1523 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 S.t1522 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 D G S.t1521 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 D G S.t1520 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 D G S.t1519 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 D G S.t1518 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 S.t1517 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 D G S.t1516 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 S.t1515 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 S.t1514 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 D G S.t1513 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 D G S.t1512 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 D G S.t1511 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 D G S.t1510 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 D G S.t1509 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 S.t1508 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 S.t1507 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 S.t1506 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 D G S.t1505 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 S.t1504 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 D G S.t1503 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 S.t1502 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 D G S.t1501 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 D G S.t1499 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 S.t1498 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 S.t1497 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 S.t1496 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 D G S.t1495 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 D G S.t1494 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 D G S.t1493 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 S.t1492 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 D G S.t1491 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 S.t1490 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 S.t1489 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 D G S.t1488 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 D G S.t1487 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 D G S.t1486 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 D G S.t1485 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 D G S.t1484 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 D G S.t1483 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 S.t1482 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 S.t1481 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 S.t1480 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 D G S.t1479 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1104 S.t1478 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1105 S.t1477 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1106 D G S.t1476 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1107 D G S.t1475 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1108 D G S.t1474 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1109 D G S.t1473 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1110 D G S.t1472 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1111 S.t1471 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1112 S.t1470 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1113 S.t1469 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1114 S.t1468 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1115 S.t1467 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1116 S.t1466 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1117 S.t1465 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1118 D G S.t1464 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1119 D G S.t1463 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1120 D G S.t1462 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1121 D G S.t1461 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1122 D G S.t1460 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1123 D G S.t1459 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1124 S.t1458 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1125 S.t1457 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1126 S.t1456 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1127 S.t1455 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1128 D G S.t1454 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1129 D G S.t1453 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1130 S.t1452 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1131 S.t1451 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1132 D G S.t1450 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1133 D G S.t1449 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1134 D G S.t1448 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1135 D G S.t1447 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1136 D G S.t1446 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1137 D G S.t1445 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1138 S.t1444 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1139 S.t1443 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1140 S.t1442 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1141 S.t1441 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1142 S.t1440 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1143 S.t1439 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1144 S.t1438 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1145 D G S.t1437 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1146 S.t1436 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1147 D G S.t1435 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1148 D G S.t1434 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1149 S.t1433 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1150 S.t1432 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1151 S.t1431 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1152 S.t1430 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1153 S.t1429 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1154 D G S.t1428 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1155 D G S.t1427 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1156 D G S.t1426 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1157 D G S.t1425 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1158 S.t1424 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1159 S.t1423 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1160 S.t1422 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1161 S.t1421 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1162 D G S.t1420 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1163 D G S.t1419 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1164 D G S.t1418 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1165 S.t1417 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1166 S.t1416 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1167 S.t1415 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1168 D G S.t1414 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1169 S.t1413 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1170 S.t1412 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1171 S.t1411 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1172 D G S.t1410 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1173 D G S.t1409 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1174 D G S.t1408 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1175 S.t1407 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1176 S.t1406 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1177 S.t1405 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1178 S.t1404 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1179 D G S.t1403 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1180 D G S.t1402 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1181 D G S.t1401 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1182 D G S.t1400 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1183 D G S.t1399 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1184 D G S.t1398 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1185 S.t1397 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1186 S.t1396 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1187 D G S.t1395 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1188 D G S.t1394 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1189 D G S.t1393 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1190 D G S.t1392 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1191 D G S.t1391 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1192 D G S.t1390 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1193 D G S.t1389 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1194 S.t1388 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1195 S.t1387 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1196 D G S.t1386 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1197 S.t1385 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1198 D G S.t1384 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1199 S.t1383 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1200 D G S.t1382 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1201 D G S.t1381 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1202 D G S.t1380 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1203 S.t1379 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1204 S.t1378 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1205 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1206 D G S.t1376 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1207 D G S.t1375 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1208 D G S.t1374 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1209 D G S.t1373 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1210 S.t1372 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1211 D G S.t1371 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1212 S.t1370 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1213 D G S.t1369 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1214 D G S.t1368 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1215 D G S.t1367 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1216 D G S.t1366 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1217 D G S.t1365 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1218 D G S.t1364 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1219 D G S.t1363 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1220 S.t1362 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1221 S.t1361 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1222 S.t1360 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1223 S.t1359 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1224 S.t1358 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1225 D G S.t1357 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1226 D G S.t1356 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1227 D G S.t1355 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1228 D G S.t1354 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1229 D G S.t1353 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1230 D G S.t1352 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1231 S.t1351 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1232 S.t1350 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1233 S.t1349 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1234 S.t1348 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1235 D G S.t1347 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1236 D G S.t1346 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1237 D G S.t1345 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1238 S.t1344 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1239 S.t1343 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1240 S.t1342 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1241 S.t1341 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1242 S.t1340 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1243 S.t1339 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1244 D G S.t1338 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1245 D G S.t1337 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1246 S.t1336 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1247 D G S.t1335 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1248 D G S.t1334 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1249 S.t1333 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1250 S.t1332 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1251 S.t1331 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1252 S.t1330 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1253 S.t1329 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1254 D G S.t1328 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1255 S.t1327 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1256 D G S.t1326 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1257 S.t1325 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1258 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1259 S.t1323 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1260 S.t1322 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1261 S.t1321 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1262 S.t1320 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1263 S.t1319 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1264 S.t1318 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1265 D G S.t1317 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1266 D G S.t1316 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1267 D G S.t1315 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1268 S.t1314 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1269 S.t1313 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1270 S.t1312 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1271 S.t1311 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1272 S.t1310 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1273 S.t1309 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1274 S.t1308 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1275 D G S.t1307 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1276 D G S.t1306 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1277 D G S.t1305 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1278 D G S.t1304 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1279 D G S.t1303 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1280 S.t1302 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1281 S.t1301 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1282 S.t1300 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1283 S.t1299 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1284 D G S.t1298 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1285 D G S.t1297 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1286 D G S.t1296 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1287 D G S.t1295 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1288 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1289 S.t1293 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1290 D G S.t1292 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1291 S.t1291 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1292 S.t1290 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1293 S.t1289 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1294 D G S.t1288 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1295 S.t1287 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1296 D G S.t1286 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1297 S.t1285 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1298 S.t1284 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1299 D G S.t1283 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1300 D G S.t1282 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1301 S.t1281 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1302 D G S.t1280 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1303 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1304 D G S.t1278 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1305 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1306 D G S.t1276 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1307 S.t1275 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1308 S.t1274 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1309 S.t1273 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1310 D G S.t1272 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1311 D G S.t1271 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1312 D G S.t1270 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1313 D G S.t1269 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1314 D G S.t1268 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1315 S.t1267 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1316 S.t1266 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1317 S.t1265 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1318 S.t1264 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1319 D G S.t1263 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1320 D G S.t1262 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1321 D G S.t1261 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1322 D G S.t1260 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1323 D G S.t1259 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1324 D G S.t1258 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1325 D G S.t1257 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1326 S.t1256 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1327 S.t1255 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1328 S.t1254 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1329 D G S.t1253 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1330 D G S.t1252 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1331 D G S.t1251 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1332 D G S.t1250 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1333 D G S.t1249 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1334 D G S.t1248 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1335 S.t1247 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1336 S.t1246 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1337 S.t1245 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1338 D G S.t1244 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1339 D G S.t1243 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1340 D G S.t1242 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1341 D G S.t1241 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1342 S.t1240 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1343 S.t1239 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1344 S.t1238 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1345 S.t1237 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1346 D G S.t1236 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1347 D G S.t1235 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1348 D G S.t1234 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1349 S.t1233 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1350 S.t1232 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1351 S.t1231 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1352 D G S.t1230 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1353 D G S.t1229 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1354 S.t1228 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1355 S.t1227 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1356 S.t1226 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1357 D G S.t1225 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1358 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1359 S.t1223 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1360 D G S.t1222 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1361 D G S.t1221 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1362 S.t1220 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1363 D G S.t1219 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1364 S.t1218 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1365 D G S.t1217 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1366 S.t1216 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1367 S.t1215 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1368 S.t1214 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1369 D G S.t1213 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1370 S.t1212 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1371 D G S.t1211 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1372 D G S.t1210 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1373 S.t1209 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1374 S.t1208 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1375 D G S.t1207 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1376 S.t1206 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1377 S.t1205 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1378 D G S.t1204 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1379 S.t1203 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1380 D G S.t1202 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1381 D G S.t1201 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1382 D G S.t1200 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1383 D G S.t1199 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1384 D G S.t1198 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1385 S.t1197 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1386 S.t1196 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1387 S.t1195 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1388 S.t1194 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1389 S.t1193 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1390 D G S.t1192 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1391 D G S.t1191 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1392 D G S.t1190 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1393 D G S.t1189 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1394 D G S.t1188 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1395 S.t1187 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1396 S.t1186 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1397 S.t1185 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1398 S.t1184 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1399 D G S.t1183 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1400 D G S.t1182 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1401 S.t1181 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1402 S.t1180 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1403 S.t1179 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1404 S.t1178 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1405 D G S.t1177 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1406 D G S.t1176 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1407 S.t1175 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1408 D G S.t1174 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1409 D G S.t1173 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1410 S.t1172 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1411 S.t1171 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1412 D G S.t1170 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1413 S.t1169 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1414 D G S.t1168 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1415 D G S.t1167 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1416 D G S.t1166 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1417 S.t1165 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1418 D G S.t1164 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1419 S.t1163 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1420 D G S.t1162 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1421 D G S.t1161 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1422 D G S.t1160 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1423 D G S.t1159 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1424 D G S.t1158 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1425 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1426 S.t1156 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1427 S.t1155 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1428 D G S.t1154 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1429 D G S.t1153 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1430 D G S.t1152 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1431 D G S.t1151 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1432 D G S.t1150 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1433 D G S.t1149 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1434 D G S.t1148 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1435 S.t1147 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1436 S.t1146 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1437 S.t1145 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1438 S.t1144 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1439 D G S.t1143 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1440 D G S.t1142 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1441 D G S.t1141 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1442 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1443 S.t1139 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1444 D G S.t1138 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1445 S.t1137 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1446 S.t1136 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1447 D G S.t1135 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1448 D G S.t1134 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1449 D G S.t1133 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1450 D G S.t1132 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1451 S.t1131 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1452 D G S.t1130 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1453 S.t1129 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1454 D G S.t1128 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1455 D G S.t1127 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1456 S.t1126 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1457 S.t1125 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1458 S.t1124 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1459 D G S.t1123 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1460 S.t1122 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1461 S.t1121 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1462 D G S.t1120 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1463 S.t1119 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1464 S.t1118 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1465 D G S.t1117 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1466 S.t1116 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1467 S.t1115 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1468 S.t1114 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1469 D G S.t1113 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1470 D G S.t1112 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1471 S.t1111 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1472 S.t1110 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1473 S.t1109 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1474 S.t1108 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1475 S.t1107 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1476 S.t1106 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1477 D G S.t1105 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1478 D G S.t1104 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1479 D G S.t1103 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1480 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1481 D G S.t1101 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1482 S.t1100 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1483 D G S.t1099 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1484 S.t1098 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1485 S.t1097 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1486 S.t1096 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1487 S.t1095 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1488 S.t1094 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1489 S.t1093 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1490 S.t1092 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1491 S.t1091 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1492 S.t1090 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1493 S.t1089 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1494 D G S.t1088 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1495 D G S.t1087 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1496 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1497 S.t1085 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1498 D G S.t1084 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1499 S.t1083 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1500 S.t1082 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1501 S.t1081 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1502 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1503 D G S.t1079 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1504 D G S.t1078 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1505 D G S.t1077 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1506 S.t1076 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1507 S.t1075 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1508 S.t1074 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1509 D G S.t1073 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1510 S.t1072 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1511 D G S.t1071 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1512 D G S.t1070 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1513 D G S.t1069 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1514 D G S.t1068 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1515 S.t1067 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1516 S.t1066 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1517 S.t1065 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1518 S.t1064 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1519 D G S.t1063 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1520 S.t1062 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1521 S.t1061 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1522 D G S.t1060 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1523 D G S.t1059 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1524 D G S.t1058 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1525 D G S.t1057 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1526 D G S.t1056 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1527 S.t1055 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1528 S.t1054 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1529 S.t1053 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1530 S.t1052 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1531 D G S.t1051 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1532 D G S.t1050 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1533 D G S.t1049 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1534 S.t1048 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1535 D G S.t1047 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1536 S.t1046 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1537 D G S.t1045 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1538 S.t1044 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1539 S.t1043 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1540 D G S.t1042 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1541 D G S.t1041 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1542 D G S.t1040 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1543 D G S.t1039 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1544 D G S.t1038 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1545 S.t1037 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1546 D G S.t1036 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1547 D G S.t1035 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1548 S.t1034 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1549 S.t1033 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1550 D G S.t1032 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1551 S.t1031 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1552 D G S.t1030 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1553 D G S.t1029 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1554 D G S.t1028 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1555 D G S.t1027 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1556 D G S.t1026 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1557 S.t1025 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1558 S.t1024 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1559 S.t1023 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1560 S.t1022 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1561 D G S.t1021 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1562 D G S.t1020 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1563 D G S.t1019 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1564 D G S.t1018 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1565 S.t1017 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1566 S.t1016 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1567 S.t1015 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1568 S.t1014 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1569 S.t1013 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1570 D G S.t1012 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1571 S.t1011 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1572 D G S.t1010 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1573 D G S.t1009 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1574 D G S.t1008 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1575 D G S.t1007 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1576 D G S.t1006 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1577 D G S.t1005 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1578 S.t1004 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1579 D G S.t1003 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1580 S.t1002 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1581 S.t1001 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1582 D G S.t1000 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1583 S.t999 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1584 S.t998 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1585 D G S.t997 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1586 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1587 S.t995 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1588 S.t994 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1589 D G S.t993 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1590 S.t992 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1591 S.t991 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1592 D G S.t990 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1593 S.t989 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1594 S.t988 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1595 D G S.t987 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1596 S.t986 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1597 S.t985 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1598 S.t984 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1599 S.t983 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1600 S.t982 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1601 D G S.t981 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1602 D G S.t980 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1603 D G S.t979 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1604 D G S.t978 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1605 S.t977 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1606 D G S.t976 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1607 D G S.t975 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1608 S.t974 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1609 S.t973 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1610 S.t972 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1611 S.t971 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1612 D G S.t970 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1613 S.t969 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1614 S.t968 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1615 S.t967 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1616 D G S.t966 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1617 D G S.t965 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1618 D G S.t964 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1619 D G S.t963 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1620 S.t962 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1621 S.t961 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1622 S.t960 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1623 S.t959 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1624 S.t958 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1625 S.t957 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1626 S.t956 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1627 S.t955 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1628 D G S.t954 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1629 D G S.t953 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1630 D G S.t952 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1631 S.t951 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1632 S.t950 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1633 S.t949 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1634 S.t948 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1635 D G S.t947 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1636 S.t946 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1637 D G S.t945 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1638 D G S.t944 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1639 D G S.t943 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1640 S.t942 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1641 D G S.t941 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1642 S.t940 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1643 D G S.t939 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1644 D G S.t938 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1645 D G S.t937 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1646 D G S.t936 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1647 D G S.t935 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1648 S.t934 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1649 S.t933 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1650 S.t932 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1651 D G S.t931 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1652 S.t930 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1653 D G S.t929 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1654 D G S.t928 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1655 D G S.t927 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1656 S.t926 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1657 S.t925 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1658 S.t924 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1659 S.t923 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1660 S.t922 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1661 S.t921 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1662 S.t920 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1663 S.t919 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1664 D G S.t918 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1665 D G S.t917 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1666 D G S.t916 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1667 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1668 D G S.t914 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1669 D G S.t913 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1670 D G S.t912 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1671 S.t911 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1672 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1673 S.t909 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1674 D G S.t908 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1675 S.t907 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1676 D G S.t906 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1677 D G S.t905 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1678 D G S.t904 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1679 D G S.t903 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1680 S.t902 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1681 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1682 S.t900 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1683 S.t899 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1684 D G S.t898 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1685 D G S.t897 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1686 S.t896 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1687 D G S.t895 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1688 S.t894 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1689 D G S.t893 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1690 S.t892 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1691 S.t891 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1692 D G S.t890 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1693 D G S.t889 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1694 S.t888 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1695 D G S.t887 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1696 D G S.t886 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1697 S.t885 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1698 D G S.t884 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1699 D G S.t883 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1700 S.t882 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1701 S.t881 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1702 S.t880 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1703 S.t879 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1704 D G S.t878 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1705 S.t877 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1706 D G S.t876 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1707 S.t875 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1708 S.t874 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1709 D G S.t873 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1710 D G S.t872 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1711 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1712 D G S.t870 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1713 D G S.t869 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1714 D G S.t868 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1715 S.t867 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1716 S.t866 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1717 S.t865 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1718 D G S.t864 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1719 S.t863 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1720 S.t862 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1721 S.t861 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1722 S.t860 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1723 D G S.t859 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1724 S.t858 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1725 S.t857 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1726 D G S.t856 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1727 D G S.t855 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1728 S.t854 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1729 D G S.t853 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1730 D G S.t852 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1731 S.t851 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1732 S.t850 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1733 S.t849 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1734 S.t848 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1735 S.t847 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1736 D G S.t846 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1737 D G S.t845 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1738 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1739 D G S.t843 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1740 D G S.t842 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1741 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1742 S.t840 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1743 D G S.t839 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1744 S.t838 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1745 D G S.t837 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1746 D G S.t836 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1747 D G S.t835 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1748 D G S.t834 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1749 D G S.t833 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1750 S.t832 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1751 S.t831 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1752 S.t830 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1753 S.t829 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1754 S.t828 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1755 S.t827 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1756 D G S.t826 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1757 D G S.t825 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1758 D G S.t824 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1759 D G S.t823 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1760 D G S.t822 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1761 D G S.t821 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1762 S.t820 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1763 D G S.t819 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1764 S.t818 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1765 S.t817 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1766 D G S.t816 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1767 S.t815 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1768 D G S.t814 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1769 D G S.t813 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1770 D G S.t812 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1771 D G S.t811 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1772 D G S.t810 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1773 D G S.t809 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1774 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1775 S.t807 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1776 D G S.t806 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1777 D G S.t805 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1778 D G S.t804 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1779 S.t803 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1780 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1781 D G S.t801 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1782 S.t800 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1783 S.t799 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1784 S.t798 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1785 D G S.t797 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1786 S.t796 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1787 D G S.t795 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1788 D G S.t794 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1789 D G S.t793 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1790 D G S.t792 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1791 D G S.t791 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1792 S.t790 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1793 D G S.t789 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1794 D G S.t788 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1795 D G S.t787 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1796 S.t786 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1797 S.t785 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1798 D G S.t784 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1799 S.t783 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1800 D G S.t782 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1801 D G S.t781 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1802 D G S.t780 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1803 D G S.t779 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1804 D G S.t778 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1805 S.t777 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1806 S.t776 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1807 D G S.t775 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1808 D G S.t774 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1809 S.t773 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1810 D G S.t772 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1811 D G S.t771 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1812 D G S.t770 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1813 D G S.t769 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1814 S.t768 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1815 S.t767 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1816 S.t766 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1817 S.t765 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1818 D G S.t764 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1819 S.t763 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1820 S.t762 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1821 D G S.t761 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1822 S.t760 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1823 S.t759 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1824 D G S.t758 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1825 D G S.t757 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1826 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1827 D G S.t755 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1828 S.t754 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1829 S.t753 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1830 S.t752 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1831 S.t751 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1832 S.t750 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1833 D G S.t749 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1834 D G S.t748 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1835 S.t747 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1836 S.t746 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1837 S.t745 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1838 S.t744 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1839 S.t743 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1840 S.t742 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1841 S.t741 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1842 D G S.t740 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1843 D G S.t739 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1844 S.t738 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1845 S.t737 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1846 S.t736 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1847 S.t735 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1848 S.t734 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1849 S.t733 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1850 D G S.t732 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1851 D G S.t731 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1852 S.t730 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1853 D G S.t729 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1854 D G S.t728 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1855 D G S.t727 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1856 S.t726 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1857 S.t725 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1858 S.t724 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1859 S.t723 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1860 S.t722 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1861 S.t721 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1862 D G S.t720 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1863 D G S.t719 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1864 S.t718 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1865 D G S.t717 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1866 S.t716 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1867 D G S.t715 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1868 S.t714 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1869 S.t713 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1870 D G S.t712 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1871 D G S.t711 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1872 S.t710 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1873 S.t709 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1874 D G S.t708 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1875 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1876 S.t706 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1877 S.t705 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1878 D G S.t704 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1879 D G S.t703 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1880 S.t702 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1881 S.t701 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1882 D G S.t700 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1883 D G S.t699 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1884 S.t698 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1885 S.t697 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1886 S.t696 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1887 D G S.t695 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1888 D G S.t694 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1889 D G S.t693 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1890 S.t692 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1891 S.t691 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1892 S.t690 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1893 D G S.t689 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1894 D G S.t688 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1895 S.t687 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1896 D G S.t686 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1897 D G S.t685 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1898 D G S.t684 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1899 D G S.t683 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1900 D G S.t682 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1901 S.t681 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1902 S.t680 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1903 S.t679 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1904 S.t678 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1905 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1906 D G S.t676 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1907 D G S.t675 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1908 D G S.t674 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1909 D G S.t673 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1910 D G S.t672 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1911 S.t671 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1912 S.t670 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1913 S.t669 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1914 D G S.t668 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1915 D G S.t667 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1916 D G S.t666 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1917 D G S.t665 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1918 D G S.t664 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1919 D G S.t663 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1920 S.t662 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1921 S.t661 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1922 D G S.t660 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1923 S.t659 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1924 D G S.t658 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1925 D G S.t657 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1926 D G S.t656 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1927 D G S.t655 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1928 S.t654 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1929 S.t653 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1930 D G S.t652 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1931 S.t651 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1932 S.t650 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1933 D G S.t649 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1934 S.t648 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1935 S.t647 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1936 D G S.t646 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1937 S.t645 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1938 S.t644 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1939 S.t643 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1940 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1941 D G S.t641 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1942 D G S.t640 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1943 S.t639 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1944 D G S.t638 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1945 D G S.t637 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1946 S.t636 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1947 S.t635 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1948 D G S.t634 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1949 D G S.t633 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1950 S.t632 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1951 D G S.t631 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1952 D G S.t630 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1953 D G S.t629 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1954 D G S.t628 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1955 S.t627 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1956 D G S.t626 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1957 D G S.t625 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1958 S.t624 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1959 S.t623 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1960 S.t622 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1961 S.t621 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1962 D G S.t620 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1963 S.t619 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1964 S.t618 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1965 D G S.t617 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1966 S.t616 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1967 S.t615 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1968 S.t614 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1969 D G S.t613 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1970 D G S.t612 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1971 D G S.t611 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1972 D G S.t610 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1973 D G S.t609 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1974 D G S.t608 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1975 S.t607 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1976 S.t606 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1977 S.t605 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1978 S.t604 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1979 D G S.t603 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1980 S.t602 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1981 D G S.t601 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1982 D G S.t600 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1983 D G S.t599 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1984 D G S.t598 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1985 D G S.t597 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1986 S.t596 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1987 S.t595 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1988 S.t594 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1989 S.t593 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1990 D G S.t592 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1991 S.t591 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1992 D G S.t590 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1993 D G S.t589 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1994 D G S.t588 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1995 S.t587 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1996 S.t586 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1997 S.t585 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1998 S.t584 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1999 D G S.t583 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2000 D G S.t582 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2001 D G S.t581 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2002 S.t580 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2003 D G S.t579 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2004 D G S.t578 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2005 D G S.t577 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2006 D G S.t576 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2007 D G S.t575 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2008 D G S.t574 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2009 S.t573 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2010 S.t572 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2011 S.t571 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2012 D G S.t570 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2013 D G S.t569 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2014 D G S.t568 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2015 D G S.t567 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2016 D G S.t566 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2017 D G S.t565 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2018 D G S.t564 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2019 S.t563 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2020 S.t562 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2021 S.t561 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2022 S.t560 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2023 S.t559 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2024 D G S.t558 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2025 D G S.t557 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2026 S.t556 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2027 S.t555 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2028 S.t554 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2029 S.t553 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2030 S.t552 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2031 D G S.t551 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2032 D G S.t550 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2033 S.t549 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2034 D G S.t548 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2035 D G S.t547 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2036 D G S.t546 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2037 S.t545 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2038 S.t544 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2039 S.t543 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2040 S.t542 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2041 S.t541 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2042 D G S.t540 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2043 D G S.t539 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2044 S.t538 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2045 S.t537 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2046 D G S.t536 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2047 S.t535 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2048 S.t534 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2049 S.t533 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2050 S.t532 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2051 S.t531 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2052 D G S.t530 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2053 S.t529 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2054 S.t528 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2055 S.t527 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2056 S.t526 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2057 S.t525 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2058 S.t524 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2059 S.t523 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2060 S.t522 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2061 S.t521 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2062 D G S.t520 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2063 D G S.t519 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2064 D G S.t518 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2065 D G S.t517 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2066 S.t516 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2067 S.t515 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2068 S.t514 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2069 S.t513 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2070 D G S.t512 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2071 D G S.t511 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2072 S.t510 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2073 S.t509 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2074 S.t508 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2075 S.t507 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2076 D G S.t506 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2077 S.t505 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2078 S.t504 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2079 D G S.t503 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2080 D G S.t502 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2081 S.t501 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2082 S.t500 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2083 S.t499 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2084 S.t498 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2085 S.t497 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2086 S.t496 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2087 S.t495 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2088 D G S.t494 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2089 D G S.t493 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2090 D G S.t492 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2091 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2092 D G S.t490 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2093 S.t489 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2094 S.t488 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2095 S.t487 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2096 S.t486 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2097 S.t485 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2098 D G S.t484 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2099 D G S.t483 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2100 D G S.t482 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2101 D G S.t481 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2102 S.t480 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2103 S.t479 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2104 S.t478 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2105 S.t477 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2106 D G S.t476 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2107 D G S.t475 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2108 D G S.t474 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2109 D G S.t473 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2110 D G S.t472 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2111 D G S.t471 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2112 S.t470 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2113 D G S.t469 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2114 S.t468 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2115 S.t467 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2116 D G S.t466 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2117 D G S.t465 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2118 D G S.t464 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2119 D G S.t463 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2120 S.t462 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2121 D G S.t461 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2122 S.t460 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2123 S.t459 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2124 D G S.t458 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2125 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2126 D G S.t456 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2127 D G S.t455 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2128 D G S.t454 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2129 D G S.t453 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2130 D G S.t452 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2131 D G S.t451 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2132 S.t450 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2133 S.t449 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2134 S.t448 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2135 D G S.t447 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2136 D G S.t446 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2137 D G S.t445 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2138 D G S.t444 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2139 D G S.t443 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2140 D G S.t442 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2141 D G S.t441 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2142 S.t440 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2143 S.t439 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2144 S.t438 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2145 S.t437 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2146 D G S.t436 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2147 D G S.t435 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2148 D G S.t434 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2149 S.t433 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2150 D G S.t432 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2151 S.t431 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2152 S.t430 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2153 D G S.t429 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2154 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2155 S.t427 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2156 D G S.t426 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2157 D G S.t425 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2158 S.t424 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2159 S.t423 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2160 D G S.t422 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2161 S.t421 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2162 D G S.t420 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2163 D G S.t419 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2164 D G S.t418 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2165 S.t417 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2166 S.t416 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2167 S.t415 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2168 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2169 S.t413 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2170 S.t412 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2171 S.t411 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2172 D G S.t410 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2173 D G S.t409 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2174 D G S.t408 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2175 D G S.t407 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2176 S.t406 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2177 S.t405 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2178 S.t404 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2179 S.t403 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2180 D G S.t402 S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2181 S.t401 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2182 D G S.t400 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2183 D G S.t399 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2184 D G S.t398 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2185 D G S.t397 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2186 S.t396 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2187 S.t395 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2188 S.t394 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2189 S.t393 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2190 S.t392 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2191 D G S.t391 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2192 D G S.t390 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2193 S.t389 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2194 D G S.t388 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2195 S.t387 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2196 S.t386 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2197 S.t385 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2198 S.t384 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2199 S.t383 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2200 D G S.t382 S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2201 D G S.t381 S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2202 D G S.t380 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2203 D G S.t379 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2204 S.t378 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2205 S.t377 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2206 S.t376 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2207 D G S.t375 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2208 D G S.t374 S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2209 D G S.t373 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2210 D G S.t372 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2211 D G S.t371 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2212 S.t370 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2213 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2214 S.t368 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2215 D G S.t367 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2216 D G S.t366 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2217 D G S.t365 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2218 D G S.t364 S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2219 D G S.t363 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2220 S.t362 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2221 S.t361 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2222 S.t360 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2223 S.t359 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2224 S.t358 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2225 D G S.t357 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2226 D G S.t356 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2227 D G S.t355 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2228 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2229 D G S.t353 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2230 S.t352 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2231 S.t351 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2232 D G S.t350 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2233 S.t349 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2234 D G S.t348 S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2235 D G S.t347 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2236 D G S.t346 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2237 D G S.t345 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2238 D G S.t344 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2239 S.t343 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2240 S.t342 G D S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2241 D G S.t341 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2242 S.t340 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2243 S.t339 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2244 S.t338 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2245 D G S.t337 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2246 D G S.t336 S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2247 S.t335 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2248 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2249 D G S.t333 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2250 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2251 S.t331 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2252 D G S.t330 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2253 S.t329 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2254 S.t328 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2255 S.t327 G D S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2256 S.t326 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2257 D G S.t325 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2258 D G S.t324 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2259 D G S.t323 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2260 S.t322 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2261 S.t321 G D S.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2262 D G S.t319 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2263 S.t318 G D S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2264 S.t317 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2265 D G S.t316 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2266 D G S.t315 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2267 D G S.t314 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2268 D G S.t313 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2269 S.t312 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2270 S.t311 G D S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2271 S.t310 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2272 D G S.t309 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2273 S.t308 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2274 S.t307 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2275 S.t306 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2276 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2277 D G S.t304 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2278 S.t303 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2279 S.t302 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2280 S.t301 G D S.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2281 D G S.t299 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2282 S.t298 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2283 D G S.t297 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2284 D G S.t296 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2285 S.t295 G D S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2286 S.t294 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2287 S.t293 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2288 S.t292 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2289 S.t291 G D S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2290 S.t290 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2291 D G S.t289 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2292 D G S.t288 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2293 D G S.t287 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2294 S.t286 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2295 S.t285 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2296 S.t284 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2297 S.t283 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2298 D G S.t282 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2299 S.t281 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2300 D G S.t280 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2301 D G S.t279 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2302 D G S.t278 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2303 D G S.t277 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2304 D G S.t276 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2305 S.t275 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2306 S.t274 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2307 S.t273 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2308 S.t272 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2309 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2310 D G S.t270 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2311 D G S.t269 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2312 S.t268 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2313 D G S.t267 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2314 D G S.t266 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2315 S.t265 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2316 S.t264 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2317 S.t263 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2318 D G S.t262 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2319 S.t261 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2320 D G S.t260 S.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2321 S.t258 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2322 S.t257 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2323 D G S.t256 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2324 D G S.t255 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2325 D G S.t254 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2326 S.t253 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2327 D G S.t252 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2328 D G S.t251 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2329 D G S.t250 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2330 D G S.t249 S.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2331 S.t247 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2332 D G S.t246 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2333 D G S.t245 S.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2334 D G S.t243 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2335 D G S.t242 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2336 D G S.t241 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2337 S.t240 G D S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2338 S.t239 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2339 S.t238 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2340 S.t237 G D S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2341 D G S.t236 S.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2342 D G S.t234 S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2343 D G S.t233 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2344 D G S.t232 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2345 S.t231 G D S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2346 S.t230 G D S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2347 S.t229 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2348 S.t228 G D S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2349 S.t227 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2350 D G S.t226 S.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2351 S.t224 G D S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2352 D G S.t223 S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2353 D G S.t222 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2354 D G S.t221 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2355 D G S.t220 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2356 D G S.t219 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2357 D G S.t218 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2358 D G S.t217 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2359 D G S.t216 S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2360 D G S.t215 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2361 S.t214 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2362 S.t213 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2363 S.t212 G D S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2364 D G S.t211 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2365 S.t210 G D S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2366 D G S.t209 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2367 D G S.t208 S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2368 D G S.t207 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2369 D G S.t206 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2370 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2371 S.t204 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2372 S.t203 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2373 S.t202 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2374 D G S.t201 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2375 D G S.t200 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2376 D G S.t199 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2377 S.t198 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2378 S.t197 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2379 S.t196 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2380 S.t195 G D S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2381 D G S.t194 S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2382 D G S.t193 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2383 D G S.t192 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2384 D G S.t191 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2385 D G S.t190 S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2386 S.t189 G D S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2387 D G S.t188 S.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2388 S.t186 G D S.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2389 S.t184 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2390 S.t183 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2391 S.t182 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2392 D G S.t181 S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2393 S.t180 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2394 D G S.t179 S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2395 D G S.t178 S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2396 S.t177 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2397 S.t176 G D S.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2398 S.t174 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2399 D G S.t173 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2400 S.t172 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2401 S.t171 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2402 S.t170 G D S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2403 S.t169 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2404 D G S.t168 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2405 S.t167 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2406 D G S.t165 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2407 D G S.t164 S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2408 S.t163 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2409 S.t162 G D S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2410 S.t161 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2411 S.t160 G D S.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2412 S.t158 G D S.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2413 D G S.t156 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2414 S.t155 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2415 S.t154 G D S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2416 D G S.t153 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2417 D G S.t152 S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2418 S.t151 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2419 D G S.t150 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2420 S.t149 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2421 S.t148 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2422 S.t147 G D S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2423 S.t146 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2424 S.t145 G D S.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2425 D G S.t143 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2426 D G S.t142 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2427 D G S.t141 S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2428 D G S.t140 S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2429 D G S.t139 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2430 D G S.t138 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2431 S.t137 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2432 S.t136 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2433 S.t135 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2434 D G S.t134 S.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2435 D G S.t132 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2436 D G S.t131 S.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2437 D G S.t129 S.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2438 D G S.t127 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2439 S.t126 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2440 D G S.t125 S.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2441 S.t123 G D S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2442 S.t122 G D S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2443 S.t121 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2444 S.t120 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2445 S.t119 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2446 S.t118 G D S.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2447 S.t116 G D S.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2448 D G S.t114 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2449 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2450 D G S.t112 S.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2451 D G S.t110 S.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2452 D G S.t108 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2453 D G S.t107 S.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2454 D G S.t105 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2455 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2456 S.t103 G D S.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2457 D G S.t101 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2458 S.t100 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2459 D G S.t99 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2460 D G S.t98 S.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2461 S.t96 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2462 D G S.t95 S.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2463 D G S.t93 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2464 S.t92 G D S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2465 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2466 S.t90 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2467 D G S.t89 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2468 D G S.t88 S.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2469 D G S.t86 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2470 D G S.t85 S.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2471 S.t83 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2472 S.t82 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2473 D G S.t81 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2474 S.t80 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2475 D G S.t78 S.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2476 S.t76 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2477 S.t75 G D S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2478 S.t74 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2479 D G S.t73 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2480 D G S.t71 S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2481 S.t70 G D S.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2482 D G S.t68 S.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2483 D G S.t66 S.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2484 S.t64 G D S.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2485 S.t62 G D S.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2486 S.t60 G D S.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2487 S.t58 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2488 S.t57 G D S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2489 D G S.t56 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2490 D G S.t54 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2491 D G S.t52 S.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2492 D G S.t50 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2493 D G S.t49 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2494 D G S.t48 S.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2495 D G S.t46 S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2496 D G S.t45 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2497 S.t43 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2498 S.t41 G D S.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2499 S.t39 G D S.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2500 D G S.t37 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2501 D G S.t36 S.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2502 D G S.t34 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2503 S.t32 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2504 S.t30 G D S.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2505 S.t28 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2506 S.t26 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2507 D G S.t24 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2508 S.t22 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2509 S.t20 G D S.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2510 D G S.t18 S.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2511 S.t16 G D S.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2512 S.t14 G D S.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2513 S.t12 G D S.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2514 D G S.t10 S.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2515 S.t8 G D S.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2516 D G S.t6 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2517 S.t5 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2518 S.t3 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2519 D G S.t1 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 S.n972 S.n970 169.035
R1 S.n985 S.n984 169.035
R2 S.n2670 S.n2669 169.035
R3 S.n3512 S.n3511 169.035
R4 S.n4343 S.n4342 169.035
R5 S.n5149 S.n5148 169.035
R6 S.n5946 S.n5945 169.035
R7 S.n6717 S.n6716 169.035
R8 S.n7479 S.n7478 169.035
R9 S.n8215 S.n8214 169.035
R10 S.n8942 S.n8941 169.035
R11 S.n9643 S.n9642 169.035
R12 S.n10335 S.n10334 169.035
R13 S.n10999 S.n10998 169.035
R14 S.n972 S.n971 169.035
R15 S.n10997 S.n10996 138.167
R16 S.n10333 S.n10332 138.167
R17 S.n9641 S.n9640 138.167
R18 S.n8940 S.n8939 138.167
R19 S.n8213 S.n8212 138.167
R20 S.n7477 S.n7476 138.167
R21 S.n6715 S.n6714 138.167
R22 S.n5944 S.n5943 138.167
R23 S.n5147 S.n5146 138.167
R24 S.n4341 S.n4340 138.167
R25 S.n3510 S.n3509 138.167
R26 S.n2668 S.n2667 138.167
R27 S.n983 S.n982 138.167
R28 S.n969 S.n968 138.167
R29 S.n526 S.n525 135.791
R30 S.n1473 S.n1472 135.791
R31 S.n2347 S.n2346 135.791
R32 S.n3129 S.n3128 135.791
R33 S.n4031 S.n4030 135.791
R34 S.n4848 S.n4847 135.791
R35 S.n5647 S.n5646 135.791
R36 S.n6420 S.n6419 135.791
R37 S.n7184 S.n7183 135.791
R38 S.n7755 S.n7754 135.791
R39 S.n8469 S.n8468 135.791
R40 S.n9354 S.n9353 135.791
R41 S.n10048 S.n10047 135.791
R42 S.n11919 S.n11918 91.519
R43 S.n12590 S.n12589 91.519
R44 S.n537 S.n536 91.519
R45 S.n9366 S.n9365 91.519
R46 S.n10059 S.n10058 91.519
R47 S.n10728 S.n10727 91.519
R48 S.n11366 S.n11365 91.519
R49 S.n12288 S.n12287 91.519
R50 S.n7767 S.n7766 91.519
R51 S.n8480 S.n8479 91.519
R52 S.n6432 S.n6431 91.519
R53 S.n7195 S.n7194 91.519
R54 S.n4860 S.n4859 91.519
R55 S.n5658 S.n5657 91.519
R56 S.n3141 S.n3140 91.519
R57 S.n4042 S.n4041 91.519
R58 S.n1485 S.n1484 91.519
R59 S.n2358 S.n2357 91.519
R60 S.n958 S.n957 91.519
R61 S.n1816 S.n1815 91.519
R62 S.n2659 S.n2658 91.519
R63 S.n3500 S.n3499 91.519
R64 S.n4332 S.n4331 91.519
R65 S.n5138 S.n5137 91.519
R66 S.n5935 S.n5934 91.519
R67 S.n6706 S.n6705 91.519
R68 S.n7468 S.n7467 91.519
R69 S.n8204 S.n8203 91.519
R70 S.n8931 S.n8930 91.519
R71 S.n9632 S.n9631 91.519
R72 S.n10324 S.n10323 91.519
R73 S.n10990 S.n10989 91.519
R74 S.n11625 S.n11624 91.519
R75 S.n11993 S.n11992 87.091
R76 S.n211 S.n210 87.091
R77 S.n208 S.n207 87.091
R78 S.n160 S.n159 87.091
R79 S.n235 S.n234 87.091
R80 S.n175 S.n174 87.091
R81 S.n189 S.n188 87.091
R82 S.n199 S.n198 87.091
R83 S.n148 S.n147 87.091
R84 S.n231 S.n230 87.091
R85 S.n136 S.n135 87.091
R86 S.n227 S.n226 87.091
R87 S.n123 S.n122 87.091
R88 S.n223 S.n222 87.091
R89 S.n110 S.n109 87.091
R90 S.n219 S.n218 87.091
R91 S.n97 S.n96 87.091
R92 S.n215 S.n214 87.091
R93 S.n11933 S.n11932 87.091
R94 S.n11937 S.n11936 87.091
R95 S.n11941 S.n11940 87.091
R96 S.n11945 S.n11944 87.091
R97 S.n11949 S.n11948 87.091
R98 S.n11953 S.n11952 87.091
R99 S.n11957 S.n11956 87.091
R100 S.n11961 S.n11960 87.091
R101 S.n11965 S.n11964 87.091
R102 S.n11969 S.n11968 87.091
R103 S.n11973 S.n11972 87.091
R104 S.n11977 S.n11976 87.091
R105 S.n11981 S.n11980 87.091
R106 S.n11985 S.n11984 87.091
R107 S.n11989 S.n11988 87.091
R108 S.n11928 S.n11927 87.091
R109 S.n974 S.t87 50.39
R110 S.n528 S.t185 50.39
R111 S.n987 S.t51 50.39
R112 S.n1475 S.t97 50.39
R113 S.n2672 S.t21 50.39
R114 S.n2349 S.t117 50.39
R115 S.n3514 S.t128 50.39
R116 S.n3131 S.t111 50.39
R117 S.n4345 S.t19 50.39
R118 S.n4033 S.t2 50.39
R119 S.n5151 S.t133 50.39
R120 S.n4850 S.t9 50.39
R121 S.n5948 S.t29 50.39
R122 S.n5649 S.t13 50.39
R123 S.n6719 S.t44 50.39
R124 S.n6422 S.t59 50.39
R125 S.n7481 S.t42 50.39
R126 S.n7186 S.t235 50.39
R127 S.n8217 S.t79 50.39
R128 S.n7757 S.t63 50.39
R129 S.n8944 S.t248 50.39
R130 S.n8471 S.t320 50.39
R131 S.n9645 S.t55 50.39
R132 S.n9356 S.t166 50.39
R133 S.n10337 S.t23 50.39
R134 S.n10050 S.t67 50.39
R135 S.n11001 S.t17 50.39
R136 S.n10718 S.t15 50.39
R137 S.t244 S.n794 48.609
R138 S.t72 S.n1438 48.609
R139 S.t175 S.n1769 48.609
R140 S.t259 S.n2257 48.609
R141 S.t187 S.n2620 48.609
R142 S.t84 S.n3092 48.609
R143 S.t38 S.n3384 48.609
R144 S.t53 S.n3904 48.609
R145 S.t94 S.n4268 48.609
R146 S.t33 S.n4704 48.609
R147 S.t77 S.n5067 48.609
R148 S.t109 S.n5481 48.609
R149 S.t25 S.n5848 48.609
R150 S.t69 S.n6246 48.609
R151 S.t4 S.n6603 48.609
R152 S.t130 S.n6988 48.609
R153 S.t102 S.n7349 48.609
R154 S.t27 S.n7718 48.609
R155 S.t11 S.n7902 48.609
R156 S.t300 S.n8425 48.609
R157 S.t40 S.n8598 48.609
R158 S.t31 S.n9120 48.609
R159 S.t225 S.n9465 48.609
R160 S.t61 S.n9792 48.609
R161 S.t124 S.n10141 48.609
R162 S.t35 S.n10452 48.609
R163 S.t144 S.n10791 48.609
R164 S.t115 S.n11082 48.609
R165 S.n11925 S.t266 3.773
R166 S.n11924 S.t379 3.773
R167 S.n11919 S.t1598 3.773
R168 S.n11645 S.t926 3.773
R169 S.n11877 S.t1225 3.773
R170 S.n11993 S.t1509 3.773
R171 S.n11990 S.t322 3.773
R172 S.n11991 S.t1191 3.773
R173 S.n11905 S.n11904 3.773
R174 S.n11905 S.t1806 3.773
R175 S.n11913 S.t143 3.773
R176 S.n11913 S.n11912 3.773
R177 S.n11916 S.t2438 3.773
R178 S.n11916 S.n11915 3.773
R179 S.n11908 S.n11907 3.773
R180 S.n11908 S.t1596 3.773
R181 S.n12314 S.n12313 3.773
R182 S.n12314 S.t459 3.773
R183 S.n12332 S.t107 3.773
R184 S.n12332 S.n12331 3.773
R185 S.n12329 S.t1646 3.773
R186 S.n12329 S.n12328 3.773
R187 S.n12317 S.n12316 3.773
R188 S.n12317 S.t265 3.773
R189 S.n12590 S.t1825 3.773
R190 S.n12592 S.t1782 3.773
R191 S.n12594 S.t1492 3.773
R192 S.n537 S.t2126 3.773
R193 S.n538 S.t693 3.773
R194 S.n518 S.t421 3.773
R195 S.n937 S.n936 3.773
R196 S.n937 S.t1534 3.773
R197 S.n952 S.t2402 3.773
R198 S.n952 S.n951 3.773
R199 S.n955 S.t93 3.773
R200 S.n955 S.n954 3.773
R201 S.n940 S.n939 3.773
R202 S.n940 S.t2350 3.773
R203 S.n211 S.t1773 3.773
R204 S.n212 S.t956 3.773
R205 S.n209 S.t1829 3.773
R206 S.n208 S.t1266 3.773
R207 S.n204 S.t1585 3.773
R208 S.n205 S.t353 3.773
R209 S.n914 S.n913 3.773
R210 S.n914 S.t2025 3.773
R211 S.n925 S.t375 3.773
R212 S.n925 S.n924 3.773
R213 S.n922 S.t127 3.773
R214 S.n922 S.n921 3.773
R215 S.n917 S.n916 3.773
R216 S.n917 S.t1823 3.773
R217 S.n1419 S.n1418 3.773
R218 S.n1419 S.t2075 3.773
R219 S.n1436 S.t422 3.773
R220 S.n1436 S.n1435 3.773
R221 S.n1433 S.t194 3.773
R222 S.n1433 S.n1432 3.773
R223 S.n1416 S.n1415 3.773
R224 S.n1416 S.t1876 3.773
R225 S.n11885 S.n11884 3.773
R226 S.n11885 S.t1750 3.773
R227 S.n11896 S.t66 3.773
R228 S.n11896 S.n11895 3.773
R229 S.n11893 S.t345 3.773
R230 S.n11893 S.n11892 3.773
R231 S.n11882 S.n11881 3.773
R232 S.n11882 S.t2563 3.773
R233 S.n12297 S.n12296 3.773
R234 S.n12297 S.t1185 3.773
R235 S.n12308 S.t2046 3.773
R236 S.n12308 S.n12307 3.773
R237 S.n12305 S.t2268 3.773
R238 S.n12305 S.n12304 3.773
R239 S.n12294 S.n12293 3.773
R240 S.n12294 S.t1993 3.773
R241 S.n12013 S.n12012 3.773
R242 S.n12013 S.t584 3.773
R243 S.n12028 S.t1453 3.773
R244 S.n12028 S.n12027 3.773
R245 S.n12025 S.t1683 3.773
R246 S.n12025 S.n12024 3.773
R247 S.n12010 S.n12009 3.773
R248 S.n12010 S.t1406 3.773
R249 S.n11395 S.n11394 3.773
R250 S.n11395 S.t120 3.773
R251 S.n11406 S.t869 3.773
R252 S.n11406 S.n11405 3.773
R253 S.n11403 S.t1120 3.773
R254 S.n11403 S.n11402 3.773
R255 S.n11392 S.n11391 3.773
R256 S.n11392 S.t817 3.773
R257 S.n11065 S.n11064 3.773
R258 S.n11065 S.t2080 3.773
R259 S.n11080 S.t426 3.773
R260 S.n11080 S.n11079 3.773
R261 S.n11077 S.t646 3.773
R262 S.n11077 S.n11076 3.773
R263 S.n11062 S.n11061 3.773
R264 S.n11062 S.t377 3.773
R265 S.n10778 S.n10777 3.773
R266 S.n10778 S.t1489 3.773
R267 S.n10789 S.t2353 3.773
R268 S.n10789 S.n10788 3.773
R269 S.n10786 S.t18 3.773
R270 S.n10786 S.n10785 3.773
R271 S.n10775 S.n10774 3.773
R272 S.n10775 S.t2302 3.773
R273 S.n10435 S.n10434 3.773
R274 S.n10435 S.t2253 3.773
R275 S.n10450 S.t1780 3.773
R276 S.n10450 S.n10449 3.773
R277 S.n10447 S.t833 3.773
R278 S.n10447 S.n10446 3.773
R279 S.n10432 S.n10431 3.773
R280 S.n10432 S.t553 3.773
R281 S.n10128 S.n10127 3.773
R282 S.n10128 S.t1667 3.773
R283 S.n10139 S.t2537 3.773
R284 S.n10139 S.n10138 3.773
R285 S.n10136 S.t267 3.773
R286 S.n10136 S.n10135 3.773
R287 S.n10125 S.n10124 3.773
R288 S.n10125 S.t2487 3.773
R289 S.n9775 S.n9774 3.773
R290 S.n9775 S.t880 3.773
R291 S.n9790 S.t1747 3.773
R292 S.n9790 S.n9789 3.773
R293 S.n9787 S.t1991 3.773
R294 S.n9787 S.n9786 3.773
R295 S.n9772 S.n9771 3.773
R296 S.n9772 S.t1918 3.773
R297 S.n9452 S.n9451 3.773
R298 S.n9452 S.t311 3.773
R299 S.n9463 S.t1182 3.773
R300 S.n9463 S.n9462 3.773
R301 S.n9460 S.t1403 3.773
R302 S.n9460 S.n9459 3.773
R303 S.n9449 S.n9448 3.773
R304 S.n9449 S.t1131 3.773
R305 S.n9103 S.n9102 3.773
R306 S.n9103 S.t2241 3.773
R307 S.n9118 S.t582 3.773
R308 S.n9118 S.n9117 3.773
R309 S.n9115 S.t816 3.773
R310 S.n9115 S.n9114 3.773
R311 S.n9100 S.n9099 3.773
R312 S.n9100 S.t538 3.773
R313 S.n8585 S.n8584 3.773
R314 S.n8585 S.t1651 3.773
R315 S.n8596 S.t2520 3.773
R316 S.n8596 S.n8595 3.773
R317 S.n8593 S.t249 3.773
R318 S.n8593 S.n8592 3.773
R319 S.n8582 S.n8581 3.773
R320 S.n8582 S.t2470 3.773
R321 S.n8408 S.n8407 3.773
R322 S.n8408 S.t1085 3.773
R323 S.n8423 S.t1953 3.773
R324 S.n8423 S.n8422 3.773
R325 S.n8420 S.t2182 3.773
R326 S.n8420 S.n8419 3.773
R327 S.n8405 S.n8404 3.773
R328 S.n8405 S.t1899 3.773
R329 S.n7889 S.n7888 3.773
R330 S.n7889 S.t619 3.773
R331 S.n7900 S.t1367 3.773
R332 S.n7900 S.n7899 3.773
R333 S.n7897 S.t1587 3.773
R334 S.n7897 S.n7896 3.773
R335 S.n7886 S.n7885 3.773
R336 S.n7886 S.t1313 3.773
R337 S.n7701 S.n7700 3.773
R338 S.n7701 S.t2553 3.773
R339 S.n7716 S.t906 3.773
R340 S.n7716 S.n7715 3.773
R341 S.n7713 S.t1153 3.773
R342 S.n7713 S.n7712 3.773
R343 S.n7698 S.n7697 3.773
R344 S.n7698 S.t850 3.773
R345 S.n7336 S.n7335 3.773
R346 S.n7336 S.t796 3.773
R347 S.n7347 S.t336 3.773
R348 S.n7347 S.n7346 3.773
R349 S.n7344 S.t1915 3.773
R350 S.n7344 S.n7343 3.773
R351 S.n7333 S.n7332 3.773
R352 S.n7333 S.t1613 3.773
R353 S.n6971 S.n6970 3.773
R354 S.n6971 S.t230 3.773
R355 S.n6986 S.t1103 3.773
R356 S.n6986 S.n6985 3.773
R357 S.n6983 S.t1326 3.773
R358 S.n6983 S.n6982 3.773
R359 S.n6968 S.n6967 3.773
R360 S.n6968 S.t1046 3.773
R361 S.n6590 S.n6589 3.773
R362 S.n6590 S.t2163 3.773
R363 S.n6601 S.t511 3.773
R364 S.n6601 S.n6600 3.773
R365 S.n6598 S.t2186 3.773
R366 S.n6598 S.n6597 3.773
R367 S.n6587 S.n6586 3.773
R368 S.n6587 S.t460 3.773
R369 S.n6229 S.n6228 3.773
R370 S.n6229 S.t777 3.773
R371 S.n6244 S.t1647 3.773
R372 S.n6244 S.n6243 3.773
R373 S.n6241 S.t1892 3.773
R374 S.n6241 S.n6240 3.773
R375 S.n6226 S.n6225 3.773
R376 S.n6226 S.t1318 3.773
R377 S.n5835 S.n5834 3.773
R378 S.n5835 S.t204 3.773
R379 S.n5846 S.t1079 3.773
R380 S.n5846 S.n5845 3.773
R381 S.n5843 S.t1307 3.773
R382 S.n5843 S.n5842 3.773
R383 S.n5832 S.n5831 3.773
R384 S.n5832 S.t1024 3.773
R385 S.n5464 S.n5463 3.773
R386 S.n5464 S.t2147 3.773
R387 S.n5479 S.t493 3.773
R388 S.n5479 S.n5478 3.773
R389 S.n5476 S.t712 3.773
R390 S.n5476 S.n5475 3.773
R391 S.n5461 S.n5460 3.773
R392 S.n5461 S.t440 3.773
R393 S.n5054 S.n5053 3.773
R394 S.n5054 S.t1556 3.773
R395 S.n5065 S.t2423 3.773
R396 S.n5065 S.n5064 3.773
R397 S.n5062 S.t134 3.773
R398 S.n5062 S.n5061 3.773
R399 S.n5051 S.n5050 3.773
R400 S.n5051 S.t2371 3.773
R401 S.n4687 S.n4686 3.773
R402 S.n4687 S.t985 3.773
R403 S.n4702 S.t1856 3.773
R404 S.n4702 S.n4701 3.773
R405 S.n4699 S.t2086 3.773
R406 S.n4699 S.n4698 3.773
R407 S.n4684 S.n4683 3.773
R408 S.n4684 S.t1795 3.773
R409 S.n4255 S.n4254 3.773
R410 S.n4255 S.t528 3.773
R411 S.n4266 S.t1271 3.773
R412 S.n4266 S.n4265 3.773
R413 S.n4263 S.t1495 3.773
R414 S.n4263 S.n4262 3.773
R415 S.n4252 S.n4251 3.773
R416 S.n4252 S.t1228 3.773
R417 S.n3887 S.n3886 3.773
R418 S.n3887 S.t286 3.773
R419 S.n3902 S.t809 3.773
R420 S.n3902 S.n3901 3.773
R421 S.n3899 S.t916 3.773
R422 S.n3899 S.n3898 3.773
R423 S.n3884 S.n3883 3.773
R424 S.n3884 S.t20 3.773
R425 S.n3371 S.n3370 3.773
R426 S.n3371 S.t261 3.773
R427 S.n3382 S.t1130 3.773
R428 S.n3382 S.n3381 3.773
R429 S.n3379 S.t887 3.773
R430 S.n3379 S.n3378 3.773
R431 S.n3368 S.n3367 3.773
R432 S.n3368 S.t2564 3.773
R433 S.n3075 S.n3074 3.773
R434 S.n3075 S.t229 3.773
R435 S.n3090 S.t1104 3.773
R436 S.n3090 S.n3089 3.773
R437 S.n3087 S.t1159 3.773
R438 S.n3087 S.n3086 3.773
R439 S.n3072 S.n3071 3.773
R440 S.n3072 S.t2538 3.773
R441 S.n2607 S.n2606 3.773
R442 S.n2607 S.t485 3.773
R443 S.n2618 S.t1352 3.773
R444 S.n2618 S.n2617 3.773
R445 S.n2615 S.t1138 3.773
R446 S.n2615 S.n2614 3.773
R447 S.n2604 S.n2603 3.773
R448 S.n2604 S.t293 3.773
R449 S.n2240 S.n2239 3.773
R450 S.n2240 S.t2127 3.773
R451 S.n2255 S.t472 3.773
R452 S.n2255 S.n2254 3.773
R453 S.n2252 S.t251 3.773
R454 S.n2252 S.n2251 3.773
R455 S.n2237 S.n2236 3.773
R456 S.n2237 S.t268 3.773
R457 S.n1756 S.n1755 3.773
R458 S.n1756 S.t2100 3.773
R459 S.n1767 S.t447 3.773
R460 S.n1767 S.n1766 3.773
R461 S.n1764 S.t220 3.773
R462 S.n1764 S.n1763 3.773
R463 S.n1753 S.n1752 3.773
R464 S.n1753 S.t1904 3.773
R465 S.n781 S.n780 3.773
R466 S.n781 S.t2053 3.773
R467 S.n792 S.t398 3.773
R468 S.n792 S.n791 3.773
R469 S.n789 S.t165 3.773
R470 S.n789 S.n788 3.773
R471 S.n784 S.n783 3.773
R472 S.n784 S.t1852 3.773
R473 S.n160 S.t746 3.773
R474 S.n153 S.t8 3.773
R475 S.n154 S.t805 3.773
R476 S.n478 S.n477 3.773
R477 S.n478 S.t525 3.773
R478 S.n489 S.t1392 3.773
R479 S.n489 S.n488 3.773
R480 S.n486 S.t1619 3.773
R481 S.n486 S.n485 3.773
R482 S.n481 S.n480 3.773
R483 S.n481 S.t1344 3.773
R484 S.n1274 S.n1273 3.773
R485 S.n1274 S.t1680 3.773
R486 S.n1287 S.t2547 3.773
R487 S.n1287 S.n1286 3.773
R488 S.n1284 S.t280 3.773
R489 S.n1284 S.n1283 3.773
R490 S.n1271 S.n1270 3.773
R491 S.n1271 S.t2498 3.773
R492 S.n9366 S.t2460 3.773
R493 S.n9367 S.t1051 3.773
R494 S.n9347 S.t747 3.773
R495 S.n9127 S.n9126 3.773
R496 S.n9127 S.t1887 3.773
R497 S.n9141 S.t233 3.773
R498 S.n9141 S.n9140 3.773
R499 S.n9144 S.t466 3.773
R500 S.n9144 S.n9143 3.773
R501 S.n9124 S.n9123 3.773
R502 S.n9124 S.t177 3.773
R503 S.n8489 S.n8488 3.773
R504 S.n8489 S.t1302 3.773
R505 S.n8500 S.t2168 3.773
R506 S.n8500 S.n8499 3.773
R507 S.n8497 S.t2396 3.773
R508 S.n8497 S.n8496 3.773
R509 S.n8486 S.n8485 3.773
R510 S.n8486 S.t2118 3.773
R511 S.n8261 S.n8260 3.773
R512 S.n8261 S.t705 3.773
R513 S.n8276 S.t1573 3.773
R514 S.n8276 S.n8275 3.773
R515 S.n8273 S.t1822 3.773
R516 S.n8273 S.n8272 3.773
R517 S.n8258 S.n8257 3.773
R518 S.n8258 S.t1528 3.773
R519 S.n7793 S.n7792 3.773
R520 S.n7793 S.t274 3.773
R521 S.n7804 S.t1009 3.773
R522 S.n7804 S.n7803 3.773
R523 S.n7801 S.t1244 3.773
R524 S.n7801 S.n7800 3.773
R525 S.n7790 S.n7789 3.773
R526 S.n7790 S.t951 3.773
R527 S.n7554 S.n7553 3.773
R528 S.n7554 S.t2203 3.773
R529 S.n7569 S.t551 3.773
R530 S.n7569 S.n7568 3.773
R531 S.n7566 S.t775 3.773
R532 S.n7566 S.n7565 3.773
R533 S.n7551 S.n7550 3.773
R534 S.n7551 S.t500 3.773
R535 S.n7240 S.n7239 3.773
R536 S.n7240 S.t1612 3.773
R537 S.n7251 S.t2484 3.773
R538 S.n7251 S.n7250 3.773
R539 S.n7248 S.t200 3.773
R540 S.n7248 S.n7247 3.773
R541 S.n7237 S.n7236 3.773
R542 S.n7237 S.t2429 3.773
R543 S.n6824 S.n6823 3.773
R544 S.n6824 S.t2378 3.773
R545 S.n6839 S.t1916 3.773
R546 S.n6839 S.n6838 3.773
R547 S.n6836 S.t965 3.773
R548 S.n6836 S.n6835 3.773
R549 S.n6821 S.n6820 3.773
R550 S.n6821 S.t670 3.773
R551 S.n6494 S.n6493 3.773
R552 S.n6494 S.t1800 3.773
R553 S.n6505 S.t138 3.773
R554 S.n6505 S.n6504 3.773
R555 S.n6502 S.t1828 3.773
R556 S.n6502 S.n6501 3.773
R557 S.n6491 S.n6490 3.773
R558 S.n6491 S.t60 3.773
R559 S.n6082 S.n6081 3.773
R560 S.n6082 S.t431 3.773
R561 S.n6097 S.t1297 3.773
R562 S.n6097 S.n6096 3.773
R563 S.n6094 S.t1519 3.773
R564 S.n6094 S.n6093 3.773
R565 S.n6079 S.n6078 3.773
R566 S.n6079 S.t955 3.773
R567 S.n5739 S.n5738 3.773
R568 S.n5739 S.t2357 3.773
R569 S.n5750 S.t699 3.773
R570 S.n5750 S.n5749 3.773
R571 S.n5747 S.t944 3.773
R572 S.n5747 S.n5746 3.773
R573 S.n5736 S.n5735 3.773
R574 S.n5736 S.t650 3.773
R575 S.n5317 S.n5316 3.773
R576 S.n5317 S.t1785 3.773
R577 S.n5332 S.t110 3.773
R578 S.n5332 S.n5331 3.773
R579 S.n5329 S.t373 3.773
R580 S.n5329 S.n5328 3.773
R581 S.n5314 S.n5313 3.773
R582 S.n5314 S.t30 3.773
R583 S.n4958 S.n4957 3.773
R584 S.n4958 S.t1218 3.773
R585 S.n4969 S.t2076 3.773
R586 S.n4969 S.n4968 3.773
R587 S.n4966 S.t2297 3.773
R588 S.n4966 S.n4965 3.773
R589 S.n4955 S.n4954 3.773
R590 S.n4955 S.t2022 3.773
R591 S.n4540 S.n4539 3.773
R592 S.n4540 S.t618 3.773
R593 S.n4555 S.t1486 3.773
R594 S.n4555 S.n4554 3.773
R595 S.n4552 S.t1717 3.773
R596 S.n4552 S.n4551 3.773
R597 S.n4537 S.n4536 3.773
R598 S.n4537 S.t1430 3.773
R599 S.n4159 S.n4158 3.773
R600 S.n4159 S.t161 3.773
R601 S.n4170 S.t908 3.773
R602 S.n4170 S.n4169 3.773
R603 S.n4167 S.t1151 3.773
R604 S.n4167 S.n4166 3.773
R605 S.n4156 S.n4155 3.773
R606 S.n4156 S.t849 3.773
R607 S.n3740 S.n3739 3.773
R608 S.n3740 S.t2110 3.773
R609 S.n3755 S.t454 3.773
R610 S.n3755 S.n3754 3.773
R611 S.n3752 S.t676 3.773
R612 S.n3752 S.n3751 3.773
R613 S.n3737 S.n3736 3.773
R614 S.n3737 S.t406 3.773
R615 S.n3275 S.n3274 3.773
R616 S.n3275 S.t360 3.773
R617 S.n3286 S.t2384 3.773
R618 S.n3286 S.n3285 3.773
R619 S.n3283 S.t1446 3.773
R620 S.n3283 S.n3282 3.773
R621 S.n3272 S.n3271 3.773
R622 S.n3272 S.t1172 3.773
R623 S.n2928 S.n2927 3.773
R624 S.n2928 S.t2283 3.773
R625 S.n2943 S.t629 3.773
R626 S.n2943 S.n2942 3.773
R627 S.n2940 S.t2304 3.773
R628 S.n2940 S.n2939 3.773
R629 S.n2925 S.n2924 3.773
R630 S.n2925 S.t580 3.773
R631 S.n2511 S.n2510 3.773
R632 S.n2511 S.t622 3.773
R633 S.n2522 S.t1491 3.773
R634 S.n2522 S.n2521 3.773
R635 S.n2519 S.t1723 3.773
R636 S.n2519 S.n2518 3.773
R637 S.n2508 S.n2507 3.773
R638 S.n2508 S.t1436 3.773
R639 S.n2091 S.n2090 3.773
R640 S.n2091 S.t342 3.773
R641 S.n2106 S.t1211 3.773
R642 S.n2106 S.n2105 3.773
R643 S.n2103 S.t1428 3.773
R644 S.n2103 S.n2102 3.773
R645 S.n2088 S.n2087 3.773
R646 S.n2088 S.t857 3.773
R647 S.n1655 S.n1654 3.773
R648 S.n1655 S.t2264 3.773
R649 S.n1666 S.t612 3.773
R650 S.n1666 S.n1665 3.773
R651 S.n1663 S.t843 3.773
R652 S.n1663 S.n1662 3.773
R653 S.n1652 S.n1651 3.773
R654 S.n1652 S.t563 3.773
R655 S.n235 S.t1184 3.773
R656 S.n236 S.t1372 3.773
R657 S.n233 S.t2238 3.773
R658 S.n501 S.n500 3.773
R659 S.n501 S.t1397 3.773
R660 S.n512 S.t2299 3.773
R661 S.n512 S.n511 3.773
R662 S.n509 S.t2045 3.773
R663 S.n509 S.n508 3.773
R664 S.n504 S.n503 3.773
R665 S.n504 S.t1212 3.773
R666 S.n10059 S.t2103 3.773
R667 S.n10060 S.t672 3.773
R668 S.n10039 S.t401 3.773
R669 S.n9803 S.n9802 3.773
R670 S.n9803 S.t1312 3.773
R671 S.n9818 S.t2180 3.773
R672 S.n9818 S.n9817 3.773
R673 S.n9821 S.t2406 3.773
R674 S.n9821 S.n9820 3.773
R675 S.n9806 S.n9805 3.773
R676 S.n9806 S.t2329 3.773
R677 S.n9373 S.n9372 3.773
R678 S.n9373 S.t718 3.773
R679 S.n9384 S.t1586 3.773
R680 S.n9384 S.n9383 3.773
R681 S.n9381 S.t1834 3.773
R682 S.n9381 S.n9380 3.773
R683 S.n9376 S.n9375 3.773
R684 S.n9376 S.t1539 3.773
R685 S.n8980 S.n8979 3.773
R686 S.n8980 S.t136 3.773
R687 S.n9000 S.t1020 3.773
R688 S.n9000 S.n8999 3.773
R689 S.n8997 S.t1253 3.773
R690 S.n8997 S.n8996 3.773
R691 S.n8983 S.n8982 3.773
R692 S.n8983 S.t961 3.773
R693 S.n8506 S.n8505 3.773
R694 S.n8506 S.t2212 3.773
R695 S.n8517 S.t436 3.773
R696 S.n8517 S.n8516 3.773
R697 S.n8514 S.t658 3.773
R698 S.n8514 S.n8513 3.773
R699 S.n8509 S.n8508 3.773
R700 S.n8509 S.t387 3.773
R701 S.n8285 S.n8284 3.773
R702 S.n8285 S.t1621 3.773
R703 S.n8305 S.t2492 3.773
R704 S.n8305 S.n8304 3.773
R705 S.n8302 S.t211 3.773
R706 S.n8302 S.n8301 3.773
R707 S.n8288 S.n8287 3.773
R708 S.n8288 S.t2434 3.773
R709 S.n7810 S.n7809 3.773
R710 S.n7810 S.t1052 3.773
R711 S.n7821 S.t1923 3.773
R712 S.n7821 S.n7820 3.773
R713 S.n7818 S.t2152 3.773
R714 S.n7818 S.n7817 3.773
R715 S.n7813 S.n7812 3.773
R716 S.n7813 S.t1865 3.773
R717 S.n7578 S.n7577 3.773
R718 S.n7578 S.t1813 3.773
R719 S.n7598 S.t1337 3.773
R720 S.n7598 S.n7597 3.773
R721 S.n7595 S.t399 3.773
R722 S.n7595 S.n7594 3.773
R723 S.n7581 S.n7580 3.773
R724 S.n7581 S.t80 3.773
R725 S.n7257 S.n7256 3.773
R726 S.n7257 S.t1237 3.773
R727 S.n7268 S.t2102 3.773
R728 S.n7268 S.n7267 3.773
R729 S.n7265 S.t2326 3.773
R730 S.n7265 S.n7264 3.773
R731 S.n7260 S.n7259 3.773
R732 S.n7260 S.t2054 3.773
R733 S.n6848 S.n6847 3.773
R734 S.n6848 S.t643 3.773
R735 S.n6868 S.t1510 3.773
R736 S.n6868 S.n6867 3.773
R737 S.n6865 S.t1746 3.773
R738 S.n6865 S.n6864 3.773
R739 S.n6851 S.n6850 3.773
R740 S.n6851 S.t1457 3.773
R741 S.n6511 S.n6510 3.773
R742 S.n6511 S.t5 3.773
R743 S.n6522 S.t936 3.773
R744 S.n6522 S.n6521 3.773
R745 S.n6519 S.t45 3.773
R746 S.n6519 S.n6518 3.773
R747 S.n6514 S.n6513 3.773
R748 S.n6514 S.t879 3.773
R749 S.n6106 S.n6105 3.773
R750 S.n6106 S.t1226 3.773
R751 S.n6126 S.t2084 3.773
R752 S.n6126 S.n6125 3.773
R753 S.n6123 S.t2307 3.773
R754 S.n6123 S.n6122 3.773
R755 S.n6109 S.n6108 3.773
R756 S.n6109 S.t1738 3.773
R757 S.n5756 S.n5755 3.773
R758 S.n5756 S.t627 3.773
R759 S.n5767 S.t1494 3.773
R760 S.n5767 S.n5766 3.773
R761 S.n5764 S.t1729 3.773
R762 S.n5764 S.n5763 3.773
R763 S.n5759 S.n5758 3.773
R764 S.n5759 S.t1442 3.773
R765 S.n5341 S.n5340 3.773
R766 S.n5341 S.t2567 3.773
R767 S.n5361 S.t918 3.773
R768 S.n5361 S.n5360 3.773
R769 S.n5358 S.t1160 3.773
R770 S.n5358 S.n5357 3.773
R771 S.n5344 S.n5343 3.773
R772 S.n5344 S.t862 3.773
R773 S.n4975 S.n4974 3.773
R774 S.n4975 S.t2119 3.773
R775 S.n4986 S.t347 3.773
R776 S.n4986 S.n4985 3.773
R777 S.n4983 S.t568 3.773
R778 S.n4983 S.n4982 3.773
R779 S.n4978 S.n4977 3.773
R780 S.n4978 S.t291 3.773
R781 S.n4564 S.n4563 3.773
R782 S.n4564 S.t1527 3.773
R783 S.n4584 S.t2394 3.773
R784 S.n4584 S.n4583 3.773
R785 S.n4581 S.t89 3.773
R786 S.n4581 S.n4580 3.773
R787 S.n4567 S.n4566 3.773
R788 S.n4567 S.t2344 3.773
R789 S.n4176 S.n4175 3.773
R790 S.n4176 S.t2293 3.773
R791 S.n4187 S.t1821 3.773
R792 S.n4187 S.n4186 3.773
R793 S.n4184 S.t872 3.773
R794 S.n4184 S.n4183 3.773
R795 S.n4179 S.n4178 3.773
R796 S.n4179 S.t587 3.773
R797 S.n3764 S.n3763 3.773
R798 S.n3764 S.t1710 3.773
R799 S.n3784 S.t2580 3.773
R800 S.n3784 S.n3783 3.773
R801 S.n3781 S.t304 3.773
R802 S.n3781 S.n3780 3.773
R803 S.n3767 S.n3766 3.773
R804 S.n3767 S.t2523 3.773
R805 S.n3292 S.n3291 3.773
R806 S.n3292 S.t1146 3.773
R807 S.n3303 S.t2006 3.773
R808 S.n3303 S.n3302 3.773
R809 S.n3300 S.t2236 3.773
R810 S.n3300 S.n3299 3.773
R811 S.n3295 S.n3294 3.773
R812 S.n3295 S.t1957 3.773
R813 S.n2952 S.n2951 3.773
R814 S.n2952 S.t555 3.773
R815 S.n2972 S.t1419 3.773
R816 S.n2972 S.n2971 3.773
R817 S.n2969 S.t574 3.773
R818 S.n2969 S.n2968 3.773
R819 S.n2955 S.n2954 3.773
R820 S.n2955 S.t1370 3.773
R821 S.n2528 S.n2527 3.773
R822 S.n2528 S.t1412 3.773
R823 S.n2539 S.t2275 3.773
R824 S.n2539 S.n2538 3.773
R825 S.n2536 S.t2511 3.773
R826 S.n2536 S.n2535 3.773
R827 S.n2531 S.n2530 3.773
R828 S.n2531 S.t2226 3.773
R829 S.n2115 S.n2114 3.773
R830 S.n2115 S.t1129 3.773
R831 S.n2135 S.t1990 3.773
R832 S.n2135 S.n2134 3.773
R833 S.n2132 S.t2218 3.773
R834 S.n2132 S.n2131 3.773
R835 S.n2118 S.n2117 3.773
R836 S.n2118 S.t1641 3.773
R837 S.n1672 S.n1671 3.773
R838 S.n1672 S.t537 3.773
R839 S.n1685 S.t1402 3.773
R840 S.n1685 S.n1684 3.773
R841 S.n1682 S.t1626 3.773
R842 S.n1682 S.n1681 3.773
R843 S.n1675 S.n1674 3.773
R844 S.n1675 S.t1351 3.773
R845 S.n1693 S.n1692 3.773
R846 S.n1693 S.t1440 3.773
R847 S.n1707 S.t2191 3.773
R848 S.n1707 S.n1706 3.773
R849 S.n1704 S.t2413 3.773
R850 S.n1704 S.n1703 3.773
R851 S.n1696 S.n1695 3.773
R852 S.n1696 S.t2138 3.773
R853 S.n1325 S.n1324 3.773
R854 S.n1325 S.t2235 3.773
R855 S.n1349 S.t1728 3.773
R856 S.n1349 S.n1348 3.773
R857 S.n1346 S.t366 3.773
R858 S.n1346 S.n1345 3.773
R859 S.n1328 S.n1327 3.773
R860 S.n1328 S.t2039 3.773
R861 S.n516 S.n515 3.773
R862 S.n516 S.t2211 3.773
R863 S.n813 S.t557 3.773
R864 S.n813 S.n812 3.773
R865 S.n816 S.t341 3.773
R866 S.n816 S.n815 3.773
R867 S.n819 S.n818 3.773
R868 S.n819 S.t2014 3.773
R869 S.n827 S.n826 3.773
R870 S.n827 S.t2185 3.773
R871 S.n842 S.t530 3.773
R872 S.n842 S.n841 3.773
R873 S.n839 S.t313 3.773
R874 S.n839 S.n838 3.773
R875 S.n830 S.n829 3.773
R876 S.n830 S.t1989 3.773
R877 S.n175 S.t1967 3.773
R878 S.n167 S.t2160 3.773
R879 S.n168 S.t506 3.773
R880 S.n2153 S.n2152 3.773
R881 S.n2153 S.t1911 3.773
R882 S.n2168 S.t260 3.773
R883 S.n2168 S.n2167 3.773
R884 S.n2165 S.t484 3.773
R885 S.n2165 S.n2164 3.773
R886 S.n2150 S.n2149 3.773
R887 S.n2150 S.t2425 3.773
R888 S.n2989 S.n2988 3.773
R889 S.n2989 S.t1343 3.773
R890 S.n3004 S.t2208 3.773
R891 S.n3004 S.n3003 3.773
R892 S.n3001 S.t1363 3.773
R893 S.n3001 S.n3000 3.773
R894 S.n2986 S.n2985 3.773
R895 S.n2986 S.t2155 3.773
R896 S.n3801 S.n3800 3.773
R897 S.n3801 S.t2497 3.773
R898 S.n3816 S.t842 3.773
R899 S.n3816 S.n3815 3.773
R900 S.n3813 S.t1088 3.773
R901 S.n3813 S.n3812 3.773
R902 S.n3798 S.n3797 3.773
R903 S.n3798 S.t783 3.773
R904 S.n4601 S.n4600 3.773
R905 S.n4601 S.t1156 3.773
R906 S.n4616 S.t2015 3.773
R907 S.n4616 S.n4615 3.773
R908 S.n4613 S.t2242 3.773
R909 S.n4613 S.n4612 3.773
R910 S.n4598 S.n4597 3.773
R911 S.n4598 S.t1969 3.773
R912 S.n5378 S.n5377 3.773
R913 S.n5378 S.t962 3.773
R914 S.n5393 S.t1835 3.773
R915 S.n5393 S.n5392 3.773
R916 S.n5390 S.t2069 3.773
R917 S.n5390 S.n5389 3.773
R918 S.n5375 S.n5374 3.773
R919 S.n5375 S.t1777 3.773
R920 S.n6143 S.n6142 3.773
R921 S.n6143 S.t2004 3.773
R922 S.n6158 S.t356 3.773
R923 S.n6158 S.n6157 3.773
R924 S.n6155 S.t578 3.773
R925 S.n6155 S.n6154 3.773
R926 S.n6140 S.n6139 3.773
R927 S.n6140 S.t2522 3.773
R928 S.n6885 S.n6884 3.773
R929 S.n6885 S.t1431 3.773
R930 S.n6900 S.t2298 3.773
R931 S.n6900 S.n6899 3.773
R932 S.n6897 S.t2528 3.773
R933 S.n6897 S.n6896 3.773
R934 S.n6882 S.n6881 3.773
R935 S.n6882 S.t2246 3.773
R936 S.n7615 S.n7614 3.773
R937 S.n7615 S.t28 3.773
R938 S.n7630 S.t945 3.773
R939 S.n7630 S.n7629 3.773
R940 S.n7627 S.t1190 3.773
R941 S.n7627 S.n7626 3.773
R942 S.n7612 S.n7611 3.773
R943 S.n7612 S.t892 3.773
R944 S.n8322 S.n8321 3.773
R945 S.n8322 S.t1245 3.773
R946 S.n8337 S.t749 3.773
R947 S.n8337 S.n8336 3.773
R948 S.n8334 S.t2337 3.773
R949 S.n8334 S.n8333 3.773
R950 S.n8319 S.n8318 3.773
R951 S.n8319 S.t2063 3.773
R952 S.n9017 S.n9016 3.773
R953 S.n9017 S.t1065 3.773
R954 S.n9032 S.t1934 3.773
R955 S.n9032 S.n9031 3.773
R956 S.n9029 S.t2161 3.773
R957 S.n9029 S.n9028 3.773
R958 S.n9014 S.n9013 3.773
R959 S.n9014 S.t1880 3.773
R960 S.n9689 S.n9688 3.773
R961 S.n9689 S.t2099 3.773
R962 S.n9704 S.t446 3.773
R963 S.n9704 S.n9703 3.773
R964 S.n9701 S.t667 3.773
R965 S.n9701 S.n9700 3.773
R966 S.n9686 S.n9685 3.773
R967 S.n9686 S.t593 3.773
R968 S.n10462 S.n10461 3.773
R969 S.n10462 S.t946 3.773
R970 S.n10476 S.t1815 3.773
R971 S.n10476 S.n10475 3.773
R972 S.n10479 S.t2056 3.773
R973 S.n10479 S.n10478 3.773
R974 S.n10459 S.n10458 3.773
R975 S.n10459 S.t1762 3.773
R976 S.n10728 S.t1522 3.773
R977 S.n10729 S.t81 3.773
R978 S.n10712 S.t2339 3.773
R979 S.n10068 S.n10067 3.773
R980 S.n10068 S.t376 3.773
R981 S.n10079 S.t1241 3.773
R982 S.n10079 S.n10078 3.773
R983 S.n10076 S.t1459 3.773
R984 S.n10076 S.n10075 3.773
R985 S.n10065 S.n10064 3.773
R986 S.n10065 S.t1193 3.773
R987 S.n9392 S.n9391 3.773
R988 S.n9392 S.t1632 3.773
R989 S.n9403 S.t2376 3.773
R990 S.n9403 S.n9402 3.773
R991 S.n9400 S.t56 3.773
R992 S.n9400 S.n9399 3.773
R993 S.n9389 S.n9388 3.773
R994 S.n9389 S.t2324 3.773
R995 S.n8525 S.n8524 3.773
R996 S.n8525 S.t480 3.773
R997 S.n8536 S.t1347 3.773
R998 S.n8536 S.n8535 3.773
R999 S.n8533 S.t1565 3.773
R1000 S.n8533 S.n8532 3.773
R1001 S.n8522 S.n8521 3.773
R1002 S.n8522 S.t1293 3.773
R1003 S.n7829 S.n7828 3.773
R1004 S.n7829 S.t651 3.773
R1005 S.n7840 S.t1518 3.773
R1006 S.n7840 S.n7839 3.773
R1007 S.n7837 S.t1761 3.773
R1008 S.n7837 S.n7836 3.773
R1009 S.n7826 S.n7825 3.773
R1010 S.n7826 S.t1470 3.773
R1011 S.n7276 S.n7275 3.773
R1012 S.n7276 S.t2020 3.773
R1013 S.n7287 S.t372 3.773
R1014 S.n7287 S.n7286 3.773
R1015 S.n7284 S.t590 3.773
R1016 S.n7284 S.n7283 3.773
R1017 S.n7273 S.n7272 3.773
R1018 S.n7273 S.t318 3.773
R1019 S.n6530 S.n6529 3.773
R1020 S.n6530 S.t847 3.773
R1021 S.n6541 S.t1714 3.773
R1022 S.n6541 S.n6540 3.773
R1023 S.n6538 S.t868 3.773
R1024 S.n6538 S.n6537 3.773
R1025 S.n6527 S.n6526 3.773
R1026 S.n6527 S.t1660 3.773
R1027 S.n5775 S.n5774 3.773
R1028 S.n5775 S.t1537 3.773
R1029 S.n5786 S.t2281 3.773
R1030 S.n5786 S.n5785 3.773
R1031 S.n5783 S.t2514 3.773
R1032 S.n5783 S.n5782 3.773
R1033 S.n5772 S.n5771 3.773
R1034 S.n5772 S.t2232 3.773
R1035 S.n4994 S.n4993 3.773
R1036 S.n4994 S.t1721 3.773
R1037 S.n5005 S.t1252 3.773
R1038 S.n5005 S.n5004 3.773
R1039 S.n5002 S.t316 3.773
R1040 S.n5002 S.n5001 3.773
R1041 S.n4991 S.n4990 3.773
R1042 S.n4991 S.t2535 3.773
R1043 S.n4195 S.n4194 3.773
R1044 S.n4195 S.t562 3.773
R1045 S.n4206 S.t1427 3.773
R1046 S.n4206 S.n4205 3.773
R1047 S.n4203 S.t1653 3.773
R1048 S.n4203 S.n4202 3.773
R1049 S.n4192 S.n4191 3.773
R1050 S.n4192 S.t1379 3.773
R1051 S.n3311 S.n3310 3.773
R1052 S.n3311 S.t1928 3.773
R1053 S.n3322 S.t279 3.773
R1054 S.n3322 S.n3321 3.773
R1055 S.n3319 S.t503 3.773
R1056 S.n3319 S.n3318 3.773
R1057 S.n3308 S.n3307 3.773
R1058 S.n3308 S.t214 3.773
R1059 S.n2547 S.n2546 3.773
R1060 S.n2547 S.t2202 3.773
R1061 S.n2558 S.t547 3.773
R1062 S.n2558 S.n2557 3.773
R1063 S.n2555 S.t771 3.773
R1064 S.n2555 S.n2554 3.773
R1065 S.n2544 S.n2543 3.773
R1066 S.n2544 S.t496 3.773
R1067 S.n1364 S.n1363 3.773
R1068 S.n1364 S.t504 3.773
R1069 S.n1383 S.t1369 3.773
R1070 S.n1383 S.n1382 3.773
R1071 S.n1380 S.t1154 3.773
R1072 S.n1380 S.n1379 3.773
R1073 S.n1367 S.n1366 3.773
R1074 S.n1367 S.t308 3.773
R1075 S.n741 S.n740 3.773
R1076 S.n741 S.t477 3.773
R1077 S.n756 S.t1346 3.773
R1078 S.n756 S.n755 3.773
R1079 S.n753 S.t1127 3.773
R1080 S.n753 S.n752 3.773
R1081 S.n744 S.n743 3.773
R1082 S.n744 S.t285 3.773
R1083 S.n859 S.n858 3.773
R1084 S.n859 S.t450 3.773
R1085 S.n875 S.t1317 3.773
R1086 S.n875 S.n874 3.773
R1087 S.n872 S.t1101 3.773
R1088 S.n872 S.n871 3.773
R1089 S.n862 S.n861 3.773
R1090 S.n862 S.t257 3.773
R1091 S.n189 S.t227 3.773
R1092 S.n178 S.t427 3.773
R1093 S.n179 S.t1292 3.773
R1094 S.n11366 S.t957 3.773
R1095 S.n11367 S.t2064 3.773
R1096 S.n11355 S.t1772 3.773
R1097 S.n11096 S.n11095 3.773
R1098 S.n11096 S.t383 3.773
R1099 S.n11104 S.t1249 3.773
R1100 S.n11104 S.n11103 3.773
R1101 S.n11107 S.t1472 3.773
R1102 S.n11107 S.n11106 3.773
R1103 S.n11093 S.n11092 3.773
R1104 S.n11093 S.t1203 3.773
R1105 S.n10742 S.n10741 3.773
R1106 S.n10742 S.t2310 3.773
R1107 S.n10750 S.t652 3.773
R1108 S.n10750 S.n10749 3.773
R1109 S.n10747 S.t893 3.773
R1110 S.n10747 S.n10746 3.773
R1111 S.n10739 S.n10738 3.773
R1112 S.n10739 S.t602 3.773
R1113 S.n10380 S.n10379 3.773
R1114 S.n10380 S.t1732 3.773
R1115 S.n10398 S.t36 3.773
R1116 S.n10398 S.n10397 3.773
R1117 S.n10395 S.t323 3.773
R1118 S.n10395 S.n10394 3.773
R1119 S.n10377 S.n10376 3.773
R1120 S.n10377 S.t2544 3.773
R1121 S.n10092 S.n10091 3.773
R1122 S.n10092 S.t1281 3.773
R1123 S.n10100 S.t2024 3.773
R1124 S.n10100 S.n10099 3.773
R1125 S.n10097 S.t2248 3.773
R1126 S.n10097 S.n10096 3.773
R1127 S.n10089 S.n10088 3.773
R1128 S.n10089 S.t1974 3.773
R1129 S.n9720 S.n9719 3.773
R1130 S.n9720 S.t488 3.773
R1131 S.n9738 S.t1356 3.773
R1132 S.n9738 S.n9737 3.773
R1133 S.n9735 S.t1574 3.773
R1134 S.n9735 S.n9734 3.773
R1135 S.n9717 S.n9716 3.773
R1136 S.n9717 S.t1506 3.773
R1137 S.n9416 S.n9415 3.773
R1138 S.n9416 S.t2416 3.773
R1139 S.n9424 S.t761 3.773
R1140 S.n9424 S.n9423 3.773
R1141 S.n9421 S.t1012 3.773
R1142 S.n9421 S.n9420 3.773
R1143 S.n9413 S.n9412 3.773
R1144 S.n9413 S.t706 3.773
R1145 S.n9048 S.n9047 3.773
R1146 S.n9048 S.t661 3.773
R1147 S.n9066 S.t191 3.773
R1148 S.n9066 S.n9065 3.773
R1149 S.n9063 S.t1771 3.773
R1150 S.n9063 S.n9062 3.773
R1151 S.n9045 S.n9044 3.773
R1152 S.n9045 S.t1482 3.773
R1153 S.n8549 S.n8548 3.773
R1154 S.n8549 S.t41 3.773
R1155 S.n8557 S.t953 3.773
R1156 S.n8557 S.n8556 3.773
R1157 S.n8554 S.t1201 3.773
R1158 S.n8554 S.n8553 3.773
R1159 S.n8546 S.n8545 3.773
R1160 S.n8546 S.t902 3.773
R1161 S.n8353 S.n8352 3.773
R1162 S.n8353 S.t2030 3.773
R1163 S.n8371 S.t380 3.773
R1164 S.n8371 S.n8370 3.773
R1165 S.n8368 S.t601 3.773
R1166 S.n8368 S.n8367 3.773
R1167 S.n8350 S.n8349 3.773
R1168 S.n8350 S.t328 3.773
R1169 S.n7853 S.n7852 3.773
R1170 S.n7853 S.t1439 3.773
R1171 S.n7861 S.t2308 3.773
R1172 S.n7861 S.n7860 3.773
R1173 S.n7858 S.t2542 3.773
R1174 S.n7858 S.n7857 3.773
R1175 S.n7850 S.n7849 3.773
R1176 S.n7850 S.t2257 3.773
R1177 S.n7646 S.n7645 3.773
R1178 S.n7646 S.t861 3.773
R1179 S.n7664 S.t1727 3.773
R1180 S.n7664 S.n7663 3.773
R1181 S.n7661 S.t1971 3.773
R1182 S.n7661 S.n7660 3.773
R1183 S.n7643 S.n7642 3.773
R1184 S.n7643 S.t1672 3.773
R1185 S.n7300 S.n7299 3.773
R1186 S.n7300 S.t294 3.773
R1187 S.n7308 S.t1161 3.773
R1188 S.n7308 S.n7307 3.773
R1189 S.n7305 S.t1384 3.773
R1190 S.n7305 S.n7304 3.773
R1191 S.n7297 S.n7296 3.773
R1192 S.n7297 S.t1109 3.773
R1193 S.n6916 S.n6915 3.773
R1194 S.n6916 S.t2222 3.773
R1195 S.n6934 S.t567 3.773
R1196 S.n6934 S.n6933 3.773
R1197 S.n6931 S.t792 3.773
R1198 S.n6931 S.n6930 3.773
R1199 S.n6913 S.n6912 3.773
R1200 S.n6913 S.t516 3.773
R1201 S.n6554 S.n6553 3.773
R1202 S.n6554 S.t1767 3.773
R1203 S.n6562 S.t2502 3.773
R1204 S.n6562 S.n6561 3.773
R1205 S.n6559 S.t1652 3.773
R1206 S.n6559 S.n6558 3.773
R1207 S.n6551 S.n6550 3.773
R1208 S.n6551 S.t2443 3.773
R1209 S.n6174 S.n6173 3.773
R1210 S.n6174 S.t396 3.773
R1211 S.n6192 S.t1262 3.773
R1212 S.n6192 S.n6191 3.773
R1213 S.n6189 S.t1487 3.773
R1214 S.n6189 S.n6188 3.773
R1215 S.n6171 S.n6170 3.773
R1216 S.n6171 S.t920 3.773
R1217 S.n5799 S.n5798 3.773
R1218 S.n5799 S.t1163 3.773
R1219 S.n5807 S.t668 3.773
R1220 S.n5807 S.n5806 3.773
R1221 S.n5804 S.t2252 3.773
R1222 S.n5804 S.n5803 3.773
R1223 S.n5796 S.n5795 3.773
R1224 S.n5796 S.t1976 3.773
R1225 S.n5409 S.n5408 3.773
R1226 S.n5409 S.t572 3.773
R1227 S.n5427 S.t1434 3.773
R1228 S.n5427 S.n5426 3.773
R1229 S.n5424 S.t1665 3.773
R1230 S.n5424 S.n5423 3.773
R1231 S.n5406 S.n5405 3.773
R1232 S.n5406 S.t1388 3.773
R1233 S.n5018 S.n5017 3.773
R1234 S.n5018 S.t2508 3.773
R1235 S.n5026 S.t856 3.773
R1236 S.n5026 S.n5025 3.773
R1237 S.n5023 S.t1105 3.773
R1238 S.n5023 S.n5022 3.773
R1239 S.n5015 S.n5014 3.773
R1240 S.n5015 S.t799 3.773
R1241 S.n4632 S.n4631 3.773
R1242 S.n4632 S.t1940 3.773
R1243 S.n4650 S.t288 3.773
R1244 S.n4650 S.n4649 3.773
R1245 S.n4647 S.t512 3.773
R1246 S.n4647 S.n4646 3.773
R1247 S.n4629 S.n4628 3.773
R1248 S.n4629 S.t231 3.773
R1249 S.n4219 S.n4218 3.773
R1250 S.n4219 S.t1350 3.773
R1251 S.n4227 S.t2217 3.773
R1252 S.n4227 S.n4226 3.773
R1253 S.n4224 S.t2440 3.773
R1254 S.n4224 S.n4223 3.773
R1255 S.n4216 S.n4215 3.773
R1256 S.n4216 S.t2164 3.773
R1257 S.n3832 S.n3831 3.773
R1258 S.n3832 S.t753 3.773
R1259 S.n3850 S.t1625 3.773
R1260 S.n3850 S.n3849 3.773
R1261 S.n3847 S.t1868 3.773
R1262 S.n3847 S.n3846 3.773
R1263 S.n3829 S.n3828 3.773
R1264 S.n3829 S.t1568 3.773
R1265 S.n3335 S.n3334 3.773
R1266 S.n3335 S.t184 3.773
R1267 S.n3343 S.t1059 3.773
R1268 S.n3343 S.n3342 3.773
R1269 S.n3340 S.t1286 3.773
R1270 S.n3340 S.n3339 3.773
R1271 S.n3332 S.n3331 3.773
R1272 S.n3332 S.t1002 3.773
R1273 S.n3020 S.n3019 3.773
R1274 S.n3020 S.t2130 3.773
R1275 S.n3038 S.t475 3.773
R1276 S.n3038 S.n3037 3.773
R1277 S.n3035 S.t2150 3.773
R1278 S.n3035 S.n3034 3.773
R1279 S.n3017 S.n3016 3.773
R1280 S.n3017 S.t424 3.773
R1281 S.n2571 S.n2570 3.773
R1282 S.n2571 S.t585 3.773
R1283 S.n2579 S.t1335 3.773
R1284 S.n2579 S.n2578 3.773
R1285 S.n2576 S.t1558 3.773
R1286 S.n2576 S.n2575 3.773
R1287 S.n2568 S.n2567 3.773
R1288 S.n2568 S.t1284 3.773
R1289 S.n2184 S.n2183 3.773
R1290 S.n2184 S.t552 3.773
R1291 S.n2202 S.t1168 3.773
R1292 S.n2202 S.n2201 3.773
R1293 S.n2199 S.t1207 3.773
R1294 S.n2199 S.n2198 3.773
R1295 S.n2181 S.n2180 3.773
R1296 S.n2181 S.t1220 3.773
R1297 S.n1720 S.n1719 3.773
R1298 S.n1720 S.t526 3.773
R1299 S.n1728 S.t1393 3.773
R1300 S.n1728 S.n1727 3.773
R1301 S.n1725 S.t1177 3.773
R1302 S.n1725 S.n1724 3.773
R1303 S.n1717 S.n1716 3.773
R1304 S.n1717 S.t335 3.773
R1305 S.n1392 S.n1391 3.773
R1306 S.n1392 S.t1287 3.773
R1307 S.n1411 S.t2156 3.773
R1308 S.n1411 S.n1410 3.773
R1309 S.n1408 S.t1935 3.773
R1310 S.n1408 S.n1407 3.773
R1311 S.n1395 S.n1394 3.773
R1312 S.n1395 S.t1092 3.773
R1313 S.n761 S.n760 3.773
R1314 S.n761 S.t1264 3.773
R1315 S.n775 S.t2132 3.773
R1316 S.n775 S.n774 3.773
R1317 S.n772 S.t1910 3.773
R1318 S.n772 S.n771 3.773
R1319 S.n764 S.n763 3.773
R1320 S.n764 S.t1066 3.773
R1321 S.n1739 S.n1738 3.773
R1322 S.n1739 S.t1314 3.773
R1323 S.n1748 S.t2183 3.773
R1324 S.n1748 S.n1747 3.773
R1325 S.n1745 S.t1960 3.773
R1326 S.n1745 S.n1744 3.773
R1327 S.n1736 S.n1735 3.773
R1328 S.n1736 S.t1121 3.773
R1329 S.n2211 S.n2210 3.773
R1330 S.n2211 S.t1341 3.773
R1331 S.n2223 S.t2206 3.773
R1332 S.n2223 S.n2222 3.773
R1333 S.n2220 S.t1985 3.773
R1334 S.n2220 S.n2219 3.773
R1335 S.n2214 S.n2213 3.773
R1336 S.n2214 S.t1997 3.773
R1337 S.n2585 S.n2584 3.773
R1338 S.n2585 S.t2219 3.773
R1339 S.n2599 S.t564 3.773
R1340 S.n2599 S.n2598 3.773
R1341 S.n2596 S.t350 3.773
R1342 S.n2596 S.n2595 3.773
R1343 S.n2588 S.n2587 3.773
R1344 S.n2588 S.t2019 3.773
R1345 S.n3047 S.n3046 3.773
R1346 S.n3047 S.t1968 3.773
R1347 S.n3058 S.t1382 3.773
R1348 S.n3058 S.n3057 3.773
R1349 S.n3055 S.t371 3.773
R1350 S.n3055 S.n3054 3.773
R1351 S.n3050 S.n3049 3.773
R1352 S.n3050 S.t1757 3.773
R1353 S.n3349 S.n3348 3.773
R1354 S.n3349 S.t1108 3.773
R1355 S.n3363 S.t1844 3.773
R1356 S.n3363 S.n3362 3.773
R1357 S.n3360 S.t2077 3.773
R1358 S.n3360 S.n3359 3.773
R1359 S.n3352 S.n3351 3.773
R1360 S.n3352 S.t1786 3.773
R1361 S.n3859 S.n3858 3.773
R1362 S.n3859 S.t1546 3.773
R1363 S.n3870 S.t2412 3.773
R1364 S.n3870 S.n3869 3.773
R1365 S.n3867 S.t112 3.773
R1366 S.n3867 S.n3866 3.773
R1367 S.n3862 S.n3861 3.773
R1368 S.n3862 S.t2358 3.773
R1369 S.n4233 S.n4232 3.773
R1370 S.n4233 S.t2137 3.773
R1371 S.n4247 S.t483 3.773
R1372 S.n4247 S.n4246 3.773
R1373 S.n4244 S.t700 3.773
R1374 S.n4244 S.n4243 3.773
R1375 S.n4236 S.n4235 3.773
R1376 S.n4236 S.t433 3.773
R1377 S.n4659 S.n4658 3.773
R1378 S.n4659 S.t198 3.773
R1379 S.n4670 S.t1071 3.773
R1380 S.n4670 S.n4669 3.773
R1381 S.n4667 S.t1298 3.773
R1382 S.n4667 S.n4666 3.773
R1383 S.n4662 S.n4661 3.773
R1384 S.n4662 S.t1017 3.773
R1385 S.n5032 S.n5031 3.773
R1386 S.n5032 S.t768 3.773
R1387 S.n5046 S.t1639 3.773
R1388 S.n5046 S.n5045 3.773
R1389 S.n5043 S.t1885 3.773
R1390 S.n5043 S.n5042 3.773
R1391 S.n5035 S.n5034 3.773
R1392 S.n5035 S.t1580 3.773
R1393 S.n5436 S.n5435 3.773
R1394 S.n5436 S.t1361 3.773
R1395 S.n5447 S.t2225 3.773
R1396 S.n5447 S.n5446 3.773
R1397 S.n5444 S.t2455 3.773
R1398 S.n5444 S.n5443 3.773
R1399 S.n5439 S.n5438 3.773
R1400 S.n5439 S.t2175 3.773
R1401 S.n5813 S.n5812 3.773
R1402 S.n5813 S.t1947 3.773
R1403 S.n5827 S.t297 3.773
R1404 S.n5827 S.n5826 3.773
R1405 S.n5824 S.t520 3.773
R1406 S.n5824 S.n5823 3.773
R1407 S.n5816 S.n5815 3.773
R1408 S.n5816 S.t239 3.773
R1409 S.n6201 S.n6200 3.773
R1410 S.n6201 S.t2518 3.773
R1411 S.n6212 S.t864 3.773
R1412 S.n6212 S.n6211 3.773
R1413 S.n6209 S.t1112 3.773
R1414 S.n6209 S.n6208 3.773
R1415 S.n6204 S.n6203 3.773
R1416 S.n6204 S.t532 3.773
R1417 S.n6568 S.n6567 3.773
R1418 S.n6568 S.t1378 3.773
R1419 S.n6582 S.t897 3.773
R1420 S.n6582 S.n6581 3.773
R1421 S.n6579 S.t1398 3.773
R1422 S.n6579 S.n6578 3.773
R1423 S.n6571 S.n6570 3.773
R1424 S.n6571 S.t2194 3.773
R1425 S.n6943 S.n6942 3.773
R1426 S.n6943 S.t607 3.773
R1427 S.n6954 S.t1476 3.773
R1428 S.n6954 S.n6953 3.773
R1429 S.n6951 S.t1706 3.773
R1430 S.n6951 S.n6950 3.773
R1431 S.n6946 S.n6945 3.773
R1432 S.n6946 S.t1424 3.773
R1433 S.n7314 S.n7313 3.773
R1434 S.n7314 S.t1206 3.773
R1435 S.n7328 S.t1945 3.773
R1436 S.n7328 S.n7327 3.773
R1437 S.n7325 S.t2169 3.773
R1438 S.n7325 S.n7324 3.773
R1439 S.n7317 S.n7316 3.773
R1440 S.n7317 S.t1888 3.773
R1441 S.n7673 S.n7672 3.773
R1442 S.n7673 S.t1645 3.773
R1443 S.n7684 S.t2516 3.773
R1444 S.n7684 S.n7683 3.773
R1445 S.n7681 S.t236 3.773
R1446 S.n7681 S.n7680 3.773
R1447 S.n7676 S.n7675 3.773
R1448 S.n7676 S.t2461 3.773
R1449 S.n7867 S.n7866 3.773
R1450 S.n7867 S.t2231 3.773
R1451 S.n7881 S.t576 3.773
R1452 S.n7881 S.n7880 3.773
R1453 S.n7878 S.t806 3.773
R1454 S.n7878 S.n7877 3.773
R1455 S.n7870 S.n7869 3.773
R1456 S.n7870 S.t527 3.773
R1457 S.n8380 S.n8379 3.773
R1458 S.n8380 S.t301 3.773
R1459 S.n8391 S.t1166 3.773
R1460 S.n8391 S.n8390 3.773
R1461 S.n8388 S.t1394 3.773
R1462 S.n8388 S.n8387 3.773
R1463 S.n8383 S.n8382 3.773
R1464 S.n8383 S.t1118 3.773
R1465 S.n8563 S.n8562 3.773
R1466 S.n8563 S.t867 3.773
R1467 S.n8577 S.t1736 3.773
R1468 S.n8577 S.n8576 3.773
R1469 S.n8574 S.t1981 3.773
R1470 S.n8574 S.n8573 3.773
R1471 S.n8566 S.n8565 3.773
R1472 S.n8566 S.t1681 3.773
R1473 S.n9075 S.n9074 3.773
R1474 S.n9075 S.t1451 3.773
R1475 S.n9086 S.t2316 3.773
R1476 S.n9086 S.n9085 3.773
R1477 S.n9083 S.t2548 3.773
R1478 S.n9083 S.n9082 3.773
R1479 S.n9078 S.n9077 3.773
R1480 S.n9078 S.t2265 3.773
R1481 S.n9430 S.n9429 3.773
R1482 S.n9430 S.t2043 3.773
R1483 S.n9444 S.t390 3.773
R1484 S.n9444 S.n9443 3.773
R1485 S.n9441 S.t613 3.773
R1486 S.n9441 S.n9440 3.773
R1487 S.n9433 S.n9432 3.773
R1488 S.n9433 S.t343 3.773
R1489 S.n9747 S.n9746 3.773
R1490 S.n9747 S.t62 3.773
R1491 S.n9758 S.t2141 3.773
R1492 S.n9758 S.n9757 3.773
R1493 S.n9755 S.t1213 3.773
R1494 S.n9755 S.n9754 3.773
R1495 S.n9750 S.n9749 3.773
R1496 S.n9750 S.t1136 3.773
R1497 S.n10106 S.n10105 3.773
R1498 S.n10106 S.t2071 3.773
R1499 S.n10120 S.t418 3.773
R1500 S.n10120 S.n10119 3.773
R1501 S.n10117 S.t640 3.773
R1502 S.n10117 S.n10116 3.773
R1503 S.n10109 S.n10108 3.773
R1504 S.n10109 S.t368 3.773
R1505 S.n10407 S.n10406 3.773
R1506 S.n10407 S.t100 3.773
R1507 S.n10418 S.t997 3.773
R1508 S.n10418 S.n10417 3.773
R1509 S.n10415 S.t1234 3.773
R1510 S.n10415 S.n10414 3.773
R1511 S.n10410 S.n10409 3.773
R1512 S.n10410 S.t940 3.773
R1513 S.n10756 S.n10755 3.773
R1514 S.n10756 S.t696 3.773
R1515 S.n10770 S.t1445 3.773
R1516 S.n10770 S.n10769 3.773
R1517 S.n10767 S.t1676 3.773
R1518 S.n10767 S.n10766 3.773
R1519 S.n10759 S.n10758 3.773
R1520 S.n10759 S.t1396 3.773
R1521 S.n11037 S.n11036 3.773
R1522 S.n11037 S.t1169 3.773
R1523 S.n11048 S.t2032 3.773
R1524 S.n11048 S.n11047 3.773
R1525 S.n11045 S.t2259 3.773
R1526 S.n11045 S.n11044 3.773
R1527 S.n11040 S.n11039 3.773
R1528 S.n11040 S.t1983 3.773
R1529 S.n11373 S.n11372 3.773
R1530 S.n11373 S.t1739 3.773
R1531 S.n11387 S.t48 3.773
R1532 S.n11387 S.n11386 3.773
R1533 S.n11384 S.t330 3.773
R1534 S.n11384 S.n11383 3.773
R1535 S.n11376 S.n11375 3.773
R1536 S.n11376 S.t2551 3.773
R1537 S.n12041 S.n12040 3.773
R1538 S.n12041 S.t2321 3.773
R1539 S.n12049 S.t663 3.773
R1540 S.n12049 S.n12048 3.773
R1541 S.n12052 S.t904 3.773
R1542 S.n12052 S.n12051 3.773
R1543 S.n12044 S.n12043 3.773
R1544 S.n12044 S.t615 3.773
R1545 S.n12288 S.t392 3.773
R1546 S.n12289 S.t1484 3.773
R1547 S.n12279 S.t1215 3.773
R1548 S.n199 S.t1015 3.773
R1549 S.n191 S.t1223 3.773
R1550 S.n192 S.t2081 3.773
R1551 S.n885 S.n884 3.773
R1552 S.n885 S.t1240 3.773
R1553 S.n904 S.t2105 3.773
R1554 S.n904 S.n903 3.773
R1555 S.n901 S.t1883 3.773
R1556 S.n901 S.n900 3.773
R1557 S.n888 S.n887 3.773
R1558 S.n888 S.t1044 3.773
R1559 S.n1296 S.n1295 3.773
R1560 S.n1296 S.t2466 3.773
R1561 S.n1315 S.t813 3.773
R1562 S.n1315 S.n1314 3.773
R1563 S.n1312 S.t1060 3.773
R1564 S.n1312 S.n1311 3.773
R1565 S.n1299 S.n1298 3.773
R1566 S.n1299 S.t754 3.773
R1567 S.n725 S.n724 3.773
R1568 S.n725 S.t2021 3.773
R1569 S.n736 S.t245 3.773
R1570 S.n736 S.n735 3.773
R1571 S.n733 S.t476 3.773
R1572 S.n733 S.n732 3.773
R1573 S.n728 S.n727 3.773
R1574 S.n728 S.t186 3.773
R1575 S.n708 S.n707 3.773
R1576 S.n708 S.t1116 3.773
R1577 S.n719 S.t1980 3.773
R1578 S.n719 S.n718 3.773
R1579 S.n716 S.t2209 3.773
R1580 S.n716 S.n715 3.773
R1581 S.n711 S.n710 3.773
R1582 S.n711 S.t1929 3.773
R1583 S.n148 S.t1702 3.773
R1584 S.n141 S.t891 3.773
R1585 S.n142 S.t1760 3.773
R1586 S.n434 S.n433 3.773
R1587 S.n434 S.t1468 3.773
R1588 S.n445 S.t2335 3.773
R1589 S.n445 S.n444 3.773
R1590 S.n442 S.t2571 3.773
R1591 S.n442 S.n441 3.773
R1592 S.n437 S.n436 3.773
R1593 S.n437 S.t2284 3.773
R1594 S.n1215 S.n1214 3.773
R1595 S.n1215 S.t90 3.773
R1596 S.n1228 S.t987 3.773
R1597 S.n1228 S.n1227 3.773
R1598 S.n1225 S.t1230 3.773
R1599 S.n1225 S.n1224 3.773
R1600 S.n1212 S.n1211 3.773
R1601 S.n1212 S.t933 3.773
R1602 S.n7767 S.t1097 3.773
R1603 S.n7768 S.t2190 3.773
R1604 S.n7748 S.t1908 3.773
R1605 S.n7725 S.n7724 3.773
R1606 S.n7725 S.t508 3.773
R1607 S.n7739 S.t1374 3.773
R1608 S.n7739 S.n7738 3.773
R1609 S.n7742 S.t1592 3.773
R1610 S.n7742 S.n7741 3.773
R1611 S.n7722 S.n7721 3.773
R1612 S.n7722 S.t1322 3.773
R1613 S.n7204 S.n7203 3.773
R1614 S.n7204 S.t2432 3.773
R1615 S.n7215 S.t779 3.773
R1616 S.n7215 S.n7214 3.773
R1617 S.n7212 S.t1027 3.773
R1618 S.n7212 S.n7211 3.773
R1619 S.n7201 S.n7200 3.773
R1620 S.n7201 S.t722 3.773
R1621 S.n6763 S.n6762 3.773
R1622 S.n6763 S.t1864 3.773
R1623 S.n6778 S.t207 3.773
R1624 S.n6778 S.n6777 3.773
R1625 S.n6775 S.t445 3.773
R1626 S.n6775 S.n6774 3.773
R1627 S.n6760 S.n6759 3.773
R1628 S.n6760 S.t148 3.773
R1629 S.n6458 S.n6457 3.773
R1630 S.n6458 S.t1404 3.773
R1631 S.n6469 S.t2151 3.773
R1632 S.n6469 S.n6468 3.773
R1633 S.n6466 S.t1303 3.773
R1634 S.n6466 S.n6465 3.773
R1635 S.n6455 S.n6454 3.773
R1636 S.n6455 S.t2098 3.773
R1637 S.n6021 S.n6020 3.773
R1638 S.n6021 S.t2545 3.773
R1639 S.n6036 S.t898 3.773
R1640 S.n6036 S.n6035 3.773
R1641 S.n6033 S.t1142 3.773
R1642 S.n6033 S.n6032 3.773
R1643 S.n6018 S.n6017 3.773
R1644 S.n6018 S.t560 3.773
R1645 S.n5703 S.n5702 3.773
R1646 S.n5703 S.t1975 3.773
R1647 S.n5714 S.t324 3.773
R1648 S.n5714 S.n5713 3.773
R1649 S.n5711 S.t550 3.773
R1650 S.n5711 S.n5710 3.773
R1651 S.n5700 S.n5699 3.773
R1652 S.n5700 S.t273 3.773
R1653 S.n5256 S.n5255 3.773
R1654 S.n5256 S.t213 3.773
R1655 S.n5271 S.t2251 3.773
R1656 S.n5271 S.n5270 3.773
R1657 S.n5268 S.t1315 3.773
R1658 S.n5268 S.n5267 3.773
R1659 S.n5253 S.n5252 3.773
R1660 S.n5253 S.t1033 3.773
R1661 S.n4922 S.n4921 3.773
R1662 S.n4922 S.t2154 3.773
R1663 S.n4933 S.t502 3.773
R1664 S.n4933 S.n4932 3.773
R1665 S.n4930 S.t719 3.773
R1666 S.n4930 S.n4929 3.773
R1667 S.n4919 S.n4918 3.773
R1668 S.n4919 S.t448 3.773
R1669 S.n4479 S.n4478 3.773
R1670 S.n4479 S.t1560 3.773
R1671 S.n4494 S.t2430 3.773
R1672 S.n4494 S.n4493 3.773
R1673 S.n4491 S.t139 3.773
R1674 S.n4491 S.n4490 3.773
R1675 S.n4476 S.n4475 3.773
R1676 S.n4476 S.t2379 3.773
R1677 S.n4123 S.n4122 3.773
R1678 S.n4123 S.t992 3.773
R1679 S.n4134 S.t1859 3.773
R1680 S.n4134 S.n4133 3.773
R1681 S.n4131 S.t2092 3.773
R1682 S.n4131 S.n4130 3.773
R1683 S.n4120 S.n4119 3.773
R1684 S.n4120 S.t1801 3.773
R1685 S.n3679 S.n3678 3.773
R1686 S.n3679 S.t413 3.773
R1687 S.n3694 S.t1276 3.773
R1688 S.n3694 S.n3693 3.773
R1689 S.n3691 S.t1501 3.773
R1690 S.n3691 S.n3690 3.773
R1691 S.n3676 S.n3675 3.773
R1692 S.n3676 S.t1231 3.773
R1693 S.n3239 S.n3238 3.773
R1694 S.n3239 S.t2342 3.773
R1695 S.n3250 S.t685 3.773
R1696 S.n3250 S.n3249 3.773
R1697 S.n3247 S.t927 3.773
R1698 S.n3247 S.n3246 3.773
R1699 S.n3236 S.n3235 3.773
R1700 S.n3236 S.t635 3.773
R1701 S.n2867 S.n2866 3.773
R1702 S.n2867 S.t1764 3.773
R1703 S.n2882 S.t85 3.773
R1704 S.n2882 S.n2881 3.773
R1705 S.n2879 S.t1787 3.773
R1706 S.n2879 S.n2878 3.773
R1707 S.n2864 S.n2863 3.773
R1708 S.n2864 S.t2574 3.773
R1709 S.n2475 S.n2474 3.773
R1710 S.n2475 S.t237 3.773
R1711 S.n2486 S.t975 3.773
R1712 S.n2486 S.n2485 3.773
R1713 S.n2483 S.t1219 3.773
R1714 S.n2483 S.n2482 3.773
R1715 S.n2472 S.n2471 3.773
R1716 S.n2472 S.t919 3.773
R1717 S.n2030 S.n2029 3.773
R1718 S.n2030 S.t2444 3.773
R1719 S.n2045 S.t788 3.773
R1720 S.n2045 S.n2044 3.773
R1721 S.n2042 S.t1042 3.773
R1722 S.n2042 S.n2041 3.773
R1723 S.n2027 S.n2026 3.773
R1724 S.n2027 S.t468 3.773
R1725 S.n1619 S.n1618 3.773
R1726 S.n1619 S.t692 3.773
R1727 S.n1630 S.t223 3.773
R1728 S.n1630 S.n1629 3.773
R1729 S.n1627 S.t1797 3.773
R1730 S.n1627 S.n1626 3.773
R1731 S.n1616 S.n1615 3.773
R1732 S.n1616 S.t1508 3.773
R1733 S.n231 S.t2491 3.773
R1734 S.n232 S.t1671 3.773
R1735 S.n229 S.t2541 3.773
R1736 S.n457 S.n456 3.773
R1737 S.n457 S.t2256 3.773
R1738 S.n460 S.t600 3.773
R1739 S.n460 S.n459 3.773
R1740 S.n468 S.t837 3.773
R1741 S.n468 S.n467 3.773
R1742 S.n463 S.n462 3.773
R1743 S.n463 S.t556 3.773
R1744 S.n8480 S.t515 3.773
R1745 S.n8481 S.t1607 3.773
R1746 S.n8460 S.t1333 3.773
R1747 S.n8436 S.n8435 3.773
R1748 S.n8436 S.t2442 3.773
R1749 S.n8451 S.t787 3.773
R1750 S.n8451 S.n8450 3.773
R1751 S.n8454 S.t1041 3.773
R1752 S.n8454 S.n8453 3.773
R1753 S.n8439 S.n8438 3.773
R1754 S.n8439 S.t735 3.773
R1755 S.n7774 S.n7773 3.773
R1756 S.n7774 S.t1878 3.773
R1757 S.n7785 S.t222 3.773
R1758 S.n7785 S.n7784 3.773
R1759 S.n7782 S.t456 3.773
R1760 S.n7782 S.n7781 3.773
R1761 S.n7777 S.n7776 3.773
R1762 S.n7777 S.t163 3.773
R1763 S.n7517 S.n7516 3.773
R1764 S.n7517 S.t1290 3.773
R1765 S.n7537 S.t2158 3.773
R1766 S.n7537 S.n7536 3.773
R1767 S.n7534 S.t2382 3.773
R1768 S.n7534 S.n7533 3.773
R1769 S.n7520 S.n7519 3.773
R1770 S.n7520 S.t2108 3.773
R1771 S.n7221 S.n7220 3.773
R1772 S.n7221 S.t830 3.773
R1773 S.n7232 S.t1563 3.773
R1774 S.n7232 S.n7231 3.773
R1775 S.n7229 S.t1808 3.773
R1776 S.n7229 S.n7228 3.773
R1777 S.n7224 S.n7223 3.773
R1778 S.n7224 S.t1515 3.773
R1779 S.n6787 S.n6786 3.773
R1780 S.n6787 S.t263 3.773
R1781 S.n6807 S.t1132 3.773
R1782 S.n6807 S.n6806 3.773
R1783 S.n6804 S.t1354 3.773
R1784 S.n6804 S.n6803 3.773
R1785 S.n6790 S.n6789 3.773
R1786 S.n6790 S.t1074 3.773
R1787 S.n6475 S.n6474 3.773
R1788 S.n6475 S.t2195 3.773
R1789 S.n6486 S.t540 3.773
R1790 S.n6486 S.n6485 3.773
R1791 S.n6483 S.t2215 3.773
R1792 S.n6483 S.n6482 3.773
R1793 S.n6478 S.n6477 3.773
R1794 S.n6478 S.t487 3.773
R1795 S.n6045 S.n6044 3.773
R1796 S.n6045 S.t2165 3.773
R1797 S.n6065 S.t1677 3.773
R1798 S.n6065 S.n6064 3.773
R1799 S.n6062 S.t728 3.773
R1800 S.n6062 S.n6061 3.773
R1801 S.n6048 S.n6047 3.773
R1802 S.n6048 S.t169 3.773
R1803 S.n5720 S.n5719 3.773
R1804 S.n5720 S.t1567 3.773
R1805 S.n5731 S.t2439 3.773
R1806 S.n5731 S.n5730 3.773
R1807 S.n5728 S.t152 3.773
R1808 S.n5728 S.n5727 3.773
R1809 S.n5723 S.n5722 3.773
R1810 S.n5723 S.t2387 3.773
R1811 S.n5280 S.n5279 3.773
R1812 S.n5280 S.t1001 3.773
R1813 S.n5300 S.t1867 3.773
R1814 S.n5300 S.n5299 3.773
R1815 S.n5297 S.t2101 3.773
R1816 S.n5297 S.n5296 3.773
R1817 S.n5283 S.n5282 3.773
R1818 S.n5283 S.t1812 3.773
R1819 S.n4939 S.n4938 3.773
R1820 S.n4939 S.t423 3.773
R1821 S.n4950 S.t1288 3.773
R1822 S.n4950 S.n4949 3.773
R1823 S.n4947 S.t1511 3.773
R1824 S.n4947 S.n4946 3.773
R1825 S.n4942 S.n4941 3.773
R1826 S.n4942 S.t1238 3.773
R1827 S.n4503 S.n4502 3.773
R1828 S.n4503 S.t2351 3.773
R1829 S.n4523 S.t694 3.773
R1830 S.n4523 S.n4522 3.773
R1831 S.n4520 S.t935 3.773
R1832 S.n4520 S.n4519 3.773
R1833 S.n4506 S.n4505 3.773
R1834 S.n4506 S.t644 3.773
R1835 S.n4140 S.n4139 3.773
R1836 S.n4140 S.t1774 3.773
R1837 S.n4151 S.t95 3.773
R1838 S.n4151 S.n4150 3.773
R1839 S.n4148 S.t364 3.773
R1840 S.n4148 S.n4147 3.773
R1841 S.n4143 S.n4142 3.773
R1842 S.n4143 S.t3 3.773
R1843 S.n3703 S.n3702 3.773
R1844 S.n3703 S.t1205 3.773
R1845 S.n3723 S.t2066 3.773
R1846 S.n3723 S.n3722 3.773
R1847 S.n3720 S.t2288 3.773
R1848 S.n3720 S.n3719 3.773
R1849 S.n3706 S.n3705 3.773
R1850 S.n3706 S.t2012 3.773
R1851 S.n3256 S.n3255 3.773
R1852 S.n3256 S.t723 3.773
R1853 S.n3267 S.t1473 3.773
R1854 S.n3267 S.n3266 3.773
R1855 S.n3264 S.t1704 3.773
R1856 S.n3264 S.n3263 3.773
R1857 S.n3259 S.n3258 3.773
R1858 S.n3259 S.t1422 3.773
R1859 S.n2891 S.n2890 3.773
R1860 S.n2891 S.t147 3.773
R1861 S.n2911 S.t1028 3.773
R1862 S.n2911 S.n2910 3.773
R1863 S.n2908 S.t178 3.773
R1864 S.n2908 S.n2907 3.773
R1865 S.n2894 S.n2893 3.773
R1866 S.n2894 S.t972 3.773
R1867 S.n2492 S.n2491 3.773
R1868 S.n2492 S.t2355 3.773
R1869 S.n2503 S.t1889 3.773
R1870 S.n2503 S.n2502 3.773
R1871 S.n2500 S.t941 3.773
R1872 S.n2500 S.n2499 3.773
R1873 S.n2495 S.n2494 3.773
R1874 S.n2495 S.t648 3.773
R1875 S.n2054 S.n2053 3.773
R1876 S.n2054 S.t2072 3.773
R1877 S.n2074 S.t419 3.773
R1878 S.n2074 S.n2073 3.773
R1879 S.n2071 S.t641 3.773
R1880 S.n2071 S.n2070 3.773
R1881 S.n2057 S.n2056 3.773
R1882 S.n2057 S.t22 3.773
R1883 S.n1636 S.n1635 3.773
R1884 S.n1636 S.t1481 3.773
R1885 S.n1647 S.t2348 3.773
R1886 S.n1647 S.n1646 3.773
R1887 S.n1644 S.t2581 3.773
R1888 S.n1644 S.n1643 3.773
R1889 S.n1639 S.n1638 3.773
R1890 S.n1639 S.t2294 3.773
R1891 S.n1237 S.n1236 3.773
R1892 S.n1237 S.t900 3.773
R1893 S.n1257 S.t1769 3.773
R1894 S.n1257 S.n1256 3.773
R1895 S.n1254 S.t2008 3.773
R1896 S.n1254 S.n1253 3.773
R1897 S.n1240 S.n1239 3.773
R1898 S.n1240 S.t1711 3.773
R1899 S.n692 S.n691 3.773
R1900 S.n692 S.t327 3.773
R1901 S.n703 S.t1200 3.773
R1902 S.n703 S.n702 3.773
R1903 S.n700 S.t1420 3.773
R1904 S.n700 S.n699 3.773
R1905 S.n695 S.n694 3.773
R1906 S.n695 S.t1147 3.773
R1907 S.n675 S.n674 3.773
R1908 S.n675 S.t2062 3.773
R1909 S.n686 S.t408 3.773
R1910 S.n686 S.n685 3.773
R1911 S.n683 S.t631 3.773
R1912 S.n683 S.n682 3.773
R1913 S.n678 S.n677 3.773
R1914 S.n678 S.t362 3.773
R1915 S.n136 S.t121 3.773
R1916 S.n128 S.t1847 3.773
R1917 S.n129 S.t1366 3.773
R1918 S.n390 S.n389 3.773
R1919 S.n390 S.t1082 3.773
R1920 S.n401 S.t1950 3.773
R1921 S.n401 S.n400 3.773
R1922 S.n398 S.t2178 3.773
R1923 S.n398 S.n397 3.773
R1924 S.n393 S.n392 3.773
R1925 S.n393 S.t1896 3.773
R1926 S.n1156 S.n1155 3.773
R1927 S.n1156 S.t2116 3.773
R1928 S.n1169 S.t465 3.773
R1929 S.n1169 S.n1168 3.773
R1930 S.n1166 S.t684 3.773
R1931 S.n1166 S.n1165 3.773
R1932 S.n1153 S.n1152 3.773
R1933 S.n1153 S.t412 3.773
R1934 S.n6432 S.t2228 3.773
R1935 S.n6433 S.t2247 3.773
R1936 S.n6413 S.t522 3.773
R1937 S.n6253 S.n6252 3.773
R1938 S.n6253 S.t848 3.773
R1939 S.n6267 S.t1716 3.773
R1940 S.n6267 S.n6266 3.773
R1941 S.n6270 S.t1963 3.773
R1942 S.n6270 S.n6269 3.773
R1943 S.n6250 S.n6249 3.773
R1944 S.n6250 S.t1385 3.773
R1945 S.n5667 S.n5666 3.773
R1946 S.n5667 S.t284 3.773
R1947 S.n5678 S.t1150 3.773
R1948 S.n5678 S.n5677 3.773
R1949 S.n5675 S.t1373 3.773
R1950 S.n5675 S.n5674 3.773
R1951 S.n5664 S.n5663 3.773
R1952 S.n5664 S.t1096 3.773
R1953 S.n5195 S.n5194 3.773
R1954 S.n5195 S.t2213 3.773
R1955 S.n5210 S.t558 3.773
R1956 S.n5210 S.n5209 3.773
R1957 S.n5207 S.t781 3.773
R1958 S.n5207 S.n5206 3.773
R1959 S.n5192 S.n5191 3.773
R1960 S.n5192 S.t507 3.773
R1961 S.n4886 S.n4885 3.773
R1962 S.n4886 S.t1754 3.773
R1963 S.n4897 S.t2493 3.773
R1964 S.n4897 S.n4896 3.773
R1965 S.n4894 S.t209 3.773
R1966 S.n4894 S.n4893 3.773
R1967 S.n4883 S.n4882 3.773
R1968 S.n4883 S.t2435 3.773
R1969 S.n4418 S.n4417 3.773
R1970 S.n4418 S.t1187 3.773
R1971 S.n4433 S.t2051 3.773
R1972 S.n4433 S.n4432 3.773
R1973 S.n4430 S.t2270 3.773
R1974 S.n4430 S.n4429 3.773
R1975 S.n4415 S.n4414 3.773
R1976 S.n4415 S.t1995 3.773
R1977 S.n4087 S.n4086 3.773
R1978 S.n4087 S.t586 3.773
R1979 S.n4098 S.t1454 3.773
R1980 S.n4098 S.n4097 3.773
R1981 S.n4095 S.t1684 3.773
R1982 S.n4095 S.n4094 3.773
R1983 S.n4084 S.n4083 3.773
R1984 S.n4084 S.t1407 3.773
R1985 S.n3618 S.n3617 3.773
R1986 S.n3618 S.t1359 3.773
R1987 S.n3633 S.t870 3.773
R1988 S.n3633 S.n3632 3.773
R1989 S.n3630 S.t2451 3.773
R1990 S.n3630 S.n3629 3.773
R1991 S.n3615 S.n3614 3.773
R1992 S.n3615 S.t2173 3.773
R1993 S.n3203 S.n3202 3.773
R1994 S.n3203 S.t765 3.773
R1995 S.n3214 S.t1636 3.773
R1996 S.n3214 S.n3213 3.773
R1997 S.n3211 S.t1881 3.773
R1998 S.n3211 S.n3210 3.773
R1999 S.n3200 S.n3199 3.773
R2000 S.n3200 S.t1577 3.773
R2001 S.n2806 S.n2805 3.773
R2002 S.n2806 S.t196 3.773
R2003 S.n2821 S.t1068 3.773
R2004 S.n2821 S.n2820 3.773
R2005 S.n2818 S.t217 3.773
R2006 S.n2818 S.n2817 3.773
R2007 S.n2803 S.n2802 3.773
R2008 S.n2803 S.t1013 3.773
R2009 S.n2439 S.n2438 3.773
R2010 S.n2439 S.t1062 3.773
R2011 S.n2450 S.t1930 3.773
R2012 S.n2450 S.n2449 3.773
R2013 S.n2447 S.t2157 3.773
R2014 S.n2447 S.n2446 3.773
R2015 S.n2436 S.n2435 3.773
R2016 S.n2436 S.t1872 3.773
R2017 S.n1969 S.n1968 3.773
R2018 S.n1969 S.t744 3.773
R2019 S.n1984 S.t1617 3.773
R2020 S.n1984 S.n1983 3.773
R2021 S.n1981 S.t1858 3.773
R2022 S.n1981 S.n1980 3.773
R2023 S.n1966 S.n1965 3.773
R2024 S.n1966 S.t1289 3.773
R2025 S.n1583 S.n1582 3.773
R2026 S.n1583 S.t176 3.773
R2027 S.n1594 S.t1050 3.773
R2028 S.n1594 S.n1593 3.773
R2029 S.n1591 S.t1278 3.773
R2030 S.n1591 S.n1590 3.773
R2031 S.n1580 S.n1579 3.773
R2032 S.n1580 S.t994 3.773
R2033 S.n227 S.t924 3.773
R2034 S.n228 S.t76 3.773
R2035 S.n225 S.t976 3.773
R2036 S.n413 S.n412 3.773
R2037 S.n413 S.t678 3.773
R2038 S.n424 S.t1549 3.773
R2039 S.n424 S.n423 3.773
R2040 S.n421 S.t1789 3.773
R2041 S.n421 S.n420 3.773
R2042 S.n416 S.n415 3.773
R2043 S.n416 S.t1498 3.773
R2044 S.n7195 S.t1649 3.773
R2045 S.n7196 S.t242 3.773
R2046 S.n7175 S.t2464 3.773
R2047 S.n6999 S.n6998 3.773
R2048 S.n6999 S.t1081 3.773
R2049 S.n7014 S.t1949 3.773
R2050 S.n7014 S.n7013 3.773
R2051 S.n7017 S.t2177 3.773
R2052 S.n7017 S.n7016 3.773
R2053 S.n7002 S.n7001 3.773
R2054 S.n7002 S.t1895 3.773
R2055 S.n6439 S.n6438 3.773
R2056 S.n6439 S.t498 3.773
R2057 S.n6450 S.t1365 3.773
R2058 S.n6450 S.n6449 3.773
R2059 S.n6447 S.t517 3.773
R2060 S.n6447 S.n6446 3.773
R2061 S.n6442 S.n6441 3.773
R2062 S.n6442 S.t1310 3.773
R2063 S.n5984 S.n5983 3.773
R2064 S.n5984 S.t1631 3.773
R2065 S.n6004 S.t2503 3.773
R2066 S.n6004 S.n6003 3.773
R2067 S.n6001 S.t221 3.773
R2068 S.n6001 S.n6000 3.773
R2069 S.n5987 S.n5986 3.773
R2070 S.n5987 S.t2170 3.773
R2071 S.n5684 S.n5683 3.773
R2072 S.n5684 S.t1196 3.773
R2073 S.n5695 S.t1933 3.773
R2074 S.n5695 S.n5694 3.773
R2075 S.n5692 S.t2162 3.773
R2076 S.n5692 S.n5691 3.773
R2077 S.n5687 S.n5686 3.773
R2078 S.n5687 S.t1877 3.773
R2079 S.n5219 S.n5218 3.773
R2080 S.n5219 S.t596 3.773
R2081 S.n5239 S.t1463 3.773
R2082 S.n5239 S.n5238 3.773
R2083 S.n5236 S.t1696 3.773
R2084 S.n5236 S.n5235 3.773
R2085 S.n5222 S.n5221 3.773
R2086 S.n5222 S.t1415 3.773
R2087 S.n4903 S.n4902 3.773
R2088 S.n4903 S.t2536 3.773
R2089 S.n4914 S.t886 3.773
R2090 S.n4914 S.n4913 3.773
R2091 S.n4911 S.t1135 3.773
R2092 S.n4911 S.n4910 3.773
R2093 S.n4906 S.n4905 3.773
R2094 S.n4906 S.t832 3.773
R2095 S.n4442 S.n4441 3.773
R2096 S.n4442 S.t776 3.773
R2097 S.n4462 S.t315 3.773
R2098 S.n4462 S.n4461 3.773
R2099 S.n4459 S.t1890 3.773
R2100 S.n4459 S.n4458 3.773
R2101 S.n4445 S.n4444 3.773
R2102 S.n4445 S.t1588 3.773
R2103 S.n4104 S.n4103 3.773
R2104 S.n4104 S.t203 3.773
R2105 S.n4115 S.t1078 3.773
R2106 S.n4115 S.n4114 3.773
R2107 S.n4112 S.t1305 3.773
R2108 S.n4112 S.n4111 3.773
R2109 S.n4107 S.n4106 3.773
R2110 S.n4107 S.t1022 3.773
R2111 S.n3642 S.n3641 3.773
R2112 S.n3642 S.t2143 3.773
R2113 S.n3662 S.t490 3.773
R2114 S.n3662 S.n3661 3.773
R2115 S.n3659 S.t708 3.773
R2116 S.n3659 S.n3658 3.773
R2117 S.n3645 S.n3644 3.773
R2118 S.n3645 S.t438 3.773
R2119 S.n3220 S.n3219 3.773
R2120 S.n3220 S.t1554 3.773
R2121 S.n3231 S.t2420 3.773
R2122 S.n3231 S.n3230 3.773
R2123 S.n3228 S.t129 3.773
R2124 S.n3228 S.n3227 3.773
R2125 S.n3223 S.n3222 3.773
R2126 S.n3223 S.t2366 3.773
R2127 S.n2830 S.n2829 3.773
R2128 S.n2830 S.t983 3.773
R2129 S.n2850 S.t1854 3.773
R2130 S.n2850 S.n2849 3.773
R2131 S.n2847 S.t1006 3.773
R2132 S.n2847 S.n2846 3.773
R2133 S.n2833 S.n2832 3.773
R2134 S.n2833 S.t1791 3.773
R2135 S.n2456 S.n2455 3.773
R2136 S.n2456 S.t1846 3.773
R2137 S.n2467 S.t188 3.773
R2138 S.n2467 S.n2466 3.773
R2139 S.n2464 S.t425 3.773
R2140 S.n2464 S.n2463 3.773
R2141 S.n2459 S.n2458 3.773
R2142 S.n2459 S.t118 3.773
R2143 S.n1993 S.n1992 3.773
R2144 S.n1993 S.t1536 3.773
R2145 S.n2013 S.t2405 3.773
R2146 S.n2013 S.n2012 3.773
R2147 S.n2010 S.t98 3.773
R2148 S.n2010 S.n2009 3.773
R2149 S.n1996 S.n1995 3.773
R2150 S.n1996 S.t2079 3.773
R2151 S.n1600 S.n1599 3.773
R2152 S.n1600 S.t1098 3.773
R2153 S.n1611 S.t1832 3.773
R2154 S.n1611 S.n1610 3.773
R2155 S.n1608 S.t2065 3.773
R2156 S.n1608 S.n1607 3.773
R2157 S.n1603 S.n1602 3.773
R2158 S.n1603 S.t1775 3.773
R2159 S.n1178 S.n1177 3.773
R2160 S.n1178 S.t509 3.773
R2161 S.n1198 S.t1375 3.773
R2162 S.n1198 S.n1197 3.773
R2163 S.n1195 S.t1593 3.773
R2164 S.n1195 S.n1194 3.773
R2165 S.n1181 S.n1180 3.773
R2166 S.n1181 S.t1323 3.773
R2167 S.n659 S.n658 3.773
R2168 S.n659 S.t1274 3.773
R2169 S.n670 S.t780 3.773
R2170 S.n670 S.n669 3.773
R2171 S.n667 S.t2362 3.773
R2172 S.n667 S.n666 3.773
R2173 S.n662 S.n661 3.773
R2174 S.n662 S.t2088 3.773
R2175 S.n642 S.n641 3.773
R2176 S.n642 S.t1650 3.773
R2177 S.n653 S.t2392 3.773
R2178 S.n653 S.n652 3.773
R2179 S.n650 S.t88 3.773
R2180 S.n650 S.n649 3.773
R2181 S.n645 S.n644 3.773
R2182 S.n645 S.t2340 3.773
R2183 S.n123 S.t2136 3.773
R2184 S.n115 S.t1321 3.773
R2185 S.n116 S.t2187 3.773
R2186 S.n346 S.n345 3.773
R2187 S.n346 S.t1906 3.773
R2188 S.n357 S.t256 3.773
R2189 S.n357 S.n356 3.773
R2190 S.n354 S.t481 3.773
R2191 S.n354 S.n353 3.773
R2192 S.n349 S.n348 3.773
R2193 S.n349 S.t195 3.773
R2194 S.n1097 S.n1096 3.773
R2195 S.n1097 S.t543 3.773
R2196 S.n1110 S.t1409 3.773
R2197 S.n1110 S.n1109 3.773
R2198 S.n1107 S.t1638 3.773
R2199 S.n1107 S.n1106 3.773
R2200 S.n1094 S.n1093 3.773
R2201 S.n1094 S.t1358 3.773
R2202 S.n4860 S.t2573 3.773
R2203 S.n4861 S.t1164 3.773
R2204 S.n4841 S.t865 3.773
R2205 S.n4711 S.n4710 3.773
R2206 S.n4711 S.t2002 3.773
R2207 S.n4725 S.t355 3.773
R2208 S.n4725 S.n4724 3.773
R2209 S.n4728 S.t575 3.773
R2210 S.n4728 S.n4727 3.773
R2211 S.n4708 S.n4707 3.773
R2212 S.n4708 S.t298 3.773
R2213 S.n4051 S.n4050 3.773
R2214 S.n4051 S.t1413 3.773
R2215 S.n4062 S.t2277 3.773
R2216 S.n4062 S.n4061 3.773
R2217 S.n4059 S.t2513 3.773
R2218 S.n4059 S.n4058 3.773
R2219 S.n4048 S.n4047 3.773
R2220 S.n4048 S.t2230 3.773
R2221 S.n3557 S.n3556 3.773
R2222 S.n3557 S.t828 3.773
R2223 S.n3572 S.t1693 3.773
R2224 S.n3572 S.n3571 3.773
R2225 S.n3569 S.t1943 3.773
R2226 S.n3569 S.n3568 3.773
R2227 S.n3554 S.n3553 3.773
R2228 S.n3554 S.t1644 3.773
R2229 S.n3167 S.n3166 3.773
R2230 S.n3167 S.t384 3.773
R2231 S.n3178 S.t1133 3.773
R2232 S.n3178 S.n3177 3.773
R2233 S.n3175 S.t1355 3.773
R2234 S.n3175 S.n3174 3.773
R2235 S.n3164 S.n3163 3.773
R2236 S.n3164 S.t1075 3.773
R2237 S.n2745 S.n2744 3.773
R2238 S.n2745 S.t2313 3.773
R2239 S.n2760 S.t655 3.773
R2240 S.n2760 S.n2759 3.773
R2241 S.n2757 S.t2333 3.773
R2242 S.n2757 S.n2756 3.773
R2243 S.n2742 S.n2741 3.773
R2244 S.n2742 S.t604 3.773
R2245 S.n2403 S.n2402 3.773
R2246 S.n2403 S.t647 3.773
R2247 S.n2414 S.t1516 3.773
R2248 S.n2414 S.n2413 3.773
R2249 S.n2411 S.t1756 3.773
R2250 S.n2411 S.n2410 3.773
R2251 S.n2400 S.n2399 3.773
R2252 S.n2400 S.t1465 3.773
R2253 S.n1908 S.n1907 3.773
R2254 S.n1908 S.t1701 3.773
R2255 S.n1923 S.t1235 3.773
R2256 S.n1923 S.n1922 3.773
R2257 S.n1920 S.t296 3.773
R2258 S.n1920 S.n1919 3.773
R2259 S.n1905 S.n1904 3.773
R2260 S.n1905 S.t2237 3.773
R2261 S.n1547 S.n1546 3.773
R2262 S.n1547 S.t1139 3.773
R2263 S.n1558 S.t1999 3.773
R2264 S.n1558 S.n1557 3.773
R2265 S.n1555 S.t2224 3.773
R2266 S.n1555 S.n1554 3.773
R2267 S.n1544 S.n1543 3.773
R2268 S.n1544 S.t1946 3.773
R2269 S.n223 S.t405 3.773
R2270 S.n224 S.t2229 3.773
R2271 S.n221 S.t453 3.773
R2272 S.n369 S.n368 3.773
R2273 S.n369 S.t160 3.773
R2274 S.n380 S.t1038 3.773
R2275 S.n380 S.n379 3.773
R2276 S.n377 S.t1270 3.773
R2277 S.n377 S.n376 3.773
R2278 S.n372 S.n371 3.773
R2279 S.n372 S.t982 3.773
R2280 S.n5658 S.t2011 3.773
R2281 S.n5659 S.t581 3.773
R2282 S.n5638 S.t310 3.773
R2283 S.n5492 S.n5491 3.773
R2284 S.n5492 S.t1421 3.773
R2285 S.n5507 S.t2286 3.773
R2286 S.n5507 S.n5506 3.773
R2287 S.n5510 S.t2519 3.773
R2288 S.n5510 S.n5509 3.773
R2289 S.n5495 S.n5494 3.773
R2290 S.n5495 S.t2239 3.773
R2291 S.n4867 S.n4866 3.773
R2292 S.n4867 S.t838 3.773
R2293 S.n4878 S.t1703 3.773
R2294 S.n4878 S.n4877 3.773
R2295 S.n4875 S.t1951 3.773
R2296 S.n4875 S.n4874 3.773
R2297 S.n4870 S.n4869 3.773
R2298 S.n4870 S.t1648 3.773
R2299 S.n4381 S.n4380 3.773
R2300 S.n4381 S.t272 3.773
R2301 S.n4401 S.t1141 3.773
R2302 S.n4401 S.n4400 3.773
R2303 S.n4398 S.t1364 3.773
R2304 S.n4398 S.n4397 3.773
R2305 S.n4384 S.n4383 3.773
R2306 S.n4384 S.t1083 3.773
R2307 S.n4068 S.n4067 3.773
R2308 S.n4068 S.t2323 3.773
R2309 S.n4079 S.t548 3.773
R2310 S.n4079 S.n4078 3.773
R2311 S.n4076 S.t774 3.773
R2312 S.n4076 S.n4075 3.773
R2313 S.n4071 S.n4070 3.773
R2314 S.n4071 S.t497 3.773
R2315 S.n3581 S.n3580 3.773
R2316 S.n3581 S.t1741 3.773
R2317 S.n3601 S.t54 3.773
R2318 S.n3601 S.n3600 3.773
R2319 S.n3598 S.t333 3.773
R2320 S.n3598 S.n3597 3.773
R2321 S.n3584 S.n3583 3.773
R2322 S.n3584 S.t2552 3.773
R2323 S.n3184 S.n3183 3.773
R2324 S.n3184 S.t1175 3.773
R2325 S.n3195 S.t2034 3.773
R2326 S.n3195 S.n3194 3.773
R2327 S.n3192 S.t2261 3.773
R2328 S.n3192 S.n3191 3.773
R2329 S.n3187 S.n3186 3.773
R2330 S.n3187 S.t1984 3.773
R2331 S.n2769 S.n2768 3.773
R2332 S.n2769 S.t1937 3.773
R2333 S.n2789 S.t1447 3.773
R2334 S.n2789 S.n2788 3.773
R2335 S.n2786 S.t1959 3.773
R2336 S.n2786 S.n2785 3.773
R2337 S.n2772 S.n2771 3.773
R2338 S.n2772 S.t228 3.773
R2339 S.n2420 S.n2419 3.773
R2340 S.n2420 S.t281 3.773
R2341 S.n2431 S.t1148 3.773
R2342 S.n2431 S.n2430 3.773
R2343 S.n2428 S.t1371 3.773
R2344 S.n2428 S.n2427 3.773
R2345 S.n2423 S.n2422 3.773
R2346 S.n2423 S.t1091 3.773
R2347 S.n1932 S.n1931 3.773
R2348 S.n1932 S.t2490 3.773
R2349 S.n1952 S.t836 3.773
R2350 S.n1952 S.n1951 3.773
R2351 S.n1935 S.t1077 3.773
R2352 S.n1935 S.n1934 3.773
R2353 S.n1938 S.n1937 3.773
R2354 S.n1938 S.t505 3.773
R2355 S.n1564 S.n1563 3.773
R2356 S.n1564 S.t1920 3.773
R2357 S.n1575 S.t269 3.773
R2358 S.n1575 S.n1574 3.773
R2359 S.n1572 S.t492 3.773
R2360 S.n1572 S.n1571 3.773
R2361 S.n1567 S.n1566 3.773
R2362 S.n1567 S.t202 3.773
R2363 S.n1119 S.n1118 3.773
R2364 S.n1119 S.t1332 3.773
R2365 S.n1139 S.t2199 3.773
R2366 S.n1139 S.n1138 3.773
R2367 S.n1136 S.t2422 3.773
R2368 S.n1136 S.n1135 3.773
R2369 S.n1122 S.n1121 3.773
R2370 S.n1122 S.t2145 3.773
R2371 S.n626 S.n625 3.773
R2372 S.n626 S.t733 3.773
R2373 S.n637 S.t1606 3.773
R2374 S.n637 S.n636 3.773
R2375 S.n634 S.t1853 3.773
R2376 S.n634 S.n633 3.773
R2377 S.n629 S.n628 3.773
R2378 S.n629 S.t1553 3.773
R2379 S.n609 S.n608 3.773
R2380 S.n609 S.t2477 3.773
R2381 S.n620 S.t824 3.773
R2382 S.n620 S.n619 3.773
R2383 S.n617 S.t1070 3.773
R2384 S.n617 S.n616 3.773
R2385 S.n612 S.n611 3.773
R2386 S.n612 S.t767 3.773
R2387 S.n110 S.t561 3.773
R2388 S.n102 S.t2263 3.773
R2389 S.n103 S.t610 3.773
R2390 S.n302 S.n301 3.773
R2391 S.n302 S.t340 3.773
R2392 S.n313 S.t2361 3.773
R2393 S.n313 S.n312 3.773
R2394 S.n310 S.t1426 3.773
R2395 S.n310 S.n309 3.773
R2396 S.n305 S.n304 3.773
R2397 S.n305 S.t1155 3.773
R2398 S.n1038 S.n1037 3.773
R2399 S.n1038 S.t135 3.773
R2400 S.n1051 S.t1018 3.773
R2401 S.n1051 S.n1050 3.773
R2402 S.n1048 S.t1251 3.773
R2403 S.n1048 S.n1047 3.773
R2404 S.n1035 S.n1034 3.773
R2405 S.n1035 S.t960 3.773
R2406 S.n3141 S.t1214 3.773
R2407 S.n3142 S.t2296 3.773
R2408 S.n3122 S.t2018 3.773
R2409 S.n3099 S.n3098 3.773
R2410 S.n3099 S.t614 3.773
R2411 S.n3113 S.t1483 3.773
R2412 S.n3113 S.n3112 3.773
R2413 S.n3116 S.t638 3.773
R2414 S.n3116 S.n3115 3.773
R2415 S.n3096 S.n3095 3.773
R2416 S.n3096 S.t1429 3.773
R2417 S.n2367 S.n2366 3.773
R2418 S.n2367 S.t1477 3.773
R2419 S.n2378 S.t2345 3.773
R2420 S.n2378 S.n2377 3.773
R2421 S.n2375 S.t2576 3.773
R2422 S.n2375 S.n2374 3.773
R2423 S.n2364 S.n2363 3.773
R2424 S.n2364 S.t2291 3.773
R2425 S.n1847 S.n1846 3.773
R2426 S.n1847 S.t1194 3.773
R2427 S.n1862 S.t2059 3.773
R2428 S.n1862 S.n1861 3.773
R2429 S.n1859 S.t2276 3.773
R2430 S.n1859 S.n1858 3.773
R2431 S.n1844 S.n1843 3.773
R2432 S.n1844 S.t1707 3.773
R2433 S.n1511 S.n1510 3.773
R2434 S.n1511 S.t716 3.773
R2435 S.n1522 S.t1464 3.773
R2436 S.n1522 S.n1521 3.773
R2437 S.n1519 S.t1697 3.773
R2438 S.n1519 S.n1518 3.773
R2439 S.n1508 S.n1507 3.773
R2440 S.n1508 S.t1416 3.773
R2441 S.n219 S.t1348 3.773
R2442 S.n220 S.t533 3.773
R2443 S.n217 S.t1400 3.773
R2444 S.n325 S.n324 3.773
R2445 S.n325 S.t1126 3.773
R2446 S.n336 S.t1988 3.773
R2447 S.n336 S.n335 3.773
R2448 S.n333 S.t2216 3.773
R2449 S.n333 S.n332 3.773
R2450 S.n328 S.n327 3.773
R2451 S.n328 S.t1939 3.773
R2452 S.n4042 S.t624 3.773
R2453 S.n4043 S.t1726 3.773
R2454 S.n4022 S.t1438 3.773
R2455 S.n3915 S.n3914 3.773
R2456 S.n3915 S.t2562 3.773
R2457 S.n3930 S.t914 3.773
R2458 S.n3930 S.n3929 3.773
R2459 S.n3933 S.t1158 3.773
R2460 S.n3933 S.n3932 3.773
R2461 S.n3918 S.n3917 3.773
R2462 S.n3918 S.t860 3.773
R2463 S.n3148 S.n3147 3.773
R2464 S.n3148 S.t1992 3.773
R2465 S.n3159 S.t344 3.773
R2466 S.n3159 S.n3158 3.773
R2467 S.n3156 S.t565 3.773
R2468 S.n3156 S.n3155 3.773
R2469 S.n3151 S.n3150 3.773
R2470 S.n3151 S.t290 3.773
R2471 S.n2708 S.n2707 3.773
R2472 S.n2708 S.t1405 3.773
R2473 S.n2728 S.t2267 3.773
R2474 S.n2728 S.n2727 3.773
R2475 S.n2725 S.t1425 3.773
R2476 S.n2725 S.n2724 3.773
R2477 S.n2711 S.n2710 3.773
R2478 S.n2711 S.t2221 3.773
R2479 S.n2384 S.n2383 3.773
R2480 S.n2384 S.t2385 3.773
R2481 S.n2395 S.t608 3.773
R2482 S.n2395 S.n2394 3.773
R2483 S.n2392 S.t839 3.773
R2484 S.n2392 S.n2391 3.773
R2485 S.n2387 S.n2386 3.773
R2486 S.n2387 S.t559 3.773
R2487 S.n1871 S.n1870 3.773
R2488 S.n1871 S.t2097 3.773
R2489 S.n1891 S.t444 3.773
R2490 S.n1891 S.n1890 3.773
R2491 S.n1888 S.t666 3.773
R2492 S.n1888 S.n1887 3.773
R2493 S.n1874 S.n1873 3.773
R2494 S.n1874 S.t74 3.773
R2495 S.n1528 S.n1527 3.773
R2496 S.n1528 S.t1507 3.773
R2497 S.n1539 S.t2373 3.773
R2498 S.n1539 S.n1538 3.773
R2499 S.n1536 S.t52 3.773
R2500 S.n1536 S.n1535 3.773
R2501 S.n1531 S.n1530 3.773
R2502 S.n1531 S.t2322 3.773
R2503 S.n1060 S.n1059 3.773
R2504 S.n1060 S.t2273 3.773
R2505 S.n1080 S.t1798 3.773
R2506 S.n1080 S.n1079 3.773
R2507 S.n1077 S.t855 3.773
R2508 S.n1077 S.n1076 3.773
R2509 S.n1063 S.n1062 3.773
R2510 S.n1063 S.t571 3.773
R2511 S.n593 S.n592 3.773
R2512 S.n593 S.t1689 3.773
R2513 S.n604 S.t2558 3.773
R2514 S.n604 S.n603 3.773
R2515 S.n601 S.t287 3.773
R2516 S.n601 S.n600 3.773
R2517 S.n596 S.n595 3.773
R2518 S.n596 S.t2507 3.773
R2519 S.n576 S.n575 3.773
R2520 S.n576 S.t2089 3.773
R2521 S.n587 S.t435 3.773
R2522 S.n587 S.n586 3.773
R2523 S.n584 S.t657 3.773
R2524 S.n584 S.n583 3.773
R2525 S.n579 S.n578 3.773
R2526 S.n579 S.t386 3.773
R2527 S.n97 S.t2550 3.773
R2528 S.n89 S.t1874 3.773
R2529 S.n90 S.t46 3.773
R2530 S.n258 S.n257 3.773
R2531 S.n258 S.t2320 3.773
R2532 S.n269 S.t665 3.773
R2533 S.n269 S.n268 3.773
R2534 S.n266 S.t903 3.773
R2535 S.n266 S.n265 3.773
R2536 S.n261 S.n260 3.773
R2537 S.n261 S.t616 3.773
R2538 S.n1445 S.n1444 3.773
R2539 S.n1445 S.t968 3.773
R2540 S.n1457 S.t1838 3.773
R2541 S.n1457 S.n1456 3.773
R2542 S.n1460 S.t2073 3.773
R2543 S.n1460 S.n1459 3.773
R2544 S.n1442 S.n1441 3.773
R2545 S.n1442 S.t1783 3.773
R2546 S.n1485 S.t1542 3.773
R2547 S.n1486 S.t108 3.773
R2548 S.n1466 S.t2356 3.773
R2549 S.n215 S.t950 3.773
R2550 S.n216 S.t119 3.773
R2551 S.n213 S.t1007 3.773
R2552 S.n281 S.n280 3.773
R2553 S.n281 S.t702 3.773
R2554 S.n292 S.t1570 3.773
R2555 S.n292 S.n291 3.773
R2556 S.n289 S.t1820 3.773
R2557 S.n289 S.n288 3.773
R2558 S.n284 S.n283 3.773
R2559 S.n284 S.t1526 3.773
R2560 S.n2358 S.t687 3.773
R2561 S.n2359 S.t1794 3.773
R2562 S.n2338 S.t1502 3.773
R2563 S.n2268 S.n2267 3.773
R2564 S.n2268 S.t404 3.773
R2565 S.n2283 S.t1269 3.773
R2566 S.n2283 S.n2282 3.773
R2567 S.n2286 S.t1493 3.773
R2568 S.n2286 S.n2285 3.773
R2569 S.n2271 S.n2270 3.773
R2570 S.n2271 S.t930 3.773
R2571 S.n1492 S.n1491 3.773
R2572 S.n1492 S.t2330 3.773
R2573 S.n1503 S.t674 3.773
R2574 S.n1503 S.n1502 3.773
R2575 S.n1500 S.t913 3.773
R2576 S.n1500 S.n1499 3.773
R2577 S.n1495 S.n1494 3.773
R2578 S.n1495 S.t623 3.773
R2579 S.n1001 S.n1000 3.773
R2580 S.n1001 S.t1755 3.773
R2581 S.n1021 S.t73 3.773
R2582 S.n1021 S.n1020 3.773
R2583 S.n1018 S.t346 3.773
R2584 S.n1018 S.n1017 3.773
R2585 S.n1004 S.n1003 3.773
R2586 S.n1004 S.t2565 3.773
R2587 S.n560 S.n559 3.773
R2588 S.n560 S.t1299 3.773
R2589 S.n571 S.t2049 3.773
R2590 S.n571 S.n570 3.773
R2591 S.n568 S.t2266 3.773
R2592 S.n568 S.n567 3.773
R2593 S.n563 S.n562 3.773
R2594 S.n563 S.t1994 3.773
R2595 S.n543 S.n542 3.773
R2596 S.n543 S.t395 3.773
R2597 S.n554 S.t1261 3.773
R2598 S.n554 S.n553 3.773
R2599 S.n551 S.t1485 3.773
R2600 S.n551 S.n550 3.773
R2601 S.n546 S.n545 3.773
R2602 S.n546 S.t1216 3.773
R2603 S.n84 S.t172 3.773
R2604 S.n61 S.t991 3.773
R2605 S.n958 S.t234 3.773
R2606 S.n960 S.t1000 3.773
R2607 S.n962 S.t698 3.773
R2608 S.n798 S.n797 3.773
R2609 S.n798 S.t1383 3.773
R2610 S.n807 S.t1189 3.773
R2611 S.n807 S.n806 3.773
R2612 S.n810 S.t2377 3.773
R2613 S.n810 S.n809 3.773
R2614 S.n801 S.n800 3.773
R2615 S.n801 S.t989 3.773
R2616 S.n1801 S.n1800 3.773
R2617 S.n1801 S.t349 3.773
R2618 S.n1810 S.t1217 3.773
R2619 S.n1810 S.n1809 3.773
R2620 S.n1813 S.t980 3.773
R2621 S.n1813 S.n1812 3.773
R2622 S.n1804 S.n1803 3.773
R2623 S.n1804 S.t122 3.773
R2624 S.n1464 S.n1463 3.773
R2625 S.n1464 S.t370 3.773
R2626 S.n1787 S.t1236 3.773
R2627 S.n1787 S.n1786 3.773
R2628 S.n1790 S.t1008 3.773
R2629 S.n1790 S.n1789 3.773
R2630 S.n1793 S.n1792 3.773
R2631 S.n1793 S.t154 3.773
R2632 S.n2308 S.n2307 3.773
R2633 S.n2308 S.t393 3.773
R2634 S.n2320 S.t1259 3.773
R2635 S.n2320 S.n2319 3.773
R2636 S.n2323 S.t1036 3.773
R2637 S.n2323 S.n2322 3.773
R2638 S.n2311 S.n2310 3.773
R2639 S.n2311 S.t1048 3.773
R2640 S.n2290 S.n2289 3.773
R2641 S.n2290 S.t1273 3.773
R2642 S.n2293 S.t2139 3.773
R2643 S.n2293 S.n2292 3.773
R2644 S.n2296 S.t1919 3.773
R2645 S.n2296 S.n2295 3.773
R2646 S.n2299 S.n2298 3.773
R2647 S.n2299 S.t1076 3.773
R2648 S.n3436 S.n3435 3.773
R2649 S.n3436 S.t1014 3.773
R2650 S.n3448 S.t1882 3.773
R2651 S.n3448 S.n3447 3.773
R2652 S.n3451 S.t1944 3.773
R2653 S.n3451 S.n3450 3.773
R2654 S.n3439 S.n3438 3.773
R2655 S.n3439 S.t803 3.773
R2656 S.n3120 S.n3119 3.773
R2657 S.n3120 S.t1043 3.773
R2658 S.n3421 S.t1912 3.773
R2659 S.n3421 S.n3420 3.773
R2660 S.n3424 S.t1669 3.773
R2661 S.n3424 S.n3423 3.773
R2662 S.n3427 S.n3426 3.773
R2663 S.n3427 S.t831 3.773
R2664 S.n3955 S.n3954 3.773
R2665 S.n3955 S.t1067 3.773
R2666 S.n3967 S.t1936 3.773
R2667 S.n3967 S.n3966 3.773
R2668 S.n3970 S.t1695 3.773
R2669 S.n3970 S.n3969 3.773
R2670 S.n3958 S.n3957 3.773
R2671 S.n3958 S.t858 3.773
R2672 S.n3937 S.n3936 3.773
R2673 S.n3937 S.t1094 3.773
R2674 S.n3940 S.t1962 3.773
R2675 S.n3940 S.n3939 3.773
R2676 S.n3943 S.t1722 3.773
R2677 S.n3943 S.n3942 3.773
R2678 S.n3946 S.n3945 3.773
R2679 S.n3946 S.t882 3.773
R2680 S.n4750 S.n4749 3.773
R2681 S.n4750 S.t1122 3.773
R2682 S.n4762 S.t246 3.773
R2683 S.n4762 S.n4761 3.773
R2684 S.n4765 S.t1749 3.773
R2685 S.n4765 S.n4764 3.773
R2686 S.n4753 S.n4752 3.773
R2687 S.n4753 S.t911 3.773
R2688 S.n4732 S.n4731 3.773
R2689 S.n4732 S.t2467 3.773
R2690 S.n4735 S.t688 3.773
R2691 S.n4735 S.n4734 3.773
R2692 S.n4738 S.t931 3.773
R2693 S.n4738 S.n4737 3.773
R2694 S.n4741 S.n4740 3.773
R2695 S.n4741 S.t639 3.773
R2696 S.n5532 S.n5531 3.773
R2697 S.n5532 S.t415 3.773
R2698 S.n5544 S.t1280 3.773
R2699 S.n5544 S.n5543 3.773
R2700 S.n5547 S.t1505 3.773
R2701 S.n5547 S.n5546 3.773
R2702 S.n5535 S.n5534 3.773
R2703 S.n5535 S.t1233 3.773
R2704 S.n5514 S.n5513 3.773
R2705 S.n5514 S.t995 3.773
R2706 S.n5517 S.t1860 3.773
R2707 S.n5517 S.n5516 3.773
R2708 S.n5520 S.t2094 3.773
R2709 S.n5520 S.n5519 3.773
R2710 S.n5523 S.n5522 3.773
R2711 S.n5523 S.t1803 3.773
R2712 S.n6292 S.n6291 3.773
R2713 S.n6292 S.t1562 3.773
R2714 S.n6304 S.t2431 3.773
R2715 S.n6304 S.n6303 3.773
R2716 S.n6307 S.t141 3.773
R2717 S.n6307 S.n6306 3.773
R2718 S.n6295 S.n6294 3.773
R2719 S.n6295 S.t2107 3.773
R2720 S.n6274 S.n6273 3.773
R2721 S.n6274 S.t430 3.773
R2722 S.n6277 S.t1295 3.773
R2723 S.n6277 S.n6276 3.773
R2724 S.n6280 S.t451 3.773
R2725 S.n6280 S.n6279 3.773
R2726 S.n6283 S.n6282 3.773
R2727 S.n6283 S.t1246 3.773
R2728 S.n7039 S.n7038 3.773
R2729 S.n7039 S.t1016 3.773
R2730 S.n7051 S.t1884 3.773
R2731 S.n7051 S.n7050 3.773
R2732 S.n7054 S.t2113 3.773
R2733 S.n7054 S.n7053 3.773
R2734 S.n7042 S.n7041 3.773
R2735 S.n7042 S.t1826 3.773
R2736 S.n7021 S.n7020 3.773
R2737 S.n7021 S.t1578 3.773
R2738 S.n7024 S.t2452 3.773
R2739 S.n7024 S.n7023 3.773
R2740 S.n7027 S.t168 3.773
R2741 S.n7027 S.n7026 3.773
R2742 S.n7030 S.n7029 3.773
R2743 S.n7030 S.t2399 3.773
R2744 S.n8050 S.n8049 3.773
R2745 S.n8050 S.t2174 3.773
R2746 S.n8062 S.t519 3.773
R2747 S.n8062 S.n8061 3.773
R2748 S.n8065 S.t739 3.773
R2749 S.n8065 S.n8064 3.773
R2750 S.n8053 S.n8052 3.773
R2751 S.n8053 S.t470 3.773
R2752 S.n7746 S.n7745 3.773
R2753 S.n7746 S.t238 3.773
R2754 S.n8035 S.t2271 3.773
R2755 S.n8035 S.n8034 3.773
R2756 S.n8038 S.t1338 3.773
R2757 S.n8038 S.n8037 3.773
R2758 S.n8041 S.n8040 3.773
R2759 S.n8041 S.t1053 3.773
R2760 S.n8762 S.n8761 3.773
R2761 S.n8762 S.t1996 3.773
R2762 S.n8774 S.t348 3.773
R2763 S.n8774 S.n8773 3.773
R2764 S.n8777 S.t569 3.773
R2765 S.n8777 S.n8776 3.773
R2766 S.n8765 S.n8764 3.773
R2767 S.n8765 S.t295 3.773
R2768 S.n8458 S.n8457 3.773
R2769 S.n8458 S.t2568 3.773
R2770 S.n8747 S.t782 3.773
R2771 S.n8747 S.n8746 3.773
R2772 S.n8750 S.t1029 3.773
R2773 S.n8750 S.n8749 3.773
R2774 S.n8753 S.n8752 3.773
R2775 S.n8753 S.t725 3.773
R2776 S.n9166 S.n9165 3.773
R2777 S.n9166 S.t510 3.773
R2778 S.n9178 S.t1376 3.773
R2779 S.n9178 S.n9177 3.773
R2780 S.n9181 S.t1597 3.773
R2781 S.n9181 S.n9180 3.773
R2782 S.n9169 S.n9168 3.773
R2783 S.n9169 S.t1325 3.773
R2784 S.n9148 S.n9147 3.773
R2785 S.n9148 S.t1100 3.773
R2786 S.n9151 S.t1965 3.773
R2787 S.n9151 S.n9150 3.773
R2788 S.n9154 S.t2193 3.773
R2789 S.n9154 S.n9153 3.773
R2790 S.n9157 S.n9156 3.773
R2791 S.n9157 S.t1913 3.773
R2792 S.n9843 S.n9842 3.773
R2793 S.n9843 S.t1661 3.773
R2794 S.n9855 S.t2530 3.773
R2795 S.n9855 S.n9854 3.773
R2796 S.n9858 S.t262 3.773
R2797 S.n9858 S.n9857 3.773
R2798 S.n9846 S.n9845 3.773
R2799 S.n9846 S.t171 3.773
R2800 S.n9825 S.n9824 3.773
R2801 S.n9825 S.t2456 3.773
R2802 S.n9828 S.t801 3.773
R2803 S.n9828 S.n9827 3.773
R2804 S.n9831 S.t1047 3.773
R2805 S.n9831 S.n9830 3.773
R2806 S.n9834 S.n9833 3.773
R2807 S.n9834 S.t742 3.773
R2808 S.n10501 S.n10500 3.773
R2809 S.n10501 S.t521 3.773
R2810 S.n10513 S.t1389 3.773
R2811 S.n10513 S.n10512 3.773
R2812 S.n10516 S.t1615 3.773
R2813 S.n10516 S.n10515 3.773
R2814 S.n10504 S.n10503 3.773
R2815 S.n10504 S.t1340 3.773
R2816 S.n10483 S.n10482 3.773
R2817 S.n10483 S.t1114 3.773
R2818 S.n10486 S.t1978 3.773
R2819 S.n10486 S.n10485 3.773
R2820 S.n10489 S.t2205 3.773
R2821 S.n10489 S.n10488 3.773
R2822 S.n10492 S.n10491 3.773
R2823 S.n10492 S.t1925 3.773
R2824 S.n11129 S.n11128 3.773
R2825 S.n11129 S.t1678 3.773
R2826 S.n11141 S.t1221 3.773
R2827 S.n11141 S.n11140 3.773
R2828 S.n11144 S.t276 3.773
R2829 S.n11144 S.n11143 3.773
R2830 S.n11132 S.n11131 3.773
R2831 S.n11132 S.t2495 3.773
R2832 S.n11111 S.n11110 3.773
R2833 S.n11111 S.t922 3.773
R2834 S.n11114 S.t1788 3.773
R2835 S.n11114 S.n11113 3.773
R2836 S.n11117 S.t2026 3.773
R2837 S.n11117 S.n11116 3.773
R2838 S.n11120 S.n11119 3.773
R2839 S.n11120 S.t1733 3.773
R2840 S.n12057 S.n12056 3.773
R2841 S.n12057 S.t1497 3.773
R2842 S.n12069 S.t2360 3.773
R2843 S.n12069 S.n12068 3.773
R2844 S.n12072 S.t37 3.773
R2845 S.n12072 S.n12071 3.773
R2846 S.n12060 S.n12059 3.773
R2847 S.n12060 S.t2314 3.773
R2848 S.n12336 S.n12335 3.773
R2849 S.n12336 S.t2087 3.773
R2850 S.n12346 S.t314 3.773
R2851 S.n12346 S.n12345 3.773
R2852 S.n12349 S.t539 3.773
R2853 S.n12349 S.n12348 3.773
R2854 S.n12339 S.n12338 3.773
R2855 S.n12339 S.t264 3.773
R2856 S.n11861 S.n11860 3.773
R2857 S.n11861 S.t2534 3.773
R2858 S.n11875 S.t883 3.773
R2859 S.n11875 S.n11874 3.773
R2860 S.n11872 S.t1134 3.773
R2861 S.n11872 S.n11871 3.773
R2862 S.n11864 S.n11863 3.773
R2863 S.n11864 S.t829 3.773
R2864 S.n11933 S.t2017 3.773
R2865 S.n11930 S.t2540 3.773
R2866 S.n11931 S.t890 3.773
R2867 S.n1816 S.t2529 3.773
R2868 S.n1818 S.t429 3.773
R2869 S.n1820 S.t126 3.773
R2870 S.n1773 S.n1772 3.773
R2871 S.n1773 S.t1180 3.773
R2872 S.n1781 S.t2016 3.773
R2873 S.n1781 S.n1780 3.773
R2874 S.n1784 S.t2112 3.773
R2875 S.n1784 S.n1783 3.773
R2876 S.n1776 S.n1775 3.773
R2877 S.n1776 S.t697 3.773
R2878 S.n2331 S.n2330 3.773
R2879 S.n2331 S.t1186 3.773
R2880 S.n2653 S.t2050 3.773
R2881 S.n2653 S.n2652 3.773
R2882 S.n2656 S.t1814 3.773
R2883 S.n2656 S.n2655 3.773
R2884 S.n2328 S.n2327 3.773
R2885 S.n2328 S.t1831 3.773
R2886 S.n11937 S.t289 3.773
R2887 S.n11935 S.t807 3.773
R2888 S.n11934 S.t1673 3.773
R2889 S.n11850 S.n11849 3.773
R2890 S.n11850 S.t932 3.773
R2891 S.n11857 S.t1796 3.773
R2892 S.n11857 S.n11856 3.773
R2893 S.n11854 S.t2035 3.773
R2894 S.n11854 S.n11853 3.773
R2895 S.n11847 S.n11846 3.773
R2896 S.n11847 S.t1742 3.773
R2897 S.n12357 S.n12356 3.773
R2898 S.n12357 S.t361 3.773
R2899 S.n12361 S.t1229 3.773
R2900 S.n12361 S.n12360 3.773
R2901 S.n12364 S.t1448 3.773
R2902 S.n12364 S.n12363 3.773
R2903 S.n12354 S.n12353 3.773
R2904 S.n12354 S.t1171 3.773
R2905 S.n12080 S.n12079 3.773
R2906 S.n12080 S.t1124 3.773
R2907 S.n12085 S.t630 3.773
R2908 S.n12085 S.n12084 3.773
R2909 S.n12088 S.t2214 3.773
R2910 S.n12088 S.n12087 3.773
R2911 S.n12077 S.n12076 3.773
R2912 S.n12077 S.t1938 3.773
R2913 S.n11166 S.n11165 3.773
R2914 S.n11166 S.t534 3.773
R2915 S.n11163 S.t1401 3.773
R2916 S.n11163 S.n11162 3.773
R2917 S.n11160 S.t1623 3.773
R2918 S.n11160 S.n11159 3.773
R2919 S.n11157 S.n11156 3.773
R2920 S.n11157 S.t1349 3.773
R2921 S.n11152 S.n11151 3.773
R2922 S.n11152 S.t2463 3.773
R2923 S.n11172 S.t811 3.773
R2924 S.n11172 S.n11171 3.773
R2925 S.n11175 S.t1056 3.773
R2926 S.n11175 S.n11174 3.773
R2927 S.n11149 S.n11148 3.773
R2928 S.n11149 S.t751 3.773
R2929 S.n10538 S.n10537 3.773
R2930 S.n10538 S.t1894 3.773
R2931 S.n10535 S.t241 3.773
R2932 S.n10535 S.n10534 3.773
R2933 S.n10532 S.t473 3.773
R2934 S.n10532 S.n10531 3.773
R2935 S.n10529 S.n10528 3.773
R2936 S.n10529 S.t180 3.773
R2937 S.n10524 S.n10523 3.773
R2938 S.n10524 S.t1308 3.773
R2939 S.n10544 S.t2176 3.773
R2940 S.n10544 S.n10543 3.773
R2941 S.n10547 S.t2401 3.773
R2942 S.n10547 S.n10546 3.773
R2943 S.n10521 S.n10520 3.773
R2944 S.n10521 S.t2128 3.773
R2945 S.n9880 S.n9879 3.773
R2946 S.n9880 S.t713 3.773
R2947 S.n9877 S.t1581 3.773
R2948 S.n9877 S.n9876 3.773
R2949 S.n9874 S.t1827 3.773
R2950 S.n9874 S.n9873 3.773
R2951 S.n9871 S.n9870 3.773
R2952 S.n9871 S.t1533 3.773
R2953 S.n9866 S.n9865 3.773
R2954 S.n9866 S.t2448 3.773
R2955 S.n9886 S.t793 3.773
R2956 S.n9886 S.n9885 3.773
R2957 S.n9889 S.t1045 3.773
R2958 S.n9889 S.n9888 3.773
R2959 S.n9863 S.n9862 3.773
R2960 S.n9863 S.t959 3.773
R2961 S.n9203 S.n9202 3.773
R2962 S.n9203 S.t2003 3.773
R2963 S.n9200 S.t226 3.773
R2964 S.n9200 S.n9199 3.773
R2965 S.n9197 S.t458 3.773
R2966 S.n9197 S.n9196 3.773
R2967 S.n9194 S.n9193 3.773
R2968 S.n9194 S.t167 3.773
R2969 S.n9189 S.n9188 3.773
R2970 S.n9189 S.t1417 3.773
R2971 S.n9209 S.t2279 3.773
R2972 S.n9209 S.n9208 3.773
R2973 S.n9212 S.t2517 3.773
R2974 S.n9212 S.n9211 3.773
R2975 S.n9186 S.n9185 3.773
R2976 S.n9186 S.t2233 3.773
R2977 S.n8799 S.n8798 3.773
R2978 S.n8799 S.t2184 3.773
R2979 S.n8796 S.t1698 3.773
R2980 S.n8796 S.n8795 3.773
R2981 S.n8793 S.t748 3.773
R2982 S.n8793 S.n8792 3.773
R2983 S.n8790 S.n8789 3.773
R2984 S.n8790 S.t479 3.773
R2985 S.n8785 S.n8784 3.773
R2986 S.n8785 S.t1589 3.773
R2987 S.n8805 S.t2462 3.773
R2988 S.n8805 S.n8804 3.773
R2989 S.n8808 S.t179 3.773
R2990 S.n8808 S.n8807 3.773
R2991 S.n8782 S.n8781 3.773
R2992 S.n8782 S.t2407 3.773
R2993 S.n8087 S.n8086 3.773
R2994 S.n8087 S.t1023 3.773
R2995 S.n8084 S.t1891 3.773
R2996 S.n8084 S.n8083 3.773
R2997 S.n8081 S.t2123 3.773
R2998 S.n8081 S.n8080 3.773
R2999 S.n8078 S.n8077 3.773
R3000 S.n8078 S.t1837 3.773
R3001 S.n8073 S.n8072 3.773
R3002 S.n8073 S.t439 3.773
R3003 S.n8093 S.t1306 3.773
R3004 S.n8093 S.n8092 3.773
R3005 S.n8096 S.t1531 3.773
R3006 S.n8096 S.n8095 3.773
R3007 S.n8070 S.n8069 3.773
R3008 S.n8070 S.t1256 3.773
R3009 S.n7076 S.n7075 3.773
R3010 S.n7076 S.t2370 3.773
R3011 S.n7073 S.t711 3.773
R3012 S.n7073 S.n7072 3.773
R3013 S.n7070 S.t954 3.773
R3014 S.n7070 S.n7069 3.773
R3015 S.n7067 S.n7066 3.773
R3016 S.n7067 S.t662 3.773
R3017 S.n7062 S.n7061 3.773
R3018 S.n7062 S.t1792 3.773
R3019 S.n7082 S.t131 3.773
R3020 S.n7082 S.n7081 3.773
R3021 S.n7085 S.t381 3.773
R3022 S.n7085 S.n7084 3.773
R3023 S.n7059 S.n7058 3.773
R3024 S.n7059 S.t43 3.773
R3025 S.n6329 S.n6328 3.773
R3026 S.n6329 S.t1227 3.773
R3027 S.n6326 S.t2083 3.773
R3028 S.n6326 S.n6325 3.773
R3029 S.n6323 S.t1242 3.773
R3030 S.n6323 S.n6322 3.773
R3031 S.n6320 S.n6319 3.773
R3032 S.n6320 S.t2031 3.773
R3033 S.n6315 S.n6314 3.773
R3034 S.n6315 S.t2352 3.773
R3035 S.n6335 S.t695 3.773
R3036 S.n6335 S.n6334 3.773
R3037 S.n6338 S.t938 3.773
R3038 S.n6338 S.n6337 3.773
R3039 S.n6312 S.n6311 3.773
R3040 S.n6312 S.t378 3.773
R3041 S.n5569 S.n5568 3.773
R3042 S.n5569 S.t1914 3.773
R3043 S.n5566 S.t99 3.773
R3044 S.n5566 S.n5565 3.773
R3045 S.n5563 S.t367 3.773
R3046 S.n5563 S.n5562 3.773
R3047 S.n5560 S.n5559 3.773
R3048 S.n5560 S.t14 3.773
R3049 S.n5555 S.n5554 3.773
R3050 S.n5555 S.t1956 3.773
R3051 S.n5575 S.t2192 3.773
R3052 S.n5575 S.n5574 3.773
R3053 S.n5578 S.t10 3.773
R3054 S.n5578 S.n5577 3.773
R3055 S.n5552 S.n5551 3.773
R3056 S.n5552 S.t1743 3.773
R3057 S.n4787 S.n4786 3.773
R3058 S.n4787 S.t1931 3.773
R3059 S.n4784 S.t282 3.773
R3060 S.n4784 S.n4783 3.773
R3061 S.n4781 S.t2560 3.773
R3062 S.n4781 S.n4780 3.773
R3063 S.n4778 S.n4777 3.773
R3064 S.n4778 S.t1719 3.773
R3065 S.n4773 S.n4772 3.773
R3066 S.n4773 S.t1903 3.773
R3067 S.n4793 S.t252 3.773
R3068 S.n4793 S.n4792 3.773
R3069 S.n4796 S.t2532 3.773
R3070 S.n4796 S.n4795 3.773
R3071 S.n4770 S.n4769 3.773
R3072 S.n4770 S.t1691 3.773
R3073 S.n3992 S.n3991 3.773
R3074 S.n3992 S.t1875 3.773
R3075 S.n3989 S.t219 3.773
R3076 S.n3989 S.n3988 3.773
R3077 S.n3986 S.t2510 3.773
R3078 S.n3986 S.n3985 3.773
R3079 S.n3983 S.n3982 3.773
R3080 S.n3983 S.t1664 3.773
R3081 S.n3978 S.n3977 3.773
R3082 S.n3978 S.t1851 3.773
R3083 S.n3998 S.t193 3.773
R3084 S.n3998 S.n3997 3.773
R3085 S.n4001 S.t2486 3.773
R3086 S.n4001 S.n4000 3.773
R3087 S.n3975 S.n3974 3.773
R3088 S.n3975 S.t1640 3.773
R3089 S.n3473 S.n3472 3.773
R3090 S.n3473 S.t1824 3.773
R3091 S.n3470 S.t164 3.773
R3092 S.n3470 S.n3469 3.773
R3093 S.n3467 S.t2457 3.773
R3094 S.n3467 S.n3466 3.773
R3095 S.n3464 S.n3463 3.773
R3096 S.n3464 S.t1614 3.773
R3097 S.n3459 S.n3458 3.773
R3098 S.n3459 S.t1793 3.773
R3099 S.n3479 S.t132 3.773
R3100 S.n3479 S.n3478 3.773
R3101 S.n3482 S.t201 3.773
R3102 S.n3482 S.n3481 3.773
R3103 S.n3456 S.n3455 3.773
R3104 S.n3456 S.t1582 3.773
R3105 S.n2648 S.n2647 3.773
R3106 S.n2648 S.t2060 3.773
R3107 S.n2645 S.t407 3.773
R3108 S.n2645 S.n2644 3.773
R3109 S.n2642 S.t173 3.773
R3110 S.n2642 S.n2641 3.773
R3111 S.n2336 S.n2335 3.773
R3112 S.n2336 S.t1857 3.773
R3113 S.n2659 S.t2318 3.773
R3114 S.n2661 S.t2367 3.773
R3115 S.n2663 S.t1805 3.773
R3116 S.n2624 S.n2623 3.773
R3117 S.n2624 S.t331 3.773
R3118 S.n2636 S.t1198 3.773
R3119 S.n2636 S.n2635 3.773
R3120 S.n2639 S.t2479 3.773
R3121 S.n2639 S.n2638 3.773
R3122 S.n2627 S.n2626 3.773
R3123 S.n2627 S.t1090 3.773
R3124 S.n3490 S.n3489 3.773
R3125 S.n3490 S.t2575 3.773
R3126 S.n3494 S.t929 3.773
R3127 S.n3494 S.n3493 3.773
R3128 S.n3497 S.t990 3.773
R3129 S.n3497 S.n3496 3.773
R3130 S.n3487 S.n3486 3.773
R3131 S.n3487 S.t2375 3.773
R3132 S.n11941 S.t1204 3.773
R3133 S.n11939 S.t1715 3.773
R3134 S.n11938 S.t6 3.773
R3135 S.n11835 S.n11834 3.773
R3136 S.n11835 S.t544 3.773
R3137 S.n11842 S.t2578 3.773
R3138 S.n11842 S.n11841 3.773
R3139 S.n11839 S.t1637 3.773
R3140 S.n11839 S.n11838 3.773
R3141 S.n11832 S.n11831 3.773
R3142 S.n11832 S.t1360 3.773
R3143 S.n12372 S.n12371 3.773
R3144 S.n12372 S.t2475 3.773
R3145 S.n12377 S.t822 3.773
R3146 S.n12377 S.n12376 3.773
R3147 S.n12380 S.t1069 3.773
R3148 S.n12380 S.n12379 3.773
R3149 S.n12369 S.n12368 3.773
R3150 S.n12369 S.t766 3.773
R3151 S.n12096 S.n12095 3.773
R3152 S.n12096 S.t1907 3.773
R3153 S.n12100 S.t254 3.773
R3154 S.n12100 S.n12099 3.773
R3155 S.n12103 S.t482 3.773
R3156 S.n12103 S.n12102 3.773
R3157 S.n12093 S.n12092 3.773
R3158 S.n12093 S.t197 3.773
R3159 S.n11414 S.n11413 3.773
R3160 S.n11414 S.t1319 3.773
R3161 S.n11419 S.t2188 3.773
R3162 S.n11419 S.n11418 3.773
R3163 S.n11422 S.t2410 3.773
R3164 S.n11422 S.n11421 3.773
R3165 S.n11411 S.n11410 3.773
R3166 S.n11411 S.t2135 3.773
R3167 S.n11183 S.n11182 3.773
R3168 S.n11183 S.t721 3.773
R3169 S.n11187 S.t1590 3.773
R3170 S.n11187 S.n11186 3.773
R3171 S.n11190 S.t1841 3.773
R3172 S.n11190 S.n11189 3.773
R3173 S.n11180 S.n11179 3.773
R3174 S.n11180 S.t1541 3.773
R3175 S.n10798 S.n10797 3.773
R3176 S.n10798 S.t145 3.773
R3177 S.n10803 S.t1026 3.773
R3178 S.n10803 S.n10802 3.773
R3179 S.n10806 S.t1260 3.773
R3180 S.n10806 S.n10805 3.773
R3181 S.n10795 S.n10794 3.773
R3182 S.n10795 S.t971 3.773
R3183 S.n10555 S.n10554 3.773
R3184 S.n10555 S.t2095 3.773
R3185 S.n10559 S.t441 3.773
R3186 S.n10559 S.n10558 3.773
R3187 S.n10562 S.t664 3.773
R3188 S.n10562 S.n10561 3.773
R3189 S.n10552 S.n10551 3.773
R3190 S.n10552 S.t394 3.773
R3191 S.n10148 S.n10147 3.773
R3192 S.n10148 S.t1628 3.773
R3193 S.n10153 S.t2372 3.773
R3194 S.n10153 S.n10152 3.773
R3195 S.n10156 S.t49 3.773
R3196 S.n10156 S.n10155 3.773
R3197 S.n10145 S.n10144 3.773
R3198 S.n10145 S.t2319 3.773
R3199 S.n9897 S.n9896 3.773
R3200 S.n9897 S.t840 3.773
R3201 S.n9901 S.t1708 3.773
R3202 S.n9901 S.n9900 3.773
R3203 S.n9904 S.t1954 3.773
R3204 S.n9904 S.n9903 3.773
R3205 S.n9894 S.n9893 3.773
R3206 S.n9894 S.t1873 3.773
R3207 S.n9472 S.n9471 3.773
R3208 S.n9472 S.t1600 3.773
R3209 S.n9477 S.t1143 3.773
R3210 S.n9477 S.n9476 3.773
R3211 S.n9480 S.t192 3.773
R3212 S.n9480 S.n9479 3.773
R3213 S.n9469 S.n9468 3.773
R3214 S.n9469 S.t2417 3.773
R3215 S.n9220 S.n9219 3.773
R3216 S.n9220 S.t1034 3.773
R3217 S.n9224 S.t1902 3.773
R3218 S.n9224 S.n9223 3.773
R3219 S.n9227 S.t2133 3.773
R3220 S.n9227 S.n9226 3.773
R3221 S.n9217 S.n9216 3.773
R3222 S.n9217 S.t1850 3.773
R3223 S.n8605 S.n8604 3.773
R3224 S.n8605 S.t449 3.773
R3225 S.n8610 S.t1316 3.773
R3226 S.n8610 S.n8609 3.773
R3227 S.n8613 S.t1540 3.773
R3228 S.n8613 S.n8612 3.773
R3229 S.n8602 S.n8601 3.773
R3230 S.n8602 S.t1267 3.773
R3231 S.n8816 S.n8815 3.773
R3232 S.n8816 S.t2380 3.773
R3233 S.n8820 S.t720 3.773
R3234 S.n8820 S.n8819 3.773
R3235 S.n8823 S.t966 3.773
R3236 S.n8823 S.n8822 3.773
R3237 S.n8813 S.n8812 3.773
R3238 S.n8813 S.t671 3.773
R3239 S.n7909 S.n7908 3.773
R3240 S.n7909 S.t1802 3.773
R3241 S.n7914 S.t140 3.773
R3242 S.n7914 S.n7913 3.773
R3243 S.n7917 S.t391 3.773
R3244 S.n7917 S.n7916 3.773
R3245 S.n7906 S.n7905 3.773
R3246 S.n7906 S.t64 3.773
R3247 S.n8104 S.n8103 3.773
R3248 S.n8104 S.t1232 3.773
R3249 S.n8108 S.t2093 3.773
R3250 S.n8108 S.n8107 3.773
R3251 S.n8111 S.t2317 3.773
R3252 S.n8111 S.n8110 3.773
R3253 S.n8101 S.n8100 3.773
R3254 S.n8101 S.t2044 3.773
R3255 S.n7356 S.n7355 3.773
R3256 S.n7356 S.t636 3.773
R3257 S.n7361 S.t1503 3.773
R3258 S.n7361 S.n7360 3.773
R3259 S.n7364 S.t1737 3.773
R3260 S.n7364 S.n7363 3.773
R3261 S.n7353 S.n7352 3.773
R3262 S.n7353 S.t1452 3.773
R3263 S.n7093 S.n7092 3.773
R3264 S.n7093 S.t2577 3.773
R3265 S.n7097 S.t928 3.773
R3266 S.n7097 S.n7096 3.773
R3267 S.n7100 S.t1167 3.773
R3268 S.n7100 S.n7099 3.773
R3269 S.n7090 S.n7089 3.773
R3270 S.n7090 S.t866 3.773
R3271 S.n6610 S.n6609 3.773
R3272 S.n6610 S.t2131 3.773
R3273 S.n6615 S.t357 3.773
R3274 S.n6615 S.n6614 3.773
R3275 S.n6618 S.t2027 3.773
R3276 S.n6618 S.n6617 3.773
R3277 S.n6607 S.n6606 3.773
R3278 S.n6607 S.t302 3.773
R3279 S.n6346 S.n6345 3.773
R3280 S.n6346 S.t275 3.773
R3281 S.n6350 S.t1611 3.773
R3282 S.n6350 S.n6349 3.773
R3283 S.n6353 S.t905 3.773
R3284 S.n6353 S.n6352 3.773
R3285 S.n6343 S.n6342 3.773
R3286 S.n6343 S.t921 3.773
R3287 S.n5855 S.n5854 3.773
R3288 S.n5855 S.t247 3.773
R3289 S.n5860 S.t1117 3.773
R3290 S.n5860 S.n5859 3.773
R3291 S.n5863 S.t876 3.773
R3292 S.n5863 S.n5862 3.773
R3293 S.n5852 S.n5851 3.773
R3294 S.n5852 S.t2555 3.773
R3295 S.n5586 S.n5585 3.773
R3296 S.n5586 S.t212 3.773
R3297 S.n5590 S.t1087 3.773
R3298 S.n5590 S.n5589 3.773
R3299 S.n5593 S.t853 3.773
R3300 S.n5593 S.n5592 3.773
R3301 S.n5583 S.n5582 3.773
R3302 S.n5583 S.t2526 3.773
R3303 S.n5074 S.n5073 3.773
R3304 S.n5074 S.t189 3.773
R3305 S.n5079 S.t1063 3.773
R3306 S.n5079 S.n5078 3.773
R3307 S.n5082 S.t826 3.773
R3308 S.n5082 S.n5081 3.773
R3309 S.n5071 S.n5070 3.773
R3310 S.n5071 S.t2504 3.773
R3311 S.n4804 S.n4803 3.773
R3312 S.n4804 S.t155 3.773
R3313 S.n4808 S.t1035 3.773
R3314 S.n4808 S.n4807 3.773
R3315 S.n4811 S.t795 3.773
R3316 S.n4811 S.n4810 3.773
R3317 S.n4801 S.n4800 3.773
R3318 S.n4801 S.t2478 3.773
R3319 S.n4275 S.n4274 3.773
R3320 S.n4275 S.t123 3.773
R3321 S.n4280 S.t1010 3.773
R3322 S.n4280 S.n4279 3.773
R3323 S.n4283 S.t769 3.773
R3324 S.n4283 S.n4282 3.773
R3325 S.n4272 S.n4271 3.773
R3326 S.n4272 S.t2449 3.773
R3327 S.n4009 S.n4008 3.773
R3328 S.n4009 S.t83 3.773
R3329 S.n4013 S.t981 3.773
R3330 S.n4013 S.n4012 3.773
R3331 S.n4016 S.t740 3.773
R3332 S.n4016 S.n4015 3.773
R3333 S.n4006 S.n4005 3.773
R3334 S.n4006 S.t2424 3.773
R3335 S.n3391 S.n3390 3.773
R3336 S.n3391 S.t39 3.773
R3337 S.n3395 S.t952 3.773
R3338 S.n3395 S.n3394 3.773
R3339 S.n3398 S.t715 3.773
R3340 S.n3398 S.n3397 3.773
R3341 S.n3388 S.n3387 3.773
R3342 S.n3388 S.t2400 3.773
R3343 S.n11945 S.t794 3.773
R3344 S.n11943 S.t1336 3.773
R3345 S.n11942 S.t852 3.773
R3346 S.n11816 S.n11815 3.773
R3347 S.n11816 S.t1330 3.773
R3348 S.n11827 S.t2197 3.773
R3349 S.n11827 S.n11826 3.773
R3350 S.n11824 S.t2421 3.773
R3351 S.n11824 S.n11823 3.773
R3352 S.n11819 S.n11818 3.773
R3353 S.n11819 S.t2144 3.773
R3354 S.n12385 S.n12384 3.773
R3355 S.n12385 S.t734 3.773
R3356 S.n12393 S.t1604 3.773
R3357 S.n12393 S.n12392 3.773
R3358 S.n12396 S.t1855 3.773
R3359 S.n12396 S.n12395 3.773
R3360 S.n12388 S.n12387 3.773
R3361 S.n12388 S.t1555 3.773
R3362 S.n12107 S.n12106 3.773
R3363 S.n12107 S.t158 3.773
R3364 S.n12115 S.t1039 3.773
R3365 S.n12115 S.n12114 3.773
R3366 S.n12118 S.t1268 3.773
R3367 S.n12118 S.n12117 3.773
R3368 S.n12110 S.n12109 3.773
R3369 S.n12110 S.t984 3.773
R3370 S.n11427 S.n11426 3.773
R3371 S.n11427 S.t2106 3.773
R3372 S.n11435 S.t452 3.773
R3373 S.n11435 S.n11434 3.773
R3374 S.n11438 S.t673 3.773
R3375 S.n11438 S.n11437 3.773
R3376 S.n11430 S.n11429 3.773
R3377 S.n11430 S.t403 3.773
R3378 S.n11194 S.n11193 3.773
R3379 S.n11194 S.t1514 3.773
R3380 S.n11202 S.t2381 3.773
R3381 S.n11202 S.n11201 3.773
R3382 S.n11205 S.t71 3.773
R3383 S.n11205 S.n11204 3.773
R3384 S.n11197 S.n11196 3.773
R3385 S.n11197 S.t2332 3.773
R3386 S.n10811 S.n10810 3.773
R3387 S.n10811 S.t1072 3.773
R3388 S.n10819 S.t1807 3.773
R3389 S.n10819 S.n10818 3.773
R3390 S.n10822 S.t2047 3.773
R3391 S.n10822 S.n10821 3.773
R3392 S.n10814 S.n10813 3.773
R3393 S.n10814 S.t1751 3.773
R3394 S.n10566 S.n10565 3.773
R3395 S.n10566 S.t486 3.773
R3396 S.n10574 S.t1353 3.773
R3397 S.n10574 S.n10573 3.773
R3398 S.n10577 S.t1569 3.773
R3399 S.n10577 S.n10576 3.773
R3400 S.n10569 S.n10568 3.773
R3401 S.n10569 S.t1300 3.773
R3402 S.n10161 S.n10160 3.773
R3403 S.n10161 S.t1255 3.773
R3404 S.n10169 S.t757 3.773
R3405 S.n10169 S.n10168 3.773
R3406 S.n10172 S.t2346 3.773
R3407 S.n10172 S.n10171 3.773
R3408 S.n10164 S.n10163 3.773
R3409 S.n10164 S.t2070 3.773
R3410 S.n9908 S.n9907 3.773
R3411 S.n9908 S.t462 3.773
R3412 S.n9916 S.t1328 3.773
R3413 S.n9916 S.n9915 3.773
R3414 S.n9919 S.t1550 3.773
R3415 S.n9919 S.n9918 3.773
R3416 S.n9911 S.n9910 3.773
R3417 S.n9911 S.t1478 3.773
R3418 S.n9485 S.n9484 3.773
R3419 S.n9485 S.t2388 3.773
R3420 S.n9493 S.t729 3.773
R3421 S.n9493 S.n9492 3.773
R3422 S.n9496 S.t979 3.773
R3423 S.n9496 S.n9495 3.773
R3424 S.n9488 S.n9487 3.773
R3425 S.n9488 S.t680 3.773
R3426 S.n9231 S.n9230 3.773
R3427 S.n9231 S.t1816 3.773
R3428 S.n9239 S.t153 3.773
R3429 S.n9239 S.n9238 3.773
R3430 S.n9242 S.t402 3.773
R3431 S.n9242 S.n9241 3.773
R3432 S.n9234 S.n9233 3.773
R3433 S.n9234 S.t82 3.773
R3434 S.n8618 S.n8617 3.773
R3435 S.n8618 S.t1239 3.773
R3436 S.n8626 S.t2104 3.773
R3437 S.n8626 S.n8625 3.773
R3438 S.n8629 S.t2328 3.773
R3439 S.n8629 S.n8628 3.773
R3440 S.n8621 S.n8620 3.773
R3441 S.n8621 S.t2057 3.773
R3442 S.n8827 S.n8826 3.773
R3443 S.n8827 S.t645 3.773
R3444 S.n8835 S.t1512 3.773
R3445 S.n8835 S.n8834 3.773
R3446 S.n8838 S.t1748 3.773
R3447 S.n8838 S.n8837 3.773
R3448 S.n8830 S.n8829 3.773
R3449 S.n8830 S.t1458 3.773
R3450 S.n7922 S.n7921 3.773
R3451 S.n7922 S.t12 3.773
R3452 S.n7930 S.t937 3.773
R3453 S.n7930 S.n7929 3.773
R3454 S.n7933 S.t1183 3.773
R3455 S.n7933 S.n7932 3.773
R3456 S.n7925 S.n7924 3.773
R3457 S.n7925 S.t881 3.773
R3458 S.n8115 S.n8114 3.773
R3459 S.n8115 S.t2013 3.773
R3460 S.n8123 S.t365 3.773
R3461 S.n8123 S.n8122 3.773
R3462 S.n8126 S.t583 3.773
R3463 S.n8126 S.n8125 3.773
R3464 S.n8118 S.n8117 3.773
R3465 S.n8118 S.t312 3.773
R3466 S.n7369 S.n7368 3.773
R3467 S.n7369 S.t1547 3.773
R3468 S.n7377 S.t2289 3.773
R3469 S.n7377 S.n7376 3.773
R3470 S.n7380 S.t2521 3.773
R3471 S.n7380 S.n7379 3.773
R3472 S.n7372 S.n7371 3.773
R3473 S.n7372 S.t2240 3.773
R3474 S.n7104 S.n7103 3.773
R3475 S.n7104 S.t1663 3.773
R3476 S.n7112 S.t1845 3.773
R3477 S.n7112 S.n7111 3.773
R3478 S.n7115 S.t2309 3.773
R3479 S.n7115 S.n7114 3.773
R3480 S.n7107 S.n7106 3.773
R3481 S.n7107 S.t1466 3.773
R3482 S.n6623 S.n6622 3.773
R3483 S.n6623 S.t1642 3.773
R3484 S.n6631 S.t2509 3.773
R3485 S.n6631 S.n6630 3.773
R3486 S.n6634 S.t2569 3.773
R3487 S.n6634 S.n6633 3.773
R3488 S.n6626 S.n6625 3.773
R3489 S.n6626 S.t1441 3.773
R3490 S.n6357 S.n6356 3.773
R3491 S.n6357 S.t1054 3.773
R3492 S.n6365 S.t1924 3.773
R3493 S.n6365 S.n6364 3.773
R3494 S.n6368 S.t1685 3.773
R3495 S.n6368 S.n6367 3.773
R3496 S.n6360 S.n6359 3.773
R3497 S.n6360 S.t1699 3.773
R3498 S.n5868 S.n5867 3.773
R3499 S.n5868 S.t1031 3.773
R3500 S.n5876 S.t1898 3.773
R3501 S.n5876 S.n5875 3.773
R3502 S.n5879 S.t1657 3.773
R3503 S.n5879 S.n5878 3.773
R3504 S.n5871 S.n5870 3.773
R3505 S.n5871 S.t818 3.773
R3506 S.n5597 S.n5596 3.773
R3507 S.n5597 S.t1004 3.773
R3508 S.n5605 S.t1870 3.773
R3509 S.n5605 S.n5604 3.773
R3510 S.n5608 S.t1633 3.773
R3511 S.n5608 S.n5607 3.773
R3512 S.n5600 S.n5599 3.773
R3513 S.n5600 S.t786 3.773
R3514 S.n5087 S.n5086 3.773
R3515 S.n5087 S.t977 3.773
R3516 S.n5095 S.t1848 3.773
R3517 S.n5095 S.n5094 3.773
R3518 S.n5098 S.t1608 3.773
R3519 S.n5098 S.n5097 3.773
R3520 S.n5090 S.n5089 3.773
R3521 S.n5090 S.t762 3.773
R3522 S.n4815 S.n4814 3.773
R3523 S.n4815 S.t948 3.773
R3524 S.n4823 S.t1817 3.773
R3525 S.n4823 S.n4822 3.773
R3526 S.n4826 S.t1575 3.773
R3527 S.n4826 S.n4825 3.773
R3528 S.n4818 S.n4817 3.773
R3529 S.n4818 S.t737 3.773
R3530 S.n4020 S.n4019 3.773
R3531 S.n4020 S.t925 3.773
R3532 S.n4306 S.t1790 3.773
R3533 S.n4306 S.n4305 3.773
R3534 S.n4309 S.t1557 3.773
R3535 S.n4309 S.n4308 3.773
R3536 S.n4312 S.n4311 3.773
R3537 S.n4312 S.t710 3.773
R3538 S.n4318 S.n4317 3.773
R3539 S.n4318 S.t896 3.773
R3540 S.n4326 S.t1765 3.773
R3541 S.n4326 S.n4325 3.773
R3542 S.n4329 S.t1532 3.773
R3543 S.n4329 S.n4328 3.773
R3544 S.n4321 S.n4320 3.773
R3545 S.n4321 S.t690 3.773
R3546 S.n3403 S.n3402 3.773
R3547 S.n3403 S.t967 3.773
R3548 S.n3415 S.t1734 3.773
R3549 S.n3415 S.n3414 3.773
R3550 S.n3418 S.t1561 3.773
R3551 S.n3418 S.n3417 3.773
R3552 S.n3406 S.n3405 3.773
R3553 S.n3406 S.t170 3.773
R3554 S.n3500 S.t2327 3.773
R3555 S.n3502 S.t1513 3.773
R3556 S.n3504 S.t2306 3.773
R3557 S.n4332 S.t2124 3.773
R3558 S.n4334 S.t2029 3.773
R3559 S.n4336 S.t1735 3.773
R3560 S.n4288 S.n4287 3.773
R3561 S.n4288 S.t741 3.773
R3562 S.n4300 S.t2572 3.773
R3563 S.n4300 S.n4299 3.773
R3564 S.n4303 S.t1296 3.773
R3565 S.n4303 S.n4302 3.773
R3566 S.n4291 S.n4290 3.773
R3567 S.n4291 S.t2408 3.773
R3568 S.n4834 S.n4833 3.773
R3569 S.n4834 S.t1731 3.773
R3570 S.n5132 S.t34 3.773
R3571 S.n5132 S.n5131 3.773
R3572 S.n5135 S.t2368 3.773
R3573 S.n5135 S.n5134 3.773
R3574 S.n4831 S.n4830 3.773
R3575 S.n4831 S.t1529 3.773
R3576 S.n11949 S.t1576 3.773
R3577 S.n11947 S.t2122 3.773
R3578 S.n11946 S.t469 3.773
R3579 S.n11805 S.n11804 3.773
R3580 S.n11805 S.t2117 3.773
R3581 S.n11812 S.t463 3.773
R3582 S.n11812 S.n11811 3.773
R3583 S.n11809 S.t686 3.773
R3584 S.n11809 S.n11808 3.773
R3585 S.n11802 S.n11801 3.773
R3586 S.n11802 S.t411 3.773
R3587 S.n12404 S.n12403 3.773
R3588 S.n12404 S.t1525 3.773
R3589 S.n12409 S.t2393 3.773
R3590 S.n12409 S.n12408 3.773
R3591 S.n12412 S.t86 3.773
R3592 S.n12412 S.n12411 3.773
R3593 S.n12401 S.n12400 3.773
R3594 S.n12401 S.t2343 3.773
R3595 S.n12126 S.n12125 3.773
R3596 S.n12126 S.t949 3.773
R3597 S.n12130 S.t1819 3.773
R3598 S.n12130 S.n12129 3.773
R3599 S.n12133 S.t2058 3.773
R3600 S.n12133 S.n12132 3.773
R3601 S.n12123 S.n12122 3.773
R3602 S.n12123 S.t1766 3.773
R3603 S.n11446 S.n11445 3.773
R3604 S.n11446 S.t495 3.773
R3605 S.n11451 S.t1243 3.773
R3606 S.n11451 S.n11450 3.773
R3607 S.n11454 S.t1461 3.773
R3608 S.n11454 S.n11453 3.773
R3609 S.n11443 S.n11442 3.773
R3610 S.n11443 S.t1195 3.773
R3611 S.n11213 S.n11212 3.773
R3612 S.n11213 S.t2428 3.773
R3613 S.n11217 S.t770 3.773
R3614 S.n11217 S.n11216 3.773
R3615 S.n11220 S.t1019 3.773
R3616 S.n11220 S.n11219 3.773
R3617 S.n11210 S.n11209 3.773
R3618 S.n11210 S.t714 3.773
R3619 S.n10830 S.n10829 3.773
R3620 S.n10830 S.t669 3.773
R3621 S.n10835 S.t199 3.773
R3622 S.n10835 S.n10834 3.773
R3623 S.n10838 S.t1778 3.773
R3624 S.n10838 S.n10837 3.773
R3625 S.n10827 S.n10826 3.773
R3626 S.n10827 S.t1490 3.773
R3627 S.n10585 S.n10584 3.773
R3628 S.n10585 S.t57 3.773
R3629 S.n10589 S.t963 3.773
R3630 S.n10589 S.n10588 3.773
R3631 S.n10592 S.t1210 3.773
R3632 S.n10592 S.n10591 3.773
R3633 S.n10582 S.n10581 3.773
R3634 S.n10582 S.t909 3.773
R3635 S.n10180 S.n10179 3.773
R3636 S.n10180 S.t2038 3.773
R3637 S.n10185 S.t388 3.773
R3638 S.n10185 S.n10184 3.773
R3639 S.n10188 S.t609 3.773
R3640 S.n10188 S.n10187 3.773
R3641 S.n10177 S.n10176 3.773
R3642 S.n10177 S.t339 3.773
R3643 S.n9927 S.n9926 3.773
R3644 S.n9927 S.t1247 3.773
R3645 S.n9931 S.t2114 3.773
R3646 S.n9931 S.n9930 3.773
R3647 S.n9934 S.t2338 3.773
R3648 S.n9934 S.n9933 3.773
R3649 S.n9924 S.n9923 3.773
R3650 S.n9924 S.t2262 3.773
R3651 S.n9504 S.n9503 3.773
R3652 S.n9504 S.t653 3.773
R3653 S.n9509 S.t1520 3.773
R3654 S.n9509 S.n9508 3.773
R3655 S.n9512 S.t1763 3.773
R3656 S.n9512 S.n9511 3.773
R3657 S.n9501 S.n9500 3.773
R3658 S.n9501 S.t1471 3.773
R3659 S.n9250 S.n9249 3.773
R3660 S.n9250 S.t32 3.773
R3661 S.n9254 S.t947 3.773
R3662 S.n9254 S.n9253 3.773
R3663 S.n9257 S.t1192 3.773
R3664 S.n9257 S.n9256 3.773
R3665 S.n9247 S.n9246 3.773
R3666 S.n9247 S.t894 3.773
R3667 S.n8637 S.n8636 3.773
R3668 S.n8637 S.t2023 3.773
R3669 S.n8642 S.t374 3.773
R3670 S.n8642 S.n8641 3.773
R3671 S.n8645 S.t592 3.773
R3672 S.n8645 S.n8644 3.773
R3673 S.n8634 S.n8633 3.773
R3674 S.n8634 S.t321 3.773
R3675 S.n8846 S.n8845 3.773
R3676 S.n8846 S.t1433 3.773
R3677 S.n8850 S.t2301 3.773
R3678 S.n8850 S.n8849 3.773
R3679 S.n8853 S.t2531 3.773
R3680 S.n8853 S.n8852 3.773
R3681 S.n8843 S.n8842 3.773
R3682 S.n8843 S.t2249 3.773
R3683 S.n7941 S.n7940 3.773
R3684 S.n7941 S.t986 3.773
R3685 S.n7946 S.t1718 3.773
R3686 S.n7946 S.n7945 3.773
R3687 S.n7949 S.t1966 3.773
R3688 S.n7949 S.n7948 3.773
R3689 S.n7938 S.n7937 3.773
R3690 S.n7938 S.t1662 3.773
R3691 S.n8134 S.n8133 3.773
R3692 S.n8134 S.t2505 3.773
R3693 S.n8138 S.t1272 3.773
R3694 S.n8138 S.n8137 3.773
R3695 S.n8141 S.t625 3.773
R3696 S.n8141 S.n8140 3.773
R3697 S.n8131 S.n8130 3.773
R3698 S.n8131 S.t2303 3.773
R3699 S.n7388 S.n7387 3.773
R3700 S.n7388 S.t2481 3.773
R3701 S.n7393 S.t825 3.773
R3702 S.n7393 S.n7392 3.773
R3703 S.n7396 S.t597 3.773
R3704 S.n7396 S.n7395 3.773
R3705 S.n7385 S.n7384 3.773
R3706 S.n7385 S.t2278 3.773
R3707 S.n7123 S.n7122 3.773
R3708 S.n7123 S.t2453 3.773
R3709 S.n7127 S.t797 3.773
R3710 S.n7127 S.n7126 3.773
R3711 S.n7130 S.t577 3.773
R3712 S.n7130 S.n7129 3.773
R3713 S.n7120 S.n7119 3.773
R3714 S.n7120 S.t2254 3.773
R3715 S.n6642 S.n6641 3.773
R3716 S.n6642 S.t2426 3.773
R3717 S.n6647 S.t772 3.773
R3718 S.n6647 S.n6646 3.773
R3719 S.n6650 S.t834 3.773
R3720 S.n6650 S.n6649 3.773
R3721 S.n6639 S.n6638 3.773
R3722 S.n6639 S.t2234 3.773
R3723 S.n6376 S.n6375 3.773
R3724 S.n6376 S.t1840 3.773
R3725 S.n6380 S.t181 3.773
R3726 S.n6380 S.n6379 3.773
R3727 S.n6383 S.t2471 3.773
R3728 S.n6383 S.n6382 3.773
R3729 S.n6373 S.n6372 3.773
R3730 S.n6373 S.t2488 3.773
R3731 S.n5887 S.n5886 3.773
R3732 S.n5887 S.t1810 3.773
R3733 S.n5892 S.t150 3.773
R3734 S.n5892 S.n5891 3.773
R3735 S.n5895 S.t2441 3.773
R3736 S.n5895 S.n5894 3.773
R3737 S.n5884 S.n5883 3.773
R3738 S.n5884 S.t1599 3.773
R3739 S.n5616 S.n5615 3.773
R3740 S.n5616 S.t1784 3.773
R3741 S.n5620 S.t114 3.773
R3742 S.n5620 S.n5619 3.773
R3743 S.n5623 S.t2418 3.773
R3744 S.n5623 S.n5622 3.773
R3745 S.n5613 S.n5612 3.773
R3746 S.n5613 S.t1572 3.773
R3747 S.n5127 S.n5126 3.773
R3748 S.n5127 S.t1759 3.773
R3749 S.n5124 S.t78 3.773
R3750 S.n5124 S.n5123 3.773
R3751 S.n5121 S.t2398 3.773
R3752 S.n5121 S.n5120 3.773
R3753 S.n4839 S.n4838 3.773
R3754 S.n4839 S.t1552 3.773
R3755 S.n5138 S.t1917 3.773
R3756 S.n5140 S.t1450 3.773
R3757 S.n5142 S.t1179 3.773
R3758 S.n5103 S.n5102 3.773
R3759 S.n5103 S.t542 3.773
R3760 S.n5115 S.t889 3.773
R3761 S.n5115 S.n5114 3.773
R3762 S.n5118 S.t1021 3.773
R3763 S.n5118 S.n5117 3.773
R3764 S.n5106 S.n5105 3.773
R3765 S.n5106 S.t2140 3.773
R3766 S.n5631 S.n5630 3.773
R3767 S.n5631 S.t2566 3.773
R3768 S.n5929 S.t917 3.773
R3769 S.n5929 S.n5928 3.773
R3770 S.n5932 S.t682 3.773
R3771 S.n5932 S.n5931 3.773
R3772 S.n5628 S.n5627 3.773
R3773 S.n5628 S.t2363 3.773
R3774 S.n11953 S.t2365 3.773
R3775 S.n11951 S.t389 3.773
R3776 S.n11950 S.t1258 3.773
R3777 S.n11790 S.n11789 3.773
R3778 S.n11790 S.t385 3.773
R3779 S.n11797 S.t1250 3.773
R3780 S.n11797 S.n11796 3.773
R3781 S.n11794 S.t1475 3.773
R3782 S.n11794 S.n11793 3.773
R3783 S.n11787 S.n11786 3.773
R3784 S.n11787 S.t1208 3.773
R3785 S.n12420 S.n12419 3.773
R3786 S.n12420 S.t2433 3.773
R3787 S.n12425 S.t656 3.773
R3788 S.n12425 S.n12424 3.773
R3789 S.n12428 S.t895 3.773
R3790 S.n12428 S.n12427 3.773
R3791 S.n12417 S.n12416 3.773
R3792 S.n12417 S.t605 3.773
R3793 S.n12141 S.n12140 3.773
R3794 S.n12141 S.t1862 3.773
R3795 S.n12145 S.t208 3.773
R3796 S.n12145 S.n12144 3.773
R3797 S.n12148 S.t442 3.773
R3798 S.n12148 S.n12147 3.773
R3799 S.n12138 S.n12137 3.773
R3800 S.n12138 S.t146 3.773
R3801 S.n11462 S.n11461 3.773
R3802 S.n11462 S.t75 3.773
R3803 S.n11467 S.t2149 3.773
R3804 S.n11467 S.n11466 3.773
R3805 S.n11470 S.t1222 3.773
R3806 S.n11470 S.n11469 3.773
R3807 S.n11459 S.n11458 3.773
R3808 S.n11459 S.t923 3.773
R3809 S.n11228 S.n11227 3.773
R3810 S.n11228 S.t2052 3.773
R3811 S.n11232 S.t397 3.773
R3812 S.n11232 S.n11231 3.773
R3813 S.n11235 S.t620 3.773
R3814 S.n11235 S.n11234 3.773
R3815 S.n11225 S.n11224 3.773
R3816 S.n11225 S.t352 3.773
R3817 S.n10846 S.n10845 3.773
R3818 S.n10846 S.t1456 3.773
R3819 S.n10851 S.t2325 3.773
R3820 S.n10851 S.n10850 3.773
R3821 S.n10854 S.t2559 3.773
R3822 S.n10854 S.n10853 3.773
R3823 S.n10843 S.n10842 3.773
R3824 S.n10843 S.t2272 3.773
R3825 S.n10600 S.n10599 3.773
R3826 S.n10600 S.t875 3.773
R3827 S.n10604 S.t1744 3.773
R3828 S.n10604 S.n10603 3.773
R3829 S.n10607 S.t1987 3.773
R3830 S.n10607 S.n10606 3.773
R3831 S.n10597 S.n10596 3.773
R3832 S.n10597 S.t1690 3.773
R3833 S.n10196 S.n10195 3.773
R3834 S.n10196 S.t307 3.773
R3835 S.n10201 S.t1176 3.773
R3836 S.n10201 S.n10200 3.773
R3837 S.n10204 S.t1399 3.773
R3838 S.n10204 S.n10203 3.773
R3839 S.n10193 S.n10192 3.773
R3840 S.n10193 S.t1125 3.773
R3841 S.n9942 S.n9941 3.773
R3842 S.n9942 S.t2033 3.773
R3843 S.n9946 S.t382 3.773
R3844 S.n9946 S.n9945 3.773
R3845 S.n9949 S.t603 3.773
R3846 S.n9949 S.n9948 3.773
R3847 S.n9939 S.n9938 3.773
R3848 S.n9939 S.t535 3.773
R3849 S.n9520 S.n9519 3.773
R3850 S.n9520 S.t1443 3.773
R3851 S.n9525 S.t2311 3.773
R3852 S.n9525 S.n9524 3.773
R3853 S.n9528 S.t2543 3.773
R3854 S.n9528 S.n9527 3.773
R3855 S.n9517 S.n9516 3.773
R3856 S.n9517 S.t2260 3.773
R3857 S.n9265 S.n9264 3.773
R3858 S.n9265 S.t863 3.773
R3859 S.n9269 S.t1730 3.773
R3860 S.n9269 S.n9268 3.773
R3861 S.n9272 S.t1972 3.773
R3862 S.n9272 S.n9271 3.773
R3863 S.n9262 S.n9261 3.773
R3864 S.n9262 S.t1675 3.773
R3865 S.n8653 S.n8652 3.773
R3866 S.n8653 S.t416 3.773
R3867 S.n8658 S.t1162 3.773
R3868 S.n8658 S.n8657 3.773
R3869 S.n8661 S.t1386 3.773
R3870 S.n8661 S.n8660 3.773
R3871 S.n8650 S.n8649 3.773
R3872 S.n8650 S.t1111 3.773
R3873 S.n8861 S.n8860 3.773
R3874 S.n8861 S.t820 3.773
R3875 S.n8865 S.t689 3.773
R3876 S.n8865 S.n8864 3.773
R3877 S.n8868 S.t1460 3.773
R3878 S.n8868 S.n8867 3.773
R3879 S.n8858 S.n8857 3.773
R3880 S.n8858 S.t621 3.773
R3881 S.n7957 S.n7956 3.773
R3882 S.n7957 S.t790 3.773
R3883 S.n7962 S.t1658 3.773
R3884 S.n7962 S.n7961 3.773
R3885 S.n7965 S.t1435 3.773
R3886 S.n7965 S.n7964 3.773
R3887 S.n7954 S.n7953 3.773
R3888 S.n7954 S.t594 3.773
R3889 S.n8149 S.n8148 3.773
R3890 S.n8149 S.t763 3.773
R3891 S.n8153 S.t1634 3.773
R3892 S.n8153 S.n8152 3.773
R3893 S.n8156 S.t1414 3.773
R3894 S.n8156 S.n8155 3.773
R3895 S.n8146 S.n8145 3.773
R3896 S.n8146 S.t573 3.773
R3897 S.n7404 S.n7403 3.773
R3898 S.n7404 S.t738 3.773
R3899 S.n7409 S.t1609 3.773
R3900 S.n7409 S.n7408 3.773
R3901 S.n7412 S.t1390 3.773
R3902 S.n7412 S.n7411 3.773
R3903 S.n7401 S.n7400 3.773
R3904 S.n7401 S.t549 3.773
R3905 S.n7138 S.n7137 3.773
R3906 S.n7138 S.t709 3.773
R3907 S.n7142 S.t1579 3.773
R3908 S.n7142 S.n7141 3.773
R3909 S.n7145 S.t1368 3.773
R3910 S.n7145 S.n7144 3.773
R3911 S.n7135 S.n7134 3.773
R3912 S.n7135 S.t524 3.773
R3913 S.n6658 S.n6657 3.773
R3914 S.n6658 S.t691 3.773
R3915 S.n6663 S.t1559 3.773
R3916 S.n6663 S.n6662 3.773
R3917 S.n6666 S.t1616 3.773
R3918 S.n6666 S.n6665 3.773
R3919 S.n6655 S.n6654 3.773
R3920 S.n6655 S.t501 3.773
R3921 S.n6391 S.n6390 3.773
R3922 S.n6391 S.t70 3.773
R3923 S.n6395 S.t970 3.773
R3924 S.n6395 S.n6394 3.773
R3925 S.n6398 S.t732 3.773
R3926 S.n6398 S.n6397 3.773
R3927 S.n6388 S.n6387 3.773
R3928 S.n6388 S.t743 3.773
R3929 S.n5924 S.n5923 3.773
R3930 S.n5924 S.t26 3.773
R3931 S.n5921 S.t943 3.773
R3932 S.n5921 S.n5920 3.773
R3933 S.n5918 S.t704 3.773
R3934 S.n5918 S.n5917 3.773
R3935 S.n5636 S.n5635 3.773
R3936 S.n5636 S.t2391 3.773
R3937 S.n5935 S.t1688 3.773
R3938 S.n5937 S.t878 3.773
R3939 S.n5939 S.t591 3.773
R3940 S.n5900 S.n5899 3.773
R3941 S.n5900 S.t338 3.773
R3942 S.n5912 S.t1725 3.773
R3943 S.n5912 S.n5911 3.773
R3944 S.n5915 S.t727 3.773
R3945 S.n5915 S.n5914 3.773
R3946 S.n5903 S.n5902 3.773
R3947 S.n5903 S.t1863 3.773
R3948 S.n6406 S.n6405 3.773
R3949 S.n6406 S.t885 3.773
R3950 S.n6700 S.t1753 3.773
R3951 S.n6700 S.n6699 3.773
R3952 S.n6703 S.t1521 3.773
R3953 S.n6703 S.n6702 3.773
R3954 S.n6403 S.n6402 3.773
R3955 S.n6403 S.t1535 3.773
R3956 S.n11957 S.t633 3.773
R3957 S.n11955 S.t1181 3.773
R3958 S.n11954 S.t2042 3.773
R3959 S.n11775 S.n11774 3.773
R3960 S.n11775 S.t1291 3.773
R3961 S.n11782 S.t2159 3.773
R3962 S.n11782 S.n11781 3.773
R3963 S.n11779 S.t2383 3.773
R3964 S.n11779 S.n11778 3.773
R3965 S.n11772 S.n11771 3.773
R3966 S.n11772 S.t2109 3.773
R3967 S.n12436 S.n12435 3.773
R3968 S.n12436 S.t2061 3.773
R3969 S.n12441 S.t1564 3.773
R3970 S.n12441 S.n12440 3.773
R3971 S.n12444 S.t628 3.773
R3972 S.n12444 S.n12443 3.773
R3973 S.n12433 S.n12432 3.773
R3974 S.n12433 S.t359 3.773
R3975 S.n12156 S.n12155 3.773
R3976 S.n12156 S.t1467 3.773
R3977 S.n12160 S.t2334 3.773
R3978 S.n12160 S.n12159 3.773
R3979 S.n12163 S.t2570 3.773
R3980 S.n12163 S.n12162 3.773
R3981 S.n12153 S.n12152 3.773
R3982 S.n12153 S.t2282 3.773
R3983 S.n11478 S.n11477 3.773
R3984 S.n11478 S.t888 3.773
R3985 S.n11483 S.t1758 3.773
R3986 S.n11483 S.n11482 3.773
R3987 S.n11486 S.t1998 3.773
R3988 S.n11486 S.n11485 3.773
R3989 S.n11475 S.n11474 3.773
R3990 S.n11475 S.t1700 3.773
R3991 S.n11243 S.n11242 3.773
R3992 S.n11243 S.t317 3.773
R3993 S.n11247 S.t1188 3.773
R3994 S.n11247 S.n11246 3.773
R3995 S.n11250 S.t1410 3.773
R3996 S.n11250 S.n11249 3.773
R3997 S.n11240 S.n11239 3.773
R3998 S.n11240 S.t1137 3.773
R3999 S.n10862 S.n10861 3.773
R4000 S.n10862 S.t2244 3.773
R4001 S.n10867 S.t589 3.773
R4002 S.n10867 S.n10866 3.773
R4003 S.n10870 S.t823 3.773
R4004 S.n10870 S.n10869 3.773
R4005 S.n10859 S.n10858 3.773
R4006 S.n10859 S.t545 3.773
R4007 S.n10615 S.n10614 3.773
R4008 S.n10615 S.t1656 3.773
R4009 S.n10619 S.t2525 3.773
R4010 S.n10619 S.n10618 3.773
R4011 S.n10622 S.t255 3.773
R4012 S.n10622 S.n10621 3.773
R4013 S.n10612 S.n10611 3.773
R4014 S.n10612 S.t2476 3.773
R4015 S.n10212 S.n10211 3.773
R4016 S.n10212 S.t1093 3.773
R4017 S.n10217 S.t1961 3.773
R4018 S.n10217 S.n10216 3.773
R4019 S.n10220 S.t2189 3.773
R4020 S.n10220 S.n10219 3.773
R4021 S.n10209 S.n10208 3.773
R4022 S.n10209 S.t1909 3.773
R4023 S.n9957 S.n9956 3.773
R4024 S.n9957 S.t303 3.773
R4025 S.n9961 S.t1170 3.773
R4026 S.n9961 S.n9960 3.773
R4027 S.n9964 S.t1395 3.773
R4028 S.n9964 S.n9963 3.773
R4029 S.n9954 S.n9953 3.773
R4030 S.n9954 S.t1320 3.773
R4031 S.n9536 S.n9535 3.773
R4032 S.n9536 S.t2354 3.773
R4033 S.n9541 S.t579 3.773
R4034 S.n9541 S.n9540 3.773
R4035 S.n9544 S.t810 3.773
R4036 S.n9544 S.n9543 3.773
R4037 S.n9533 S.n9532 3.773
R4038 S.n9533 S.t529 3.773
R4039 S.n9280 S.n9279 3.773
R4040 S.n9280 S.t1654 3.773
R4041 S.n9284 S.t101 3.773
R4042 S.n9284 S.n9283 3.773
R4043 S.n9287 S.t2300 3.773
R4044 S.n9287 S.n9286 3.773
R4045 S.n9277 S.n9276 3.773
R4046 S.n9277 S.t1455 3.773
R4047 S.n8669 S.n8668 3.773
R4048 S.n8669 S.t1629 3.773
R4049 S.n8674 S.t2500 3.773
R4050 S.n8674 S.n8673 3.773
R4051 S.n8677 S.t2274 3.773
R4052 S.n8677 S.n8676 3.773
R4053 S.n8666 S.n8665 3.773
R4054 S.n8666 S.t1432 3.773
R4055 S.n8876 S.n8875 3.773
R4056 S.n8876 S.t1602 3.773
R4057 S.n8880 S.t2473 3.773
R4058 S.n8880 S.n8879 3.773
R4059 S.n8883 S.t2250 3.773
R4060 S.n8883 S.n8882 3.773
R4061 S.n8873 S.n8872 3.773
R4062 S.n8873 S.t1411 3.773
R4063 S.n7973 S.n7972 3.773
R4064 S.n7973 S.t1571 3.773
R4065 S.n7978 S.t2446 3.773
R4066 S.n7978 S.n7977 3.773
R4067 S.n7981 S.t2227 3.773
R4068 S.n7981 S.n7980 3.773
R4069 S.n7970 S.n7969 3.773
R4070 S.n7970 S.t1387 3.773
R4071 S.n8164 S.n8163 3.773
R4072 S.n8164 S.t1551 3.773
R4073 S.n8168 S.t2419 3.773
R4074 S.n8168 S.n8167 3.773
R4075 S.n8171 S.t2204 3.773
R4076 S.n8171 S.n8170 3.773
R4077 S.n8161 S.n8160 3.773
R4078 S.n8161 S.t1362 3.773
R4079 S.n7420 S.n7419 3.773
R4080 S.n7420 S.t1530 3.773
R4081 S.n7425 S.t2397 3.773
R4082 S.n7425 S.n7424 3.773
R4083 S.n7428 S.t2179 3.773
R4084 S.n7428 S.n7427 3.773
R4085 S.n7417 S.n7416 3.773
R4086 S.n7417 S.t1339 3.773
R4087 S.n7153 S.n7152 3.773
R4088 S.n7153 S.t1504 3.773
R4089 S.n7157 S.t2369 3.773
R4090 S.n7157 S.n7156 3.773
R4091 S.n7160 S.t2153 3.773
R4092 S.n7160 S.n7159 3.773
R4093 S.n7150 S.n7149 3.773
R4094 S.n7150 S.t1309 3.773
R4095 S.n6695 S.n6694 3.773
R4096 S.n6695 S.t1480 3.773
R4097 S.n6692 S.t2347 3.773
R4098 S.n6692 S.n6691 3.773
R4099 S.n6689 S.t2403 3.773
R4100 S.n6689 S.n6688 3.773
R4101 S.n6411 S.n6410 3.773
R4102 S.n6411 S.t1285 3.773
R4103 S.n6706 S.t1479 3.773
R4104 S.n6708 S.t319 3.773
R4105 S.n6710 S.t2258 3.773
R4106 S.n6671 S.n6670 3.773
R4107 S.n6671 S.t351 3.773
R4108 S.n6683 S.t611 3.773
R4109 S.n6683 S.n6682 3.773
R4110 S.n6686 S.t1128 3.773
R4111 S.n6686 S.n6685 3.773
R4112 S.n6674 S.n6673 3.773
R4113 S.n6674 S.t1591 3.773
R4114 S.n7168 S.n7167 3.773
R4115 S.n7168 S.t2290 3.773
R4116 S.n7462 S.t637 3.773
R4117 S.n7462 S.n7461 3.773
R4118 S.n7465 S.t420 3.773
R4119 S.n7465 S.n7464 3.773
R4120 S.n7165 S.n7164 3.773
R4121 S.n7165 S.t2096 3.773
R4122 S.n11961 S.t1543 3.773
R4123 S.n11959 S.t2085 3.773
R4124 S.n11958 S.t432 3.773
R4125 S.n11760 S.n11759 3.773
R4126 S.n11760 S.t899 3.773
R4127 S.n11767 S.t1768 3.773
R4128 S.n11767 S.n11766 3.773
R4129 S.n11764 S.t2005 3.773
R4130 S.n11764 S.n11763 3.773
R4131 S.n11757 S.n11756 3.773
R4132 S.n11757 S.t1709 3.773
R4133 S.n12452 S.n12451 3.773
R4134 S.n12452 S.t326 3.773
R4135 S.n12457 S.t1199 3.773
R4136 S.n12457 S.n12456 3.773
R4137 S.n12460 S.t1418 3.773
R4138 S.n12460 S.n12459 3.773
R4139 S.n12449 S.n12448 3.773
R4140 S.n12449 S.t1145 3.773
R4141 S.n12171 S.n12170 3.773
R4142 S.n12171 S.t2255 3.773
R4143 S.n12175 S.t598 3.773
R4144 S.n12175 S.n12174 3.773
R4145 S.n12178 S.t835 3.773
R4146 S.n12178 S.n12177 3.773
R4147 S.n12168 S.n12167 3.773
R4148 S.n12168 S.t554 3.773
R4149 S.n11494 S.n11493 3.773
R4150 S.n11494 S.t1670 3.773
R4151 S.n11499 S.t2539 3.773
R4152 S.n11499 S.n11498 3.773
R4153 S.n11502 S.t270 3.773
R4154 S.n11502 S.n11501 3.773
R4155 S.n11491 S.n11490 3.773
R4156 S.n11491 S.t2489 3.773
R4157 S.n11258 S.n11257 3.773
R4158 S.n11258 S.t1107 3.773
R4159 S.n11262 S.t1970 3.773
R4160 S.n11262 S.n11261 3.773
R4161 S.n11265 S.t2198 3.773
R4162 S.n11265 S.n11264 3.773
R4163 S.n11255 S.n11254 3.773
R4164 S.n11255 S.t1921 3.773
R4165 S.n10878 S.n10877 3.773
R4166 S.n10878 S.t513 3.773
R4167 S.n10883 S.t1380 3.773
R4168 S.n10883 S.n10882 3.773
R4169 S.n10886 S.t1605 3.773
R4170 S.n10886 S.n10885 3.773
R4171 S.n10875 S.n10874 3.773
R4172 S.n10875 S.t1331 3.773
R4173 S.n10630 S.n10629 3.773
R4174 S.n10630 S.t2445 3.773
R4175 S.n10634 S.t789 3.773
R4176 S.n10634 S.n10633 3.773
R4177 S.n10637 S.t1040 3.773
R4178 S.n10637 S.n10636 3.773
R4179 S.n10627 S.n10626 3.773
R4180 S.n10627 S.t736 3.773
R4181 S.n10228 S.n10227 3.773
R4182 S.n10228 S.t2001 3.773
R4183 S.n10233 S.t218 3.773
R4184 S.n10233 S.n10232 3.773
R4185 S.n10236 S.t455 3.773
R4186 S.n10236 S.n10235 3.773
R4187 S.n10225 S.n10224 3.773
R4188 S.n10225 S.t162 3.773
R4189 S.n9972 S.n9971 3.773
R4190 S.n9972 S.t2494 3.773
R4191 S.n9976 S.t2078 3.773
R4192 S.n9976 S.n9975 3.773
R4193 S.n9979 S.t617 3.773
R4194 S.n9979 S.n9978 3.773
R4195 S.n9969 S.n9968 3.773
R4196 S.n9969 S.t149 3.773
R4197 S.n9552 S.n9551 3.773
R4198 S.n9552 S.t2468 3.773
R4199 S.n9557 S.t814 3.773
R4200 S.n9557 S.n9556 3.773
R4201 S.n9560 S.t588 3.773
R4202 S.n9560 S.n9559 3.773
R4203 S.n9549 S.n9548 3.773
R4204 S.n9549 S.t2269 3.773
R4205 S.n9295 S.n9294 3.773
R4206 S.n9295 S.t2436 3.773
R4207 S.n9299 S.t784 3.773
R4208 S.n9299 S.n9298 3.773
R4209 S.n9302 S.t570 3.773
R4210 S.n9302 S.n9301 3.773
R4211 S.n9292 S.n9291 3.773
R4212 S.n9292 S.t2245 3.773
R4213 S.n8685 S.n8684 3.773
R4214 S.n8685 S.t2415 3.773
R4215 S.n8690 S.t758 3.773
R4216 S.n8690 S.n8689 3.773
R4217 S.n8693 S.t546 3.773
R4218 S.n8693 S.n8692 3.773
R4219 S.n8682 S.n8681 3.773
R4220 S.n8682 S.t2223 3.773
R4221 S.n8891 S.n8890 3.773
R4222 S.n8891 S.t2390 3.773
R4223 S.n8895 S.t731 3.773
R4224 S.n8895 S.n8894 3.773
R4225 S.n8898 S.t518 3.773
R4226 S.n8898 S.n8897 3.773
R4227 S.n8888 S.n8887 3.773
R4228 S.n8888 S.t2200 3.773
R4229 S.n7989 S.n7988 3.773
R4230 S.n7989 S.t2364 3.773
R4231 S.n7994 S.t703 3.773
R4232 S.n7994 S.n7993 3.773
R4233 S.n7997 S.t494 3.773
R4234 S.n7997 S.n7996 3.773
R4235 S.n7986 S.n7985 3.773
R4236 S.n7986 S.t2172 3.773
R4237 S.n8179 S.n8178 3.773
R4238 S.n8179 S.t2341 3.773
R4239 S.n8183 S.t683 3.773
R4240 S.n8183 S.n8182 3.773
R4241 S.n8186 S.t471 3.773
R4242 S.n8186 S.n8185 3.773
R4243 S.n8176 S.n8175 3.773
R4244 S.n8176 S.t2148 3.773
R4245 S.n7457 S.n7456 3.773
R4246 S.n7457 S.t2315 3.773
R4247 S.n7454 S.t660 3.773
R4248 S.n7454 S.n7453 3.773
R4249 S.n7451 S.t443 3.773
R4250 S.n7451 S.n7450 3.773
R4251 S.n7173 S.n7172 3.773
R4252 S.n7173 S.t2125 3.773
R4253 S.n7468 S.t1488 3.773
R4254 S.n7470 S.t536 3.773
R4255 S.n7472 S.t258 3.773
R4256 S.n7433 S.n7432 3.773
R4257 S.n7433 S.t103 3.773
R4258 S.n7445 S.t1449 3.773
R4259 S.n7445 S.n7444 3.773
R4260 S.n7448 S.t206 3.773
R4261 S.n7448 S.n7447 3.773
R4262 S.n7436 S.n7435 3.773
R4263 S.n7436 S.t1329 3.773
R4264 S.n8194 S.n8193 3.773
R4265 S.n8194 S.t606 3.773
R4266 S.n8198 S.t1474 3.773
R4267 S.n8198 S.n8197 3.773
R4268 S.n8201 S.t1257 3.773
R4269 S.n8201 S.n8200 3.773
R4270 S.n8191 S.n8190 3.773
R4271 S.n8191 S.t417 3.773
R4272 S.n11965 S.t1173 3.773
R4273 S.n11963 S.t1686 3.773
R4274 S.n11962 S.t2554 3.773
R4275 S.n11745 S.n11744 3.773
R4276 S.n11745 S.t1679 3.773
R4277 S.n11752 S.t2546 3.773
R4278 S.n11752 S.n11751 3.773
R4279 S.n11749 S.t278 3.773
R4280 S.n11749 S.n11748 3.773
R4281 S.n11742 S.n11741 3.773
R4282 S.n11742 S.t2496 3.773
R4283 S.n12468 S.n12467 3.773
R4284 S.n12468 S.t1115 3.773
R4285 S.n12473 S.t1979 3.773
R4286 S.n12473 S.n12472 3.773
R4287 S.n12476 S.t2207 3.773
R4288 S.n12476 S.n12475 3.773
R4289 S.n12465 S.n12464 3.773
R4290 S.n12465 S.t1927 3.773
R4291 S.n12186 S.n12185 3.773
R4292 S.n12186 S.t523 3.773
R4293 S.n12190 S.t1391 3.773
R4294 S.n12190 S.n12189 3.773
R4295 S.n12193 S.t1618 3.773
R4296 S.n12193 S.n12192 3.773
R4297 S.n12183 S.n12182 3.773
R4298 S.n12183 S.t1342 3.773
R4299 S.n11510 S.n11509 3.773
R4300 S.n11510 S.t2458 3.773
R4301 S.n11515 S.t804 3.773
R4302 S.n11515 S.n11514 3.773
R4303 S.n11518 S.t1049 3.773
R4304 S.n11518 S.n11517 3.773
R4305 S.n11507 S.n11506 3.773
R4306 S.n11507 S.t745 3.773
R4307 S.n11273 S.n11272 3.773
R4308 S.n11273 S.t1886 3.773
R4309 S.n11277 S.t232 3.773
R4310 S.n11277 S.n11276 3.773
R4311 S.n11280 S.t464 3.773
R4312 S.n11280 S.n11279 3.773
R4313 S.n11270 S.n11269 3.773
R4314 S.n11270 S.t174 3.773
R4315 S.n10894 S.n10893 3.773
R4316 S.n10894 S.t1423 3.773
R4317 S.n10899 S.t2166 3.773
R4318 S.n10899 S.n10898 3.773
R4319 S.n10902 S.t2395 3.773
R4320 S.n10902 S.n10901 3.773
R4321 S.n10891 S.n10890 3.773
R4322 S.n10891 S.t2120 3.773
R4323 S.n10645 S.n10644 3.773
R4324 S.n10645 S.t1209 3.773
R4325 S.n10649 S.t1705 3.773
R4326 S.n10649 S.n10648 3.773
R4327 S.n10652 S.t1839 3.773
R4328 S.n10652 S.n10651 3.773
R4329 S.n10642 S.n10641 3.773
R4330 S.n10642 S.t998 3.773
R4331 S.n10244 S.n10243 3.773
R4332 S.n10244 S.t1178 3.773
R4333 S.n10249 S.t2041 3.773
R4334 S.n10249 S.n10248 3.773
R4335 S.n10252 S.t1809 3.773
R4336 S.n10252 S.n10251 3.773
R4337 S.n10241 S.n10240 3.773
R4338 S.n10241 S.t969 3.773
R4339 S.n9987 S.n9986 3.773
R4340 S.n9987 S.t750 3.773
R4341 S.n9991 S.t1622 3.773
R4342 S.n9991 S.n9990 3.773
R4343 S.n9994 S.t1408 3.773
R4344 S.n9994 S.n9993 3.773
R4345 S.n9984 S.n9983 3.773
R4346 S.n9984 S.t942 3.773
R4347 S.n9568 S.n9567 3.773
R4348 S.n9568 S.t726 3.773
R4349 S.n9573 S.t1595 3.773
R4350 S.n9573 S.n9572 3.773
R4351 S.n9576 S.t1381 3.773
R4352 S.n9576 S.n9575 3.773
R4353 S.n9565 S.n9564 3.773
R4354 S.n9565 S.t541 3.773
R4355 S.n9310 S.n9309 3.773
R4356 S.n9310 S.t701 3.773
R4357 S.n9314 S.t1566 3.773
R4358 S.n9314 S.n9313 3.773
R4359 S.n9317 S.t1357 3.773
R4360 S.n9317 S.n9316 3.773
R4361 S.n9307 S.n9306 3.773
R4362 S.n9307 S.t514 3.773
R4363 S.n8701 S.n8700 3.773
R4364 S.n8701 S.t679 3.773
R4365 S.n8706 S.t1548 3.773
R4366 S.n8706 S.n8705 3.773
R4367 S.n8709 S.t1334 3.773
R4368 S.n8709 S.n8708 3.773
R4369 S.n8698 S.n8697 3.773
R4370 S.n8698 S.t489 3.773
R4371 S.n8906 S.n8905 3.773
R4372 S.n8906 S.t654 3.773
R4373 S.n8910 S.t1524 3.773
R4374 S.n8910 S.n8909 3.773
R4375 S.n8913 S.t1304 3.773
R4376 S.n8913 S.n8912 3.773
R4377 S.n8903 S.n8902 3.773
R4378 S.n8903 S.t467 3.773
R4379 S.n8005 S.n8004 3.773
R4380 S.n8005 S.t632 3.773
R4381 S.n8009 S.t1499 3.773
R4382 S.n8009 S.n8008 3.773
R4383 S.n8012 S.t1283 3.773
R4384 S.n8012 S.n8011 3.773
R4385 S.n8002 S.n8001 3.773
R4386 S.n8002 S.t437 3.773
R4387 S.n8204 S.t1282 3.773
R4388 S.n8206 S.t2480 3.773
R4389 S.n8208 S.t2201 3.773
R4390 S.n8017 S.n8016 3.773
R4391 S.n8017 S.t2427 3.773
R4392 S.n8029 S.t2285 3.773
R4393 S.n8029 S.n8028 3.773
R4394 S.n8032 S.t2437 3.773
R4395 S.n8032 S.n8031 3.773
R4396 S.n8020 S.n8019 3.773
R4397 S.n8020 S.t1055 3.773
R4398 S.n8921 S.n8920 3.773
R4399 S.n8921 S.t1444 3.773
R4400 S.n8925 S.t2312 3.773
R4401 S.n8925 S.n8924 3.773
R4402 S.n8928 S.t2091 3.773
R4403 S.n8928 S.n8927 3.773
R4404 S.n8918 S.n8917 3.773
R4405 S.n8918 S.t1254 3.773
R4406 S.n11969 S.t1955 3.773
R4407 S.n11967 S.t2472 3.773
R4408 S.n11966 S.t819 3.773
R4409 S.n11730 S.n11729 3.773
R4410 S.n11730 S.t2465 3.773
R4411 S.n11737 S.t812 3.773
R4412 S.n11737 S.n11736 3.773
R4413 S.n11734 S.t1058 3.773
R4414 S.n11734 S.n11733 3.773
R4415 S.n11727 S.n11726 3.773
R4416 S.n11727 S.t752 3.773
R4417 S.n12484 S.n12483 3.773
R4418 S.n12484 S.t1897 3.773
R4419 S.n12489 S.t243 3.773
R4420 S.n12489 S.n12488 3.773
R4421 S.n12492 S.t474 3.773
R4422 S.n12492 S.n12491 3.773
R4423 S.n12481 S.n12480 3.773
R4424 S.n12481 S.t183 3.773
R4425 S.n12201 S.n12200 3.773
R4426 S.n12201 S.t1311 3.773
R4427 S.n12205 S.t2181 3.773
R4428 S.n12205 S.n12204 3.773
R4429 S.n12208 S.t2404 3.773
R4430 S.n12208 S.n12207 3.773
R4431 S.n12198 S.n12197 3.773
R4432 S.n12198 S.t2129 3.773
R4433 S.n11526 S.n11525 3.773
R4434 S.n11526 S.t851 3.773
R4435 S.n11531 S.t1583 3.773
R4436 S.n11531 S.n11530 3.773
R4437 S.n11534 S.t1833 3.773
R4438 S.n11534 S.n11533 3.773
R4439 S.n11523 S.n11522 3.773
R4440 S.n11523 S.t1538 3.773
R4441 S.n11288 S.n11287 3.773
R4442 S.n11288 S.t2037 3.773
R4443 S.n11292 S.t1152 3.773
R4444 S.n11292 S.n11291 3.773
R4445 S.n11295 S.t142 3.773
R4446 S.n11295 S.n11294 3.773
R4447 S.n11285 S.n11284 3.773
R4448 S.n11285 S.t1836 3.773
R4449 S.n10910 S.n10909 3.773
R4450 S.n10910 S.t2009 3.773
R4451 S.n10915 S.t363 3.773
R4452 S.n10915 S.n10914 3.773
R4453 S.n10918 S.t105 3.773
R4454 S.n10918 S.n10917 3.773
R4455 S.n10907 S.n10906 3.773
R4456 S.n10907 S.t1804 3.773
R4457 S.n10660 S.n10659 3.773
R4458 S.n10660 S.t1986 3.773
R4459 S.n10664 S.t337 3.773
R4460 S.n10664 S.n10663 3.773
R4461 S.n10667 S.t68 3.773
R4462 S.n10667 S.n10666 3.773
R4463 S.n10657 S.n10656 3.773
R4464 S.n10657 S.t1781 3.773
R4465 S.n10260 S.n10259 3.773
R4466 S.n10260 S.t1964 3.773
R4467 S.n10265 S.t309 3.773
R4468 S.n10265 S.n10264 3.773
R4469 S.n10268 S.t24 3.773
R4470 S.n10268 S.n10267 3.773
R4471 S.n10257 S.n10256 3.773
R4472 S.n10257 S.t1752 3.773
R4473 S.n10002 S.n10001 3.773
R4474 S.n10002 S.t1544 3.773
R4475 S.n10006 S.t2409 3.773
R4476 S.n10006 S.n10005 3.773
R4477 S.n10009 S.t2196 3.773
R4478 S.n10009 S.n10008 3.773
R4479 S.n9999 S.n9998 3.773
R4480 S.n9999 S.t1724 3.773
R4481 S.n9584 S.n9583 3.773
R4482 S.n9584 S.t1517 3.773
R4483 S.n9589 S.t2386 3.773
R4484 S.n9589 S.n9588 3.773
R4485 S.n9592 S.t2167 3.773
R4486 S.n9592 S.n9591 3.773
R4487 S.n9581 S.n9580 3.773
R4488 S.n9581 S.t1327 3.773
R4489 S.n9325 S.n9324 3.773
R4490 S.n9325 S.t1496 3.773
R4491 S.n9329 S.t2359 3.773
R4492 S.n9329 S.n9328 3.773
R4493 S.n9332 S.t2142 3.773
R4494 S.n9332 S.n9331 3.773
R4495 S.n9322 S.n9321 3.773
R4496 S.n9322 S.t1301 3.773
R4497 S.n8717 S.n8716 3.773
R4498 S.n8717 S.t1469 3.773
R4499 S.n8721 S.t2336 3.773
R4500 S.n8721 S.n8720 3.773
R4501 S.n8724 S.t2121 3.773
R4502 S.n8724 S.n8723 3.773
R4503 S.n8714 S.n8713 3.773
R4504 S.n8714 S.t1275 3.773
R4505 S.n8931 S.t1073 3.773
R4506 S.n8933 S.t1922 3.773
R4507 S.n8935 S.t1620 3.773
R4508 S.n8729 S.n8728 3.773
R4509 S.n8729 S.t2220 3.773
R4510 S.n8741 S.t599 3.773
R4511 S.n8741 S.n8740 3.773
R4512 S.n8744 S.t2171 3.773
R4513 S.n8744 S.n8743 3.773
R4514 S.n8732 S.n8731 3.773
R4515 S.n8732 S.t760 3.773
R4516 S.n9340 S.n9339 3.773
R4517 S.n9340 S.t2280 3.773
R4518 S.n9626 S.t626 3.773
R4519 S.n9626 S.n9625 3.773
R4520 S.n9629 S.t410 3.773
R4521 S.n9629 S.n9628 3.773
R4522 S.n9337 S.n9336 3.773
R4523 S.n9337 S.t2090 3.773
R4524 S.n11973 S.t215 3.773
R4525 S.n11971 S.t730 3.773
R4526 S.n11970 S.t1601 3.773
R4527 S.n11715 S.n11714 3.773
R4528 S.n11715 S.t724 3.773
R4529 S.n11722 S.t1594 3.773
R4530 S.n11722 S.n11721 3.773
R4531 S.n11719 S.t1843 3.773
R4532 S.n11719 S.n11718 3.773
R4533 S.n11712 S.n11711 3.773
R4534 S.n11712 S.t1545 3.773
R4535 S.n12500 S.n12499 3.773
R4536 S.n12500 S.t292 3.773
R4537 S.n12505 S.t1030 3.773
R4538 S.n12505 S.n12504 3.773
R4539 S.n12508 S.t1263 3.773
R4540 S.n12508 S.n12507 3.773
R4541 S.n12497 S.n12496 3.773
R4542 S.n12497 S.t974 3.773
R4543 S.n12216 S.n12215 3.773
R4544 S.n12216 S.t358 3.773
R4545 S.n12220 S.t566 3.773
R4546 S.n12220 S.n12219 3.773
R4547 S.n12223 S.t993 3.773
R4548 S.n12223 S.n12222 3.773
R4549 S.n12213 S.n12212 3.773
R4550 S.n12213 S.t137 3.773
R4551 S.n11542 S.n11541 3.773
R4552 S.n11542 S.t329 3.773
R4553 S.n11547 S.t1202 3.773
R4554 S.n11547 S.n11546 3.773
R4555 S.n11550 S.t964 3.773
R4556 S.n11550 S.n11549 3.773
R4557 S.n11539 S.n11538 3.773
R4558 S.n11539 S.t96 3.773
R4559 S.n11303 S.n11302 3.773
R4560 S.n11303 S.t306 3.773
R4561 S.n11307 S.t1174 3.773
R4562 S.n11307 S.n11306 3.773
R4563 S.n11310 S.t939 3.773
R4564 S.n11310 S.n11309 3.773
R4565 S.n11300 S.n11299 3.773
R4566 S.n11300 S.t58 3.773
R4567 S.n10926 S.n10925 3.773
R4568 S.n10926 S.t283 3.773
R4569 S.n10931 S.t1149 3.773
R4570 S.n10931 S.n10930 3.773
R4571 S.n10934 S.t912 3.773
R4572 S.n10934 S.n10933 3.773
R4573 S.n10923 S.n10922 3.773
R4574 S.n10923 S.t16 3.773
R4575 S.n10675 S.n10674 3.773
R4576 S.n10675 S.t253 3.773
R4577 S.n10679 S.t1123 3.773
R4578 S.n10679 S.n10678 3.773
R4579 S.n10682 S.t884 3.773
R4580 S.n10682 S.n10681 3.773
R4581 S.n10672 S.n10671 3.773
R4582 S.n10672 S.t2561 3.773
R4583 S.n10276 S.n10275 3.773
R4584 S.n10276 S.t224 3.773
R4585 S.n10281 S.t1099 3.773
R4586 S.n10281 S.n10280 3.773
R4587 S.n10284 S.t859 3.773
R4588 S.n10284 S.n10283 3.773
R4589 S.n10273 S.n10272 3.773
R4590 S.n10273 S.t2533 3.773
R4591 S.n10017 S.n10016 3.773
R4592 S.n10017 S.t2331 3.773
R4593 S.n10021 S.t675 3.773
R4594 S.n10021 S.n10020 3.773
R4595 S.n10024 S.t461 3.773
R4596 S.n10024 S.n10023 3.773
R4597 S.n10014 S.n10013 3.773
R4598 S.n10014 S.t2512 3.773
R4599 S.n9621 S.n9620 3.773
R4600 S.n9621 S.t2305 3.773
R4601 S.n9618 S.t649 3.773
R4602 S.n9618 S.n9617 3.773
R4603 S.n9615 S.t434 3.773
R4604 S.n9615 S.n9614 3.773
R4605 S.n9345 S.n9344 3.773
R4606 S.n9345 S.t2115 3.773
R4607 S.n9632 S.t846 3.773
R4608 S.n9634 S.t1345 3.773
R4609 S.n9636 S.t1061 3.773
R4610 S.n9597 S.n9596 3.773
R4611 S.n9597 S.t2010 3.773
R4612 S.n9609 S.t1437 3.773
R4613 S.n9609 S.n9608 3.773
R4614 S.n9612 S.t1900 3.773
R4615 S.n9612 S.n9611 3.773
R4616 S.n9600 S.n9599 3.773
R4617 S.n9600 S.t499 3.773
R4618 S.n10032 S.n10031 3.773
R4619 S.n10032 S.t595 3.773
R4620 S.n10318 S.t1462 3.773
R4621 S.n10318 S.n10317 3.773
R4622 S.n10321 S.t1248 3.773
R4623 S.n10321 S.n10320 3.773
R4624 S.n10029 S.n10028 3.773
R4625 S.n10029 S.t773 3.773
R4626 S.n11977 S.t1003 3.773
R4627 S.n11975 S.t1523 3.773
R4628 S.n11974 S.t2389 3.773
R4629 S.n11700 S.n11699 3.773
R4630 S.n11700 S.t1197 3.773
R4631 S.n11707 S.t2515 3.773
R4632 S.n11707 S.n11706 3.773
R4633 S.n11704 S.t1830 3.773
R4634 S.n11704 S.n11703 3.773
R4635 S.n11697 S.n11696 3.773
R4636 S.n11697 S.t988 3.773
R4637 S.n12516 S.n12515 3.773
R4638 S.n12516 S.t1165 3.773
R4639 S.n12521 S.t2028 3.773
R4640 S.n12521 S.n12520 3.773
R4641 S.n12524 S.t1799 3.773
R4642 S.n12524 S.n12523 3.773
R4643 S.n12513 S.n12512 3.773
R4644 S.n12513 S.t958 3.773
R4645 S.n12231 S.n12230 3.773
R4646 S.n12231 S.t1144 3.773
R4647 S.n12235 S.t2007 3.773
R4648 S.n12235 S.n12234 3.773
R4649 S.n12238 S.t1776 3.773
R4650 S.n12238 S.n12237 3.773
R4651 S.n12228 S.n12227 3.773
R4652 S.n12228 S.t934 3.773
R4653 S.n11558 S.n11557 3.773
R4654 S.n11558 S.t1119 3.773
R4655 S.n11563 S.t1982 3.773
R4656 S.n11563 S.n11562 3.773
R4657 S.n11566 S.t1745 3.773
R4658 S.n11566 S.n11565 3.773
R4659 S.n11555 S.n11554 3.773
R4660 S.n11555 S.t907 3.773
R4661 S.n11318 S.n11317 3.773
R4662 S.n11318 S.t1089 3.773
R4663 S.n11322 S.t1958 3.773
R4664 S.n11322 S.n11321 3.773
R4665 S.n11325 S.t1720 3.773
R4666 S.n11325 S.n11324 3.773
R4667 S.n11315 S.n11314 3.773
R4668 S.n11315 S.t877 3.773
R4669 S.n10942 S.n10941 3.773
R4670 S.n10942 S.t1064 3.773
R4671 S.n10947 S.t1932 3.773
R4672 S.n10947 S.n10946 3.773
R4673 S.n10950 S.t1692 3.773
R4674 S.n10950 S.n10949 3.773
R4675 S.n10939 S.n10938 3.773
R4676 S.n10939 S.t854 3.773
R4677 S.n10690 S.n10689 3.773
R4678 S.n10690 S.t1037 3.773
R4679 S.n10694 S.t1905 3.773
R4680 S.n10694 S.n10693 3.773
R4681 S.n10697 S.t1666 3.773
R4682 S.n10697 S.n10696 3.773
R4683 S.n10687 S.n10686 3.773
R4684 S.n10687 S.t827 3.773
R4685 S.n10313 S.n10312 3.773
R4686 S.n10313 S.t1011 3.773
R4687 S.n10310 S.t1879 3.773
R4688 S.n10310 S.n10309 3.773
R4689 S.n10307 S.t1643 3.773
R4690 S.n10307 S.n10306 3.773
R4691 S.n10037 S.n10036 3.773
R4692 S.n10037 S.t798 3.773
R4693 S.n10324 S.t634 3.773
R4694 S.n10326 S.t755 3.773
R4695 S.n10328 S.t681 3.773
R4696 S.n10289 S.n10288 3.773
R4697 S.n10289 S.t1106 3.773
R4698 S.n10301 S.t125 3.773
R4699 S.n10301 S.n10300 3.773
R4700 S.n10304 S.t2483 3.773
R4701 S.n10304 S.n10303 3.773
R4702 S.n10292 S.n10291 3.773
R4703 S.n10292 S.t1095 3.773
R4704 S.n10705 S.n10704 3.773
R4705 S.n10705 S.t1818 3.773
R4706 S.n10984 S.t156 3.773
R4707 S.n10984 S.n10983 3.773
R4708 S.n10987 S.t2454 3.773
R4709 S.n10987 S.n10986 3.773
R4710 S.n10702 S.n10701 3.773
R4711 S.n10702 S.t1610 3.773
R4712 S.n11981 S.t1668 3.773
R4713 S.n11979 S.t478 3.773
R4714 S.n11978 S.t778 3.773
R4715 S.n11685 S.n11684 3.773
R4716 S.n11685 S.t1977 3.773
R4717 S.n11692 S.t325 3.773
R4718 S.n11692 S.n11691 3.773
R4719 S.n11689 S.t50 3.773
R4720 S.n11689 S.n11688 3.773
R4721 S.n11682 S.n11681 3.773
R4722 S.n11682 S.t1770 3.773
R4723 S.n12532 S.n12531 3.773
R4724 S.n12532 S.t1952 3.773
R4725 S.n12537 S.t299 3.773
R4726 S.n12537 S.n12536 3.773
R4727 S.n12540 S.t1 3.773
R4728 S.n12540 S.n12539 3.773
R4729 S.n12529 S.n12528 3.773
R4730 S.n12529 S.t1740 3.773
R4731 S.n12246 S.n12245 3.773
R4732 S.n12246 S.t1926 3.773
R4733 S.n12250 S.t277 3.773
R4734 S.n12250 S.n12249 3.773
R4735 S.n12253 S.t2556 3.773
R4736 S.n12253 S.n12252 3.773
R4737 S.n12243 S.n12242 3.773
R4738 S.n12243 S.t1713 3.773
R4739 S.n11574 S.n11573 3.773
R4740 S.n11574 S.t1901 3.773
R4741 S.n11579 S.t250 3.773
R4742 S.n11579 S.n11578 3.773
R4743 S.n11582 S.t2527 3.773
R4744 S.n11582 S.n11581 3.773
R4745 S.n11571 S.n11570 3.773
R4746 S.n11571 S.t1687 3.773
R4747 S.n11333 S.n11332 3.773
R4748 S.n11333 S.t1871 3.773
R4749 S.n11337 S.t216 3.773
R4750 S.n11337 S.n11336 3.773
R4751 S.n11340 S.t2506 3.773
R4752 S.n11340 S.n11339 3.773
R4753 S.n11330 S.n11329 3.773
R4754 S.n11330 S.t1659 3.773
R4755 S.n10979 S.n10978 3.773
R4756 S.n10979 S.t1849 3.773
R4757 S.n10976 S.t190 3.773
R4758 S.n10976 S.n10975 3.773
R4759 S.n10973 S.t2482 3.773
R4760 S.n10973 S.n10972 3.773
R4761 S.n10710 S.n10709 3.773
R4762 S.n10710 S.t1635 3.773
R4763 S.n10990 S.t2243 3.773
R4764 S.n10992 S.t409 3.773
R4765 S.n10994 S.t92 3.773
R4766 S.n10955 S.n10954 3.773
R4767 S.n10955 S.t874 3.773
R4768 S.n10967 S.t978 3.773
R4769 S.n10967 S.n10966 3.773
R4770 S.n10970 S.t2210 3.773
R4771 S.n10970 S.n10969 3.773
R4772 S.n10958 S.n10957 3.773
R4773 S.n10958 S.t800 3.773
R4774 S.n11348 S.n11347 3.773
R4775 S.n11348 S.t116 3.773
R4776 S.n11619 S.t1005 3.773
R4777 S.n11619 S.n11618 3.773
R4778 S.n11622 S.t764 3.773
R4779 S.n11622 S.n11621 3.773
R4780 S.n11345 S.n11344 3.773
R4781 S.n11345 S.t2447 3.773
R4782 S.n11985 S.t2459 3.773
R4783 S.n11983 S.t1265 3.773
R4784 S.n11982 S.t2134 3.773
R4785 S.n11670 S.n11669 3.773
R4786 S.n11670 S.t240 3.773
R4787 S.n11677 S.t1113 3.773
R4788 S.n11677 S.n11676 3.773
R4789 S.n11674 S.t873 3.773
R4790 S.n11674 S.n11673 3.773
R4791 S.n11667 S.n11666 3.773
R4792 S.n11667 S.t2549 3.773
R4793 S.n12548 S.n12547 3.773
R4794 S.n12548 S.t210 3.773
R4795 S.n12553 S.t1084 3.773
R4796 S.n12553 S.n12552 3.773
R4797 S.n12556 S.t845 3.773
R4798 S.n12556 S.n12555 3.773
R4799 S.n12545 S.n12544 3.773
R4800 S.n12545 S.t2524 3.773
R4801 S.n12261 S.n12260 3.773
R4802 S.n12261 S.t182 3.773
R4803 S.n12265 S.t1057 3.773
R4804 S.n12265 S.n12264 3.773
R4805 S.n12268 S.t821 3.773
R4806 S.n12268 S.n12267 3.773
R4807 S.n12258 S.n12257 3.773
R4808 S.n12258 S.t2501 3.773
R4809 S.n11614 S.n11613 3.773
R4810 S.n11614 S.t151 3.773
R4811 S.n11611 S.t1032 3.773
R4812 S.n11611 S.n11610 3.773
R4813 S.n11608 S.t791 3.773
R4814 S.n11608 S.n11607 3.773
R4815 S.n11353 S.n11352 3.773
R4816 S.n11353 S.t2474 3.773
R4817 S.n11625 S.t2040 3.773
R4818 S.n11627 S.t2349 3.773
R4819 S.n11629 S.t2074 3.773
R4820 S.n11585 S.n11584 3.773
R4821 S.n11585 S.t659 3.773
R4822 S.n11602 S.t1811 3.773
R4823 S.n11602 S.n11601 3.773
R4824 S.n11605 S.t1941 3.773
R4825 S.n11605 S.n11604 3.773
R4826 S.n11588 S.n11587 3.773
R4827 S.n11588 S.t531 3.773
R4828 S.n12575 S.n12574 3.773
R4829 S.n12575 S.t973 3.773
R4830 S.n12584 S.t1842 3.773
R4831 S.n12584 S.n12583 3.773
R4832 S.n12587 S.t1603 3.773
R4833 S.n12587 S.n12586 3.773
R4834 S.n12578 S.n12577 3.773
R4835 S.n12578 S.t759 3.773
R4836 S.n11989 S.t717 3.773
R4837 S.n11986 S.t2055 3.773
R4838 S.n11987 S.t400 3.773
R4839 S.n11651 S.n11650 3.773
R4840 S.n11651 S.t1025 3.773
R4841 S.n11662 S.t1893 3.773
R4842 S.n11662 S.n11661 3.773
R4843 S.n11659 S.t1655 3.773
R4844 S.n11659 S.n11658 3.773
R4845 S.n11654 S.n11653 3.773
R4846 S.n11654 S.t815 3.773
R4847 S.n12277 S.n12276 3.773
R4848 S.n12277 S.t999 3.773
R4849 S.n12559 S.t1866 3.773
R4850 S.n12559 S.n12558 3.773
R4851 S.n12562 S.t1630 3.773
R4852 S.n12562 S.n12561 3.773
R4853 S.n12565 S.n12564 3.773
R4854 S.n12565 S.t785 3.773
R4855 S.n11928 S.t2295 3.773
R4856 S.n11929 S.t1110 3.773
R4857 S.n11926 S.t1973 3.773
R4858 S.n528 S.n526 2.808
R4859 S.n1475 S.n1473 2.808
R4860 S.n2349 S.n2347 2.808
R4861 S.n3131 S.n3129 2.808
R4862 S.n4033 S.n4031 2.808
R4863 S.n4850 S.n4848 2.808
R4864 S.n5649 S.n5647 2.808
R4865 S.n6422 S.n6420 2.808
R4866 S.n7186 S.n7184 2.808
R4867 S.n7757 S.n7755 2.808
R4868 S.n8471 S.n8469 2.808
R4869 S.n9356 S.n9354 2.808
R4870 S.n10050 S.n10048 2.808
R4871 S.n10718 S.n10716 2.808
R4872 S.n65 S.n64 2.645
R4873 S.n522 S.n521 2.645
R4874 S.n1469 S.n1468 2.645
R4875 S.n2343 S.n2342 2.645
R4876 S.n3125 S.n3124 2.645
R4877 S.n4027 S.n4026 2.645
R4878 S.n4844 S.n4843 2.645
R4879 S.n5643 S.n5642 2.645
R4880 S.n6416 S.n6415 2.645
R4881 S.n7180 S.n7179 2.645
R4882 S.n7751 S.n7750 2.645
R4883 S.n8465 S.n8464 2.645
R4884 S.n9350 S.n9349 2.645
R4885 S.n10044 S.n10043 2.645
R4886 S.n11642 S.n11641 0.21
R4887 S.n976 S.n975 0.172
R4888 S.n67 S.n63 0.164
R4889 S.n11996 S.n11995 0.143
R4890 S.n2217 S.n2216 0.133
R4891 S.n1807 S.n1806 0.133
R4892 S.n245 S.n237 0.123
R4893 S.n131 S.n130 0.123
R4894 S.n118 S.n117 0.123
R4895 S.n105 S.n104 0.123
R4896 S.n92 S.n91 0.123
R4897 S.n57 S.n56 0.12
R4898 S.n20 S.n19 0.12
R4899 S.n29 S.n28 0.12
R4900 S.n38 S.n37 0.12
R4901 S.n47 S.n46 0.12
R4902 S.n12626 S.n1827 0.114
R4903 S.n12627 S.n980 0.111
R4904 S.n12625 S.n2696 0.111
R4905 S.n12623 S.n4369 0.111
R4906 S.n12622 S.n5175 0.111
R4907 S.n12621 S.n5972 0.111
R4908 S.n12620 S.n6743 0.111
R4909 S.n12619 S.n7505 0.111
R4910 S.n12618 S.n8241 0.111
R4911 S.n12617 S.n8968 0.111
R4912 S.n12616 S.n9669 0.111
R4913 S.n12615 S.n10361 0.111
R4914 S.n12614 S.n11025 0.111
R4915 S.n12613 S.n11644 0.111
R4916 S.n12612 S.n12611 0.11
R4917 S.n12624 S.n3537 0.11
R4918 S.n11996 S.n11923 0.11
R4919 S.n11381 S.n11379 0.109
R4920 S.n10764 S.n10762 0.109
R4921 S.n10114 S.n10112 0.109
R4922 S.n9438 S.n9436 0.109
R4923 S.n8571 S.n8569 0.109
R4924 S.n7875 S.n7873 0.109
R4925 S.n7322 S.n7320 0.109
R4926 S.n6576 S.n6574 0.109
R4927 S.n5821 S.n5819 0.109
R4928 S.n5040 S.n5038 0.109
R4929 S.n4241 S.n4239 0.109
R4930 S.n3357 S.n3355 0.109
R4931 S.n2593 S.n2591 0.109
R4932 S.n2632 S.n2629 0.106
R4933 S.n3411 S.n3408 0.106
R4934 S.n4296 S.n4293 0.106
R4935 S.n5111 S.n5108 0.106
R4936 S.n5908 S.n5905 0.106
R4937 S.n6679 S.n6676 0.106
R4938 S.n7441 S.n7438 0.106
R4939 S.n8025 S.n8022 0.106
R4940 S.n8737 S.n8734 0.106
R4941 S.n9605 S.n9602 0.106
R4942 S.n10297 S.n10294 0.106
R4943 S.n10963 S.n10960 0.106
R4944 S.n12325 S.n12320 0.106
R4945 S.n2177 S.n2176 0.097
R4946 S.n3013 S.n3012 0.097
R4947 S.n3825 S.n3824 0.097
R4948 S.n4625 S.n4624 0.097
R4949 S.n5402 S.n5401 0.097
R4950 S.n6167 S.n6166 0.097
R4951 S.n6909 S.n6908 0.097
R4952 S.n7639 S.n7638 0.097
R4953 S.n8346 S.n8345 0.097
R4954 S.n9041 S.n9040 0.097
R4955 S.n9713 S.n9712 0.097
R4956 S.n10373 S.n10372 0.097
R4957 S.n11090 S.n11089 0.097
R4958 S.n1374 S.n1373 0.097
R4959 S.n1402 S.n1401 0.097
R4960 S.n12604 S.n12603 0.095
R4961 S.n12282 S.n12281 0.093
R4962 S.n1331 S.n1330 0.087
R4963 S.n977 S.n974 0.081
R4964 S.n990 S.n987 0.081
R4965 S.n2675 S.n2672 0.081
R4966 S.n3516 S.n3514 0.081
R4967 S.n4348 S.n4345 0.081
R4968 S.n5154 S.n5151 0.081
R4969 S.n5951 S.n5948 0.081
R4970 S.n6722 S.n6719 0.081
R4971 S.n7484 S.n7481 0.081
R4972 S.n8220 S.n8217 0.081
R4973 S.n8947 S.n8944 0.081
R4974 S.n9648 S.n9645 0.081
R4975 S.n10340 S.n10337 0.081
R4976 S.n11004 S.n11001 0.081
R4977 S.n11085 S.n11084 0.08
R4978 S.n10368 S.n10367 0.08
R4979 S.n9708 S.n9707 0.08
R4980 S.n9036 S.n9035 0.08
R4981 S.n8341 S.n8340 0.08
R4982 S.n7634 S.n7633 0.08
R4983 S.n6904 S.n6903 0.08
R4984 S.n6162 S.n6161 0.08
R4985 S.n5397 S.n5396 0.08
R4986 S.n4620 S.n4619 0.08
R4987 S.n3820 S.n3819 0.08
R4988 S.n3008 S.n3007 0.08
R4989 S.n2172 S.n2171 0.08
R4990 S.n1404 S.n1403 0.08
R4991 S.n1376 S.n1375 0.08
R4992 S.n2689 S.n2688 0.079
R4993 S.n3530 S.n3529 0.079
R4994 S.n4362 S.n4361 0.079
R4995 S.n5168 S.n5167 0.079
R4996 S.n5965 S.n5964 0.079
R4997 S.n6736 S.n6735 0.079
R4998 S.n7498 S.n7497 0.079
R4999 S.n8234 S.n8233 0.079
R5000 S.n8961 S.n8960 0.079
R5001 S.n9662 S.n9661 0.079
R5002 S.n10354 S.n10353 0.079
R5003 S.n11018 S.n11017 0.079
R5004 S.n1712 S.n1711 0.077
R5005 S.n2563 S.n2562 0.077
R5006 S.n3327 S.n3326 0.077
R5007 S.n4211 S.n4210 0.077
R5008 S.n5010 S.n5009 0.077
R5009 S.n5791 S.n5790 0.077
R5010 S.n6546 S.n6545 0.077
R5011 S.n7292 S.n7291 0.077
R5012 S.n7845 S.n7844 0.077
R5013 S.n8541 S.n8540 0.077
R5014 S.n9408 S.n9407 0.077
R5015 S.n10084 S.n10083 0.077
R5016 S.n10734 S.n10733 0.077
R5017 S.n750 S.n749 0.077
R5018 S.n769 S.n768 0.077
R5019 S.n2692 S.n2691 0.075
R5020 S.n3533 S.n3532 0.075
R5021 S.n4365 S.n4364 0.075
R5022 S.n5171 S.n5170 0.075
R5023 S.n5968 S.n5967 0.075
R5024 S.n6739 S.n6738 0.075
R5025 S.n7501 S.n7500 0.075
R5026 S.n8237 S.n8236 0.075
R5027 S.n8964 S.n8963 0.075
R5028 S.n9665 S.n9664 0.075
R5029 S.n10357 S.n10356 0.075
R5030 S.n11021 S.n11020 0.075
R5031 S.n10723 S.n10722 0.074
R5032 S.n10055 S.n10054 0.074
R5033 S.n9361 S.n9360 0.074
R5034 S.n8476 S.n8475 0.074
R5035 S.n7762 S.n7761 0.074
R5036 S.n7191 S.n7190 0.074
R5037 S.n6427 S.n6426 0.074
R5038 S.n5654 S.n5653 0.074
R5039 S.n4855 S.n4854 0.074
R5040 S.n4038 S.n4037 0.074
R5041 S.n3136 S.n3135 0.074
R5042 S.n2354 S.n2353 0.074
R5043 S.n1480 S.n1479 0.074
R5044 S.n533 S.n532 0.074
R5045 S.n10375 S.n10374 0.071
R5046 S.n9715 S.n9714 0.071
R5047 S.n9043 S.n9042 0.071
R5048 S.n8348 S.n8347 0.071
R5049 S.n7641 S.n7640 0.071
R5050 S.n6911 S.n6910 0.071
R5051 S.n6169 S.n6168 0.071
R5052 S.n5404 S.n5403 0.071
R5053 S.n4627 S.n4626 0.071
R5054 S.n3827 S.n3826 0.071
R5055 S.n3015 S.n3014 0.071
R5056 S.n2179 S.n2178 0.071
R5057 S.n1370 S.n1369 0.071
R5058 S.n1398 S.n1397 0.071
R5059 S.n12323 S.n12322 0.07
R5060 S.n202 S.n200 0.067
R5061 S.n202 S.n201 0.067
R5062 S.n164 S.n162 0.067
R5063 S.n164 S.n163 0.067
R5064 S.n183 S.n181 0.067
R5065 S.n183 S.n182 0.067
R5066 S.n196 S.n194 0.067
R5067 S.n196 S.n195 0.067
R5068 S.n6 S.n4 0.067
R5069 S.n6 S.n5 0.067
R5070 S.n151 S.n149 0.067
R5071 S.n151 S.n150 0.067
R5072 S.n14 S.n12 0.067
R5073 S.n14 S.n13 0.067
R5074 S.n139 S.n137 0.067
R5075 S.n139 S.n138 0.067
R5076 S.n23 S.n21 0.067
R5077 S.n23 S.n22 0.067
R5078 S.n126 S.n124 0.067
R5079 S.n126 S.n125 0.067
R5080 S.n32 S.n30 0.067
R5081 S.n32 S.n31 0.067
R5082 S.n113 S.n111 0.067
R5083 S.n113 S.n112 0.067
R5084 S.n41 S.n39 0.067
R5085 S.n41 S.n40 0.067
R5086 S.n100 S.n98 0.067
R5087 S.n100 S.n99 0.067
R5088 S.n50 S.n48 0.067
R5089 S.n50 S.n49 0.067
R5090 S.n87 S.n85 0.067
R5091 S.n87 S.n86 0.067
R5092 S.n54 S.n53 0.067
R5093 S.n54 S.n52 0.067
R5094 S.n977 S.n967 0.067
R5095 S.n977 S.n965 0.067
R5096 S.n2675 S.n2666 0.067
R5097 S.n2675 S.n2665 0.067
R5098 S.n3516 S.n3515 0.067
R5099 S.n4348 S.n4339 0.067
R5100 S.n4348 S.n4338 0.067
R5101 S.n5154 S.n5145 0.067
R5102 S.n5154 S.n5144 0.067
R5103 S.n5951 S.n5942 0.067
R5104 S.n5951 S.n5941 0.067
R5105 S.n6722 S.n6713 0.067
R5106 S.n6722 S.n6712 0.067
R5107 S.n7484 S.n7475 0.067
R5108 S.n7484 S.n7474 0.067
R5109 S.n8220 S.n8211 0.067
R5110 S.n8220 S.n8210 0.067
R5111 S.n8947 S.n8938 0.067
R5112 S.n8947 S.n8937 0.067
R5113 S.n9648 S.n9639 0.067
R5114 S.n9648 S.n9638 0.067
R5115 S.n10340 S.n10331 0.067
R5116 S.n10340 S.n10330 0.067
R5117 S.n3516 S.n3506 0.067
R5118 S.n80 S.n79 0.066
R5119 S.n870 S.n869 0.066
R5120 S.n979 S.n978 0.065
R5121 S.n197 S.n196 0.063
R5122 S.n1431 S.n1430 0.063
R5123 S.n1762 S.n1761 0.063
R5124 S.n2250 S.n2249 0.063
R5125 S.n2613 S.n2612 0.063
R5126 S.n3085 S.n3084 0.063
R5127 S.n3377 S.n3376 0.063
R5128 S.n3897 S.n3896 0.063
R5129 S.n4261 S.n4260 0.063
R5130 S.n4697 S.n4696 0.063
R5131 S.n5060 S.n5059 0.063
R5132 S.n5474 S.n5473 0.063
R5133 S.n5841 S.n5840 0.063
R5134 S.n6239 S.n6238 0.063
R5135 S.n6596 S.n6595 0.063
R5136 S.n6981 S.n6980 0.063
R5137 S.n7342 S.n7341 0.063
R5138 S.n7711 S.n7710 0.063
R5139 S.n7895 S.n7894 0.063
R5140 S.n8418 S.n8417 0.063
R5141 S.n8591 S.n8590 0.063
R5142 S.n9113 S.n9112 0.063
R5143 S.n9458 S.n9457 0.063
R5144 S.n9785 S.n9784 0.063
R5145 S.n10134 S.n10133 0.063
R5146 S.n10445 S.n10444 0.063
R5147 S.n10784 S.n10783 0.063
R5148 S.n11075 S.n11074 0.063
R5149 S.n11401 S.n11400 0.063
R5150 S.n12023 S.n12022 0.063
R5151 S.n12303 S.n12302 0.063
R5152 S.n920 S.n907 0.063
R5153 S.n1344 S.n1320 0.063
R5154 S.n1702 S.n1688 0.063
R5155 S.n2163 S.n2162 0.063
R5156 S.n2553 S.n2552 0.063
R5157 S.n2999 S.n2998 0.063
R5158 S.n3317 S.n3316 0.063
R5159 S.n3811 S.n3810 0.063
R5160 S.n4201 S.n4200 0.063
R5161 S.n4611 S.n4610 0.063
R5162 S.n5000 S.n4999 0.063
R5163 S.n5388 S.n5387 0.063
R5164 S.n5781 S.n5780 0.063
R5165 S.n6153 S.n6152 0.063
R5166 S.n6536 S.n6535 0.063
R5167 S.n6895 S.n6894 0.063
R5168 S.n7282 S.n7281 0.063
R5169 S.n7625 S.n7624 0.063
R5170 S.n7835 S.n7834 0.063
R5171 S.n8332 S.n8331 0.063
R5172 S.n8531 S.n8530 0.063
R5173 S.n9027 S.n9026 0.063
R5174 S.n9398 S.n9397 0.063
R5175 S.n9699 S.n9698 0.063
R5176 S.n10074 S.n10073 0.063
R5177 S.n1406 S.n1386 0.063
R5178 S.n2218 S.n2205 0.063
R5179 S.n3053 S.n3041 0.063
R5180 S.n3865 S.n3853 0.063
R5181 S.n4665 S.n4653 0.063
R5182 S.n5442 S.n5430 0.063
R5183 S.n6207 S.n6195 0.063
R5184 S.n6949 S.n6937 0.063
R5185 S.n7679 S.n7667 0.063
R5186 S.n8386 S.n8374 0.063
R5187 S.n9081 S.n9069 0.063
R5188 S.n9753 S.n9741 0.063
R5189 S.n10413 S.n10401 0.063
R5190 S.n11043 S.n11031 0.063
R5191 S.n899 S.n879 0.063
R5192 S.n8995 S.n8974 0.063
R5193 S.n8300 S.n8279 0.063
R5194 S.n7593 S.n7572 0.063
R5195 S.n6863 S.n6842 0.063
R5196 S.n6121 S.n6100 0.063
R5197 S.n5356 S.n5335 0.063
R5198 S.n4579 S.n4558 0.063
R5199 S.n3779 S.n3758 0.063
R5200 S.n2967 S.n2946 0.063
R5201 S.n2130 S.n2109 0.063
R5202 S.n1310 S.n1291 0.063
R5203 S.n507 S.n492 0.063
R5204 S.n1282 S.n1281 0.063
R5205 S.n1661 S.n1660 0.063
R5206 S.n2101 S.n2100 0.063
R5207 S.n2517 S.n2516 0.063
R5208 S.n2938 S.n2937 0.063
R5209 S.n3281 S.n3280 0.063
R5210 S.n3750 S.n3749 0.063
R5211 S.n4165 S.n4164 0.063
R5212 S.n4550 S.n4549 0.063
R5213 S.n4964 S.n4963 0.063
R5214 S.n5327 S.n5326 0.063
R5215 S.n5745 S.n5744 0.063
R5216 S.n6092 S.n6091 0.063
R5217 S.n6500 S.n6499 0.063
R5218 S.n6834 S.n6833 0.063
R5219 S.n7246 S.n7245 0.063
R5220 S.n7564 S.n7563 0.063
R5221 S.n7799 S.n7798 0.063
R5222 S.n8271 S.n8270 0.063
R5223 S.n8495 S.n8494 0.063
R5224 S.n7532 S.n7511 0.063
R5225 S.n6802 S.n6781 0.063
R5226 S.n6060 S.n6039 0.063
R5227 S.n5295 S.n5274 0.063
R5228 S.n4518 S.n4497 0.063
R5229 S.n3718 S.n3697 0.063
R5230 S.n2906 S.n2885 0.063
R5231 S.n2069 S.n2048 0.063
R5232 S.n1252 S.n1232 0.063
R5233 S.n466 S.n448 0.063
R5234 S.n1223 S.n1222 0.063
R5235 S.n1625 S.n1624 0.063
R5236 S.n2040 S.n2039 0.063
R5237 S.n2481 S.n2480 0.063
R5238 S.n2877 S.n2876 0.063
R5239 S.n3245 S.n3244 0.063
R5240 S.n3689 S.n3688 0.063
R5241 S.n4129 S.n4128 0.063
R5242 S.n4489 S.n4488 0.063
R5243 S.n4928 S.n4927 0.063
R5244 S.n5266 S.n5265 0.063
R5245 S.n5709 S.n5708 0.063
R5246 S.n6031 S.n6030 0.063
R5247 S.n6464 S.n6463 0.063
R5248 S.n6773 S.n6772 0.063
R5249 S.n7210 S.n7209 0.063
R5250 S.n5999 S.n5978 0.063
R5251 S.n5234 S.n5213 0.063
R5252 S.n4457 S.n4436 0.063
R5253 S.n3657 S.n3636 0.063
R5254 S.n2845 S.n2824 0.063
R5255 S.n2008 S.n1987 0.063
R5256 S.n1193 S.n1173 0.063
R5257 S.n419 S.n404 0.063
R5258 S.n1164 S.n1163 0.063
R5259 S.n1589 S.n1588 0.063
R5260 S.n1979 S.n1978 0.063
R5261 S.n2445 S.n2444 0.063
R5262 S.n2816 S.n2815 0.063
R5263 S.n3209 S.n3208 0.063
R5264 S.n3628 S.n3627 0.063
R5265 S.n4093 S.n4092 0.063
R5266 S.n4428 S.n4427 0.063
R5267 S.n4892 S.n4891 0.063
R5268 S.n5205 S.n5204 0.063
R5269 S.n5673 S.n5672 0.063
R5270 S.n4396 S.n4375 0.063
R5271 S.n3596 S.n3575 0.063
R5272 S.n2784 S.n2763 0.063
R5273 S.n1950 S.n1926 0.063
R5274 S.n1134 S.n1114 0.063
R5275 S.n375 S.n360 0.063
R5276 S.n1105 S.n1104 0.063
R5277 S.n1553 S.n1552 0.063
R5278 S.n1918 S.n1917 0.063
R5279 S.n2409 S.n2408 0.063
R5280 S.n2755 S.n2754 0.063
R5281 S.n3173 S.n3172 0.063
R5282 S.n3567 S.n3566 0.063
R5283 S.n4057 S.n4056 0.063
R5284 S.n2723 S.n2702 0.063
R5285 S.n1886 S.n1865 0.063
R5286 S.n1075 S.n1055 0.063
R5287 S.n331 S.n316 0.063
R5288 S.n1046 S.n1045 0.063
R5289 S.n1517 S.n1516 0.063
R5290 S.n1857 S.n1856 0.063
R5291 S.n2373 S.n2372 0.063
R5292 S.n1016 S.n996 0.063
R5293 S.n287 S.n272 0.063
R5294 S.n950 S.n949 0.063
R5295 S.n203 S.n202 0.062
R5296 S.n152 S.n151 0.062
R5297 S.n140 S.n139 0.062
R5298 S.n127 S.n126 0.062
R5299 S.n114 S.n113 0.062
R5300 S.n101 S.n100 0.062
R5301 S.n88 S.n87 0.062
R5302 S.n184 S.n183 0.061
R5303 S.n7 S.n6 0.06
R5304 S.n15 S.n14 0.06
R5305 S.n24 S.n23 0.06
R5306 S.n33 S.n32 0.06
R5307 S.n42 S.n41 0.06
R5308 S.n51 S.n50 0.06
R5309 S.n55 S.n54 0.06
R5310 S.n12031 S.n12030 0.059
R5311 S.n2148 S.n2138 0.059
R5312 S.n165 S.n164 0.059
R5313 S.n2678 S.n2677 0.058
R5314 S.n3519 S.n3518 0.058
R5315 S.n4351 S.n4350 0.058
R5316 S.n5157 S.n5156 0.058
R5317 S.n5954 S.n5953 0.058
R5318 S.n6725 S.n6724 0.058
R5319 S.n7487 S.n7486 0.058
R5320 S.n8223 S.n8222 0.058
R5321 S.n8950 S.n8949 0.058
R5322 S.n9651 S.n9650 0.058
R5323 S.n10343 S.n10342 0.058
R5324 S.n11007 S.n11006 0.058
R5325 S.n979 S.n977 0.058
R5326 S.n83 S.n61 0.055
R5327 S.n11920 S.n11645 0.054
R5328 S.n535 S.n518 0.054
R5329 S.n9364 S.n9347 0.054
R5330 S.n10057 S.n10039 0.054
R5331 S.n10726 S.n10712 0.054
R5332 S.n11364 S.n11355 0.054
R5333 S.n12286 S.n12279 0.054
R5334 S.n7765 S.n7748 0.054
R5335 S.n8478 S.n8460 0.054
R5336 S.n6430 S.n6413 0.054
R5337 S.n7193 S.n7175 0.054
R5338 S.n4858 S.n4841 0.054
R5339 S.n5656 S.n5638 0.054
R5340 S.n3139 S.n3122 0.054
R5341 S.n4040 S.n4022 0.054
R5342 S.n1483 S.n1466 0.054
R5343 S.n2356 S.n2338 0.054
R5344 S S.n12627 0.054
R5345 S.n12593 S.n12592 0.054
R5346 S.n961 S.n960 0.054
R5347 S.n1819 S.n1818 0.054
R5348 S.n2662 S.n2661 0.054
R5349 S.n3503 S.n3502 0.054
R5350 S.n4335 S.n4334 0.054
R5351 S.n5141 S.n5140 0.054
R5352 S.n5938 S.n5937 0.054
R5353 S.n6709 S.n6708 0.054
R5354 S.n7471 S.n7470 0.054
R5355 S.n8207 S.n8206 0.054
R5356 S.n8934 S.n8933 0.054
R5357 S.n9635 S.n9634 0.054
R5358 S.n10327 S.n10326 0.054
R5359 S.n10993 S.n10992 0.054
R5360 S.n11628 S.n11627 0.054
R5361 S S.n245 0.053
R5362 S.n531 S.n530 0.053
R5363 S.n1478 S.n1477 0.053
R5364 S.n2352 S.n2351 0.053
R5365 S.n3134 S.n3133 0.053
R5366 S.n4036 S.n4035 0.053
R5367 S.n4853 S.n4852 0.053
R5368 S.n5652 S.n5651 0.053
R5369 S.n6425 S.n6424 0.053
R5370 S.n7189 S.n7188 0.053
R5371 S.n7760 S.n7759 0.053
R5372 S.n8474 S.n8473 0.053
R5373 S.n9359 S.n9358 0.053
R5374 S.n10053 S.n10052 0.053
R5375 S.n10721 S.n10720 0.053
R5376 S.n11917 S.n11916 0.053
R5377 S.n12330 S.n12329 0.053
R5378 S.n956 S.n955 0.053
R5379 S.n923 S.n922 0.053
R5380 S.n1434 S.n1433 0.053
R5381 S.n11894 S.n11893 0.053
R5382 S.n12306 S.n12305 0.053
R5383 S.n12026 S.n12025 0.053
R5384 S.n11404 S.n11403 0.053
R5385 S.n11078 S.n11077 0.053
R5386 S.n10787 S.n10786 0.053
R5387 S.n10448 S.n10447 0.053
R5388 S.n10137 S.n10136 0.053
R5389 S.n9788 S.n9787 0.053
R5390 S.n9461 S.n9460 0.053
R5391 S.n9116 S.n9115 0.053
R5392 S.n8594 S.n8593 0.053
R5393 S.n8421 S.n8420 0.053
R5394 S.n7898 S.n7897 0.053
R5395 S.n7714 S.n7713 0.053
R5396 S.n7345 S.n7344 0.053
R5397 S.n6984 S.n6983 0.053
R5398 S.n6599 S.n6598 0.053
R5399 S.n6242 S.n6241 0.053
R5400 S.n5844 S.n5843 0.053
R5401 S.n5477 S.n5476 0.053
R5402 S.n5063 S.n5062 0.053
R5403 S.n4700 S.n4699 0.053
R5404 S.n4264 S.n4263 0.053
R5405 S.n3900 S.n3899 0.053
R5406 S.n3380 S.n3379 0.053
R5407 S.n3088 S.n3087 0.053
R5408 S.n2616 S.n2615 0.053
R5409 S.n2253 S.n2252 0.053
R5410 S.n1765 S.n1764 0.053
R5411 S.n790 S.n789 0.053
R5412 S.n487 S.n486 0.053
R5413 S.n1285 S.n1284 0.053
R5414 S.n9145 S.n9144 0.053
R5415 S.n8498 S.n8497 0.053
R5416 S.n8274 S.n8273 0.053
R5417 S.n7802 S.n7801 0.053
R5418 S.n7567 S.n7566 0.053
R5419 S.n7249 S.n7248 0.053
R5420 S.n6837 S.n6836 0.053
R5421 S.n6503 S.n6502 0.053
R5422 S.n6095 S.n6094 0.053
R5423 S.n5748 S.n5747 0.053
R5424 S.n5330 S.n5329 0.053
R5425 S.n4967 S.n4966 0.053
R5426 S.n4553 S.n4552 0.053
R5427 S.n4168 S.n4167 0.053
R5428 S.n3753 S.n3752 0.053
R5429 S.n3284 S.n3283 0.053
R5430 S.n2941 S.n2940 0.053
R5431 S.n2520 S.n2519 0.053
R5432 S.n2104 S.n2103 0.053
R5433 S.n1664 S.n1663 0.053
R5434 S.n510 S.n509 0.053
R5435 S.n9822 S.n9821 0.053
R5436 S.n9382 S.n9381 0.053
R5437 S.n8998 S.n8997 0.053
R5438 S.n8515 S.n8514 0.053
R5439 S.n8303 S.n8302 0.053
R5440 S.n7819 S.n7818 0.053
R5441 S.n7596 S.n7595 0.053
R5442 S.n7266 S.n7265 0.053
R5443 S.n6866 S.n6865 0.053
R5444 S.n6520 S.n6519 0.053
R5445 S.n6124 S.n6123 0.053
R5446 S.n5765 S.n5764 0.053
R5447 S.n5359 S.n5358 0.053
R5448 S.n4984 S.n4983 0.053
R5449 S.n4582 S.n4581 0.053
R5450 S.n4185 S.n4184 0.053
R5451 S.n3782 S.n3781 0.053
R5452 S.n3301 S.n3300 0.053
R5453 S.n2970 S.n2969 0.053
R5454 S.n2537 S.n2536 0.053
R5455 S.n2133 S.n2132 0.053
R5456 S.n1683 S.n1682 0.053
R5457 S.n1705 S.n1704 0.053
R5458 S.n1347 S.n1346 0.053
R5459 S.n817 S.n816 0.053
R5460 S.n840 S.n839 0.053
R5461 S.n2166 S.n2165 0.053
R5462 S.n3002 S.n3001 0.053
R5463 S.n3814 S.n3813 0.053
R5464 S.n4614 S.n4613 0.053
R5465 S.n5391 S.n5390 0.053
R5466 S.n6156 S.n6155 0.053
R5467 S.n6898 S.n6897 0.053
R5468 S.n7628 S.n7627 0.053
R5469 S.n8335 S.n8334 0.053
R5470 S.n9030 S.n9029 0.053
R5471 S.n9702 S.n9701 0.053
R5472 S.n10480 S.n10479 0.053
R5473 S.n10077 S.n10076 0.053
R5474 S.n9401 S.n9400 0.053
R5475 S.n8534 S.n8533 0.053
R5476 S.n7838 S.n7837 0.053
R5477 S.n7285 S.n7284 0.053
R5478 S.n6539 S.n6538 0.053
R5479 S.n5784 S.n5783 0.053
R5480 S.n5003 S.n5002 0.053
R5481 S.n4204 S.n4203 0.053
R5482 S.n3320 S.n3319 0.053
R5483 S.n2556 S.n2555 0.053
R5484 S.n1381 S.n1380 0.053
R5485 S.n754 S.n753 0.053
R5486 S.n873 S.n872 0.053
R5487 S.n11108 S.n11107 0.053
R5488 S.n10748 S.n10747 0.053
R5489 S.n10396 S.n10395 0.053
R5490 S.n10098 S.n10097 0.053
R5491 S.n9736 S.n9735 0.053
R5492 S.n9422 S.n9421 0.053
R5493 S.n9064 S.n9063 0.053
R5494 S.n8555 S.n8554 0.053
R5495 S.n8369 S.n8368 0.053
R5496 S.n7859 S.n7858 0.053
R5497 S.n7662 S.n7661 0.053
R5498 S.n7306 S.n7305 0.053
R5499 S.n6932 S.n6931 0.053
R5500 S.n6560 S.n6559 0.053
R5501 S.n6190 S.n6189 0.053
R5502 S.n5805 S.n5804 0.053
R5503 S.n5425 S.n5424 0.053
R5504 S.n5024 S.n5023 0.053
R5505 S.n4648 S.n4647 0.053
R5506 S.n4225 S.n4224 0.053
R5507 S.n3848 S.n3847 0.053
R5508 S.n3341 S.n3340 0.053
R5509 S.n3036 S.n3035 0.053
R5510 S.n2577 S.n2576 0.053
R5511 S.n2200 S.n2199 0.053
R5512 S.n1726 S.n1725 0.053
R5513 S.n1409 S.n1408 0.053
R5514 S.n773 S.n772 0.053
R5515 S.n1746 S.n1745 0.053
R5516 S.n2221 S.n2220 0.053
R5517 S.n2597 S.n2596 0.053
R5518 S.n3056 S.n3055 0.053
R5519 S.n3361 S.n3360 0.053
R5520 S.n3868 S.n3867 0.053
R5521 S.n4245 S.n4244 0.053
R5522 S.n4668 S.n4667 0.053
R5523 S.n5044 S.n5043 0.053
R5524 S.n5445 S.n5444 0.053
R5525 S.n5825 S.n5824 0.053
R5526 S.n6210 S.n6209 0.053
R5527 S.n6580 S.n6579 0.053
R5528 S.n6952 S.n6951 0.053
R5529 S.n7326 S.n7325 0.053
R5530 S.n7682 S.n7681 0.053
R5531 S.n7879 S.n7878 0.053
R5532 S.n8389 S.n8388 0.053
R5533 S.n8575 S.n8574 0.053
R5534 S.n9084 S.n9083 0.053
R5535 S.n9442 S.n9441 0.053
R5536 S.n9756 S.n9755 0.053
R5537 S.n10118 S.n10117 0.053
R5538 S.n10416 S.n10415 0.053
R5539 S.n10768 S.n10767 0.053
R5540 S.n11046 S.n11045 0.053
R5541 S.n11385 S.n11384 0.053
R5542 S.n12053 S.n12052 0.053
R5543 S.n902 S.n901 0.053
R5544 S.n1313 S.n1312 0.053
R5545 S.n734 S.n733 0.053
R5546 S.n717 S.n716 0.053
R5547 S.n443 S.n442 0.053
R5548 S.n1226 S.n1225 0.053
R5549 S.n7743 S.n7742 0.053
R5550 S.n7213 S.n7212 0.053
R5551 S.n6776 S.n6775 0.053
R5552 S.n6467 S.n6466 0.053
R5553 S.n6034 S.n6033 0.053
R5554 S.n5712 S.n5711 0.053
R5555 S.n5269 S.n5268 0.053
R5556 S.n4931 S.n4930 0.053
R5557 S.n4492 S.n4491 0.053
R5558 S.n4132 S.n4131 0.053
R5559 S.n3692 S.n3691 0.053
R5560 S.n3248 S.n3247 0.053
R5561 S.n2880 S.n2879 0.053
R5562 S.n2484 S.n2483 0.053
R5563 S.n2043 S.n2042 0.053
R5564 S.n1628 S.n1627 0.053
R5565 S.n469 S.n468 0.053
R5566 S.n8455 S.n8454 0.053
R5567 S.n7783 S.n7782 0.053
R5568 S.n7535 S.n7534 0.053
R5569 S.n7230 S.n7229 0.053
R5570 S.n6805 S.n6804 0.053
R5571 S.n6484 S.n6483 0.053
R5572 S.n6063 S.n6062 0.053
R5573 S.n5729 S.n5728 0.053
R5574 S.n5298 S.n5297 0.053
R5575 S.n4948 S.n4947 0.053
R5576 S.n4521 S.n4520 0.053
R5577 S.n4149 S.n4148 0.053
R5578 S.n3721 S.n3720 0.053
R5579 S.n3265 S.n3264 0.053
R5580 S.n2909 S.n2908 0.053
R5581 S.n2501 S.n2500 0.053
R5582 S.n2072 S.n2071 0.053
R5583 S.n1645 S.n1644 0.053
R5584 S.n1255 S.n1254 0.053
R5585 S.n701 S.n700 0.053
R5586 S.n684 S.n683 0.053
R5587 S.n399 S.n398 0.053
R5588 S.n1167 S.n1166 0.053
R5589 S.n6271 S.n6270 0.053
R5590 S.n5676 S.n5675 0.053
R5591 S.n5208 S.n5207 0.053
R5592 S.n4895 S.n4894 0.053
R5593 S.n4431 S.n4430 0.053
R5594 S.n4096 S.n4095 0.053
R5595 S.n3631 S.n3630 0.053
R5596 S.n3212 S.n3211 0.053
R5597 S.n2819 S.n2818 0.053
R5598 S.n2448 S.n2447 0.053
R5599 S.n1982 S.n1981 0.053
R5600 S.n1592 S.n1591 0.053
R5601 S.n422 S.n421 0.053
R5602 S.n7018 S.n7017 0.053
R5603 S.n6448 S.n6447 0.053
R5604 S.n6002 S.n6001 0.053
R5605 S.n5693 S.n5692 0.053
R5606 S.n5237 S.n5236 0.053
R5607 S.n4912 S.n4911 0.053
R5608 S.n4460 S.n4459 0.053
R5609 S.n4113 S.n4112 0.053
R5610 S.n3660 S.n3659 0.053
R5611 S.n3229 S.n3228 0.053
R5612 S.n2848 S.n2847 0.053
R5613 S.n2465 S.n2464 0.053
R5614 S.n2011 S.n2010 0.053
R5615 S.n1609 S.n1608 0.053
R5616 S.n1196 S.n1195 0.053
R5617 S.n668 S.n667 0.053
R5618 S.n651 S.n650 0.053
R5619 S.n355 S.n354 0.053
R5620 S.n1108 S.n1107 0.053
R5621 S.n4729 S.n4728 0.053
R5622 S.n4060 S.n4059 0.053
R5623 S.n3570 S.n3569 0.053
R5624 S.n3176 S.n3175 0.053
R5625 S.n2758 S.n2757 0.053
R5626 S.n2412 S.n2411 0.053
R5627 S.n1921 S.n1920 0.053
R5628 S.n1556 S.n1555 0.053
R5629 S.n378 S.n377 0.053
R5630 S.n5511 S.n5510 0.053
R5631 S.n4876 S.n4875 0.053
R5632 S.n4399 S.n4398 0.053
R5633 S.n4077 S.n4076 0.053
R5634 S.n3599 S.n3598 0.053
R5635 S.n3193 S.n3192 0.053
R5636 S.n2787 S.n2786 0.053
R5637 S.n2429 S.n2428 0.053
R5638 S.n1936 S.n1935 0.053
R5639 S.n1573 S.n1572 0.053
R5640 S.n1137 S.n1136 0.053
R5641 S.n635 S.n634 0.053
R5642 S.n618 S.n617 0.053
R5643 S.n311 S.n310 0.053
R5644 S.n1049 S.n1048 0.053
R5645 S.n3117 S.n3116 0.053
R5646 S.n2376 S.n2375 0.053
R5647 S.n1860 S.n1859 0.053
R5648 S.n1520 S.n1519 0.053
R5649 S.n334 S.n333 0.053
R5650 S.n3934 S.n3933 0.053
R5651 S.n3157 S.n3156 0.053
R5652 S.n2726 S.n2725 0.053
R5653 S.n2393 S.n2392 0.053
R5654 S.n1889 S.n1888 0.053
R5655 S.n1537 S.n1536 0.053
R5656 S.n1078 S.n1077 0.053
R5657 S.n602 S.n601 0.053
R5658 S.n585 S.n584 0.053
R5659 S.n267 S.n266 0.053
R5660 S.n1461 S.n1460 0.053
R5661 S.n290 S.n289 0.053
R5662 S.n2287 S.n2286 0.053
R5663 S.n1501 S.n1500 0.053
R5664 S.n1019 S.n1018 0.053
R5665 S.n569 S.n568 0.053
R5666 S.n552 S.n551 0.053
R5667 S.n811 S.n810 0.053
R5668 S.n1814 S.n1813 0.053
R5669 S.n1791 S.n1790 0.053
R5670 S.n2324 S.n2323 0.053
R5671 S.n2297 S.n2296 0.053
R5672 S.n3452 S.n3451 0.053
R5673 S.n3425 S.n3424 0.053
R5674 S.n3971 S.n3970 0.053
R5675 S.n3944 S.n3943 0.053
R5676 S.n4766 S.n4765 0.053
R5677 S.n4739 S.n4738 0.053
R5678 S.n5548 S.n5547 0.053
R5679 S.n5521 S.n5520 0.053
R5680 S.n6308 S.n6307 0.053
R5681 S.n6281 S.n6280 0.053
R5682 S.n7055 S.n7054 0.053
R5683 S.n7028 S.n7027 0.053
R5684 S.n8066 S.n8065 0.053
R5685 S.n8039 S.n8038 0.053
R5686 S.n8778 S.n8777 0.053
R5687 S.n8751 S.n8750 0.053
R5688 S.n9182 S.n9181 0.053
R5689 S.n9155 S.n9154 0.053
R5690 S.n9859 S.n9858 0.053
R5691 S.n9832 S.n9831 0.053
R5692 S.n10517 S.n10516 0.053
R5693 S.n10490 S.n10489 0.053
R5694 S.n11145 S.n11144 0.053
R5695 S.n11118 S.n11117 0.053
R5696 S.n12073 S.n12072 0.053
R5697 S.n12350 S.n12349 0.053
R5698 S.n11873 S.n11872 0.053
R5699 S.n1785 S.n1784 0.053
R5700 S.n2657 S.n2656 0.053
R5701 S.n11855 S.n11854 0.053
R5702 S.n12365 S.n12364 0.053
R5703 S.n12089 S.n12088 0.053
R5704 S.n11161 S.n11160 0.053
R5705 S.n11176 S.n11175 0.053
R5706 S.n10533 S.n10532 0.053
R5707 S.n10548 S.n10547 0.053
R5708 S.n9875 S.n9874 0.053
R5709 S.n9890 S.n9889 0.053
R5710 S.n9198 S.n9197 0.053
R5711 S.n9213 S.n9212 0.053
R5712 S.n8794 S.n8793 0.053
R5713 S.n8809 S.n8808 0.053
R5714 S.n8082 S.n8081 0.053
R5715 S.n8097 S.n8096 0.053
R5716 S.n7071 S.n7070 0.053
R5717 S.n7086 S.n7085 0.053
R5718 S.n6324 S.n6323 0.053
R5719 S.n6339 S.n6338 0.053
R5720 S.n5564 S.n5563 0.053
R5721 S.n5579 S.n5578 0.053
R5722 S.n4782 S.n4781 0.053
R5723 S.n4797 S.n4796 0.053
R5724 S.n3987 S.n3986 0.053
R5725 S.n4002 S.n4001 0.053
R5726 S.n3468 S.n3467 0.053
R5727 S.n3483 S.n3482 0.053
R5728 S.n2643 S.n2642 0.053
R5729 S.n2640 S.n2639 0.053
R5730 S.n3498 S.n3497 0.053
R5731 S.n11840 S.n11839 0.053
R5732 S.n12381 S.n12380 0.053
R5733 S.n12104 S.n12103 0.053
R5734 S.n11423 S.n11422 0.053
R5735 S.n11191 S.n11190 0.053
R5736 S.n10807 S.n10806 0.053
R5737 S.n10563 S.n10562 0.053
R5738 S.n10157 S.n10156 0.053
R5739 S.n9905 S.n9904 0.053
R5740 S.n9481 S.n9480 0.053
R5741 S.n9228 S.n9227 0.053
R5742 S.n8614 S.n8613 0.053
R5743 S.n8824 S.n8823 0.053
R5744 S.n7918 S.n7917 0.053
R5745 S.n8112 S.n8111 0.053
R5746 S.n7365 S.n7364 0.053
R5747 S.n7101 S.n7100 0.053
R5748 S.n6619 S.n6618 0.053
R5749 S.n6354 S.n6353 0.053
R5750 S.n5864 S.n5863 0.053
R5751 S.n5594 S.n5593 0.053
R5752 S.n5083 S.n5082 0.053
R5753 S.n4812 S.n4811 0.053
R5754 S.n4284 S.n4283 0.053
R5755 S.n4017 S.n4016 0.053
R5756 S.n3399 S.n3398 0.053
R5757 S.n11825 S.n11824 0.053
R5758 S.n12397 S.n12396 0.053
R5759 S.n12119 S.n12118 0.053
R5760 S.n11439 S.n11438 0.053
R5761 S.n11206 S.n11205 0.053
R5762 S.n10823 S.n10822 0.053
R5763 S.n10578 S.n10577 0.053
R5764 S.n10173 S.n10172 0.053
R5765 S.n9920 S.n9919 0.053
R5766 S.n9497 S.n9496 0.053
R5767 S.n9243 S.n9242 0.053
R5768 S.n8630 S.n8629 0.053
R5769 S.n8839 S.n8838 0.053
R5770 S.n7934 S.n7933 0.053
R5771 S.n8127 S.n8126 0.053
R5772 S.n7381 S.n7380 0.053
R5773 S.n7116 S.n7115 0.053
R5774 S.n6635 S.n6634 0.053
R5775 S.n6369 S.n6368 0.053
R5776 S.n5880 S.n5879 0.053
R5777 S.n5609 S.n5608 0.053
R5778 S.n5099 S.n5098 0.053
R5779 S.n4827 S.n4826 0.053
R5780 S.n4310 S.n4309 0.053
R5781 S.n4330 S.n4329 0.053
R5782 S.n3419 S.n3418 0.053
R5783 S.n4304 S.n4303 0.053
R5784 S.n5136 S.n5135 0.053
R5785 S.n11810 S.n11809 0.053
R5786 S.n12413 S.n12412 0.053
R5787 S.n12134 S.n12133 0.053
R5788 S.n11455 S.n11454 0.053
R5789 S.n11221 S.n11220 0.053
R5790 S.n10839 S.n10838 0.053
R5791 S.n10593 S.n10592 0.053
R5792 S.n10189 S.n10188 0.053
R5793 S.n9935 S.n9934 0.053
R5794 S.n9513 S.n9512 0.053
R5795 S.n9258 S.n9257 0.053
R5796 S.n8646 S.n8645 0.053
R5797 S.n8854 S.n8853 0.053
R5798 S.n7950 S.n7949 0.053
R5799 S.n8142 S.n8141 0.053
R5800 S.n7397 S.n7396 0.053
R5801 S.n7131 S.n7130 0.053
R5802 S.n6651 S.n6650 0.053
R5803 S.n6384 S.n6383 0.053
R5804 S.n5896 S.n5895 0.053
R5805 S.n5624 S.n5623 0.053
R5806 S.n5122 S.n5121 0.053
R5807 S.n5119 S.n5118 0.053
R5808 S.n5933 S.n5932 0.053
R5809 S.n11795 S.n11794 0.053
R5810 S.n12429 S.n12428 0.053
R5811 S.n12149 S.n12148 0.053
R5812 S.n11471 S.n11470 0.053
R5813 S.n11236 S.n11235 0.053
R5814 S.n10855 S.n10854 0.053
R5815 S.n10608 S.n10607 0.053
R5816 S.n10205 S.n10204 0.053
R5817 S.n9950 S.n9949 0.053
R5818 S.n9529 S.n9528 0.053
R5819 S.n9273 S.n9272 0.053
R5820 S.n8662 S.n8661 0.053
R5821 S.n8869 S.n8868 0.053
R5822 S.n7966 S.n7965 0.053
R5823 S.n8157 S.n8156 0.053
R5824 S.n7413 S.n7412 0.053
R5825 S.n7146 S.n7145 0.053
R5826 S.n6667 S.n6666 0.053
R5827 S.n6399 S.n6398 0.053
R5828 S.n5919 S.n5918 0.053
R5829 S.n5916 S.n5915 0.053
R5830 S.n6704 S.n6703 0.053
R5831 S.n11780 S.n11779 0.053
R5832 S.n12445 S.n12444 0.053
R5833 S.n12164 S.n12163 0.053
R5834 S.n11487 S.n11486 0.053
R5835 S.n11251 S.n11250 0.053
R5836 S.n10871 S.n10870 0.053
R5837 S.n10623 S.n10622 0.053
R5838 S.n10221 S.n10220 0.053
R5839 S.n9965 S.n9964 0.053
R5840 S.n9545 S.n9544 0.053
R5841 S.n9288 S.n9287 0.053
R5842 S.n8678 S.n8677 0.053
R5843 S.n8884 S.n8883 0.053
R5844 S.n7982 S.n7981 0.053
R5845 S.n8172 S.n8171 0.053
R5846 S.n7429 S.n7428 0.053
R5847 S.n7161 S.n7160 0.053
R5848 S.n6690 S.n6689 0.053
R5849 S.n6687 S.n6686 0.053
R5850 S.n7466 S.n7465 0.053
R5851 S.n11765 S.n11764 0.053
R5852 S.n12461 S.n12460 0.053
R5853 S.n12179 S.n12178 0.053
R5854 S.n11503 S.n11502 0.053
R5855 S.n11266 S.n11265 0.053
R5856 S.n10887 S.n10886 0.053
R5857 S.n10638 S.n10637 0.053
R5858 S.n10237 S.n10236 0.053
R5859 S.n9980 S.n9979 0.053
R5860 S.n9561 S.n9560 0.053
R5861 S.n9303 S.n9302 0.053
R5862 S.n8694 S.n8693 0.053
R5863 S.n8899 S.n8898 0.053
R5864 S.n7998 S.n7997 0.053
R5865 S.n8187 S.n8186 0.053
R5866 S.n7452 S.n7451 0.053
R5867 S.n7449 S.n7448 0.053
R5868 S.n8202 S.n8201 0.053
R5869 S.n11750 S.n11749 0.053
R5870 S.n12477 S.n12476 0.053
R5871 S.n12194 S.n12193 0.053
R5872 S.n11519 S.n11518 0.053
R5873 S.n11281 S.n11280 0.053
R5874 S.n10903 S.n10902 0.053
R5875 S.n10653 S.n10652 0.053
R5876 S.n10253 S.n10252 0.053
R5877 S.n9995 S.n9994 0.053
R5878 S.n9577 S.n9576 0.053
R5879 S.n9318 S.n9317 0.053
R5880 S.n8710 S.n8709 0.053
R5881 S.n8914 S.n8913 0.053
R5882 S.n8013 S.n8012 0.053
R5883 S.n8033 S.n8032 0.053
R5884 S.n8929 S.n8928 0.053
R5885 S.n11735 S.n11734 0.053
R5886 S.n12493 S.n12492 0.053
R5887 S.n12209 S.n12208 0.053
R5888 S.n11535 S.n11534 0.053
R5889 S.n11296 S.n11295 0.053
R5890 S.n10919 S.n10918 0.053
R5891 S.n10668 S.n10667 0.053
R5892 S.n10269 S.n10268 0.053
R5893 S.n10010 S.n10009 0.053
R5894 S.n9593 S.n9592 0.053
R5895 S.n9333 S.n9332 0.053
R5896 S.n8725 S.n8724 0.053
R5897 S.n8745 S.n8744 0.053
R5898 S.n9630 S.n9629 0.053
R5899 S.n11720 S.n11719 0.053
R5900 S.n12509 S.n12508 0.053
R5901 S.n12224 S.n12223 0.053
R5902 S.n11551 S.n11550 0.053
R5903 S.n11311 S.n11310 0.053
R5904 S.n10935 S.n10934 0.053
R5905 S.n10683 S.n10682 0.053
R5906 S.n10285 S.n10284 0.053
R5907 S.n10025 S.n10024 0.053
R5908 S.n9616 S.n9615 0.053
R5909 S.n9613 S.n9612 0.053
R5910 S.n10322 S.n10321 0.053
R5911 S.n11705 S.n11704 0.053
R5912 S.n12525 S.n12524 0.053
R5913 S.n12239 S.n12238 0.053
R5914 S.n11567 S.n11566 0.053
R5915 S.n11326 S.n11325 0.053
R5916 S.n10951 S.n10950 0.053
R5917 S.n10698 S.n10697 0.053
R5918 S.n10308 S.n10307 0.053
R5919 S.n10305 S.n10304 0.053
R5920 S.n10988 S.n10987 0.053
R5921 S.n11690 S.n11689 0.053
R5922 S.n12541 S.n12540 0.053
R5923 S.n12254 S.n12253 0.053
R5924 S.n11583 S.n11582 0.053
R5925 S.n11341 S.n11340 0.053
R5926 S.n10974 S.n10973 0.053
R5927 S.n10971 S.n10970 0.053
R5928 S.n11623 S.n11622 0.053
R5929 S.n11675 S.n11674 0.053
R5930 S.n12557 S.n12556 0.053
R5931 S.n12269 S.n12268 0.053
R5932 S.n11609 S.n11608 0.053
R5933 S.n11606 S.n11605 0.053
R5934 S.n12588 S.n12587 0.053
R5935 S.n11660 S.n11659 0.053
R5936 S.n12563 S.n12562 0.053
R5937 S.n993 S.n992 0.052
R5938 S.n2688 S.n2687 0.052
R5939 S.n1831 S.n1830 0.052
R5940 S.n3529 S.n3528 0.052
R5941 S.n4361 S.n4360 0.052
R5942 S.n3541 S.n3540 0.052
R5943 S.n5167 S.n5166 0.052
R5944 S.n4373 S.n4372 0.052
R5945 S.n5964 S.n5963 0.052
R5946 S.n5179 S.n5178 0.052
R5947 S.n6735 S.n6734 0.052
R5948 S.n5976 S.n5975 0.052
R5949 S.n7497 S.n7496 0.052
R5950 S.n6747 S.n6746 0.052
R5951 S.n8233 S.n8232 0.052
R5952 S.n7509 S.n7508 0.052
R5953 S.n8960 S.n8959 0.052
R5954 S.n8245 S.n8244 0.052
R5955 S.n9661 S.n9660 0.052
R5956 S.n8972 S.n8971 0.052
R5957 S.n10353 S.n10352 0.052
R5958 S.n9673 S.n9672 0.052
R5959 S.n11017 S.n11016 0.052
R5960 S.n10365 S.n10364 0.052
R5961 S.n11029 S.n11028 0.052
R5962 S.n12609 S.n12608 0.052
R5963 S.n12322 S.n12321 0.052
R5964 S.n2700 S.n2699 0.052
R5965 S.n11994 S.n11924 0.052
R5966 S.n824 S.n823 0.051
R5967 S.n10472 S.n10470 0.051
R5968 S.n9795 S.n9794 0.051
R5969 S.n9137 S.n9135 0.051
R5970 S.n8428 S.n8427 0.051
R5971 S.n7735 S.n7733 0.051
R5972 S.n6991 S.n6990 0.051
R5973 S.n6263 S.n6261 0.051
R5974 S.n5484 S.n5483 0.051
R5975 S.n4721 S.n4719 0.051
R5976 S.n3907 S.n3906 0.051
R5977 S.n3109 S.n3107 0.051
R5978 S.n2260 S.n2259 0.051
R5979 S.n1453 S.n1451 0.051
R5980 S.n929 S.n928 0.051
R5981 S.n967 S.n966 0.051
R5982 S.n965 S.n964 0.051
R5983 S.n10474 S.n10473 0.05
R5984 S.n12047 S.n12034 0.05
R5985 S.n891 S.n890 0.05
R5986 S.n9811 S.n9810 0.05
R5987 S.n9816 S.n9797 0.05
R5988 S.n9139 S.n9138 0.05
R5989 S.n8446 S.n8443 0.05
R5990 S.n8449 S.n8430 0.05
R5991 S.n7737 S.n7736 0.05
R5992 S.n7009 S.n7006 0.05
R5993 S.n7012 S.n6993 0.05
R5994 S.n6265 S.n6264 0.05
R5995 S.n5500 S.n5499 0.05
R5996 S.n5505 S.n5486 0.05
R5997 S.n4723 S.n4722 0.05
R5998 S.n3925 S.n3922 0.05
R5999 S.n3928 S.n3909 0.05
R6000 S.n3111 S.n3110 0.05
R6001 S.n2276 S.n2275 0.05
R6002 S.n2281 S.n2262 0.05
R6003 S.n1455 S.n1454 0.05
R6004 S.n950 S.n931 0.05
R6005 S.n910 S.n909 0.05
R6006 S.n1715 S.n1714 0.049
R6007 S.n2566 S.n2565 0.049
R6008 S.n3330 S.n3329 0.049
R6009 S.n4214 S.n4213 0.049
R6010 S.n5013 S.n5012 0.049
R6011 S.n5794 S.n5793 0.049
R6012 S.n6549 S.n6548 0.049
R6013 S.n7295 S.n7294 0.049
R6014 S.n7848 S.n7847 0.049
R6015 S.n8544 S.n8543 0.049
R6016 S.n9411 S.n9410 0.049
R6017 S.n10087 S.n10086 0.049
R6018 S.n10737 S.n10736 0.049
R6019 S.n748 S.n747 0.049
R6020 S.n767 S.n766 0.049
R6021 S.n11642 S.n11640 0.049
R6022 S.n11599 S.n11598 0.048
R6023 S.n991 S.n990 0.048
R6024 S.n2676 S.n2675 0.048
R6025 S.n3517 S.n3516 0.048
R6026 S.n4349 S.n4348 0.048
R6027 S.n5155 S.n5154 0.048
R6028 S.n5952 S.n5951 0.048
R6029 S.n6723 S.n6722 0.048
R6030 S.n7485 S.n7484 0.048
R6031 S.n8221 S.n8220 0.048
R6032 S.n8948 S.n8947 0.048
R6033 S.n9649 S.n9648 0.048
R6034 S.n10341 S.n10340 0.048
R6035 S.n11005 S.n11004 0.048
R6036 S.n11639 S.n11638 0.048
R6037 S.n11911 S.n11909 0.047
R6038 S.n12327 S.n12318 0.047
R6039 S.n12611 S.n12595 0.047
R6040 S.n950 S.n941 0.047
R6041 S.n920 S.n918 0.047
R6042 S.n1431 S.n1417 0.047
R6043 S.n11891 S.n11883 0.047
R6044 S.n12303 S.n12295 0.047
R6045 S.n12023 S.n12011 0.047
R6046 S.n11401 S.n11393 0.047
R6047 S.n11075 S.n11063 0.047
R6048 S.n10784 S.n10776 0.047
R6049 S.n10445 S.n10433 0.047
R6050 S.n10134 S.n10126 0.047
R6051 S.n9785 S.n9773 0.047
R6052 S.n9458 S.n9450 0.047
R6053 S.n9113 S.n9101 0.047
R6054 S.n8591 S.n8583 0.047
R6055 S.n8418 S.n8406 0.047
R6056 S.n7895 S.n7887 0.047
R6057 S.n7711 S.n7699 0.047
R6058 S.n7342 S.n7334 0.047
R6059 S.n6981 S.n6969 0.047
R6060 S.n6596 S.n6588 0.047
R6061 S.n6239 S.n6227 0.047
R6062 S.n5841 S.n5833 0.047
R6063 S.n5474 S.n5462 0.047
R6064 S.n5060 S.n5052 0.047
R6065 S.n4697 S.n4685 0.047
R6066 S.n4261 S.n4253 0.047
R6067 S.n3897 S.n3885 0.047
R6068 S.n3377 S.n3369 0.047
R6069 S.n3085 S.n3073 0.047
R6070 S.n2613 S.n2605 0.047
R6071 S.n2250 S.n2238 0.047
R6072 S.n1762 S.n1754 0.047
R6073 S.n787 S.n785 0.047
R6074 S.n484 S.n482 0.047
R6075 S.n1282 S.n1272 0.047
R6076 S.n9139 S.n9125 0.047
R6077 S.n8495 S.n8487 0.047
R6078 S.n8271 S.n8259 0.047
R6079 S.n7799 S.n7791 0.047
R6080 S.n7564 S.n7552 0.047
R6081 S.n7246 S.n7238 0.047
R6082 S.n6834 S.n6822 0.047
R6083 S.n6500 S.n6492 0.047
R6084 S.n6092 S.n6080 0.047
R6085 S.n5745 S.n5737 0.047
R6086 S.n5327 S.n5315 0.047
R6087 S.n4964 S.n4956 0.047
R6088 S.n4550 S.n4538 0.047
R6089 S.n4165 S.n4157 0.047
R6090 S.n3750 S.n3738 0.047
R6091 S.n3281 S.n3273 0.047
R6092 S.n2938 S.n2926 0.047
R6093 S.n2517 S.n2509 0.047
R6094 S.n2101 S.n2089 0.047
R6095 S.n1661 S.n1653 0.047
R6096 S.n507 S.n505 0.047
R6097 S.n9816 S.n9807 0.047
R6098 S.n9379 S.n9377 0.047
R6099 S.n8995 S.n8984 0.047
R6100 S.n8512 S.n8510 0.047
R6101 S.n8300 S.n8289 0.047
R6102 S.n7816 S.n7814 0.047
R6103 S.n7593 S.n7582 0.047
R6104 S.n7263 S.n7261 0.047
R6105 S.n6863 S.n6852 0.047
R6106 S.n6517 S.n6515 0.047
R6107 S.n6121 S.n6110 0.047
R6108 S.n5762 S.n5760 0.047
R6109 S.n5356 S.n5345 0.047
R6110 S.n4981 S.n4979 0.047
R6111 S.n4579 S.n4568 0.047
R6112 S.n4182 S.n4180 0.047
R6113 S.n3779 S.n3768 0.047
R6114 S.n3298 S.n3296 0.047
R6115 S.n2967 S.n2956 0.047
R6116 S.n2534 S.n2532 0.047
R6117 S.n2130 S.n2119 0.047
R6118 S.n1680 S.n1676 0.047
R6119 S.n1702 S.n1697 0.047
R6120 S.n1344 S.n1329 0.047
R6121 S.n822 S.n820 0.047
R6122 S.n837 S.n831 0.047
R6123 S.n2163 S.n2151 0.047
R6124 S.n2999 S.n2987 0.047
R6125 S.n3811 S.n3799 0.047
R6126 S.n4611 S.n4599 0.047
R6127 S.n5388 S.n5376 0.047
R6128 S.n6153 S.n6141 0.047
R6129 S.n6895 S.n6883 0.047
R6130 S.n7625 S.n7613 0.047
R6131 S.n8332 S.n8320 0.047
R6132 S.n9027 S.n9015 0.047
R6133 S.n9699 S.n9687 0.047
R6134 S.n10474 S.n10460 0.047
R6135 S.n10074 S.n10066 0.047
R6136 S.n9398 S.n9390 0.047
R6137 S.n8531 S.n8523 0.047
R6138 S.n7835 S.n7827 0.047
R6139 S.n7282 S.n7274 0.047
R6140 S.n6536 S.n6528 0.047
R6141 S.n5781 S.n5773 0.047
R6142 S.n5000 S.n4992 0.047
R6143 S.n4201 S.n4193 0.047
R6144 S.n3317 S.n3309 0.047
R6145 S.n2553 S.n2545 0.047
R6146 S.n1378 S.n1368 0.047
R6147 S.n751 S.n745 0.047
R6148 S.n870 S.n863 0.047
R6149 S.n11102 S.n11094 0.047
R6150 S.n10745 S.n10740 0.047
R6151 S.n10393 S.n10378 0.047
R6152 S.n10095 S.n10090 0.047
R6153 S.n9733 S.n9718 0.047
R6154 S.n9419 S.n9414 0.047
R6155 S.n9061 S.n9046 0.047
R6156 S.n8552 S.n8547 0.047
R6157 S.n8366 S.n8351 0.047
R6158 S.n7856 S.n7851 0.047
R6159 S.n7659 S.n7644 0.047
R6160 S.n7303 S.n7298 0.047
R6161 S.n6929 S.n6914 0.047
R6162 S.n6557 S.n6552 0.047
R6163 S.n6187 S.n6172 0.047
R6164 S.n5802 S.n5797 0.047
R6165 S.n5422 S.n5407 0.047
R6166 S.n5021 S.n5016 0.047
R6167 S.n4645 S.n4630 0.047
R6168 S.n4222 S.n4217 0.047
R6169 S.n3845 S.n3830 0.047
R6170 S.n3338 S.n3333 0.047
R6171 S.n3033 S.n3018 0.047
R6172 S.n2574 S.n2569 0.047
R6173 S.n2197 S.n2182 0.047
R6174 S.n1723 S.n1718 0.047
R6175 S.n1406 S.n1396 0.047
R6176 S.n770 S.n765 0.047
R6177 S.n1743 S.n1737 0.047
R6178 S.n2218 S.n2215 0.047
R6179 S.n2594 S.n2589 0.047
R6180 S.n3053 S.n3051 0.047
R6181 S.n3358 S.n3353 0.047
R6182 S.n3865 S.n3863 0.047
R6183 S.n4242 S.n4237 0.047
R6184 S.n4665 S.n4663 0.047
R6185 S.n5041 S.n5036 0.047
R6186 S.n5442 S.n5440 0.047
R6187 S.n5822 S.n5817 0.047
R6188 S.n6207 S.n6205 0.047
R6189 S.n6577 S.n6572 0.047
R6190 S.n6949 S.n6947 0.047
R6191 S.n7323 S.n7318 0.047
R6192 S.n7679 S.n7677 0.047
R6193 S.n7876 S.n7871 0.047
R6194 S.n8386 S.n8384 0.047
R6195 S.n8572 S.n8567 0.047
R6196 S.n9081 S.n9079 0.047
R6197 S.n9439 S.n9434 0.047
R6198 S.n9753 S.n9751 0.047
R6199 S.n10115 S.n10110 0.047
R6200 S.n10413 S.n10411 0.047
R6201 S.n10765 S.n10760 0.047
R6202 S.n11043 S.n11041 0.047
R6203 S.n11382 S.n11377 0.047
R6204 S.n12047 S.n12045 0.047
R6205 S.n899 S.n889 0.047
R6206 S.n1310 S.n1300 0.047
R6207 S.n731 S.n729 0.047
R6208 S.n714 S.n712 0.047
R6209 S.n440 S.n438 0.047
R6210 S.n1223 S.n1213 0.047
R6211 S.n7737 S.n7723 0.047
R6212 S.n7210 S.n7202 0.047
R6213 S.n6773 S.n6761 0.047
R6214 S.n6464 S.n6456 0.047
R6215 S.n6031 S.n6019 0.047
R6216 S.n5709 S.n5701 0.047
R6217 S.n5266 S.n5254 0.047
R6218 S.n4928 S.n4920 0.047
R6219 S.n4489 S.n4477 0.047
R6220 S.n4129 S.n4121 0.047
R6221 S.n3689 S.n3677 0.047
R6222 S.n3245 S.n3237 0.047
R6223 S.n2877 S.n2865 0.047
R6224 S.n2481 S.n2473 0.047
R6225 S.n2040 S.n2028 0.047
R6226 S.n1625 S.n1617 0.047
R6227 S.n466 S.n464 0.047
R6228 S.n8449 S.n8440 0.047
R6229 S.n7780 S.n7778 0.047
R6230 S.n7532 S.n7521 0.047
R6231 S.n7227 S.n7225 0.047
R6232 S.n6802 S.n6791 0.047
R6233 S.n6481 S.n6479 0.047
R6234 S.n6060 S.n6049 0.047
R6235 S.n5726 S.n5724 0.047
R6236 S.n5295 S.n5284 0.047
R6237 S.n4945 S.n4943 0.047
R6238 S.n4518 S.n4507 0.047
R6239 S.n4146 S.n4144 0.047
R6240 S.n3718 S.n3707 0.047
R6241 S.n3262 S.n3260 0.047
R6242 S.n2906 S.n2895 0.047
R6243 S.n2498 S.n2496 0.047
R6244 S.n2069 S.n2058 0.047
R6245 S.n1642 S.n1640 0.047
R6246 S.n1252 S.n1241 0.047
R6247 S.n698 S.n696 0.047
R6248 S.n681 S.n679 0.047
R6249 S.n396 S.n394 0.047
R6250 S.n1164 S.n1154 0.047
R6251 S.n6265 S.n6251 0.047
R6252 S.n5673 S.n5665 0.047
R6253 S.n5205 S.n5193 0.047
R6254 S.n4892 S.n4884 0.047
R6255 S.n4428 S.n4416 0.047
R6256 S.n4093 S.n4085 0.047
R6257 S.n3628 S.n3616 0.047
R6258 S.n3209 S.n3201 0.047
R6259 S.n2816 S.n2804 0.047
R6260 S.n2445 S.n2437 0.047
R6261 S.n1979 S.n1967 0.047
R6262 S.n1589 S.n1581 0.047
R6263 S.n419 S.n417 0.047
R6264 S.n7012 S.n7003 0.047
R6265 S.n6445 S.n6443 0.047
R6266 S.n5999 S.n5988 0.047
R6267 S.n5690 S.n5688 0.047
R6268 S.n5234 S.n5223 0.047
R6269 S.n4909 S.n4907 0.047
R6270 S.n4457 S.n4446 0.047
R6271 S.n4110 S.n4108 0.047
R6272 S.n3657 S.n3646 0.047
R6273 S.n3226 S.n3224 0.047
R6274 S.n2845 S.n2834 0.047
R6275 S.n2462 S.n2460 0.047
R6276 S.n2008 S.n1997 0.047
R6277 S.n1606 S.n1604 0.047
R6278 S.n1193 S.n1182 0.047
R6279 S.n665 S.n663 0.047
R6280 S.n648 S.n646 0.047
R6281 S.n352 S.n350 0.047
R6282 S.n1105 S.n1095 0.047
R6283 S.n4723 S.n4709 0.047
R6284 S.n4057 S.n4049 0.047
R6285 S.n3567 S.n3555 0.047
R6286 S.n3173 S.n3165 0.047
R6287 S.n2755 S.n2743 0.047
R6288 S.n2409 S.n2401 0.047
R6289 S.n1918 S.n1906 0.047
R6290 S.n1553 S.n1545 0.047
R6291 S.n375 S.n373 0.047
R6292 S.n5505 S.n5496 0.047
R6293 S.n4873 S.n4871 0.047
R6294 S.n4396 S.n4385 0.047
R6295 S.n4074 S.n4072 0.047
R6296 S.n3596 S.n3585 0.047
R6297 S.n3190 S.n3188 0.047
R6298 S.n2784 S.n2773 0.047
R6299 S.n2426 S.n2424 0.047
R6300 S.n1950 S.n1939 0.047
R6301 S.n1570 S.n1568 0.047
R6302 S.n1134 S.n1123 0.047
R6303 S.n632 S.n630 0.047
R6304 S.n615 S.n613 0.047
R6305 S.n308 S.n306 0.047
R6306 S.n1046 S.n1036 0.047
R6307 S.n3111 S.n3097 0.047
R6308 S.n2373 S.n2365 0.047
R6309 S.n1857 S.n1845 0.047
R6310 S.n1517 S.n1509 0.047
R6311 S.n331 S.n329 0.047
R6312 S.n3928 S.n3919 0.047
R6313 S.n3154 S.n3152 0.047
R6314 S.n2723 S.n2712 0.047
R6315 S.n2390 S.n2388 0.047
R6316 S.n1886 S.n1875 0.047
R6317 S.n1534 S.n1532 0.047
R6318 S.n1075 S.n1064 0.047
R6319 S.n599 S.n597 0.047
R6320 S.n582 S.n580 0.047
R6321 S.n264 S.n262 0.047
R6322 S.n1455 S.n1443 0.047
R6323 S.n287 S.n285 0.047
R6324 S.n2281 S.n2272 0.047
R6325 S.n1498 S.n1496 0.047
R6326 S.n1016 S.n1005 0.047
R6327 S.n566 S.n564 0.047
R6328 S.n549 S.n547 0.047
R6329 S.n980 S.n963 0.047
R6330 S.n805 S.n802 0.047
R6331 S.n1808 S.n1805 0.047
R6332 S.n1798 S.n1794 0.047
R6333 S.n2318 S.n2312 0.047
R6334 S.n2304 S.n2300 0.047
R6335 S.n3446 S.n3440 0.047
R6336 S.n3432 S.n3428 0.047
R6337 S.n3965 S.n3959 0.047
R6338 S.n3951 S.n3947 0.047
R6339 S.n4760 S.n4754 0.047
R6340 S.n4746 S.n4742 0.047
R6341 S.n5542 S.n5536 0.047
R6342 S.n5528 S.n5524 0.047
R6343 S.n6302 S.n6296 0.047
R6344 S.n6288 S.n6284 0.047
R6345 S.n7049 S.n7043 0.047
R6346 S.n7035 S.n7031 0.047
R6347 S.n8060 S.n8054 0.047
R6348 S.n8046 S.n8042 0.047
R6349 S.n8772 S.n8766 0.047
R6350 S.n8758 S.n8754 0.047
R6351 S.n9176 S.n9170 0.047
R6352 S.n9162 S.n9158 0.047
R6353 S.n9853 S.n9847 0.047
R6354 S.n9839 S.n9835 0.047
R6355 S.n10511 S.n10505 0.047
R6356 S.n10497 S.n10493 0.047
R6357 S.n11139 S.n11133 0.047
R6358 S.n11125 S.n11121 0.047
R6359 S.n12067 S.n12061 0.047
R6360 S.n12344 S.n12340 0.047
R6361 S.n11870 S.n11865 0.047
R6362 S.n1826 S.n1821 0.047
R6363 S.n1779 S.n1777 0.047
R6364 S.n2651 S.n2329 0.047
R6365 S.n11852 S.n11848 0.047
R6366 S.n12359 S.n12355 0.047
R6367 S.n12083 S.n12078 0.047
R6368 S.n11168 S.n11158 0.047
R6369 S.n11170 S.n11150 0.047
R6370 S.n10540 S.n10530 0.047
R6371 S.n10542 S.n10522 0.047
R6372 S.n9882 S.n9872 0.047
R6373 S.n9884 S.n9864 0.047
R6374 S.n9205 S.n9195 0.047
R6375 S.n9207 S.n9187 0.047
R6376 S.n8801 S.n8791 0.047
R6377 S.n8803 S.n8783 0.047
R6378 S.n8089 S.n8079 0.047
R6379 S.n8091 S.n8071 0.047
R6380 S.n7078 S.n7068 0.047
R6381 S.n7080 S.n7060 0.047
R6382 S.n6331 S.n6321 0.047
R6383 S.n6333 S.n6313 0.047
R6384 S.n5571 S.n5561 0.047
R6385 S.n5573 S.n5553 0.047
R6386 S.n4789 S.n4779 0.047
R6387 S.n4791 S.n4771 0.047
R6388 S.n3994 S.n3984 0.047
R6389 S.n3996 S.n3976 0.047
R6390 S.n3475 S.n3465 0.047
R6391 S.n3477 S.n3457 0.047
R6392 S.n2650 S.n2337 0.047
R6393 S.n2696 S.n2664 0.047
R6394 S.n2634 S.n2628 0.047
R6395 S.n3492 S.n3488 0.047
R6396 S.n11837 S.n11833 0.047
R6397 S.n12375 S.n12370 0.047
R6398 S.n12098 S.n12094 0.047
R6399 S.n11417 S.n11412 0.047
R6400 S.n11185 S.n11181 0.047
R6401 S.n10801 S.n10796 0.047
R6402 S.n10557 S.n10553 0.047
R6403 S.n10151 S.n10146 0.047
R6404 S.n9899 S.n9895 0.047
R6405 S.n9475 S.n9470 0.047
R6406 S.n9222 S.n9218 0.047
R6407 S.n8608 S.n8603 0.047
R6408 S.n8818 S.n8814 0.047
R6409 S.n7912 S.n7907 0.047
R6410 S.n8106 S.n8102 0.047
R6411 S.n7359 S.n7354 0.047
R6412 S.n7095 S.n7091 0.047
R6413 S.n6613 S.n6608 0.047
R6414 S.n6348 S.n6344 0.047
R6415 S.n5858 S.n5853 0.047
R6416 S.n5588 S.n5584 0.047
R6417 S.n5077 S.n5072 0.047
R6418 S.n4806 S.n4802 0.047
R6419 S.n4278 S.n4273 0.047
R6420 S.n4011 S.n4007 0.047
R6421 S.n3393 S.n3389 0.047
R6422 S.n11822 S.n11820 0.047
R6423 S.n12391 S.n12389 0.047
R6424 S.n12113 S.n12111 0.047
R6425 S.n11433 S.n11431 0.047
R6426 S.n11200 S.n11198 0.047
R6427 S.n10817 S.n10815 0.047
R6428 S.n10572 S.n10570 0.047
R6429 S.n10167 S.n10165 0.047
R6430 S.n9914 S.n9912 0.047
R6431 S.n9491 S.n9489 0.047
R6432 S.n9237 S.n9235 0.047
R6433 S.n8624 S.n8622 0.047
R6434 S.n8833 S.n8831 0.047
R6435 S.n7928 S.n7926 0.047
R6436 S.n8121 S.n8119 0.047
R6437 S.n7375 S.n7373 0.047
R6438 S.n7110 S.n7108 0.047
R6439 S.n6629 S.n6627 0.047
R6440 S.n6363 S.n6361 0.047
R6441 S.n5874 S.n5872 0.047
R6442 S.n5603 S.n5601 0.047
R6443 S.n5093 S.n5091 0.047
R6444 S.n4821 S.n4819 0.047
R6445 S.n4315 S.n4313 0.047
R6446 S.n4324 S.n4322 0.047
R6447 S.n3413 S.n3407 0.047
R6448 S.n3537 S.n3505 0.047
R6449 S.n4369 S.n4337 0.047
R6450 S.n4298 S.n4292 0.047
R6451 S.n5130 S.n4832 0.047
R6452 S.n11807 S.n11803 0.047
R6453 S.n12407 S.n12402 0.047
R6454 S.n12128 S.n12124 0.047
R6455 S.n11449 S.n11444 0.047
R6456 S.n11215 S.n11211 0.047
R6457 S.n10833 S.n10828 0.047
R6458 S.n10587 S.n10583 0.047
R6459 S.n10183 S.n10178 0.047
R6460 S.n9929 S.n9925 0.047
R6461 S.n9507 S.n9502 0.047
R6462 S.n9252 S.n9248 0.047
R6463 S.n8640 S.n8635 0.047
R6464 S.n8848 S.n8844 0.047
R6465 S.n7944 S.n7939 0.047
R6466 S.n8136 S.n8132 0.047
R6467 S.n7391 S.n7386 0.047
R6468 S.n7125 S.n7121 0.047
R6469 S.n6645 S.n6640 0.047
R6470 S.n6378 S.n6374 0.047
R6471 S.n5890 S.n5885 0.047
R6472 S.n5618 S.n5614 0.047
R6473 S.n5129 S.n4840 0.047
R6474 S.n5175 S.n5143 0.047
R6475 S.n5113 S.n5107 0.047
R6476 S.n5927 S.n5629 0.047
R6477 S.n11792 S.n11788 0.047
R6478 S.n12423 S.n12418 0.047
R6479 S.n12143 S.n12139 0.047
R6480 S.n11465 S.n11460 0.047
R6481 S.n11230 S.n11226 0.047
R6482 S.n10849 S.n10844 0.047
R6483 S.n10602 S.n10598 0.047
R6484 S.n10199 S.n10194 0.047
R6485 S.n9944 S.n9940 0.047
R6486 S.n9523 S.n9518 0.047
R6487 S.n9267 S.n9263 0.047
R6488 S.n8656 S.n8651 0.047
R6489 S.n8863 S.n8859 0.047
R6490 S.n7960 S.n7955 0.047
R6491 S.n8151 S.n8147 0.047
R6492 S.n7407 S.n7402 0.047
R6493 S.n7140 S.n7136 0.047
R6494 S.n6661 S.n6656 0.047
R6495 S.n6393 S.n6389 0.047
R6496 S.n5926 S.n5637 0.047
R6497 S.n5972 S.n5940 0.047
R6498 S.n5910 S.n5904 0.047
R6499 S.n6698 S.n6404 0.047
R6500 S.n11777 S.n11773 0.047
R6501 S.n12439 S.n12434 0.047
R6502 S.n12158 S.n12154 0.047
R6503 S.n11481 S.n11476 0.047
R6504 S.n11245 S.n11241 0.047
R6505 S.n10865 S.n10860 0.047
R6506 S.n10617 S.n10613 0.047
R6507 S.n10215 S.n10210 0.047
R6508 S.n9959 S.n9955 0.047
R6509 S.n9539 S.n9534 0.047
R6510 S.n9282 S.n9278 0.047
R6511 S.n8672 S.n8667 0.047
R6512 S.n8878 S.n8874 0.047
R6513 S.n7976 S.n7971 0.047
R6514 S.n8166 S.n8162 0.047
R6515 S.n7423 S.n7418 0.047
R6516 S.n7155 S.n7151 0.047
R6517 S.n6697 S.n6412 0.047
R6518 S.n6743 S.n6711 0.047
R6519 S.n6681 S.n6675 0.047
R6520 S.n7460 S.n7166 0.047
R6521 S.n11762 S.n11758 0.047
R6522 S.n12455 S.n12450 0.047
R6523 S.n12173 S.n12169 0.047
R6524 S.n11497 S.n11492 0.047
R6525 S.n11260 S.n11256 0.047
R6526 S.n10881 S.n10876 0.047
R6527 S.n10632 S.n10628 0.047
R6528 S.n10231 S.n10226 0.047
R6529 S.n9974 S.n9970 0.047
R6530 S.n9555 S.n9550 0.047
R6531 S.n9297 S.n9293 0.047
R6532 S.n8688 S.n8683 0.047
R6533 S.n8893 S.n8889 0.047
R6534 S.n7992 S.n7987 0.047
R6535 S.n8181 S.n8177 0.047
R6536 S.n7459 S.n7174 0.047
R6537 S.n7505 S.n7473 0.047
R6538 S.n7443 S.n7437 0.047
R6539 S.n8196 S.n8192 0.047
R6540 S.n11747 S.n11743 0.047
R6541 S.n12471 S.n12466 0.047
R6542 S.n12188 S.n12184 0.047
R6543 S.n11513 S.n11508 0.047
R6544 S.n11275 S.n11271 0.047
R6545 S.n10897 S.n10892 0.047
R6546 S.n10647 S.n10643 0.047
R6547 S.n10247 S.n10242 0.047
R6548 S.n9989 S.n9985 0.047
R6549 S.n9571 S.n9566 0.047
R6550 S.n9312 S.n9308 0.047
R6551 S.n8704 S.n8699 0.047
R6552 S.n8908 S.n8904 0.047
R6553 S.n8007 S.n8003 0.047
R6554 S.n8241 S.n8209 0.047
R6555 S.n8027 S.n8021 0.047
R6556 S.n8923 S.n8919 0.047
R6557 S.n11732 S.n11728 0.047
R6558 S.n12487 S.n12482 0.047
R6559 S.n12203 S.n12199 0.047
R6560 S.n11529 S.n11524 0.047
R6561 S.n11290 S.n11286 0.047
R6562 S.n10913 S.n10908 0.047
R6563 S.n10662 S.n10658 0.047
R6564 S.n10263 S.n10258 0.047
R6565 S.n10004 S.n10000 0.047
R6566 S.n9587 S.n9582 0.047
R6567 S.n9327 S.n9323 0.047
R6568 S.n8719 S.n8715 0.047
R6569 S.n8968 S.n8936 0.047
R6570 S.n8739 S.n8733 0.047
R6571 S.n9624 S.n9338 0.047
R6572 S.n11717 S.n11713 0.047
R6573 S.n12503 S.n12498 0.047
R6574 S.n12218 S.n12214 0.047
R6575 S.n11545 S.n11540 0.047
R6576 S.n11305 S.n11301 0.047
R6577 S.n10929 S.n10924 0.047
R6578 S.n10677 S.n10673 0.047
R6579 S.n10279 S.n10274 0.047
R6580 S.n10019 S.n10015 0.047
R6581 S.n9623 S.n9346 0.047
R6582 S.n9669 S.n9637 0.047
R6583 S.n9607 S.n9601 0.047
R6584 S.n10316 S.n10030 0.047
R6585 S.n11702 S.n11698 0.047
R6586 S.n12519 S.n12514 0.047
R6587 S.n12233 S.n12229 0.047
R6588 S.n11561 S.n11556 0.047
R6589 S.n11320 S.n11316 0.047
R6590 S.n10945 S.n10940 0.047
R6591 S.n10692 S.n10688 0.047
R6592 S.n10315 S.n10038 0.047
R6593 S.n10361 S.n10329 0.047
R6594 S.n10299 S.n10293 0.047
R6595 S.n10982 S.n10703 0.047
R6596 S.n11687 S.n11683 0.047
R6597 S.n12535 S.n12530 0.047
R6598 S.n12248 S.n12244 0.047
R6599 S.n11577 S.n11572 0.047
R6600 S.n11335 S.n11331 0.047
R6601 S.n10981 S.n10711 0.047
R6602 S.n11025 S.n10995 0.047
R6603 S.n10965 S.n10959 0.047
R6604 S.n11617 S.n11346 0.047
R6605 S.n11672 S.n11668 0.047
R6606 S.n12551 S.n12546 0.047
R6607 S.n12263 S.n12259 0.047
R6608 S.n11616 S.n11354 0.047
R6609 S.n11644 S.n11630 0.047
R6610 S.n11600 S.n11589 0.047
R6611 S.n12582 S.n12579 0.047
R6612 S.n11657 S.n11655 0.047
R6613 S.n12568 S.n12566 0.047
R6614 S.n1342 S.n1337 0.047
R6615 S.n9683 S.n9682 0.047
R6616 S.n9011 S.n9010 0.047
R6617 S.n8316 S.n8315 0.047
R6618 S.n7609 S.n7608 0.047
R6619 S.n6879 S.n6878 0.047
R6620 S.n6137 S.n6136 0.047
R6621 S.n5372 S.n5371 0.047
R6622 S.n4595 S.n4594 0.047
R6623 S.n3795 S.n3794 0.047
R6624 S.n2983 S.n2982 0.047
R6625 S.n2147 S.n2146 0.047
R6626 S.t7 S.n166 0.046
R6627 S.t7 S.n156 0.046
R6628 S.t7 S.n144 0.046
R6629 S.t7 S.n132 0.046
R6630 S.t7 S.n119 0.046
R6631 S.t7 S.n106 0.046
R6632 S.t7 S.n93 0.046
R6633 S.n1808 S.n1798 0.046
R6634 S.n2651 S.n2650 0.046
R6635 S.n5130 S.n5129 0.045
R6636 S.n5927 S.n5926 0.045
R6637 S.n6698 S.n6697 0.045
R6638 S.n7460 S.n7459 0.045
R6639 S.n9624 S.n9623 0.045
R6640 S.n10316 S.n10315 0.045
R6641 S.n10982 S.n10981 0.045
R6642 S.n11617 S.n11616 0.045
R6643 S.n4324 S.n4315 0.045
R6644 S.n173 S.n171 0.045
R6645 S.n12581 S.n12580 0.045
R6646 S.n855 S.n854 0.045
R6647 S.n1359 S.n1351 0.045
R6648 S.n2194 S.n2186 0.045
R6649 S.n3030 S.n3022 0.045
R6650 S.n3842 S.n3834 0.045
R6651 S.n4642 S.n4634 0.045
R6652 S.n5419 S.n5411 0.045
R6653 S.n6184 S.n6176 0.045
R6654 S.n6926 S.n6918 0.045
R6655 S.n7656 S.n7648 0.045
R6656 S.n8363 S.n8355 0.045
R6657 S.n9058 S.n9050 0.045
R6658 S.n9730 S.n9722 0.045
R6659 S.n10390 S.n10382 0.045
R6660 S.n2680 S.n2679 0.045
R6661 S.n3521 S.n3520 0.045
R6662 S.n4353 S.n4352 0.045
R6663 S.n5159 S.n5158 0.045
R6664 S.n5956 S.n5955 0.045
R6665 S.n6727 S.n6726 0.045
R6666 S.n7489 S.n7488 0.045
R6667 S.n8225 S.n8224 0.045
R6668 S.n8952 S.n8951 0.045
R6669 S.n9653 S.n9652 0.045
R6670 S.n10345 S.n10344 0.045
R6671 S.n11009 S.n11008 0.045
R6672 S.n12582 S.n12568 0.044
R6673 S.n2318 S.n2305 0.044
R6674 S.n3446 S.n3433 0.044
R6675 S.n3965 S.n3952 0.044
R6676 S.n4760 S.n4747 0.044
R6677 S.n5542 S.n5529 0.044
R6678 S.n6302 S.n6289 0.044
R6679 S.n7049 S.n7036 0.044
R6680 S.n8060 S.n8047 0.044
R6681 S.n8772 S.n8759 0.044
R6682 S.n9176 S.n9163 0.044
R6683 S.n9853 S.n9840 0.044
R6684 S.n10511 S.n10498 0.044
R6685 S.n11139 S.n11126 0.044
R6686 S.n12067 S.n12054 0.044
R6687 S.n3477 S.n3476 0.044
R6688 S.n3996 S.n3995 0.044
R6689 S.n4791 S.n4790 0.044
R6690 S.n5573 S.n5572 0.044
R6691 S.n6333 S.n6332 0.044
R6692 S.n7080 S.n7079 0.044
R6693 S.n8091 S.n8090 0.044
R6694 S.n8803 S.n8802 0.044
R6695 S.n9207 S.n9206 0.044
R6696 S.n9884 S.n9883 0.044
R6697 S.n10542 S.n10541 0.044
R6698 S.n11170 S.n11169 0.044
R6699 S.n12083 S.n12082 0.044
R6700 S.n497 S.n496 0.044
R6701 S.n453 S.n452 0.044
R6702 S.n409 S.n408 0.044
R6703 S.n365 S.n364 0.044
R6704 S.n321 S.n320 0.044
R6705 S.n277 S.n276 0.044
R6706 S.n834 S.n833 0.043
R6707 S.n12034 S.n12033 0.043
R6708 S.n1293 S.n1292 0.042
R6709 S.n2111 S.n2110 0.042
R6710 S.n2948 S.n2947 0.042
R6711 S.n3760 S.n3759 0.042
R6712 S.n4560 S.n4559 0.042
R6713 S.n5337 S.n5336 0.042
R6714 S.n6102 S.n6101 0.042
R6715 S.n6844 S.n6843 0.042
R6716 S.n7574 S.n7573 0.042
R6717 S.n8281 S.n8280 0.042
R6718 S.n8976 S.n8975 0.042
R6719 S.n1234 S.n1233 0.042
R6720 S.n2050 S.n2049 0.042
R6721 S.n2887 S.n2886 0.042
R6722 S.n3699 S.n3698 0.042
R6723 S.n4499 S.n4498 0.042
R6724 S.n5276 S.n5275 0.042
R6725 S.n6041 S.n6040 0.042
R6726 S.n6783 S.n6782 0.042
R6727 S.n7513 S.n7512 0.042
R6728 S.n1175 S.n1174 0.042
R6729 S.n1989 S.n1988 0.042
R6730 S.n2826 S.n2825 0.042
R6731 S.n3638 S.n3637 0.042
R6732 S.n4438 S.n4437 0.042
R6733 S.n5215 S.n5214 0.042
R6734 S.n5980 S.n5979 0.042
R6735 S.n1116 S.n1115 0.042
R6736 S.n1928 S.n1927 0.042
R6737 S.n2765 S.n2764 0.042
R6738 S.n3577 S.n3576 0.042
R6739 S.n4377 S.n4376 0.042
R6740 S.n1057 S.n1056 0.042
R6741 S.n1867 S.n1866 0.042
R6742 S.n2704 S.n2703 0.042
R6743 S.n998 S.n997 0.042
R6744 S.n12019 S.n12016 0.042
R6745 S.n11071 S.n11068 0.042
R6746 S.n10441 S.n10438 0.042
R6747 S.n9781 S.n9778 0.042
R6748 S.n9109 S.n9106 0.042
R6749 S.n8414 S.n8411 0.042
R6750 S.n7707 S.n7704 0.042
R6751 S.n6977 S.n6974 0.042
R6752 S.n6235 S.n6232 0.042
R6753 S.n5470 S.n5467 0.042
R6754 S.n4693 S.n4690 0.042
R6755 S.n3893 S.n3890 0.042
R6756 S.n3081 S.n3078 0.042
R6757 S.n2246 S.n2243 0.042
R6758 S.n1427 S.n1422 0.042
R6759 S.n8267 S.n8264 0.042
R6760 S.n7560 S.n7557 0.042
R6761 S.n6830 S.n6827 0.042
R6762 S.n6088 S.n6085 0.042
R6763 S.n5323 S.n5320 0.042
R6764 S.n4546 S.n4543 0.042
R6765 S.n3746 S.n3743 0.042
R6766 S.n2934 S.n2931 0.042
R6767 S.n2097 S.n2094 0.042
R6768 S.n9695 S.n9692 0.042
R6769 S.n9023 S.n9020 0.042
R6770 S.n8328 S.n8325 0.042
R6771 S.n7621 S.n7618 0.042
R6772 S.n6891 S.n6888 0.042
R6773 S.n6149 S.n6146 0.042
R6774 S.n5384 S.n5381 0.042
R6775 S.n4607 S.n4604 0.042
R6776 S.n3807 S.n3804 0.042
R6777 S.n2995 S.n2992 0.042
R6778 S.n2159 S.n2156 0.042
R6779 S.n6769 S.n6766 0.042
R6780 S.n6027 S.n6024 0.042
R6781 S.n5262 S.n5259 0.042
R6782 S.n4485 S.n4482 0.042
R6783 S.n3685 S.n3682 0.042
R6784 S.n2873 S.n2870 0.042
R6785 S.n2036 S.n2033 0.042
R6786 S.n5201 S.n5198 0.042
R6787 S.n4424 S.n4421 0.042
R6788 S.n3624 S.n3621 0.042
R6789 S.n2812 S.n2809 0.042
R6790 S.n1975 S.n1972 0.042
R6791 S.n3563 S.n3560 0.042
R6792 S.n2751 S.n2748 0.042
R6793 S.n1914 S.n1911 0.042
R6794 S.n1853 S.n1850 0.042
R6795 S.n11033 S.n11032 0.042
R6796 S.n10403 S.n10402 0.042
R6797 S.n9743 S.n9742 0.042
R6798 S.n9071 S.n9070 0.042
R6799 S.n8376 S.n8375 0.042
R6800 S.n7669 S.n7668 0.042
R6801 S.n6939 S.n6938 0.042
R6802 S.n6197 S.n6196 0.042
R6803 S.n5432 S.n5431 0.042
R6804 S.n4655 S.n4654 0.042
R6805 S.n3855 S.n3854 0.042
R6806 S.n3043 S.n3042 0.042
R6807 S.n2207 S.n2206 0.042
R6808 S.n1388 S.n1387 0.042
R6809 S.n882 S.n881 0.041
R6810 S.n10457 S.n10456 0.041
R6811 S.n249 S.n248 0.041
R6812 S.n531 S.n522 0.04
R6813 S.n1478 S.n1469 0.04
R6814 S.n2352 S.n2343 0.04
R6815 S.n3134 S.n3125 0.04
R6816 S.n4036 S.n4027 0.04
R6817 S.n4853 S.n4844 0.04
R6818 S.n5652 S.n5643 0.04
R6819 S.n6425 S.n6416 0.04
R6820 S.n7189 S.n7180 0.04
R6821 S.n7760 S.n7751 0.04
R6822 S.n8474 S.n8465 0.04
R6823 S.n9359 S.n9350 0.04
R6824 S.n10053 S.n10044 0.04
R6825 S.n81 S.n67 0.04
R6826 S.n66 S.n65 0.039
R6827 S.n12600 S.n12599 0.039
R6828 S.n2681 S.n2680 0.039
R6829 S.n2686 S.n2685 0.039
R6830 S.n3522 S.n3521 0.039
R6831 S.n3527 S.n3526 0.039
R6832 S.n4354 S.n4353 0.039
R6833 S.n4359 S.n4358 0.039
R6834 S.n5160 S.n5159 0.039
R6835 S.n5165 S.n5164 0.039
R6836 S.n5957 S.n5956 0.039
R6837 S.n5962 S.n5961 0.039
R6838 S.n6728 S.n6727 0.039
R6839 S.n6733 S.n6732 0.039
R6840 S.n7490 S.n7489 0.039
R6841 S.n7495 S.n7494 0.039
R6842 S.n8226 S.n8225 0.039
R6843 S.n8231 S.n8230 0.039
R6844 S.n8953 S.n8952 0.039
R6845 S.n8958 S.n8957 0.039
R6846 S.n9654 S.n9653 0.039
R6847 S.n9659 S.n9658 0.039
R6848 S.n10346 S.n10345 0.039
R6849 S.n10351 S.n10350 0.039
R6850 S.n11010 S.n11009 0.039
R6851 S.n11015 S.n11014 0.039
R6852 S.n530 S.n523 0.039
R6853 S.n1477 S.n1470 0.039
R6854 S.n2351 S.n2344 0.039
R6855 S.n3133 S.n3126 0.039
R6856 S.n4035 S.n4028 0.039
R6857 S.n4852 S.n4845 0.039
R6858 S.n5651 S.n5644 0.039
R6859 S.n6424 S.n6417 0.039
R6860 S.n7188 S.n7181 0.039
R6861 S.n7759 S.n7752 0.039
R6862 S.n8473 S.n8466 0.039
R6863 S.n9358 S.n9351 0.039
R6864 S.n10052 S.n10045 0.039
R6865 S.n10720 S.n10714 0.039
R6866 S.n12282 S.n12280 0.038
R6867 S.n12007 S.n12006 0.038
R6868 S.n11059 S.n11058 0.038
R6869 S.n10429 S.n10428 0.038
R6870 S.n9769 S.n9768 0.038
R6871 S.n9097 S.n9096 0.038
R6872 S.n8402 S.n8401 0.038
R6873 S.n7695 S.n7694 0.038
R6874 S.n6965 S.n6964 0.038
R6875 S.n6223 S.n6222 0.038
R6876 S.n5458 S.n5457 0.038
R6877 S.n4681 S.n4680 0.038
R6878 S.n3881 S.n3880 0.038
R6879 S.n3069 S.n3068 0.038
R6880 S.n2234 S.n2233 0.038
R6881 S.n8255 S.n8254 0.038
R6882 S.n7548 S.n7547 0.038
R6883 S.n6818 S.n6817 0.038
R6884 S.n6076 S.n6075 0.038
R6885 S.n5311 S.n5310 0.038
R6886 S.n4534 S.n4533 0.038
R6887 S.n3734 S.n3733 0.038
R6888 S.n2922 S.n2921 0.038
R6889 S.n2085 S.n2084 0.038
R6890 S.n1268 S.n1267 0.038
R6891 S.n8993 S.n8988 0.038
R6892 S.n8298 S.n8293 0.038
R6893 S.n7591 S.n7586 0.038
R6894 S.n6861 S.n6856 0.038
R6895 S.n6119 S.n6114 0.038
R6896 S.n5354 S.n5349 0.038
R6897 S.n4577 S.n4572 0.038
R6898 S.n3777 S.n3772 0.038
R6899 S.n2965 S.n2960 0.038
R6900 S.n2128 S.n2123 0.038
R6901 S.n1308 S.n1304 0.038
R6902 S.n6757 S.n6756 0.038
R6903 S.n6015 S.n6014 0.038
R6904 S.n5250 S.n5249 0.038
R6905 S.n4473 S.n4472 0.038
R6906 S.n3673 S.n3672 0.038
R6907 S.n2861 S.n2860 0.038
R6908 S.n2024 S.n2023 0.038
R6909 S.n1209 S.n1208 0.038
R6910 S.n7530 S.n7525 0.038
R6911 S.n6800 S.n6795 0.038
R6912 S.n6058 S.n6053 0.038
R6913 S.n5293 S.n5288 0.038
R6914 S.n4516 S.n4511 0.038
R6915 S.n3716 S.n3711 0.038
R6916 S.n2904 S.n2899 0.038
R6917 S.n2067 S.n2062 0.038
R6918 S.n1250 S.n1245 0.038
R6919 S.n5189 S.n5188 0.038
R6920 S.n4412 S.n4411 0.038
R6921 S.n3612 S.n3611 0.038
R6922 S.n2800 S.n2799 0.038
R6923 S.n1963 S.n1962 0.038
R6924 S.n1150 S.n1149 0.038
R6925 S.n5997 S.n5992 0.038
R6926 S.n5232 S.n5227 0.038
R6927 S.n4455 S.n4450 0.038
R6928 S.n3655 S.n3650 0.038
R6929 S.n2843 S.n2838 0.038
R6930 S.n2006 S.n2001 0.038
R6931 S.n1191 S.n1186 0.038
R6932 S.n3551 S.n3550 0.038
R6933 S.n2739 S.n2738 0.038
R6934 S.n1902 S.n1901 0.038
R6935 S.n1091 S.n1090 0.038
R6936 S.n4394 S.n4389 0.038
R6937 S.n3594 S.n3589 0.038
R6938 S.n2782 S.n2777 0.038
R6939 S.n1948 S.n1943 0.038
R6940 S.n1132 S.n1127 0.038
R6941 S.n1841 S.n1840 0.038
R6942 S.n1032 S.n1031 0.038
R6943 S.n2721 S.n2716 0.038
R6944 S.n1884 S.n1879 0.038
R6945 S.n1073 S.n1068 0.038
R6946 S.n1014 S.n1009 0.038
R6947 S.n944 S.n943 0.038
R6948 S.n11101 S.n11099 0.037
R6949 S.n12600 S.n12597 0.037
R6950 S.n12599 S.n12598 0.037
R6951 S.n2197 S.n2179 0.037
R6952 S.n3033 S.n3015 0.037
R6953 S.n3845 S.n3827 0.037
R6954 S.n4645 S.n4627 0.037
R6955 S.n5422 S.n5404 0.037
R6956 S.n6187 S.n6169 0.037
R6957 S.n6929 S.n6911 0.037
R6958 S.n7659 S.n7641 0.037
R6959 S.n8366 S.n8348 0.037
R6960 S.n9061 S.n9043 0.037
R6961 S.n9733 S.n9715 0.037
R6962 S.n10393 S.n10375 0.037
R6963 S.n11102 S.n11091 0.037
R6964 S.n1406 S.n1398 0.037
R6965 S.n1378 S.n1370 0.037
R6966 S.n2686 S.n2683 0.037
R6967 S.n2685 S.n2684 0.037
R6968 S.n3527 S.n3524 0.037
R6969 S.n3526 S.n3525 0.037
R6970 S.n4359 S.n4356 0.037
R6971 S.n4358 S.n4357 0.037
R6972 S.n5165 S.n5162 0.037
R6973 S.n5164 S.n5163 0.037
R6974 S.n5962 S.n5959 0.037
R6975 S.n5961 S.n5960 0.037
R6976 S.n6733 S.n6730 0.037
R6977 S.n6732 S.n6731 0.037
R6978 S.n7495 S.n7492 0.037
R6979 S.n7494 S.n7493 0.037
R6980 S.n8231 S.n8228 0.037
R6981 S.n8230 S.n8229 0.037
R6982 S.n8958 S.n8955 0.037
R6983 S.n8957 S.n8956 0.037
R6984 S.n9659 S.n9656 0.037
R6985 S.n9658 S.n9657 0.037
R6986 S.n10351 S.n10348 0.037
R6987 S.n10350 S.n10349 0.037
R6988 S.n11015 S.n11012 0.037
R6989 S.n11014 S.n11013 0.037
R6990 S.n11648 S.n11647 0.037
R6991 S.n12572 S.n12571 0.037
R6992 S.n980 S.n249 0.036
R6993 S.n1742 S.n1741 0.036
R6994 S.n2582 S.n2581 0.036
R6995 S.n3346 S.n3345 0.036
R6996 S.n4230 S.n4229 0.036
R6997 S.n5029 S.n5028 0.036
R6998 S.n5810 S.n5809 0.036
R6999 S.n6565 S.n6564 0.036
R7000 S.n7311 S.n7310 0.036
R7001 S.n7864 S.n7863 0.036
R7002 S.n8560 S.n8559 0.036
R7003 S.n9427 S.n9426 0.036
R7004 S.n10103 S.n10102 0.036
R7005 S.n10753 S.n10752 0.036
R7006 S.n11370 S.n11369 0.036
R7007 S.n9370 S.n9369 0.035
R7008 S.n8503 S.n8502 0.035
R7009 S.n7807 S.n7806 0.035
R7010 S.n7254 S.n7253 0.035
R7011 S.n6508 S.n6507 0.035
R7012 S.n5753 S.n5752 0.035
R7013 S.n4972 S.n4971 0.035
R7014 S.n4173 S.n4172 0.035
R7015 S.n3289 S.n3288 0.035
R7016 S.n2525 S.n2524 0.035
R7017 S.n1669 S.n1668 0.035
R7018 S.n7771 S.n7770 0.035
R7019 S.n7218 S.n7217 0.035
R7020 S.n6472 S.n6471 0.035
R7021 S.n5717 S.n5716 0.035
R7022 S.n4936 S.n4935 0.035
R7023 S.n4137 S.n4136 0.035
R7024 S.n3253 S.n3252 0.035
R7025 S.n2489 S.n2488 0.035
R7026 S.n1633 S.n1632 0.035
R7027 S.n6436 S.n6435 0.035
R7028 S.n5681 S.n5680 0.035
R7029 S.n4900 S.n4899 0.035
R7030 S.n4101 S.n4100 0.035
R7031 S.n3217 S.n3216 0.035
R7032 S.n2453 S.n2452 0.035
R7033 S.n1597 S.n1596 0.035
R7034 S.n4864 S.n4863 0.035
R7035 S.n4065 S.n4064 0.035
R7036 S.n3181 S.n3180 0.035
R7037 S.n2417 S.n2416 0.035
R7038 S.n1561 S.n1560 0.035
R7039 S.n3145 S.n3144 0.035
R7040 S.n2381 S.n2380 0.035
R7041 S.n1525 S.n1524 0.035
R7042 S.n1489 S.n1488 0.035
R7043 S.n11902 S.n11901 0.035
R7044 S.n12601 S.n12600 0.035
R7045 S.n12007 S.n12002 0.035
R7046 S.n11059 S.n11054 0.035
R7047 S.n10429 S.n10424 0.035
R7048 S.n9769 S.n9764 0.035
R7049 S.n9097 S.n9092 0.035
R7050 S.n8402 S.n8397 0.035
R7051 S.n7695 S.n7690 0.035
R7052 S.n6965 S.n6960 0.035
R7053 S.n6223 S.n6218 0.035
R7054 S.n5458 S.n5453 0.035
R7055 S.n4681 S.n4676 0.035
R7056 S.n3881 S.n3876 0.035
R7057 S.n3069 S.n3064 0.035
R7058 S.n2234 S.n2229 0.035
R7059 S.n8255 S.n8250 0.035
R7060 S.n7548 S.n7543 0.035
R7061 S.n6818 S.n6813 0.035
R7062 S.n6076 S.n6071 0.035
R7063 S.n5311 S.n5306 0.035
R7064 S.n4534 S.n4529 0.035
R7065 S.n3734 S.n3729 0.035
R7066 S.n2922 S.n2917 0.035
R7067 S.n2085 S.n2080 0.035
R7068 S.n1268 S.n1263 0.035
R7069 S.n10474 S.n10457 0.035
R7070 S.n1308 S.n1307 0.035
R7071 S.n2128 S.n2127 0.035
R7072 S.n2965 S.n2964 0.035
R7073 S.n3777 S.n3776 0.035
R7074 S.n4577 S.n4576 0.035
R7075 S.n5354 S.n5353 0.035
R7076 S.n6119 S.n6118 0.035
R7077 S.n6861 S.n6860 0.035
R7078 S.n7591 S.n7590 0.035
R7079 S.n8298 S.n8297 0.035
R7080 S.n8993 S.n8992 0.035
R7081 S.n6757 S.n6752 0.035
R7082 S.n6015 S.n6010 0.035
R7083 S.n5250 S.n5245 0.035
R7084 S.n4473 S.n4468 0.035
R7085 S.n3673 S.n3668 0.035
R7086 S.n2861 S.n2856 0.035
R7087 S.n2024 S.n2019 0.035
R7088 S.n1209 S.n1204 0.035
R7089 S.n1250 S.n1249 0.035
R7090 S.n2067 S.n2066 0.035
R7091 S.n2904 S.n2903 0.035
R7092 S.n3716 S.n3715 0.035
R7093 S.n4516 S.n4515 0.035
R7094 S.n5293 S.n5292 0.035
R7095 S.n6058 S.n6057 0.035
R7096 S.n6800 S.n6799 0.035
R7097 S.n7530 S.n7529 0.035
R7098 S.n5189 S.n5184 0.035
R7099 S.n4412 S.n4407 0.035
R7100 S.n3612 S.n3607 0.035
R7101 S.n2800 S.n2795 0.035
R7102 S.n1963 S.n1958 0.035
R7103 S.n1150 S.n1145 0.035
R7104 S.n1191 S.n1190 0.035
R7105 S.n2006 S.n2005 0.035
R7106 S.n2843 S.n2842 0.035
R7107 S.n3655 S.n3654 0.035
R7108 S.n4455 S.n4454 0.035
R7109 S.n5232 S.n5231 0.035
R7110 S.n5997 S.n5996 0.035
R7111 S.n3551 S.n3546 0.035
R7112 S.n2739 S.n2734 0.035
R7113 S.n1902 S.n1897 0.035
R7114 S.n1091 S.n1086 0.035
R7115 S.n1132 S.n1131 0.035
R7116 S.n1948 S.n1947 0.035
R7117 S.n2782 S.n2781 0.035
R7118 S.n3594 S.n3593 0.035
R7119 S.n4394 S.n4393 0.035
R7120 S.n1841 S.n1836 0.035
R7121 S.n1032 S.n1027 0.035
R7122 S.n1073 S.n1072 0.035
R7123 S.n1884 S.n1883 0.035
R7124 S.n2721 S.n2720 0.035
R7125 S.n1014 S.n1013 0.035
R7126 S.n2679 S.n2678 0.035
R7127 S.n2689 S.n2686 0.035
R7128 S.n3520 S.n3519 0.035
R7129 S.n3530 S.n3527 0.035
R7130 S.n4352 S.n4351 0.035
R7131 S.n4362 S.n4359 0.035
R7132 S.n5158 S.n5157 0.035
R7133 S.n5168 S.n5165 0.035
R7134 S.n5955 S.n5954 0.035
R7135 S.n5965 S.n5962 0.035
R7136 S.n6726 S.n6725 0.035
R7137 S.n6736 S.n6733 0.035
R7138 S.n7488 S.n7487 0.035
R7139 S.n7498 S.n7495 0.035
R7140 S.n8224 S.n8223 0.035
R7141 S.n8234 S.n8231 0.035
R7142 S.n8951 S.n8950 0.035
R7143 S.n8961 S.n8958 0.035
R7144 S.n9652 S.n9651 0.035
R7145 S.n9662 S.n9659 0.035
R7146 S.n10344 S.n10343 0.035
R7147 S.n10354 S.n10351 0.035
R7148 S.n11008 S.n11007 0.035
R7149 S.n11018 S.n11015 0.035
R7150 S.n11634 S.n11633 0.034
R7151 S.n11878 S.n11877 0.034
R7152 S.n539 S.n538 0.034
R7153 S.n9368 S.n9367 0.034
R7154 S.n10061 S.n10060 0.034
R7155 S.n10730 S.n10729 0.034
R7156 S.n11368 S.n11367 0.034
R7157 S.n12290 S.n12289 0.034
R7158 S.n7769 S.n7768 0.034
R7159 S.n8482 S.n8481 0.034
R7160 S.n6434 S.n6433 0.034
R7161 S.n7197 S.n7196 0.034
R7162 S.n4862 S.n4861 0.034
R7163 S.n5660 S.n5659 0.034
R7164 S.n3143 S.n3142 0.034
R7165 S.n4044 S.n4043 0.034
R7166 S.n1487 S.n1486 0.034
R7167 S.n2360 S.n2359 0.034
R7168 S.n165 S.n161 0.034
R7169 S.n158 S.n157 0.034
R7170 S.n146 S.n145 0.034
R7171 S.n134 S.n133 0.034
R7172 S.n121 S.n120 0.034
R7173 S.n108 S.n107 0.034
R7174 S.n95 S.n94 0.034
R7175 S.n11870 S.n11866 0.034
R7176 S.n12344 S.n12341 0.034
R7177 S.n12067 S.n12063 0.034
R7178 S.n11125 S.n11122 0.034
R7179 S.n11139 S.n11135 0.034
R7180 S.n10497 S.n10494 0.034
R7181 S.n10511 S.n10507 0.034
R7182 S.n9839 S.n9836 0.034
R7183 S.n9853 S.n9849 0.034
R7184 S.n9162 S.n9159 0.034
R7185 S.n9176 S.n9172 0.034
R7186 S.n8758 S.n8755 0.034
R7187 S.n8772 S.n8768 0.034
R7188 S.n8046 S.n8043 0.034
R7189 S.n8060 S.n8056 0.034
R7190 S.n7035 S.n7032 0.034
R7191 S.n7049 S.n7045 0.034
R7192 S.n6288 S.n6285 0.034
R7193 S.n6302 S.n6298 0.034
R7194 S.n5528 S.n5525 0.034
R7195 S.n5542 S.n5538 0.034
R7196 S.n4746 S.n4743 0.034
R7197 S.n4760 S.n4756 0.034
R7198 S.n3951 S.n3948 0.034
R7199 S.n3965 S.n3961 0.034
R7200 S.n3432 S.n3429 0.034
R7201 S.n3446 S.n3442 0.034
R7202 S.n2304 S.n2301 0.034
R7203 S.n2318 S.n2314 0.034
R7204 S.n1798 S.n1795 0.034
R7205 S.n1826 S.n981 0.034
R7206 S.n2696 S.n1828 0.034
R7207 S.n4369 S.n3538 0.034
R7208 S.n5175 S.n4370 0.034
R7209 S.n5972 S.n5176 0.034
R7210 S.n6743 S.n5973 0.034
R7211 S.n7505 S.n6744 0.034
R7212 S.n8241 S.n7506 0.034
R7213 S.n8968 S.n8242 0.034
R7214 S.n9669 S.n8969 0.034
R7215 S.n10361 S.n9670 0.034
R7216 S.n11025 S.n10362 0.034
R7217 S.n11644 S.n11026 0.034
R7218 S.n12611 S.n12610 0.034
R7219 S.n3537 S.n2697 0.034
R7220 S.n529 S.n524 0.034
R7221 S.n1476 S.n1471 0.034
R7222 S.n2350 S.n2345 0.034
R7223 S.n3132 S.n3127 0.034
R7224 S.n4034 S.n4029 0.034
R7225 S.n4851 S.n4846 0.034
R7226 S.n5650 S.n5645 0.034
R7227 S.n6423 S.n6418 0.034
R7228 S.n7187 S.n7182 0.034
R7229 S.n7758 S.n7753 0.034
R7230 S.n8472 S.n8467 0.034
R7231 S.n9357 S.n9352 0.034
R7232 S.n10051 S.n10046 0.034
R7233 S.n10719 S.n10715 0.034
R7234 S.n10723 S.n10713 0.034
R7235 S.n10055 S.n10042 0.034
R7236 S.n9361 S.n9348 0.034
R7237 S.n8476 S.n8463 0.034
R7238 S.n7762 S.n7749 0.034
R7239 S.n7191 S.n7178 0.034
R7240 S.n6427 S.n6414 0.034
R7241 S.n5654 S.n5641 0.034
R7242 S.n4855 S.n4842 0.034
R7243 S.n4038 S.n4025 0.034
R7244 S.n3136 S.n3123 0.034
R7245 S.n2354 S.n2341 0.034
R7246 S.n1480 S.n1467 0.034
R7247 S.n533 S.n520 0.034
R7248 S.t0 S.n11991 0.034
R7249 S.t0 S.n11990 0.034
R7250 S.t7 S.n209 0.034
R7251 S.t7 S.n212 0.034
R7252 S.t7 S.n205 0.034
R7253 S.t7 S.n204 0.034
R7254 S.t7 S.n154 0.034
R7255 S.t7 S.n153 0.034
R7256 S.t7 S.n233 0.034
R7257 S.t7 S.n236 0.034
R7258 S.t7 S.n168 0.034
R7259 S.t7 S.n167 0.034
R7260 S.t7 S.n179 0.034
R7261 S.t7 S.n178 0.034
R7262 S.t7 S.n192 0.034
R7263 S.t7 S.n191 0.034
R7264 S.t7 S.n142 0.034
R7265 S.t7 S.n141 0.034
R7266 S.t7 S.n229 0.034
R7267 S.t7 S.n232 0.034
R7268 S.t7 S.n129 0.034
R7269 S.t7 S.n128 0.034
R7270 S.t7 S.n225 0.034
R7271 S.t7 S.n228 0.034
R7272 S.t7 S.n116 0.034
R7273 S.t7 S.n115 0.034
R7274 S.t7 S.n221 0.034
R7275 S.t7 S.n224 0.034
R7276 S.t7 S.n103 0.034
R7277 S.t7 S.n102 0.034
R7278 S.t7 S.n217 0.034
R7279 S.t7 S.n220 0.034
R7280 S.t7 S.n90 0.034
R7281 S.t7 S.n89 0.034
R7282 S.t7 S.n213 0.034
R7283 S.t7 S.n216 0.034
R7284 S.t0 S.n11931 0.034
R7285 S.t0 S.n11930 0.034
R7286 S.t0 S.n11934 0.034
R7287 S.t0 S.n11935 0.034
R7288 S.t0 S.n11938 0.034
R7289 S.t0 S.n11939 0.034
R7290 S.t0 S.n11942 0.034
R7291 S.t0 S.n11943 0.034
R7292 S.t0 S.n11946 0.034
R7293 S.t0 S.n11947 0.034
R7294 S.t0 S.n11950 0.034
R7295 S.t0 S.n11951 0.034
R7296 S.t0 S.n11954 0.034
R7297 S.t0 S.n11955 0.034
R7298 S.t0 S.n11958 0.034
R7299 S.t0 S.n11959 0.034
R7300 S.t0 S.n11962 0.034
R7301 S.t0 S.n11963 0.034
R7302 S.t0 S.n11966 0.034
R7303 S.t0 S.n11967 0.034
R7304 S.t0 S.n11970 0.034
R7305 S.t0 S.n11971 0.034
R7306 S.t0 S.n11974 0.034
R7307 S.t0 S.n11975 0.034
R7308 S.t0 S.n11978 0.034
R7309 S.t0 S.n11979 0.034
R7310 S.t0 S.n11982 0.034
R7311 S.t0 S.n11983 0.034
R7312 S.t0 S.n11987 0.034
R7313 S.t0 S.n11986 0.034
R7314 S.t0 S.n11926 0.034
R7315 S.t0 S.n11929 0.034
R7316 S.n81 S.n80 0.033
R7317 S.n1701 S.n1700 0.033
R7318 S.n12283 S.n12282 0.032
R7319 S.n11357 S.n11356 0.032
R7320 S.n1448 S.n1447 0.031
R7321 S.t65 S.n11878 0.031
R7322 S.t244 S.n539 0.031
R7323 S.t225 S.n9368 0.031
R7324 S.t124 S.n10061 0.031
R7325 S.t144 S.n10730 0.031
R7326 S.t47 S.n11368 0.031
R7327 S.t106 S.n12290 0.031
R7328 S.t11 S.n7769 0.031
R7329 S.t40 S.n8482 0.031
R7330 S.t4 S.n6434 0.031
R7331 S.t102 S.n7197 0.031
R7332 S.t77 S.n4862 0.031
R7333 S.t25 S.n5660 0.031
R7334 S.t38 S.n3143 0.031
R7335 S.t94 S.n4044 0.031
R7336 S.t175 S.n1487 0.031
R7337 S.t187 S.n2360 0.031
R7338 S.n12002 S.n12001 0.031
R7339 S.n11054 S.n11053 0.031
R7340 S.n10424 S.n10423 0.031
R7341 S.n9764 S.n9763 0.031
R7342 S.n9092 S.n9091 0.031
R7343 S.n8397 S.n8396 0.031
R7344 S.n7690 S.n7689 0.031
R7345 S.n6960 S.n6959 0.031
R7346 S.n6218 S.n6217 0.031
R7347 S.n5453 S.n5452 0.031
R7348 S.n4676 S.n4675 0.031
R7349 S.n3876 S.n3875 0.031
R7350 S.n3064 S.n3063 0.031
R7351 S.n2229 S.n2228 0.031
R7352 S.n8250 S.n8249 0.031
R7353 S.n7543 S.n7542 0.031
R7354 S.n6813 S.n6812 0.031
R7355 S.n6071 S.n6070 0.031
R7356 S.n5306 S.n5305 0.031
R7357 S.n4529 S.n4528 0.031
R7358 S.n3729 S.n3728 0.031
R7359 S.n2917 S.n2916 0.031
R7360 S.n2080 S.n2079 0.031
R7361 S.n1263 S.n1262 0.031
R7362 S.n1307 S.n1306 0.031
R7363 S.n2127 S.n2126 0.031
R7364 S.n2964 S.n2963 0.031
R7365 S.n3776 S.n3775 0.031
R7366 S.n4576 S.n4575 0.031
R7367 S.n5353 S.n5352 0.031
R7368 S.n6118 S.n6117 0.031
R7369 S.n6860 S.n6859 0.031
R7370 S.n7590 S.n7589 0.031
R7371 S.n8297 S.n8296 0.031
R7372 S.n8992 S.n8991 0.031
R7373 S.n6752 S.n6751 0.031
R7374 S.n6010 S.n6009 0.031
R7375 S.n5245 S.n5244 0.031
R7376 S.n4468 S.n4467 0.031
R7377 S.n3668 S.n3667 0.031
R7378 S.n2856 S.n2855 0.031
R7379 S.n2019 S.n2018 0.031
R7380 S.n1204 S.n1203 0.031
R7381 S.n1249 S.n1248 0.031
R7382 S.n2066 S.n2065 0.031
R7383 S.n2903 S.n2902 0.031
R7384 S.n3715 S.n3714 0.031
R7385 S.n4515 S.n4514 0.031
R7386 S.n5292 S.n5291 0.031
R7387 S.n6057 S.n6056 0.031
R7388 S.n6799 S.n6798 0.031
R7389 S.n7529 S.n7528 0.031
R7390 S.n5184 S.n5183 0.031
R7391 S.n4407 S.n4406 0.031
R7392 S.n3607 S.n3606 0.031
R7393 S.n2795 S.n2794 0.031
R7394 S.n1958 S.n1957 0.031
R7395 S.n1145 S.n1144 0.031
R7396 S.n1190 S.n1189 0.031
R7397 S.n2005 S.n2004 0.031
R7398 S.n2842 S.n2841 0.031
R7399 S.n3654 S.n3653 0.031
R7400 S.n4454 S.n4453 0.031
R7401 S.n5231 S.n5230 0.031
R7402 S.n5996 S.n5995 0.031
R7403 S.n3546 S.n3545 0.031
R7404 S.n2734 S.n2733 0.031
R7405 S.n1897 S.n1896 0.031
R7406 S.n1086 S.n1085 0.031
R7407 S.n1131 S.n1130 0.031
R7408 S.n1947 S.n1946 0.031
R7409 S.n2781 S.n2780 0.031
R7410 S.n3593 S.n3592 0.031
R7411 S.n4393 S.n4392 0.031
R7412 S.n1836 S.n1835 0.031
R7413 S.n1027 S.n1026 0.031
R7414 S.n1072 S.n1071 0.031
R7415 S.n1883 S.n1882 0.031
R7416 S.n2720 S.n2719 0.031
R7417 S.n1013 S.n1012 0.031
R7418 S.n239 S.n238 0.031
R7419 S.n240 S.n239 0.031
R7420 S.n241 S.n240 0.031
R7421 S.n242 S.n241 0.031
R7422 S.n243 S.n242 0.031
R7423 S.n244 S.n243 0.031
R7424 S.n245 S.n244 0.031
R7425 S.n247 S.n246 0.031
R7426 S.n12627 S.n12626 0.031
R7427 S.n12626 S.n12625 0.031
R7428 S.n12625 S.n12624 0.031
R7429 S.n12624 S.n12623 0.031
R7430 S.n12623 S.n12622 0.031
R7431 S.n12622 S.n12621 0.031
R7432 S.n12621 S.n12620 0.031
R7433 S.n12620 S.n12619 0.031
R7434 S.n12619 S.n12618 0.031
R7435 S.n12618 S.n12617 0.031
R7436 S.n12617 S.n12616 0.031
R7437 S.n12616 S.n12615 0.031
R7438 S.n12615 S.n12614 0.031
R7439 S.n12614 S.n12613 0.031
R7440 S.n12613 S.n12612 0.031
R7441 S.n12612 S.n11996 0.031
R7442 S.n11868 S.n11867 0.031
R7443 S.n12065 S.n12064 0.031
R7444 S.n11137 S.n11136 0.031
R7445 S.n10509 S.n10508 0.031
R7446 S.n9851 S.n9850 0.031
R7447 S.n9174 S.n9173 0.031
R7448 S.n8770 S.n8769 0.031
R7449 S.n8058 S.n8057 0.031
R7450 S.n7047 S.n7046 0.031
R7451 S.n6300 S.n6299 0.031
R7452 S.n5540 S.n5539 0.031
R7453 S.n4758 S.n4757 0.031
R7454 S.n3963 S.n3962 0.031
R7455 S.n3444 S.n3443 0.031
R7456 S.n2316 S.n2315 0.031
R7457 S.n9814 S.n9813 0.031
R7458 S.n5503 S.n5502 0.031
R7459 S.n2279 S.n2278 0.031
R7460 S.n9799 S.n9798 0.03
R7461 S.n8432 S.n8431 0.03
R7462 S.n6995 S.n6994 0.03
R7463 S.n5488 S.n5487 0.03
R7464 S.n3911 S.n3910 0.03
R7465 S.n2264 S.n2263 0.03
R7466 S.n10387 S.n10386 0.03
R7467 S.n9727 S.n9726 0.03
R7468 S.n9055 S.n9054 0.03
R7469 S.n8360 S.n8359 0.03
R7470 S.n7653 S.n7652 0.03
R7471 S.n6923 S.n6922 0.03
R7472 S.n6181 S.n6180 0.03
R7473 S.n5416 S.n5415 0.03
R7474 S.n4639 S.n4638 0.03
R7475 S.n3839 S.n3838 0.03
R7476 S.n3027 S.n3026 0.03
R7477 S.n2191 S.n2190 0.03
R7478 S.n1356 S.n1355 0.03
R7479 S.n848 S.n847 0.03
R7480 S.n933 S.n932 0.03
R7481 S.n9132 S.n9129 0.029
R7482 S.n10467 S.n10464 0.029
R7483 S.n7730 S.n7727 0.029
R7484 S.n6258 S.n6255 0.029
R7485 S.n4716 S.n4713 0.029
R7486 S.n3104 S.n3101 0.029
R7487 S.n1427 S.n1426 0.029
R7488 S.n2246 S.n2245 0.029
R7489 S.n3081 S.n3080 0.029
R7490 S.n3893 S.n3892 0.029
R7491 S.n4693 S.n4692 0.029
R7492 S.n5470 S.n5469 0.029
R7493 S.n6235 S.n6234 0.029
R7494 S.n6977 S.n6976 0.029
R7495 S.n7707 S.n7706 0.029
R7496 S.n8414 S.n8413 0.029
R7497 S.n9109 S.n9108 0.029
R7498 S.n9781 S.n9780 0.029
R7499 S.n10441 S.n10440 0.029
R7500 S.n11071 S.n11070 0.029
R7501 S.n12019 S.n12018 0.029
R7502 S.n2159 S.n2158 0.029
R7503 S.n2995 S.n2994 0.029
R7504 S.n3807 S.n3806 0.029
R7505 S.n4607 S.n4606 0.029
R7506 S.n5384 S.n5383 0.029
R7507 S.n6149 S.n6148 0.029
R7508 S.n6891 S.n6890 0.029
R7509 S.n7621 S.n7620 0.029
R7510 S.n8328 S.n8327 0.029
R7511 S.n9023 S.n9022 0.029
R7512 S.n9695 S.n9694 0.029
R7513 S.n2097 S.n2096 0.029
R7514 S.n2934 S.n2933 0.029
R7515 S.n3746 S.n3745 0.029
R7516 S.n4546 S.n4545 0.029
R7517 S.n5323 S.n5322 0.029
R7518 S.n6088 S.n6087 0.029
R7519 S.n6830 S.n6829 0.029
R7520 S.n7560 S.n7559 0.029
R7521 S.n8267 S.n8266 0.029
R7522 S.n2036 S.n2035 0.029
R7523 S.n2873 S.n2872 0.029
R7524 S.n3685 S.n3684 0.029
R7525 S.n4485 S.n4484 0.029
R7526 S.n5262 S.n5261 0.029
R7527 S.n6027 S.n6026 0.029
R7528 S.n6769 S.n6768 0.029
R7529 S.n1975 S.n1974 0.029
R7530 S.n2812 S.n2811 0.029
R7531 S.n3624 S.n3623 0.029
R7532 S.n4424 S.n4423 0.029
R7533 S.n5201 S.n5200 0.029
R7534 S.n1914 S.n1913 0.029
R7535 S.n2751 S.n2750 0.029
R7536 S.n3563 S.n3562 0.029
R7537 S.n1853 S.n1852 0.029
R7538 S.n2984 S.n2983 0.029
R7539 S.n3796 S.n3795 0.029
R7540 S.n4596 S.n4595 0.029
R7541 S.n5373 S.n5372 0.029
R7542 S.n6138 S.n6137 0.029
R7543 S.n6880 S.n6879 0.029
R7544 S.n7610 S.n7609 0.029
R7545 S.n8317 S.n8316 0.029
R7546 S.n9012 S.n9011 0.029
R7547 S.n9684 S.n9683 0.029
R7548 S.n10386 S.n10385 0.029
R7549 S.n9726 S.n9725 0.029
R7550 S.n9054 S.n9053 0.029
R7551 S.n8359 S.n8358 0.029
R7552 S.n7652 S.n7651 0.029
R7553 S.n6922 S.n6921 0.029
R7554 S.n6180 S.n6179 0.029
R7555 S.n5415 S.n5414 0.029
R7556 S.n4638 S.n4637 0.029
R7557 S.n3838 S.n3837 0.029
R7558 S.n3026 S.n3025 0.029
R7559 S.n2190 S.n2189 0.029
R7560 S.n1355 S.n1354 0.029
R7561 S.n847 S.n846 0.029
R7562 S.n12002 S.n11999 0.028
R7563 S.n11054 S.n11051 0.028
R7564 S.n10424 S.n10421 0.028
R7565 S.n9764 S.n9761 0.028
R7566 S.n9092 S.n9089 0.028
R7567 S.n8397 S.n8394 0.028
R7568 S.n7690 S.n7687 0.028
R7569 S.n6960 S.n6957 0.028
R7570 S.n6218 S.n6215 0.028
R7571 S.n5453 S.n5450 0.028
R7572 S.n4676 S.n4673 0.028
R7573 S.n3876 S.n3873 0.028
R7574 S.n3064 S.n3061 0.028
R7575 S.n2229 S.n2226 0.028
R7576 S.n8250 S.n8247 0.028
R7577 S.n7543 S.n7540 0.028
R7578 S.n6813 S.n6810 0.028
R7579 S.n6071 S.n6068 0.028
R7580 S.n5306 S.n5303 0.028
R7581 S.n4529 S.n4526 0.028
R7582 S.n3729 S.n3726 0.028
R7583 S.n2917 S.n2914 0.028
R7584 S.n2080 S.n2077 0.028
R7585 S.n1263 S.n1260 0.028
R7586 S.n2127 S.n2124 0.028
R7587 S.n2964 S.n2961 0.028
R7588 S.n3776 S.n3773 0.028
R7589 S.n4576 S.n4573 0.028
R7590 S.n5353 S.n5350 0.028
R7591 S.n6118 S.n6115 0.028
R7592 S.n6860 S.n6857 0.028
R7593 S.n7590 S.n7587 0.028
R7594 S.n8297 S.n8294 0.028
R7595 S.n8992 S.n8989 0.028
R7596 S.n6752 S.n6749 0.028
R7597 S.n6010 S.n6007 0.028
R7598 S.n5245 S.n5242 0.028
R7599 S.n4468 S.n4465 0.028
R7600 S.n3668 S.n3665 0.028
R7601 S.n2856 S.n2853 0.028
R7602 S.n2019 S.n2016 0.028
R7603 S.n1204 S.n1201 0.028
R7604 S.n1249 S.n1246 0.028
R7605 S.n2066 S.n2063 0.028
R7606 S.n2903 S.n2900 0.028
R7607 S.n3715 S.n3712 0.028
R7608 S.n4515 S.n4512 0.028
R7609 S.n5292 S.n5289 0.028
R7610 S.n6057 S.n6054 0.028
R7611 S.n6799 S.n6796 0.028
R7612 S.n7529 S.n7526 0.028
R7613 S.n5184 S.n5181 0.028
R7614 S.n4407 S.n4404 0.028
R7615 S.n3607 S.n3604 0.028
R7616 S.n2795 S.n2792 0.028
R7617 S.n1958 S.n1955 0.028
R7618 S.n1145 S.n1142 0.028
R7619 S.n1190 S.n1187 0.028
R7620 S.n2005 S.n2002 0.028
R7621 S.n2842 S.n2839 0.028
R7622 S.n3654 S.n3651 0.028
R7623 S.n4454 S.n4451 0.028
R7624 S.n5231 S.n5228 0.028
R7625 S.n5996 S.n5993 0.028
R7626 S.n3546 S.n3543 0.028
R7627 S.n2734 S.n2731 0.028
R7628 S.n1897 S.n1894 0.028
R7629 S.n1086 S.n1083 0.028
R7630 S.n1131 S.n1128 0.028
R7631 S.n1947 S.n1944 0.028
R7632 S.n2781 S.n2778 0.028
R7633 S.n3593 S.n3590 0.028
R7634 S.n4393 S.n4390 0.028
R7635 S.n1836 S.n1833 0.028
R7636 S.n1027 S.n1024 0.028
R7637 S.n1072 S.n1069 0.028
R7638 S.n1883 S.n1880 0.028
R7639 S.n2720 S.n2717 0.028
R7640 S.n1013 S.n1010 0.028
R7641 S.n2175 S.n2174 0.028
R7642 S.n2177 S.n2175 0.028
R7643 S.n3011 S.n3010 0.028
R7644 S.n3013 S.n3011 0.028
R7645 S.n3823 S.n3822 0.028
R7646 S.n3825 S.n3823 0.028
R7647 S.n4623 S.n4622 0.028
R7648 S.n4625 S.n4623 0.028
R7649 S.n5400 S.n5399 0.028
R7650 S.n5402 S.n5400 0.028
R7651 S.n6165 S.n6164 0.028
R7652 S.n6167 S.n6165 0.028
R7653 S.n6907 S.n6906 0.028
R7654 S.n6909 S.n6907 0.028
R7655 S.n7637 S.n7636 0.028
R7656 S.n7639 S.n7637 0.028
R7657 S.n8344 S.n8343 0.028
R7658 S.n8346 S.n8344 0.028
R7659 S.n9039 S.n9038 0.028
R7660 S.n9041 S.n9039 0.028
R7661 S.n9711 S.n9710 0.028
R7662 S.n9713 S.n9711 0.028
R7663 S.n10371 S.n10370 0.028
R7664 S.n10373 S.n10371 0.028
R7665 S.n11088 S.n11087 0.028
R7666 S.n11090 S.n11088 0.028
R7667 S.n1372 S.n1371 0.028
R7668 S.n1374 S.n1372 0.028
R7669 S.n1400 S.n1399 0.028
R7670 S.n1402 S.n1400 0.028
R7671 S.n974 S.n969 0.028
R7672 S.n987 S.n983 0.028
R7673 S.n2672 S.n2668 0.028
R7674 S.n3514 S.n3510 0.028
R7675 S.n4345 S.n4341 0.028
R7676 S.n5151 S.n5147 0.028
R7677 S.n5948 S.n5944 0.028
R7678 S.n6719 S.n6715 0.028
R7679 S.n7481 S.n7477 0.028
R7680 S.n8217 S.n8213 0.028
R7681 S.n8944 S.n8940 0.028
R7682 S.n9645 S.n9641 0.028
R7683 S.n10337 S.n10333 0.028
R7684 S.n11001 S.n10997 0.028
R7685 S.n11889 S.n11888 0.028
R7686 S.n10467 S.n10466 0.028
R7687 S.n9132 S.n9131 0.028
R7688 S.n7730 S.n7729 0.028
R7689 S.n6258 S.n6257 0.028
R7690 S.n4716 S.n4715 0.028
R7691 S.n3104 S.n3103 0.028
R7692 S.n2148 S.n2147 0.028
R7693 S.n11648 S.n11646 0.027
R7694 S.n12572 S.n12570 0.027
R7695 S.n870 S.n865 0.027
R7696 S.n893 S.n892 0.027
R7697 S.n9813 S.n9812 0.027
R7698 S.n8445 S.n8444 0.027
R7699 S.n7008 S.n7007 0.027
R7700 S.n5502 S.n5501 0.027
R7701 S.n3924 S.n3923 0.027
R7702 S.n2278 S.n2277 0.027
R7703 S.n1826 S.n1825 0.027
R7704 S.n2314 S.n2313 0.027
R7705 S.n3442 S.n3441 0.027
R7706 S.n3961 S.n3960 0.027
R7707 S.n4756 S.n4755 0.027
R7708 S.n5538 S.n5537 0.027
R7709 S.n6298 S.n6297 0.027
R7710 S.n7045 S.n7044 0.027
R7711 S.n8056 S.n8055 0.027
R7712 S.n8768 S.n8767 0.027
R7713 S.n9172 S.n9171 0.027
R7714 S.n9849 S.n9848 0.027
R7715 S.n10507 S.n10506 0.027
R7716 S.n11135 S.n11134 0.027
R7717 S.n12063 S.n12062 0.027
R7718 S.n1678 S.n1677 0.027
R7719 S.n1431 S.n1428 0.026
R7720 S.n1762 S.n1759 0.026
R7721 S.n2250 S.n2247 0.026
R7722 S.n2613 S.n2610 0.026
R7723 S.n3085 S.n3082 0.026
R7724 S.n3377 S.n3374 0.026
R7725 S.n3897 S.n3894 0.026
R7726 S.n4261 S.n4258 0.026
R7727 S.n4697 S.n4694 0.026
R7728 S.n5060 S.n5057 0.026
R7729 S.n5474 S.n5471 0.026
R7730 S.n5841 S.n5838 0.026
R7731 S.n6239 S.n6236 0.026
R7732 S.n6596 S.n6593 0.026
R7733 S.n6981 S.n6978 0.026
R7734 S.n7342 S.n7339 0.026
R7735 S.n7711 S.n7708 0.026
R7736 S.n7895 S.n7892 0.026
R7737 S.n8418 S.n8415 0.026
R7738 S.n8591 S.n8588 0.026
R7739 S.n9113 S.n9110 0.026
R7740 S.n9458 S.n9455 0.026
R7741 S.n9785 S.n9782 0.026
R7742 S.n10134 S.n10131 0.026
R7743 S.n10445 S.n10442 0.026
R7744 S.n10784 S.n10781 0.026
R7745 S.n11075 S.n11072 0.026
R7746 S.n11401 S.n11398 0.026
R7747 S.n12023 S.n12020 0.026
R7748 S.n12303 S.n12300 0.026
R7749 S.n11891 S.n11890 0.026
R7750 S.n787 S.n779 0.026
R7751 S.n1344 S.n1322 0.026
R7752 S.n1702 S.n1690 0.026
R7753 S.n2163 S.n2160 0.026
R7754 S.n2553 S.n2550 0.026
R7755 S.n2999 S.n2996 0.026
R7756 S.n3317 S.n3314 0.026
R7757 S.n3811 S.n3808 0.026
R7758 S.n4201 S.n4198 0.026
R7759 S.n4611 S.n4608 0.026
R7760 S.n5000 S.n4997 0.026
R7761 S.n5388 S.n5385 0.026
R7762 S.n5781 S.n5778 0.026
R7763 S.n6153 S.n6150 0.026
R7764 S.n6536 S.n6533 0.026
R7765 S.n6895 S.n6892 0.026
R7766 S.n7282 S.n7279 0.026
R7767 S.n7625 S.n7622 0.026
R7768 S.n7835 S.n7832 0.026
R7769 S.n8332 S.n8329 0.026
R7770 S.n8531 S.n8528 0.026
R7771 S.n9027 S.n9024 0.026
R7772 S.n9398 S.n9395 0.026
R7773 S.n9699 S.n9696 0.026
R7774 S.n10074 S.n10071 0.026
R7775 S.n10474 S.n10468 0.026
R7776 S.n1712 S.n1710 0.026
R7777 S.n2563 S.n2561 0.026
R7778 S.n3327 S.n3325 0.026
R7779 S.n4211 S.n4209 0.026
R7780 S.n5010 S.n5008 0.026
R7781 S.n5791 S.n5789 0.026
R7782 S.n6546 S.n6544 0.026
R7783 S.n7292 S.n7290 0.026
R7784 S.n7845 S.n7843 0.026
R7785 S.n8541 S.n8539 0.026
R7786 S.n9408 S.n9406 0.026
R7787 S.n10084 S.n10082 0.026
R7788 S.n10734 S.n10732 0.026
R7789 S.n11381 S.n11380 0.026
R7790 S.n10764 S.n10763 0.026
R7791 S.n10114 S.n10113 0.026
R7792 S.n9438 S.n9437 0.026
R7793 S.n8571 S.n8570 0.026
R7794 S.n7875 S.n7874 0.026
R7795 S.n7322 S.n7321 0.026
R7796 S.n6576 S.n6575 0.026
R7797 S.n5821 S.n5820 0.026
R7798 S.n5040 S.n5039 0.026
R7799 S.n4241 S.n4240 0.026
R7800 S.n3357 S.n3356 0.026
R7801 S.n2593 S.n2592 0.026
R7802 S.n1732 S.n1731 0.026
R7803 S.n1406 S.n1389 0.026
R7804 S.n2218 S.n2208 0.026
R7805 S.n3053 S.n3044 0.026
R7806 S.n3865 S.n3856 0.026
R7807 S.n4665 S.n4656 0.026
R7808 S.n5442 S.n5433 0.026
R7809 S.n6207 S.n6198 0.026
R7810 S.n6949 S.n6940 0.026
R7811 S.n7679 S.n7670 0.026
R7812 S.n8386 S.n8377 0.026
R7813 S.n9081 S.n9072 0.026
R7814 S.n9753 S.n9744 0.026
R7815 S.n10413 S.n10404 0.026
R7816 S.n11043 S.n11034 0.026
R7817 S.n12047 S.n12038 0.026
R7818 S.n899 S.n883 0.026
R7819 S.n9816 S.n9800 0.026
R7820 S.n8995 S.n8977 0.026
R7821 S.n8300 S.n8282 0.026
R7822 S.n7593 S.n7575 0.026
R7823 S.n6863 S.n6845 0.026
R7824 S.n6121 S.n6103 0.026
R7825 S.n5356 S.n5338 0.026
R7826 S.n4579 S.n4561 0.026
R7827 S.n3779 S.n3761 0.026
R7828 S.n2967 S.n2949 0.026
R7829 S.n2130 S.n2112 0.026
R7830 S.n1310 S.n1294 0.026
R7831 S.n1282 S.n1277 0.026
R7832 S.n1661 S.n1658 0.026
R7833 S.n2101 S.n2098 0.026
R7834 S.n2517 S.n2514 0.026
R7835 S.n2938 S.n2935 0.026
R7836 S.n3281 S.n3278 0.026
R7837 S.n3750 S.n3747 0.026
R7838 S.n4165 S.n4162 0.026
R7839 S.n4550 S.n4547 0.026
R7840 S.n4964 S.n4961 0.026
R7841 S.n5327 S.n5324 0.026
R7842 S.n5745 S.n5742 0.026
R7843 S.n6092 S.n6089 0.026
R7844 S.n6500 S.n6497 0.026
R7845 S.n6834 S.n6831 0.026
R7846 S.n7246 S.n7243 0.026
R7847 S.n7564 S.n7561 0.026
R7848 S.n7799 S.n7796 0.026
R7849 S.n8271 S.n8268 0.026
R7850 S.n8495 S.n8492 0.026
R7851 S.n9139 S.n9133 0.026
R7852 S.n8449 S.n8433 0.026
R7853 S.n7532 S.n7514 0.026
R7854 S.n6802 S.n6784 0.026
R7855 S.n6060 S.n6042 0.026
R7856 S.n5295 S.n5277 0.026
R7857 S.n4518 S.n4500 0.026
R7858 S.n3718 S.n3700 0.026
R7859 S.n2906 S.n2888 0.026
R7860 S.n2069 S.n2051 0.026
R7861 S.n1252 S.n1235 0.026
R7862 S.n1223 S.n1218 0.026
R7863 S.n1625 S.n1622 0.026
R7864 S.n2040 S.n2037 0.026
R7865 S.n2481 S.n2478 0.026
R7866 S.n2877 S.n2874 0.026
R7867 S.n3245 S.n3242 0.026
R7868 S.n3689 S.n3686 0.026
R7869 S.n4129 S.n4126 0.026
R7870 S.n4489 S.n4486 0.026
R7871 S.n4928 S.n4925 0.026
R7872 S.n5266 S.n5263 0.026
R7873 S.n5709 S.n5706 0.026
R7874 S.n6031 S.n6028 0.026
R7875 S.n6464 S.n6461 0.026
R7876 S.n6773 S.n6770 0.026
R7877 S.n7210 S.n7207 0.026
R7878 S.n7737 S.n7731 0.026
R7879 S.n7012 S.n6996 0.026
R7880 S.n5999 S.n5981 0.026
R7881 S.n5234 S.n5216 0.026
R7882 S.n4457 S.n4439 0.026
R7883 S.n3657 S.n3639 0.026
R7884 S.n2845 S.n2827 0.026
R7885 S.n2008 S.n1990 0.026
R7886 S.n1193 S.n1176 0.026
R7887 S.n1164 S.n1159 0.026
R7888 S.n1589 S.n1586 0.026
R7889 S.n1979 S.n1976 0.026
R7890 S.n2445 S.n2442 0.026
R7891 S.n2816 S.n2813 0.026
R7892 S.n3209 S.n3206 0.026
R7893 S.n3628 S.n3625 0.026
R7894 S.n4093 S.n4090 0.026
R7895 S.n4428 S.n4425 0.026
R7896 S.n4892 S.n4889 0.026
R7897 S.n5205 S.n5202 0.026
R7898 S.n5673 S.n5670 0.026
R7899 S.n6265 S.n6259 0.026
R7900 S.n5505 S.n5489 0.026
R7901 S.n4396 S.n4378 0.026
R7902 S.n3596 S.n3578 0.026
R7903 S.n2784 S.n2766 0.026
R7904 S.n1950 S.n1929 0.026
R7905 S.n1134 S.n1117 0.026
R7906 S.n1105 S.n1100 0.026
R7907 S.n1553 S.n1550 0.026
R7908 S.n1918 S.n1915 0.026
R7909 S.n2409 S.n2406 0.026
R7910 S.n2755 S.n2752 0.026
R7911 S.n3173 S.n3170 0.026
R7912 S.n3567 S.n3564 0.026
R7913 S.n4057 S.n4054 0.026
R7914 S.n4723 S.n4717 0.026
R7915 S.n3928 S.n3912 0.026
R7916 S.n2723 S.n2705 0.026
R7917 S.n1886 S.n1868 0.026
R7918 S.n1075 S.n1058 0.026
R7919 S.n1046 S.n1041 0.026
R7920 S.n1517 S.n1514 0.026
R7921 S.n1857 S.n1854 0.026
R7922 S.n2373 S.n2370 0.026
R7923 S.n3111 S.n3105 0.026
R7924 S.n2281 S.n2265 0.026
R7925 S.n1016 S.n999 0.026
R7926 S.n1455 S.n1449 0.026
R7927 S.n950 S.n945 0.026
R7928 S.n950 S.n934 0.026
R7929 S.n12327 S.n12311 0.026
R7930 S.n837 S.n836 0.026
R7931 S.t7 S.n59 0.025
R7932 S.t7 S.n2 0.025
R7933 S.t7 S.n10 0.025
R7934 S.t7 S.n18 0.025
R7935 S.t7 S.n27 0.025
R7936 S.t7 S.n36 0.025
R7937 S.t7 S.n45 0.025
R7938 S.n187 S.n186 0.024
R7939 S.n989 S.n988 0.024
R7940 S.n2674 S.n2673 0.024
R7941 S.n3508 S.n3507 0.024
R7942 S.n4347 S.n4346 0.024
R7943 S.n5153 S.n5152 0.024
R7944 S.n5950 S.n5949 0.024
R7945 S.n6721 S.n6720 0.024
R7946 S.n7483 S.n7482 0.024
R7947 S.n8219 S.n8218 0.024
R7948 S.n8946 S.n8945 0.024
R7949 S.n9647 S.n9646 0.024
R7950 S.n10339 S.n10338 0.024
R7951 S.n11003 S.n11002 0.024
R7952 S.n11637 S.n11636 0.024
R7953 S.n9683 S.n9678 0.024
R7954 S.n9011 S.n9006 0.024
R7955 S.n8316 S.n8311 0.024
R7956 S.n7609 S.n7604 0.024
R7957 S.n6879 S.n6874 0.024
R7958 S.n6137 S.n6132 0.024
R7959 S.n5372 S.n5367 0.024
R7960 S.n4595 S.n4590 0.024
R7961 S.n3795 S.n3790 0.024
R7962 S.n2983 S.n2978 0.024
R7963 S.n2147 S.n2142 0.024
R7964 S.n2197 S.n2173 0.024
R7965 S.n3033 S.n3009 0.024
R7966 S.n3845 S.n3821 0.024
R7967 S.n4645 S.n4621 0.024
R7968 S.n5422 S.n5398 0.024
R7969 S.n6187 S.n6163 0.024
R7970 S.n6929 S.n6905 0.024
R7971 S.n7659 S.n7635 0.024
R7972 S.n8366 S.n8342 0.024
R7973 S.n9061 S.n9037 0.024
R7974 S.n9733 S.n9709 0.024
R7975 S.n10393 S.n10369 0.024
R7976 S.n11102 S.n11086 0.024
R7977 S.n1406 S.n1405 0.024
R7978 S.n1378 S.n1377 0.024
R7979 S.n1342 S.n1341 0.024
R7980 S.n1825 S.n1824 0.024
R7981 S.n186 S.n185 0.024
R7982 S.n2700 S.n2698 0.023
R7983 S.n12320 S.n12319 0.023
R7984 S.n12609 S.n12596 0.023
R7985 S.n945 S.n942 0.023
R7986 S.n474 S.n473 0.023
R7987 S.n498 S.n494 0.023
R7988 S.n835 S.n832 0.023
R7989 S.n1377 S.n1376 0.023
R7990 S.t7 S.n187 0.023
R7991 S.n11358 S.n11357 0.023
R7992 S.n11086 S.n11085 0.023
R7993 S.n10369 S.n10368 0.023
R7994 S.n9709 S.n9708 0.023
R7995 S.n9037 S.n9036 0.023
R7996 S.n8342 S.n8341 0.023
R7997 S.n7635 S.n7634 0.023
R7998 S.n6905 S.n6904 0.023
R7999 S.n6163 S.n6162 0.023
R8000 S.n5398 S.n5397 0.023
R8001 S.n4621 S.n4620 0.023
R8002 S.n3821 S.n3820 0.023
R8003 S.n3009 S.n3008 0.023
R8004 S.n2173 S.n2172 0.023
R8005 S.n2197 S.n2177 0.023
R8006 S.n3033 S.n3013 0.023
R8007 S.n3845 S.n3825 0.023
R8008 S.n4645 S.n4625 0.023
R8009 S.n5422 S.n5402 0.023
R8010 S.n6187 S.n6167 0.023
R8011 S.n6929 S.n6909 0.023
R8012 S.n7659 S.n7639 0.023
R8013 S.n8366 S.n8346 0.023
R8014 S.n9061 S.n9041 0.023
R8015 S.n9733 S.n9713 0.023
R8016 S.n10393 S.n10373 0.023
R8017 S.n11102 S.n11090 0.023
R8018 S.n748 S.n746 0.023
R8019 S.n1405 S.n1404 0.023
R8020 S.n894 S.n893 0.023
R8021 S.n1406 S.n1402 0.023
R8022 S.n1378 S.n1374 0.023
R8023 S.n475 S.n471 0.023
R8024 S.n430 S.n429 0.023
R8025 S.n454 S.n450 0.023
R8026 S.n8446 S.n8445 0.023
R8027 S.n431 S.n427 0.023
R8028 S.n386 S.n385 0.023
R8029 S.n410 S.n406 0.023
R8030 S.n7009 S.n7008 0.023
R8031 S.n387 S.n383 0.023
R8032 S.n342 S.n341 0.023
R8033 S.n366 S.n362 0.023
R8034 S.n343 S.n339 0.023
R8035 S.n298 S.n297 0.023
R8036 S.n322 S.n318 0.023
R8037 S.n3925 S.n3924 0.023
R8038 S.n299 S.n295 0.023
R8039 S.n254 S.n253 0.023
R8040 S.n278 S.n274 0.023
R8041 S.n255 S.n251 0.023
R8042 S.n993 S.n991 0.023
R8043 S.n1823 S.n1822 0.023
R8044 S.n1831 S.n1829 0.023
R8045 S.n2683 S.n2682 0.023
R8046 S.n3524 S.n3523 0.023
R8047 S.n3541 S.n3539 0.023
R8048 S.n4356 S.n4355 0.023
R8049 S.n4373 S.n4371 0.023
R8050 S.n5162 S.n5161 0.023
R8051 S.n5179 S.n5177 0.023
R8052 S.n5959 S.n5958 0.023
R8053 S.n5976 S.n5974 0.023
R8054 S.n6730 S.n6729 0.023
R8055 S.n6747 S.n6745 0.023
R8056 S.n7492 S.n7491 0.023
R8057 S.n7509 S.n7507 0.023
R8058 S.n8228 S.n8227 0.023
R8059 S.n8245 S.n8243 0.023
R8060 S.n8955 S.n8954 0.023
R8061 S.n8972 S.n8970 0.023
R8062 S.n9656 S.n9655 0.023
R8063 S.n9673 S.n9671 0.023
R8064 S.n10348 S.n10347 0.023
R8065 S.n10365 S.n10363 0.023
R8066 S.n11012 S.n11011 0.023
R8067 S.n11029 S.n11027 0.023
R8068 S.n9678 S.n9675 0.023
R8069 S.n9006 S.n9003 0.023
R8070 S.n8311 S.n8308 0.023
R8071 S.n7604 S.n7601 0.023
R8072 S.n6874 S.n6872 0.023
R8073 S.n6132 S.n6129 0.023
R8074 S.n5367 S.n5364 0.023
R8075 S.n4590 S.n4588 0.023
R8076 S.n3790 S.n3787 0.023
R8077 S.n2978 S.n2976 0.023
R8078 S.n2142 S.n2139 0.023
R8079 S.n1341 S.n1338 0.023
R8080 S.n1333 S.n1332 0.023
R8081 S.n1332 S.n1331 0.022
R8082 S.n10388 S.n10384 0.022
R8083 S.n9728 S.n9724 0.022
R8084 S.n9056 S.n9052 0.022
R8085 S.n8361 S.n8357 0.022
R8086 S.n7654 S.n7650 0.022
R8087 S.n6924 S.n6920 0.022
R8088 S.n6182 S.n6178 0.022
R8089 S.n5417 S.n5413 0.022
R8090 S.n4640 S.n4636 0.022
R8091 S.n3840 S.n3836 0.022
R8092 S.n3028 S.n3024 0.022
R8093 S.n2192 S.n2188 0.022
R8094 S.n1357 S.n1353 0.022
R8095 S.n849 S.n845 0.022
R8096 S.n12033 S.n12032 0.022
R8097 S.n2692 S.n2690 0.022
R8098 S.n3533 S.n3531 0.022
R8099 S.n4365 S.n4363 0.022
R8100 S.n5171 S.n5169 0.022
R8101 S.n5968 S.n5966 0.022
R8102 S.n6739 S.n6737 0.022
R8103 S.n7501 S.n7499 0.022
R8104 S.n8237 S.n8235 0.022
R8105 S.n8964 S.n8962 0.022
R8106 S.n9665 S.n9663 0.022
R8107 S.n10357 S.n10355 0.022
R8108 S.n11021 S.n11019 0.022
R8109 S.n10472 S.n10471 0.022
R8110 S.n9795 S.n9793 0.022
R8111 S.n9137 S.n9136 0.022
R8112 S.n8428 S.n8426 0.022
R8113 S.n7735 S.n7734 0.022
R8114 S.n6991 S.n6989 0.022
R8115 S.n6263 S.n6262 0.022
R8116 S.n5484 S.n5482 0.022
R8117 S.n4721 S.n4720 0.022
R8118 S.n3907 S.n3905 0.022
R8119 S.n3109 S.n3108 0.022
R8120 S.n2260 S.n2258 0.022
R8121 S.n1453 S.n1452 0.022
R8122 S.n929 S.n927 0.022
R8123 S.n12037 S.n12036 0.022
R8124 S.n1426 S.n1425 0.021
R8125 S.n1422 S.n1421 0.021
R8126 S.n2245 S.n2244 0.021
R8127 S.n2243 S.n2242 0.021
R8128 S.n3080 S.n3079 0.021
R8129 S.n3078 S.n3077 0.021
R8130 S.n3892 S.n3891 0.021
R8131 S.n3890 S.n3889 0.021
R8132 S.n4692 S.n4691 0.021
R8133 S.n4690 S.n4689 0.021
R8134 S.n5469 S.n5468 0.021
R8135 S.n5467 S.n5466 0.021
R8136 S.n6234 S.n6233 0.021
R8137 S.n6232 S.n6231 0.021
R8138 S.n6976 S.n6975 0.021
R8139 S.n6974 S.n6973 0.021
R8140 S.n7706 S.n7705 0.021
R8141 S.n7704 S.n7703 0.021
R8142 S.n8413 S.n8412 0.021
R8143 S.n8411 S.n8410 0.021
R8144 S.n9108 S.n9107 0.021
R8145 S.n9106 S.n9105 0.021
R8146 S.n9780 S.n9779 0.021
R8147 S.n9778 S.n9777 0.021
R8148 S.n10440 S.n10439 0.021
R8149 S.n10438 S.n10437 0.021
R8150 S.n11070 S.n11069 0.021
R8151 S.n11068 S.n11067 0.021
R8152 S.n12018 S.n12017 0.021
R8153 S.n12016 S.n12015 0.021
R8154 S.n11888 S.n11887 0.021
R8155 S.n909 S.n908 0.021
R8156 S.n1319 S.n1318 0.021
R8157 S.n2158 S.n2157 0.021
R8158 S.n2156 S.n2155 0.021
R8159 S.n2994 S.n2993 0.021
R8160 S.n2992 S.n2991 0.021
R8161 S.n3806 S.n3805 0.021
R8162 S.n3804 S.n3803 0.021
R8163 S.n4606 S.n4605 0.021
R8164 S.n4604 S.n4603 0.021
R8165 S.n5383 S.n5382 0.021
R8166 S.n5381 S.n5380 0.021
R8167 S.n6148 S.n6147 0.021
R8168 S.n6146 S.n6145 0.021
R8169 S.n6890 S.n6889 0.021
R8170 S.n6888 S.n6887 0.021
R8171 S.n7620 S.n7619 0.021
R8172 S.n7618 S.n7617 0.021
R8173 S.n8327 S.n8326 0.021
R8174 S.n8325 S.n8324 0.021
R8175 S.n9022 S.n9021 0.021
R8176 S.n9020 S.n9019 0.021
R8177 S.n9694 S.n9693 0.021
R8178 S.n9692 S.n9691 0.021
R8179 S.n10466 S.n10465 0.021
R8180 S.n1280 S.n1279 0.021
R8181 S.n2096 S.n2095 0.021
R8182 S.n2094 S.n2093 0.021
R8183 S.n2933 S.n2932 0.021
R8184 S.n2931 S.n2930 0.021
R8185 S.n3745 S.n3744 0.021
R8186 S.n3743 S.n3742 0.021
R8187 S.n4545 S.n4544 0.021
R8188 S.n4543 S.n4542 0.021
R8189 S.n5322 S.n5321 0.021
R8190 S.n5320 S.n5319 0.021
R8191 S.n6087 S.n6086 0.021
R8192 S.n6085 S.n6084 0.021
R8193 S.n6829 S.n6828 0.021
R8194 S.n6827 S.n6826 0.021
R8195 S.n7559 S.n7558 0.021
R8196 S.n7557 S.n7556 0.021
R8197 S.n8266 S.n8265 0.021
R8198 S.n8264 S.n8263 0.021
R8199 S.n9131 S.n9130 0.021
R8200 S.n1221 S.n1220 0.021
R8201 S.n2035 S.n2034 0.021
R8202 S.n2033 S.n2032 0.021
R8203 S.n2872 S.n2871 0.021
R8204 S.n2870 S.n2869 0.021
R8205 S.n3684 S.n3683 0.021
R8206 S.n3682 S.n3681 0.021
R8207 S.n4484 S.n4483 0.021
R8208 S.n4482 S.n4481 0.021
R8209 S.n5261 S.n5260 0.021
R8210 S.n5259 S.n5258 0.021
R8211 S.n6026 S.n6025 0.021
R8212 S.n6024 S.n6023 0.021
R8213 S.n6768 S.n6767 0.021
R8214 S.n6766 S.n6765 0.021
R8215 S.n7729 S.n7728 0.021
R8216 S.n1162 S.n1161 0.021
R8217 S.n1974 S.n1973 0.021
R8218 S.n1972 S.n1971 0.021
R8219 S.n2811 S.n2810 0.021
R8220 S.n2809 S.n2808 0.021
R8221 S.n3623 S.n3622 0.021
R8222 S.n3621 S.n3620 0.021
R8223 S.n4423 S.n4422 0.021
R8224 S.n4421 S.n4420 0.021
R8225 S.n5200 S.n5199 0.021
R8226 S.n5198 S.n5197 0.021
R8227 S.n6257 S.n6256 0.021
R8228 S.n1103 S.n1102 0.021
R8229 S.n1913 S.n1912 0.021
R8230 S.n1911 S.n1910 0.021
R8231 S.n2750 S.n2749 0.021
R8232 S.n2748 S.n2747 0.021
R8233 S.n3562 S.n3561 0.021
R8234 S.n3560 S.n3559 0.021
R8235 S.n4715 S.n4714 0.021
R8236 S.n1044 S.n1043 0.021
R8237 S.n1852 S.n1851 0.021
R8238 S.n1850 S.n1849 0.021
R8239 S.n3103 S.n3102 0.021
R8240 S.n11361 S.n11360 0.021
R8241 S.n12001 S.n12000 0.021
R8242 S.n11053 S.n11052 0.021
R8243 S.n10423 S.n10422 0.021
R8244 S.n9763 S.n9762 0.021
R8245 S.n9091 S.n9090 0.021
R8246 S.n8396 S.n8395 0.021
R8247 S.n7689 S.n7688 0.021
R8248 S.n6959 S.n6958 0.021
R8249 S.n6217 S.n6216 0.021
R8250 S.n5452 S.n5451 0.021
R8251 S.n4675 S.n4674 0.021
R8252 S.n3875 S.n3874 0.021
R8253 S.n3063 S.n3062 0.021
R8254 S.n2228 S.n2227 0.021
R8255 S.n907 S.n906 0.021
R8256 S.n8249 S.n8248 0.021
R8257 S.n7542 S.n7541 0.021
R8258 S.n6812 S.n6811 0.021
R8259 S.n6070 S.n6069 0.021
R8260 S.n5305 S.n5304 0.021
R8261 S.n4528 S.n4527 0.021
R8262 S.n3728 S.n3727 0.021
R8263 S.n2916 S.n2915 0.021
R8264 S.n2079 S.n2078 0.021
R8265 S.n1262 S.n1261 0.021
R8266 S.n10473 S.n10472 0.021
R8267 S.n11101 S.n11100 0.021
R8268 S.n1306 S.n1305 0.021
R8269 S.n2126 S.n2125 0.021
R8270 S.n2963 S.n2962 0.021
R8271 S.n3775 S.n3774 0.021
R8272 S.n4575 S.n4574 0.021
R8273 S.n5352 S.n5351 0.021
R8274 S.n6117 S.n6116 0.021
R8275 S.n6859 S.n6858 0.021
R8276 S.n7589 S.n7588 0.021
R8277 S.n8296 S.n8295 0.021
R8278 S.n8991 S.n8990 0.021
R8279 S.n9797 S.n9795 0.021
R8280 S.n492 S.n491 0.021
R8281 S.n9138 S.n9137 0.021
R8282 S.n6751 S.n6750 0.021
R8283 S.n6009 S.n6008 0.021
R8284 S.n5244 S.n5243 0.021
R8285 S.n4467 S.n4466 0.021
R8286 S.n3667 S.n3666 0.021
R8287 S.n2855 S.n2854 0.021
R8288 S.n2018 S.n2017 0.021
R8289 S.n1203 S.n1202 0.021
R8290 S.n1248 S.n1247 0.021
R8291 S.n2065 S.n2064 0.021
R8292 S.n2902 S.n2901 0.021
R8293 S.n3714 S.n3713 0.021
R8294 S.n4514 S.n4513 0.021
R8295 S.n5291 S.n5290 0.021
R8296 S.n6056 S.n6055 0.021
R8297 S.n6798 S.n6797 0.021
R8298 S.n7528 S.n7527 0.021
R8299 S.n8430 S.n8428 0.021
R8300 S.n448 S.n447 0.021
R8301 S.n7736 S.n7735 0.021
R8302 S.n5183 S.n5182 0.021
R8303 S.n4406 S.n4405 0.021
R8304 S.n3606 S.n3605 0.021
R8305 S.n2794 S.n2793 0.021
R8306 S.n1957 S.n1956 0.021
R8307 S.n1144 S.n1143 0.021
R8308 S.n1189 S.n1188 0.021
R8309 S.n2004 S.n2003 0.021
R8310 S.n2841 S.n2840 0.021
R8311 S.n3653 S.n3652 0.021
R8312 S.n4453 S.n4452 0.021
R8313 S.n5230 S.n5229 0.021
R8314 S.n5995 S.n5994 0.021
R8315 S.n6993 S.n6991 0.021
R8316 S.n404 S.n403 0.021
R8317 S.n6264 S.n6263 0.021
R8318 S.n3545 S.n3544 0.021
R8319 S.n2733 S.n2732 0.021
R8320 S.n1896 S.n1895 0.021
R8321 S.n1085 S.n1084 0.021
R8322 S.n1130 S.n1129 0.021
R8323 S.n1946 S.n1945 0.021
R8324 S.n2780 S.n2779 0.021
R8325 S.n3592 S.n3591 0.021
R8326 S.n4392 S.n4391 0.021
R8327 S.n5486 S.n5484 0.021
R8328 S.n360 S.n359 0.021
R8329 S.n4722 S.n4721 0.021
R8330 S.n1835 S.n1834 0.021
R8331 S.n1026 S.n1025 0.021
R8332 S.n1071 S.n1070 0.021
R8333 S.n1882 S.n1881 0.021
R8334 S.n2719 S.n2718 0.021
R8335 S.n3909 S.n3907 0.021
R8336 S.n316 S.n315 0.021
R8337 S.n3110 S.n3109 0.021
R8338 S.n1012 S.n1011 0.021
R8339 S.n2262 S.n2260 0.021
R8340 S.n272 S.n271 0.021
R8341 S.n1454 S.n1453 0.021
R8342 S.n931 S.n929 0.021
R8343 S.n11643 S.n11642 0.021
R8344 S.n881 S.n880 0.02
R8345 S.n496 S.n495 0.02
R8346 S.n452 S.n451 0.02
R8347 S.n408 S.n407 0.02
R8348 S.n364 S.n363 0.02
R8349 S.n320 S.n319 0.02
R8350 S.n276 S.n275 0.02
R8351 S.n948 S.n947 0.02
R8352 S.n11901 S.n11900 0.02
R8353 S.n9678 S.n9677 0.02
R8354 S.n9006 S.n9005 0.02
R8355 S.n8311 S.n8310 0.02
R8356 S.n7604 S.n7603 0.02
R8357 S.n6874 S.n6873 0.02
R8358 S.n6132 S.n6131 0.02
R8359 S.n5367 S.n5366 0.02
R8360 S.n4590 S.n4589 0.02
R8361 S.n3790 S.n3789 0.02
R8362 S.n2978 S.n2977 0.02
R8363 S.n2142 S.n2141 0.02
R8364 S.n10473 S.n10469 0.02
R8365 S.n12034 S.n12031 0.02
R8366 S.n1341 S.n1340 0.02
R8367 S.n9797 S.n9796 0.02
R8368 S.n9138 S.n9134 0.02
R8369 S.n8430 S.n8429 0.02
R8370 S.n7736 S.n7732 0.02
R8371 S.n6993 S.n6992 0.02
R8372 S.n6264 S.n6260 0.02
R8373 S.n5486 S.n5485 0.02
R8374 S.n4722 S.n4718 0.02
R8375 S.n3909 S.n3908 0.02
R8376 S.n3110 S.n3106 0.02
R8377 S.n2262 S.n2261 0.02
R8378 S.n1454 S.n1450 0.02
R8379 S.n931 S.n930 0.02
R8380 S.n898 S.n897 0.02
R8381 S.t7 S.n173 0.019
R8382 S.n1715 S.n1713 0.019
R8383 S.n2566 S.n2564 0.019
R8384 S.n3330 S.n3328 0.019
R8385 S.n4214 S.n4212 0.019
R8386 S.n5013 S.n5011 0.019
R8387 S.n5794 S.n5792 0.019
R8388 S.n6549 S.n6547 0.019
R8389 S.n7295 S.n7293 0.019
R8390 S.n7848 S.n7846 0.019
R8391 S.n8544 S.n8542 0.019
R8392 S.n9411 S.n9409 0.019
R8393 S.n10087 S.n10085 0.019
R8394 S.n10737 S.n10735 0.019
R8395 S.n856 S.n855 0.019
R8396 S.n1734 S.n1733 0.019
R8397 S.n10392 S.n10391 0.019
R8398 S.n9732 S.n9731 0.019
R8399 S.n9060 S.n9059 0.019
R8400 S.n8365 S.n8364 0.019
R8401 S.n7658 S.n7657 0.019
R8402 S.n6928 S.n6927 0.019
R8403 S.n6186 S.n6185 0.019
R8404 S.n5421 S.n5420 0.019
R8405 S.n4644 S.n4643 0.019
R8406 S.n3844 S.n3843 0.019
R8407 S.n3032 S.n3031 0.019
R8408 S.n2196 S.n2195 0.019
R8409 S.n1361 S.n1360 0.019
R8410 S.n12274 S.n12273 0.019
R8411 S.n867 S.n866 0.018
R8412 S.n974 S.n973 0.018
R8413 S.n987 S.n986 0.018
R8414 S.n2672 S.n2671 0.018
R8415 S.n3514 S.n3513 0.018
R8416 S.n4345 S.n4344 0.018
R8417 S.n5151 S.n5150 0.018
R8418 S.n5948 S.n5947 0.018
R8419 S.n6719 S.n6718 0.018
R8420 S.n7481 S.n7480 0.018
R8421 S.n8217 S.n8216 0.018
R8422 S.n8944 S.n8943 0.018
R8423 S.n9645 S.n9644 0.018
R8424 S.n10337 S.n10336 0.018
R8425 S.n11001 S.n11000 0.018
R8426 S.n173 S.n172 0.018
R8427 S.n494 S.n493 0.018
R8428 S.n471 S.n470 0.018
R8429 S.n450 S.n449 0.018
R8430 S.n427 S.n426 0.018
R8431 S.n406 S.n405 0.018
R8432 S.n383 S.n382 0.018
R8433 S.n362 S.n361 0.018
R8434 S.n339 S.n338 0.018
R8435 S.n318 S.n317 0.018
R8436 S.n295 S.n294 0.018
R8437 S.n274 S.n273 0.018
R8438 S.n251 S.n250 0.018
R8439 S.n11596 S.n11595 0.018
R8440 S.n177 S.n176 0.018
R8441 S.n1340 S.n1339 0.018
R8442 S.n9677 S.n9676 0.018
R8443 S.n9005 S.n9004 0.018
R8444 S.n8310 S.n8309 0.018
R8445 S.n7603 S.n7602 0.018
R8446 S.n6131 S.n6130 0.018
R8447 S.n5366 S.n5365 0.018
R8448 S.n3789 S.n3788 0.018
R8449 S.n2141 S.n2140 0.018
R8450 S.n11593 S.n11592 0.017
R8451 S.n11600 S.n11597 0.017
R8452 S.n12606 S.n12605 0.017
R8453 S.n12605 S.n12604 0.017
R8454 S.n2695 S.n2694 0.017
R8455 S.n3536 S.n3535 0.017
R8456 S.n4368 S.n4367 0.017
R8457 S.n5174 S.n5173 0.017
R8458 S.n5971 S.n5970 0.017
R8459 S.n6742 S.n6741 0.017
R8460 S.n7504 S.n7503 0.017
R8461 S.n8240 S.n8239 0.017
R8462 S.n8967 S.n8966 0.017
R8463 S.n9668 S.n9667 0.017
R8464 S.n10360 S.n10359 0.017
R8465 S.n11024 S.n11023 0.017
R8466 S.n1344 S.n1333 0.016
R8467 S.n1702 S.n1698 0.016
R8468 S.n9816 S.n9808 0.016
R8469 S.n8449 S.n8441 0.016
R8470 S.n7012 S.n7004 0.016
R8471 S.n5505 S.n5497 0.016
R8472 S.n3928 S.n3920 0.016
R8473 S.n2281 S.n2273 0.016
R8474 S.n2693 S.n2692 0.016
R8475 S.n3534 S.n3533 0.016
R8476 S.n4366 S.n4365 0.016
R8477 S.n5172 S.n5171 0.016
R8478 S.n5969 S.n5968 0.016
R8479 S.n6740 S.n6739 0.016
R8480 S.n7502 S.n7501 0.016
R8481 S.n8238 S.n8237 0.016
R8482 S.n8965 S.n8964 0.016
R8483 S.n9666 S.n9665 0.016
R8484 S.n10358 S.n10357 0.016
R8485 S.n11022 S.n11021 0.016
R8486 S.n6872 S.n6871 0.015
R8487 S.n4588 S.n4587 0.015
R8488 S.n2976 S.n2975 0.015
R8489 S.n12570 S.n12569 0.015
R8490 S.n1344 S.n1343 0.015
R8491 S.n10390 S.n10389 0.015
R8492 S.n10389 S.n10388 0.015
R8493 S.n10388 S.n10387 0.015
R8494 S.n9730 S.n9729 0.015
R8495 S.n9729 S.n9728 0.015
R8496 S.n9728 S.n9727 0.015
R8497 S.n9058 S.n9057 0.015
R8498 S.n9057 S.n9056 0.015
R8499 S.n9056 S.n9055 0.015
R8500 S.n8363 S.n8362 0.015
R8501 S.n8362 S.n8361 0.015
R8502 S.n8361 S.n8360 0.015
R8503 S.n7656 S.n7655 0.015
R8504 S.n7655 S.n7654 0.015
R8505 S.n7654 S.n7653 0.015
R8506 S.n6926 S.n6925 0.015
R8507 S.n6925 S.n6924 0.015
R8508 S.n6924 S.n6923 0.015
R8509 S.n6184 S.n6183 0.015
R8510 S.n6183 S.n6182 0.015
R8511 S.n6182 S.n6181 0.015
R8512 S.n5419 S.n5418 0.015
R8513 S.n5418 S.n5417 0.015
R8514 S.n5417 S.n5416 0.015
R8515 S.n4642 S.n4641 0.015
R8516 S.n4641 S.n4640 0.015
R8517 S.n4640 S.n4639 0.015
R8518 S.n3842 S.n3841 0.015
R8519 S.n3841 S.n3840 0.015
R8520 S.n3840 S.n3839 0.015
R8521 S.n3030 S.n3029 0.015
R8522 S.n3029 S.n3028 0.015
R8523 S.n3028 S.n3027 0.015
R8524 S.n2194 S.n2193 0.015
R8525 S.n2193 S.n2192 0.015
R8526 S.n2192 S.n2191 0.015
R8527 S.n1359 S.n1358 0.015
R8528 S.n1358 S.n1357 0.015
R8529 S.n1357 S.n1356 0.015
R8530 S.n850 S.n849 0.015
R8531 S.n849 S.n848 0.015
R8532 S.n12036 S.n12035 0.015
R8533 S.n896 S.n895 0.015
R8534 S.n2696 S.n2676 0.015
R8535 S.n3537 S.n3517 0.015
R8536 S.n4369 S.n4349 0.015
R8537 S.n5175 S.n5155 0.015
R8538 S.n5972 S.n5952 0.015
R8539 S.n6743 S.n6723 0.015
R8540 S.n7505 S.n7485 0.015
R8541 S.n8241 S.n8221 0.015
R8542 S.n8968 S.n8948 0.015
R8543 S.n9669 S.n9649 0.015
R8544 S.n10361 S.n10341 0.015
R8545 S.n11025 S.n11005 0.015
R8546 S.n12272 S.n12271 0.015
R8547 S.n12271 S.n12270 0.015
R8548 S.n11595 S.n11594 0.015
R8549 S.n11644 S.n11639 0.015
R8550 S.n12004 S.n12003 0.015
R8551 S.n11056 S.n11055 0.015
R8552 S.n10426 S.n10425 0.015
R8553 S.n9766 S.n9765 0.015
R8554 S.n9094 S.n9093 0.015
R8555 S.n8399 S.n8398 0.015
R8556 S.n7692 S.n7691 0.015
R8557 S.n6962 S.n6961 0.015
R8558 S.n6220 S.n6219 0.015
R8559 S.n5455 S.n5454 0.015
R8560 S.n4678 S.n4677 0.015
R8561 S.n3878 S.n3877 0.015
R8562 S.n3066 S.n3065 0.015
R8563 S.n2231 S.n2230 0.015
R8564 S.n8252 S.n8251 0.015
R8565 S.n7545 S.n7544 0.015
R8566 S.n6815 S.n6814 0.015
R8567 S.n6073 S.n6072 0.015
R8568 S.n5308 S.n5307 0.015
R8569 S.n4531 S.n4530 0.015
R8570 S.n3731 S.n3730 0.015
R8571 S.n2919 S.n2918 0.015
R8572 S.n2082 S.n2081 0.015
R8573 S.n1265 S.n1264 0.015
R8574 S.n8986 S.n8985 0.015
R8575 S.n8291 S.n8290 0.015
R8576 S.n7584 S.n7583 0.015
R8577 S.n6854 S.n6853 0.015
R8578 S.n6112 S.n6111 0.015
R8579 S.n5347 S.n5346 0.015
R8580 S.n4570 S.n4569 0.015
R8581 S.n3770 S.n3769 0.015
R8582 S.n2958 S.n2957 0.015
R8583 S.n2121 S.n2120 0.015
R8584 S.n1302 S.n1301 0.015
R8585 S.n6754 S.n6753 0.015
R8586 S.n6012 S.n6011 0.015
R8587 S.n5247 S.n5246 0.015
R8588 S.n4470 S.n4469 0.015
R8589 S.n3670 S.n3669 0.015
R8590 S.n2858 S.n2857 0.015
R8591 S.n2021 S.n2020 0.015
R8592 S.n1206 S.n1205 0.015
R8593 S.n7523 S.n7522 0.015
R8594 S.n6793 S.n6792 0.015
R8595 S.n6051 S.n6050 0.015
R8596 S.n5286 S.n5285 0.015
R8597 S.n4509 S.n4508 0.015
R8598 S.n3709 S.n3708 0.015
R8599 S.n2897 S.n2896 0.015
R8600 S.n2060 S.n2059 0.015
R8601 S.n1243 S.n1242 0.015
R8602 S.n5186 S.n5185 0.015
R8603 S.n4409 S.n4408 0.015
R8604 S.n3609 S.n3608 0.015
R8605 S.n2797 S.n2796 0.015
R8606 S.n1960 S.n1959 0.015
R8607 S.n1147 S.n1146 0.015
R8608 S.n5990 S.n5989 0.015
R8609 S.n5225 S.n5224 0.015
R8610 S.n4448 S.n4447 0.015
R8611 S.n3648 S.n3647 0.015
R8612 S.n2836 S.n2835 0.015
R8613 S.n1999 S.n1998 0.015
R8614 S.n1184 S.n1183 0.015
R8615 S.n3548 S.n3547 0.015
R8616 S.n2736 S.n2735 0.015
R8617 S.n1899 S.n1898 0.015
R8618 S.n1088 S.n1087 0.015
R8619 S.n4387 S.n4386 0.015
R8620 S.n3587 S.n3586 0.015
R8621 S.n2775 S.n2774 0.015
R8622 S.n1941 S.n1940 0.015
R8623 S.n1125 S.n1124 0.015
R8624 S.n1838 S.n1837 0.015
R8625 S.n1029 S.n1028 0.015
R8626 S.n2714 S.n2713 0.015
R8627 S.n1877 S.n1876 0.015
R8628 S.n1066 S.n1065 0.015
R8629 S.n1007 S.n1006 0.015
R8630 S.n853 S.n852 0.014
R8631 S.n11633 S.n11631 0.014
R8632 S.n1269 S.n1268 0.014
R8633 S.n2129 S.n2128 0.014
R8634 S.n2966 S.n2965 0.014
R8635 S.n3778 S.n3777 0.014
R8636 S.n4578 S.n4577 0.014
R8637 S.n5355 S.n5354 0.014
R8638 S.n6120 S.n6119 0.014
R8639 S.n6862 S.n6861 0.014
R8640 S.n7592 S.n7591 0.014
R8641 S.n8299 S.n8298 0.014
R8642 S.n8994 S.n8993 0.014
R8643 S.n1210 S.n1209 0.014
R8644 S.n2068 S.n2067 0.014
R8645 S.n2905 S.n2904 0.014
R8646 S.n3717 S.n3716 0.014
R8647 S.n4517 S.n4516 0.014
R8648 S.n5294 S.n5293 0.014
R8649 S.n6059 S.n6058 0.014
R8650 S.n6801 S.n6800 0.014
R8651 S.n7531 S.n7530 0.014
R8652 S.n1151 S.n1150 0.014
R8653 S.n2007 S.n2006 0.014
R8654 S.n2844 S.n2843 0.014
R8655 S.n3656 S.n3655 0.014
R8656 S.n4456 S.n4455 0.014
R8657 S.n5233 S.n5232 0.014
R8658 S.n5998 S.n5997 0.014
R8659 S.n1092 S.n1091 0.014
R8660 S.n1949 S.n1948 0.014
R8661 S.n2783 S.n2782 0.014
R8662 S.n3595 S.n3594 0.014
R8663 S.n4395 S.n4394 0.014
R8664 S.n1033 S.n1032 0.014
R8665 S.n1885 S.n1884 0.014
R8666 S.n2722 S.n2721 0.014
R8667 S.n11657 S.n11648 0.014
R8668 S.n12582 S.n12572 0.014
R8669 S.n1343 S.n1342 0.014
R8670 S.n1679 S.n1678 0.014
R8671 S.n2633 S.n2632 0.014
R8672 S.n4297 S.n4296 0.014
R8673 S.n5112 S.n5111 0.014
R8674 S.n5909 S.n5908 0.014
R8675 S.n6680 S.n6679 0.014
R8676 S.n7442 S.n7441 0.014
R8677 S.n8026 S.n8025 0.014
R8678 S.n8738 S.n8737 0.014
R8679 S.n9606 S.n9605 0.014
R8680 S.n10298 S.n10297 0.014
R8681 S.n10964 S.n10963 0.014
R8682 S.n12326 S.n12325 0.014
R8683 S.n3412 S.n3411 0.014
R8684 S.n12008 S.n12007 0.013
R8685 S.n11060 S.n11059 0.013
R8686 S.n10430 S.n10429 0.013
R8687 S.n9770 S.n9769 0.013
R8688 S.n9098 S.n9097 0.013
R8689 S.n8403 S.n8402 0.013
R8690 S.n7696 S.n7695 0.013
R8691 S.n6966 S.n6965 0.013
R8692 S.n6224 S.n6223 0.013
R8693 S.n5459 S.n5458 0.013
R8694 S.n4682 S.n4681 0.013
R8695 S.n3882 S.n3881 0.013
R8696 S.n3070 S.n3069 0.013
R8697 S.n2235 S.n2234 0.013
R8698 S.n8256 S.n8255 0.013
R8699 S.n7549 S.n7548 0.013
R8700 S.n6819 S.n6818 0.013
R8701 S.n6077 S.n6076 0.013
R8702 S.n5312 S.n5311 0.013
R8703 S.n4535 S.n4534 0.013
R8704 S.n3735 S.n3734 0.013
R8705 S.n2923 S.n2922 0.013
R8706 S.n2086 S.n2085 0.013
R8707 S.n1309 S.n1308 0.013
R8708 S.n6758 S.n6757 0.013
R8709 S.n6016 S.n6015 0.013
R8710 S.n5251 S.n5250 0.013
R8711 S.n4474 S.n4473 0.013
R8712 S.n3674 S.n3673 0.013
R8713 S.n2862 S.n2861 0.013
R8714 S.n2025 S.n2024 0.013
R8715 S.n1251 S.n1250 0.013
R8716 S.n5190 S.n5189 0.013
R8717 S.n4413 S.n4412 0.013
R8718 S.n3613 S.n3612 0.013
R8719 S.n2801 S.n2800 0.013
R8720 S.n1964 S.n1963 0.013
R8721 S.n1192 S.n1191 0.013
R8722 S.n3552 S.n3551 0.013
R8723 S.n2740 S.n2739 0.013
R8724 S.n1903 S.n1902 0.013
R8725 S.n1133 S.n1132 0.013
R8726 S.n1842 S.n1841 0.013
R8727 S.n1074 S.n1073 0.013
R8728 S.n1015 S.n1014 0.013
R8729 S.n11099 S.n11098 0.013
R8730 S.n2632 S.n2631 0.013
R8731 S.n3411 S.n3410 0.013
R8732 S.n4296 S.n4295 0.013
R8733 S.n5111 S.n5110 0.013
R8734 S.n5908 S.n5907 0.013
R8735 S.n6679 S.n6678 0.013
R8736 S.n7441 S.n7440 0.013
R8737 S.n8025 S.n8024 0.013
R8738 S.n8737 S.n8736 0.013
R8739 S.n9605 S.n9604 0.013
R8740 S.n10297 S.n10296 0.013
R8741 S.n10963 S.n10962 0.013
R8742 S.n12325 S.n12324 0.013
R8743 S.t7 S.n0 0.012
R8744 S.t7 S.n8 0.012
R8745 S.t7 S.n16 0.012
R8746 S.t7 S.n25 0.012
R8747 S.t7 S.n34 0.012
R8748 S.t7 S.n43 0.012
R8749 S.t7 S.n60 0.012
R8750 S.n11639 S.n11635 0.012
R8751 S.n12602 S.n12601 0.012
R8752 S.n12005 S.n12004 0.012
R8753 S.n11057 S.n11056 0.012
R8754 S.n10427 S.n10426 0.012
R8755 S.n9767 S.n9766 0.012
R8756 S.n9095 S.n9094 0.012
R8757 S.n8400 S.n8399 0.012
R8758 S.n7693 S.n7692 0.012
R8759 S.n6963 S.n6962 0.012
R8760 S.n6221 S.n6220 0.012
R8761 S.n5456 S.n5455 0.012
R8762 S.n4679 S.n4678 0.012
R8763 S.n3879 S.n3878 0.012
R8764 S.n3067 S.n3066 0.012
R8765 S.n2232 S.n2231 0.012
R8766 S.n920 S.n911 0.012
R8767 S.n8253 S.n8252 0.012
R8768 S.n7546 S.n7545 0.012
R8769 S.n6816 S.n6815 0.012
R8770 S.n6074 S.n6073 0.012
R8771 S.n5309 S.n5308 0.012
R8772 S.n4532 S.n4531 0.012
R8773 S.n3732 S.n3731 0.012
R8774 S.n2920 S.n2919 0.012
R8775 S.n2083 S.n2082 0.012
R8776 S.n1266 S.n1265 0.012
R8777 S.n8987 S.n8986 0.012
R8778 S.n8292 S.n8291 0.012
R8779 S.n7585 S.n7584 0.012
R8780 S.n6855 S.n6854 0.012
R8781 S.n6113 S.n6112 0.012
R8782 S.n5348 S.n5347 0.012
R8783 S.n4571 S.n4570 0.012
R8784 S.n3771 S.n3770 0.012
R8785 S.n2959 S.n2958 0.012
R8786 S.n2122 S.n2121 0.012
R8787 S.n1336 S.n1335 0.012
R8788 S.n9681 S.n9680 0.012
R8789 S.n9009 S.n9008 0.012
R8790 S.n8314 S.n8313 0.012
R8791 S.n7607 S.n7606 0.012
R8792 S.n6877 S.n6876 0.012
R8793 S.n6135 S.n6134 0.012
R8794 S.n5370 S.n5369 0.012
R8795 S.n4593 S.n4592 0.012
R8796 S.n3793 S.n3792 0.012
R8797 S.n2981 S.n2980 0.012
R8798 S.n2145 S.n2144 0.012
R8799 S.n1303 S.n1302 0.012
R8800 S.n507 S.n498 0.012
R8801 S.n6755 S.n6754 0.012
R8802 S.n6013 S.n6012 0.012
R8803 S.n5248 S.n5247 0.012
R8804 S.n4471 S.n4470 0.012
R8805 S.n3671 S.n3670 0.012
R8806 S.n2859 S.n2858 0.012
R8807 S.n2022 S.n2021 0.012
R8808 S.n1207 S.n1206 0.012
R8809 S.n7524 S.n7523 0.012
R8810 S.n6794 S.n6793 0.012
R8811 S.n6052 S.n6051 0.012
R8812 S.n5287 S.n5286 0.012
R8813 S.n4510 S.n4509 0.012
R8814 S.n3710 S.n3709 0.012
R8815 S.n2898 S.n2897 0.012
R8816 S.n2061 S.n2060 0.012
R8817 S.n1244 S.n1243 0.012
R8818 S.n466 S.n454 0.012
R8819 S.n5187 S.n5186 0.012
R8820 S.n4410 S.n4409 0.012
R8821 S.n3610 S.n3609 0.012
R8822 S.n2798 S.n2797 0.012
R8823 S.n1961 S.n1960 0.012
R8824 S.n1148 S.n1147 0.012
R8825 S.n5991 S.n5990 0.012
R8826 S.n5226 S.n5225 0.012
R8827 S.n4449 S.n4448 0.012
R8828 S.n3649 S.n3648 0.012
R8829 S.n2837 S.n2836 0.012
R8830 S.n2000 S.n1999 0.012
R8831 S.n1185 S.n1184 0.012
R8832 S.n419 S.n410 0.012
R8833 S.n3549 S.n3548 0.012
R8834 S.n2737 S.n2736 0.012
R8835 S.n1900 S.n1899 0.012
R8836 S.n1089 S.n1088 0.012
R8837 S.n4388 S.n4387 0.012
R8838 S.n3588 S.n3587 0.012
R8839 S.n2776 S.n2775 0.012
R8840 S.n1942 S.n1941 0.012
R8841 S.n1126 S.n1125 0.012
R8842 S.n375 S.n366 0.012
R8843 S.n1839 S.n1838 0.012
R8844 S.n1030 S.n1029 0.012
R8845 S.n2715 S.n2714 0.012
R8846 S.n1878 S.n1877 0.012
R8847 S.n1067 S.n1066 0.012
R8848 S.n331 S.n322 0.012
R8849 S.n1008 S.n1007 0.012
R8850 S.n287 S.n278 0.012
R8851 S.n2631 S.n2630 0.012
R8852 S.n2690 S.n2689 0.012
R8853 S.n3531 S.n3530 0.012
R8854 S.n3410 S.n3409 0.012
R8855 S.n4295 S.n4294 0.012
R8856 S.n4363 S.n4362 0.012
R8857 S.n5110 S.n5109 0.012
R8858 S.n5169 S.n5168 0.012
R8859 S.n5907 S.n5906 0.012
R8860 S.n5966 S.n5965 0.012
R8861 S.n6678 S.n6677 0.012
R8862 S.n6737 S.n6736 0.012
R8863 S.n7440 S.n7439 0.012
R8864 S.n7499 S.n7498 0.012
R8865 S.n8024 S.n8023 0.012
R8866 S.n8235 S.n8234 0.012
R8867 S.n8736 S.n8735 0.012
R8868 S.n8962 S.n8961 0.012
R8869 S.n9604 S.n9603 0.012
R8870 S.n9663 S.n9662 0.012
R8871 S.n10296 S.n10295 0.012
R8872 S.n10355 S.n10354 0.012
R8873 S.n10962 S.n10961 0.012
R8874 S.n11019 S.n11018 0.012
R8875 S.n12324 S.n12323 0.012
R8876 S.n11600 S.n11593 0.01
R8877 S.n722 S.n721 0.01
R8878 S.n689 S.n688 0.01
R8879 S.n656 S.n655 0.01
R8880 S.n623 S.n622 0.01
R8881 S.n590 S.n589 0.01
R8882 S.n557 S.n556 0.01
R8883 S.n10455 S.n10454 0.01
R8884 S.n837 S.n835 0.01
R8885 S.n1723 S.n1715 0.01
R8886 S.n2574 S.n2566 0.01
R8887 S.n3338 S.n3330 0.01
R8888 S.n4222 S.n4214 0.01
R8889 S.n5021 S.n5013 0.01
R8890 S.n5802 S.n5794 0.01
R8891 S.n6557 S.n6549 0.01
R8892 S.n7303 S.n7295 0.01
R8893 S.n7856 S.n7848 0.01
R8894 S.n8552 S.n8544 0.01
R8895 S.n9419 S.n9411 0.01
R8896 S.n10095 S.n10087 0.01
R8897 S.n10745 S.n10737 0.01
R8898 S.n751 S.n748 0.01
R8899 S.n11382 S.n11378 0.01
R8900 S.n10765 S.n10761 0.01
R8901 S.n10115 S.n10111 0.01
R8902 S.n9439 S.n9435 0.01
R8903 S.n8572 S.n8568 0.01
R8904 S.n7876 S.n7872 0.01
R8905 S.n7323 S.n7319 0.01
R8906 S.n6577 S.n6573 0.01
R8907 S.n5822 S.n5818 0.01
R8908 S.n5041 S.n5037 0.01
R8909 S.n4242 S.n4238 0.01
R8910 S.n3358 S.n3354 0.01
R8911 S.n2594 S.n2590 0.01
R8912 S.n1743 S.n1734 0.01
R8913 S.n899 S.n898 0.01
R8914 S.n770 S.n767 0.01
R8915 S.n475 S.n474 0.01
R8916 S.n431 S.n430 0.01
R8917 S.n387 S.n386 0.01
R8918 S.n343 S.n342 0.01
R8919 S.n299 S.n298 0.01
R8920 S.n255 S.n254 0.01
R8921 S.n805 S.n803 0.01
R8922 S.n1826 S.n1823 0.01
R8923 S.n1826 S.n993 0.01
R8924 S.n2696 S.n1831 0.01
R8925 S.n4369 S.n3541 0.01
R8926 S.n5175 S.n4373 0.01
R8927 S.n5972 S.n5179 0.01
R8928 S.n6743 S.n5976 0.01
R8929 S.n7505 S.n6747 0.01
R8930 S.n8241 S.n7509 0.01
R8931 S.n8968 S.n8245 0.01
R8932 S.n9669 S.n8972 0.01
R8933 S.n10361 S.n9673 0.01
R8934 S.n11025 S.n10365 0.01
R8935 S.n11644 S.n11029 0.01
R8936 S.n12611 S.n12609 0.01
R8937 S.n3537 S.n2700 0.01
R8938 S.n870 S.n853 0.01
R8939 S.n498 S.n497 0.01
R8940 S.n454 S.n453 0.01
R8941 S.n410 S.n409 0.01
R8942 S.n366 S.n365 0.01
R8943 S.n322 S.n321 0.01
R8944 S.n278 S.n277 0.01
R8945 S.n12604 S.n12602 0.01
R8946 S.n1701 S.n1699 0.01
R8947 S.n473 S.n472 0.01
R8948 S.n429 S.n428 0.01
R8949 S.n385 S.n384 0.01
R8950 S.n341 S.n340 0.01
R8951 S.n297 S.n296 0.01
R8952 S.n253 S.n252 0.01
R8953 S.n11363 S.n11361 0.01
R8954 S.n10056 S.n10041 0.01
R8955 S.n8477 S.n8462 0.01
R8956 S.n7192 S.n7177 0.01
R8957 S.n5655 S.n5640 0.01
R8958 S.n4039 S.n4024 0.01
R8959 S.n2355 S.n2340 0.01
R8960 S.n11923 S.n11921 0.009
R8961 S.n12607 S.n12606 0.009
R8962 S.n11102 S.n11101 0.009
R8963 S.n12611 S.n11997 0.009
R8964 S.n12006 S.n12005 0.008
R8965 S.n11058 S.n11057 0.008
R8966 S.n10428 S.n10427 0.008
R8967 S.n9768 S.n9767 0.008
R8968 S.n9096 S.n9095 0.008
R8969 S.n8401 S.n8400 0.008
R8970 S.n7694 S.n7693 0.008
R8971 S.n6964 S.n6963 0.008
R8972 S.n6222 S.n6221 0.008
R8973 S.n5457 S.n5456 0.008
R8974 S.n4680 S.n4679 0.008
R8975 S.n3880 S.n3879 0.008
R8976 S.n3068 S.n3067 0.008
R8977 S.n2233 S.n2232 0.008
R8978 S.n8254 S.n8253 0.008
R8979 S.n7547 S.n7546 0.008
R8980 S.n6817 S.n6816 0.008
R8981 S.n6075 S.n6074 0.008
R8982 S.n5310 S.n5309 0.008
R8983 S.n4533 S.n4532 0.008
R8984 S.n3733 S.n3732 0.008
R8985 S.n2921 S.n2920 0.008
R8986 S.n2084 S.n2083 0.008
R8987 S.n1267 S.n1266 0.008
R8988 S.n8988 S.n8987 0.008
R8989 S.n8293 S.n8292 0.008
R8990 S.n7586 S.n7585 0.008
R8991 S.n6856 S.n6855 0.008
R8992 S.n6114 S.n6113 0.008
R8993 S.n5349 S.n5348 0.008
R8994 S.n4572 S.n4571 0.008
R8995 S.n3772 S.n3771 0.008
R8996 S.n2960 S.n2959 0.008
R8997 S.n2123 S.n2122 0.008
R8998 S.n1304 S.n1303 0.008
R8999 S.n6756 S.n6755 0.008
R9000 S.n6014 S.n6013 0.008
R9001 S.n5249 S.n5248 0.008
R9002 S.n4472 S.n4471 0.008
R9003 S.n3672 S.n3671 0.008
R9004 S.n2860 S.n2859 0.008
R9005 S.n2023 S.n2022 0.008
R9006 S.n1208 S.n1207 0.008
R9007 S.n7525 S.n7524 0.008
R9008 S.n6795 S.n6794 0.008
R9009 S.n6053 S.n6052 0.008
R9010 S.n5288 S.n5287 0.008
R9011 S.n4511 S.n4510 0.008
R9012 S.n3711 S.n3710 0.008
R9013 S.n2899 S.n2898 0.008
R9014 S.n2062 S.n2061 0.008
R9015 S.n1245 S.n1244 0.008
R9016 S.n5188 S.n5187 0.008
R9017 S.n4411 S.n4410 0.008
R9018 S.n3611 S.n3610 0.008
R9019 S.n2799 S.n2798 0.008
R9020 S.n1962 S.n1961 0.008
R9021 S.n1149 S.n1148 0.008
R9022 S.n5992 S.n5991 0.008
R9023 S.n5227 S.n5226 0.008
R9024 S.n4450 S.n4449 0.008
R9025 S.n3650 S.n3649 0.008
R9026 S.n2838 S.n2837 0.008
R9027 S.n2001 S.n2000 0.008
R9028 S.n1186 S.n1185 0.008
R9029 S.n3550 S.n3549 0.008
R9030 S.n2738 S.n2737 0.008
R9031 S.n1901 S.n1900 0.008
R9032 S.n1090 S.n1089 0.008
R9033 S.n4389 S.n4388 0.008
R9034 S.n3589 S.n3588 0.008
R9035 S.n2777 S.n2776 0.008
R9036 S.n1943 S.n1942 0.008
R9037 S.n1127 S.n1126 0.008
R9038 S.n1840 S.n1839 0.008
R9039 S.n1031 S.n1030 0.008
R9040 S.n2716 S.n2715 0.008
R9041 S.n1879 S.n1878 0.008
R9042 S.n1068 S.n1067 0.008
R9043 S.n1009 S.n1008 0.008
R9044 S.n1430 S.n1429 0.008
R9045 S.n1761 S.n1760 0.008
R9046 S.n2249 S.n2248 0.008
R9047 S.n2612 S.n2611 0.008
R9048 S.n3084 S.n3083 0.008
R9049 S.n3376 S.n3375 0.008
R9050 S.n3896 S.n3895 0.008
R9051 S.n4260 S.n4259 0.008
R9052 S.n4696 S.n4695 0.008
R9053 S.n5059 S.n5058 0.008
R9054 S.n5473 S.n5472 0.008
R9055 S.n5840 S.n5839 0.008
R9056 S.n6238 S.n6237 0.008
R9057 S.n6595 S.n6594 0.008
R9058 S.n6980 S.n6979 0.008
R9059 S.n7341 S.n7340 0.008
R9060 S.n7710 S.n7709 0.008
R9061 S.n7894 S.n7893 0.008
R9062 S.n8417 S.n8416 0.008
R9063 S.n8590 S.n8589 0.008
R9064 S.n9112 S.n9111 0.008
R9065 S.n9457 S.n9456 0.008
R9066 S.n9784 S.n9783 0.008
R9067 S.n10133 S.n10132 0.008
R9068 S.n10444 S.n10443 0.008
R9069 S.n10783 S.n10782 0.008
R9070 S.n11074 S.n11073 0.008
R9071 S.n11400 S.n11399 0.008
R9072 S.n12022 S.n12021 0.008
R9073 S.n12302 S.n12301 0.008
R9074 S.n1424 S.n1423 0.008
R9075 S.n1320 S.n1317 0.008
R9076 S.n1688 S.n1687 0.008
R9077 S.n2162 S.n2161 0.008
R9078 S.n2552 S.n2551 0.008
R9079 S.n2998 S.n2997 0.008
R9080 S.n3316 S.n3315 0.008
R9081 S.n3810 S.n3809 0.008
R9082 S.n4200 S.n4199 0.008
R9083 S.n4610 S.n4609 0.008
R9084 S.n4999 S.n4998 0.008
R9085 S.n5387 S.n5386 0.008
R9086 S.n5780 S.n5779 0.008
R9087 S.n6152 S.n6151 0.008
R9088 S.n6535 S.n6534 0.008
R9089 S.n6894 S.n6893 0.008
R9090 S.n7281 S.n7280 0.008
R9091 S.n7624 S.n7623 0.008
R9092 S.n7834 S.n7833 0.008
R9093 S.n8331 S.n8330 0.008
R9094 S.n8530 S.n8529 0.008
R9095 S.n9026 S.n9025 0.008
R9096 S.n9397 S.n9396 0.008
R9097 S.n9698 S.n9697 0.008
R9098 S.n10073 S.n10072 0.008
R9099 S.n1723 S.n1712 0.008
R9100 S.n2574 S.n2563 0.008
R9101 S.n3338 S.n3327 0.008
R9102 S.n4222 S.n4211 0.008
R9103 S.n5021 S.n5010 0.008
R9104 S.n5802 S.n5791 0.008
R9105 S.n6557 S.n6546 0.008
R9106 S.n7303 S.n7292 0.008
R9107 S.n7856 S.n7845 0.008
R9108 S.n8552 S.n8541 0.008
R9109 S.n9419 S.n9408 0.008
R9110 S.n10095 S.n10084 0.008
R9111 S.n10745 S.n10734 0.008
R9112 S.n751 S.n750 0.008
R9113 S.n11382 S.n11381 0.008
R9114 S.n10765 S.n10764 0.008
R9115 S.n10115 S.n10114 0.008
R9116 S.n9439 S.n9438 0.008
R9117 S.n8572 S.n8571 0.008
R9118 S.n7876 S.n7875 0.008
R9119 S.n7323 S.n7322 0.008
R9120 S.n6577 S.n6576 0.008
R9121 S.n5822 S.n5821 0.008
R9122 S.n5041 S.n5040 0.008
R9123 S.n4242 S.n4241 0.008
R9124 S.n3358 S.n3357 0.008
R9125 S.n2594 S.n2593 0.008
R9126 S.n1743 S.n1732 0.008
R9127 S.n1386 S.n1385 0.008
R9128 S.n2205 S.n2204 0.008
R9129 S.n3041 S.n3040 0.008
R9130 S.n3853 S.n3852 0.008
R9131 S.n4653 S.n4652 0.008
R9132 S.n5430 S.n5429 0.008
R9133 S.n6195 S.n6194 0.008
R9134 S.n6937 S.n6936 0.008
R9135 S.n7667 S.n7666 0.008
R9136 S.n8374 S.n8373 0.008
R9137 S.n9069 S.n9068 0.008
R9138 S.n9741 S.n9740 0.008
R9139 S.n10401 S.n10400 0.008
R9140 S.n11031 S.n11030 0.008
R9141 S.n879 S.n878 0.008
R9142 S.n895 S.n891 0.008
R9143 S.n895 S.n894 0.008
R9144 S.n770 S.n769 0.008
R9145 S.n9815 S.n9811 0.008
R9146 S.n8974 S.n8973 0.008
R9147 S.n8279 S.n8278 0.008
R9148 S.n7572 S.n7571 0.008
R9149 S.n6842 S.n6841 0.008
R9150 S.n6100 S.n6099 0.008
R9151 S.n5335 S.n5334 0.008
R9152 S.n4558 S.n4557 0.008
R9153 S.n3758 S.n3757 0.008
R9154 S.n2946 S.n2945 0.008
R9155 S.n2109 S.n2108 0.008
R9156 S.n1291 S.n1290 0.008
R9157 S.n1281 S.n1278 0.008
R9158 S.n1660 S.n1659 0.008
R9159 S.n2100 S.n2099 0.008
R9160 S.n2516 S.n2515 0.008
R9161 S.n2937 S.n2936 0.008
R9162 S.n3280 S.n3279 0.008
R9163 S.n3749 S.n3748 0.008
R9164 S.n4164 S.n4163 0.008
R9165 S.n4549 S.n4548 0.008
R9166 S.n4963 S.n4962 0.008
R9167 S.n5326 S.n5325 0.008
R9168 S.n5744 S.n5743 0.008
R9169 S.n6091 S.n6090 0.008
R9170 S.n6499 S.n6498 0.008
R9171 S.n6833 S.n6832 0.008
R9172 S.n7245 S.n7244 0.008
R9173 S.n7563 S.n7562 0.008
R9174 S.n7798 S.n7797 0.008
R9175 S.n8270 S.n8269 0.008
R9176 S.n8494 S.n8493 0.008
R9177 S.n8448 S.n8446 0.008
R9178 S.n7511 S.n7510 0.008
R9179 S.n6781 S.n6780 0.008
R9180 S.n6039 S.n6038 0.008
R9181 S.n5274 S.n5273 0.008
R9182 S.n4497 S.n4496 0.008
R9183 S.n3697 S.n3696 0.008
R9184 S.n2885 S.n2884 0.008
R9185 S.n2048 S.n2047 0.008
R9186 S.n1232 S.n1231 0.008
R9187 S.n1222 S.n1219 0.008
R9188 S.n1624 S.n1623 0.008
R9189 S.n2039 S.n2038 0.008
R9190 S.n2480 S.n2479 0.008
R9191 S.n2876 S.n2875 0.008
R9192 S.n3244 S.n3243 0.008
R9193 S.n3688 S.n3687 0.008
R9194 S.n4128 S.n4127 0.008
R9195 S.n4488 S.n4487 0.008
R9196 S.n4927 S.n4926 0.008
R9197 S.n5265 S.n5264 0.008
R9198 S.n5708 S.n5707 0.008
R9199 S.n6030 S.n6029 0.008
R9200 S.n6463 S.n6462 0.008
R9201 S.n6772 S.n6771 0.008
R9202 S.n7209 S.n7208 0.008
R9203 S.n7011 S.n7009 0.008
R9204 S.n5978 S.n5977 0.008
R9205 S.n5213 S.n5212 0.008
R9206 S.n4436 S.n4435 0.008
R9207 S.n3636 S.n3635 0.008
R9208 S.n2824 S.n2823 0.008
R9209 S.n1987 S.n1986 0.008
R9210 S.n1173 S.n1172 0.008
R9211 S.n1163 S.n1160 0.008
R9212 S.n1588 S.n1587 0.008
R9213 S.n1978 S.n1977 0.008
R9214 S.n2444 S.n2443 0.008
R9215 S.n2815 S.n2814 0.008
R9216 S.n3208 S.n3207 0.008
R9217 S.n3627 S.n3626 0.008
R9218 S.n4092 S.n4091 0.008
R9219 S.n4427 S.n4426 0.008
R9220 S.n4891 S.n4890 0.008
R9221 S.n5204 S.n5203 0.008
R9222 S.n5672 S.n5671 0.008
R9223 S.n5504 S.n5500 0.008
R9224 S.n4375 S.n4374 0.008
R9225 S.n3575 S.n3574 0.008
R9226 S.n2763 S.n2762 0.008
R9227 S.n1926 S.n1925 0.008
R9228 S.n1114 S.n1113 0.008
R9229 S.n1104 S.n1101 0.008
R9230 S.n1552 S.n1551 0.008
R9231 S.n1917 S.n1916 0.008
R9232 S.n2408 S.n2407 0.008
R9233 S.n2754 S.n2753 0.008
R9234 S.n3172 S.n3171 0.008
R9235 S.n3566 S.n3565 0.008
R9236 S.n4056 S.n4055 0.008
R9237 S.n3927 S.n3925 0.008
R9238 S.n2702 S.n2701 0.008
R9239 S.n1865 S.n1864 0.008
R9240 S.n1055 S.n1054 0.008
R9241 S.n1045 S.n1042 0.008
R9242 S.n1516 S.n1515 0.008
R9243 S.n1856 S.n1855 0.008
R9244 S.n2372 S.n2371 0.008
R9245 S.n2280 S.n2276 0.008
R9246 S.n996 S.n995 0.008
R9247 S.n949 S.n946 0.008
R9248 S.n805 S.n804 0.008
R9249 S.n980 S.n247 0.008
R9250 S.n11600 S.n11599 0.008
R9251 S.n11899 S.n11898 0.008
R9252 S.n869 S.n868 0.008
R9253 S.n869 S.n867 0.007
R9254 S.t7 S.n165 0.007
R9255 S.t7 S.n158 0.007
R9256 S.t7 S.n146 0.007
R9257 S.t7 S.n134 0.007
R9258 S.t7 S.n121 0.007
R9259 S.t7 S.n108 0.007
R9260 S.t7 S.n95 0.007
R9261 S.n852 S.n851 0.007
R9262 S.n11592 S.n11591 0.007
R9263 S.n1425 S.n1424 0.006
R9264 S.n1320 S.n1319 0.006
R9265 S.n1281 S.n1280 0.006
R9266 S.n1222 S.n1221 0.006
R9267 S.n1163 S.n1162 0.006
R9268 S.n1104 S.n1103 0.006
R9269 S.n1045 S.n1044 0.006
R9270 S.n949 S.n948 0.006
R9271 S.n11900 S.n11899 0.006
R9272 S.n484 S.n475 0.006
R9273 S.n440 S.n431 0.006
R9274 S.n396 S.n387 0.006
R9275 S.n352 S.n343 0.006
R9276 S.n308 S.n299 0.006
R9277 S.n264 S.n255 0.006
R9278 S.n837 S.n824 0.005
R9279 S.n1337 S.n1336 0.005
R9280 S.n9682 S.n9681 0.005
R9281 S.n9010 S.n9009 0.005
R9282 S.n8315 S.n8314 0.005
R9283 S.n7608 S.n7607 0.005
R9284 S.n6878 S.n6877 0.005
R9285 S.n6136 S.n6135 0.005
R9286 S.n5371 S.n5370 0.005
R9287 S.n4594 S.n4593 0.005
R9288 S.n3794 S.n3793 0.005
R9289 S.n2982 S.n2981 0.005
R9290 S.n2146 S.n2145 0.005
R9291 S.t7 S.n170 0.005
R9292 S.n9810 S.n9809 0.005
R9293 S.n8443 S.n8442 0.005
R9294 S.n7006 S.n7005 0.005
R9295 S.n5499 S.n5498 0.005
R9296 S.n3922 S.n3921 0.005
R9297 S.n2275 S.n2274 0.005
R9298 S.t7 S.n184 0.005
R9299 S.n11909 S.n11908 0.004
R9300 S.n12318 S.n12317 0.004
R9301 S.n12595 S.n12594 0.004
R9302 S.n941 S.n940 0.004
R9303 S.n918 S.n917 0.004
R9304 S.n1417 S.n1416 0.004
R9305 S.n11883 S.n11882 0.004
R9306 S.n12295 S.n12294 0.004
R9307 S.n12011 S.n12010 0.004
R9308 S.n11393 S.n11392 0.004
R9309 S.n11063 S.n11062 0.004
R9310 S.n10776 S.n10775 0.004
R9311 S.n10433 S.n10432 0.004
R9312 S.n10126 S.n10125 0.004
R9313 S.n9773 S.n9772 0.004
R9314 S.n9450 S.n9449 0.004
R9315 S.n9101 S.n9100 0.004
R9316 S.n8583 S.n8582 0.004
R9317 S.n8406 S.n8405 0.004
R9318 S.n7887 S.n7886 0.004
R9319 S.n7699 S.n7698 0.004
R9320 S.n7334 S.n7333 0.004
R9321 S.n6969 S.n6968 0.004
R9322 S.n6588 S.n6587 0.004
R9323 S.n6227 S.n6226 0.004
R9324 S.n5833 S.n5832 0.004
R9325 S.n5462 S.n5461 0.004
R9326 S.n5052 S.n5051 0.004
R9327 S.n4685 S.n4684 0.004
R9328 S.n4253 S.n4252 0.004
R9329 S.n3885 S.n3884 0.004
R9330 S.n3369 S.n3368 0.004
R9331 S.n3073 S.n3072 0.004
R9332 S.n2605 S.n2604 0.004
R9333 S.n2238 S.n2237 0.004
R9334 S.n1754 S.n1753 0.004
R9335 S.n785 S.n784 0.004
R9336 S.n482 S.n481 0.004
R9337 S.n1272 S.n1271 0.004
R9338 S.n9125 S.n9124 0.004
R9339 S.n8487 S.n8486 0.004
R9340 S.n8259 S.n8258 0.004
R9341 S.n7791 S.n7790 0.004
R9342 S.n7552 S.n7551 0.004
R9343 S.n7238 S.n7237 0.004
R9344 S.n6822 S.n6821 0.004
R9345 S.n6492 S.n6491 0.004
R9346 S.n6080 S.n6079 0.004
R9347 S.n5737 S.n5736 0.004
R9348 S.n5315 S.n5314 0.004
R9349 S.n4956 S.n4955 0.004
R9350 S.n4538 S.n4537 0.004
R9351 S.n4157 S.n4156 0.004
R9352 S.n3738 S.n3737 0.004
R9353 S.n3273 S.n3272 0.004
R9354 S.n2926 S.n2925 0.004
R9355 S.n2509 S.n2508 0.004
R9356 S.n2089 S.n2088 0.004
R9357 S.n1653 S.n1652 0.004
R9358 S.n505 S.n504 0.004
R9359 S.n9807 S.n9806 0.004
R9360 S.n9377 S.n9376 0.004
R9361 S.n8984 S.n8983 0.004
R9362 S.n8510 S.n8509 0.004
R9363 S.n8289 S.n8288 0.004
R9364 S.n7814 S.n7813 0.004
R9365 S.n7582 S.n7581 0.004
R9366 S.n7261 S.n7260 0.004
R9367 S.n6852 S.n6851 0.004
R9368 S.n6515 S.n6514 0.004
R9369 S.n6110 S.n6109 0.004
R9370 S.n5760 S.n5759 0.004
R9371 S.n5345 S.n5344 0.004
R9372 S.n4979 S.n4978 0.004
R9373 S.n4568 S.n4567 0.004
R9374 S.n4180 S.n4179 0.004
R9375 S.n3768 S.n3767 0.004
R9376 S.n3296 S.n3295 0.004
R9377 S.n2956 S.n2955 0.004
R9378 S.n2532 S.n2531 0.004
R9379 S.n2119 S.n2118 0.004
R9380 S.n1676 S.n1675 0.004
R9381 S.n1697 S.n1696 0.004
R9382 S.n1329 S.n1328 0.004
R9383 S.n820 S.n819 0.004
R9384 S.n831 S.n830 0.004
R9385 S.n2151 S.n2150 0.004
R9386 S.n2987 S.n2986 0.004
R9387 S.n3799 S.n3798 0.004
R9388 S.n4599 S.n4598 0.004
R9389 S.n5376 S.n5375 0.004
R9390 S.n6141 S.n6140 0.004
R9391 S.n6883 S.n6882 0.004
R9392 S.n7613 S.n7612 0.004
R9393 S.n8320 S.n8319 0.004
R9394 S.n9015 S.n9014 0.004
R9395 S.n9687 S.n9686 0.004
R9396 S.n10460 S.n10459 0.004
R9397 S.n10066 S.n10065 0.004
R9398 S.n9390 S.n9389 0.004
R9399 S.n8523 S.n8522 0.004
R9400 S.n7827 S.n7826 0.004
R9401 S.n7274 S.n7273 0.004
R9402 S.n6528 S.n6527 0.004
R9403 S.n5773 S.n5772 0.004
R9404 S.n4992 S.n4991 0.004
R9405 S.n4193 S.n4192 0.004
R9406 S.n3309 S.n3308 0.004
R9407 S.n2545 S.n2544 0.004
R9408 S.n1368 S.n1367 0.004
R9409 S.n745 S.n744 0.004
R9410 S.n863 S.n862 0.004
R9411 S.n11094 S.n11093 0.004
R9412 S.n10740 S.n10739 0.004
R9413 S.n10378 S.n10377 0.004
R9414 S.n10090 S.n10089 0.004
R9415 S.n9718 S.n9717 0.004
R9416 S.n9414 S.n9413 0.004
R9417 S.n9046 S.n9045 0.004
R9418 S.n8547 S.n8546 0.004
R9419 S.n8351 S.n8350 0.004
R9420 S.n7851 S.n7850 0.004
R9421 S.n7644 S.n7643 0.004
R9422 S.n7298 S.n7297 0.004
R9423 S.n6914 S.n6913 0.004
R9424 S.n6552 S.n6551 0.004
R9425 S.n6172 S.n6171 0.004
R9426 S.n5797 S.n5796 0.004
R9427 S.n5407 S.n5406 0.004
R9428 S.n5016 S.n5015 0.004
R9429 S.n4630 S.n4629 0.004
R9430 S.n4217 S.n4216 0.004
R9431 S.n3830 S.n3829 0.004
R9432 S.n3333 S.n3332 0.004
R9433 S.n3018 S.n3017 0.004
R9434 S.n2569 S.n2568 0.004
R9435 S.n2182 S.n2181 0.004
R9436 S.n1718 S.n1717 0.004
R9437 S.n1396 S.n1395 0.004
R9438 S.n765 S.n764 0.004
R9439 S.n1737 S.n1736 0.004
R9440 S.n2215 S.n2214 0.004
R9441 S.n2589 S.n2588 0.004
R9442 S.n3051 S.n3050 0.004
R9443 S.n3353 S.n3352 0.004
R9444 S.n3863 S.n3862 0.004
R9445 S.n4237 S.n4236 0.004
R9446 S.n4663 S.n4662 0.004
R9447 S.n5036 S.n5035 0.004
R9448 S.n5440 S.n5439 0.004
R9449 S.n5817 S.n5816 0.004
R9450 S.n6205 S.n6204 0.004
R9451 S.n6572 S.n6571 0.004
R9452 S.n6947 S.n6946 0.004
R9453 S.n7318 S.n7317 0.004
R9454 S.n7677 S.n7676 0.004
R9455 S.n7871 S.n7870 0.004
R9456 S.n8384 S.n8383 0.004
R9457 S.n8567 S.n8566 0.004
R9458 S.n9079 S.n9078 0.004
R9459 S.n9434 S.n9433 0.004
R9460 S.n9751 S.n9750 0.004
R9461 S.n10110 S.n10109 0.004
R9462 S.n10411 S.n10410 0.004
R9463 S.n10760 S.n10759 0.004
R9464 S.n11041 S.n11040 0.004
R9465 S.n11377 S.n11376 0.004
R9466 S.n12045 S.n12044 0.004
R9467 S.n889 S.n888 0.004
R9468 S.n1300 S.n1299 0.004
R9469 S.n729 S.n728 0.004
R9470 S.n712 S.n711 0.004
R9471 S.n438 S.n437 0.004
R9472 S.n1213 S.n1212 0.004
R9473 S.n7723 S.n7722 0.004
R9474 S.n7202 S.n7201 0.004
R9475 S.n6761 S.n6760 0.004
R9476 S.n6456 S.n6455 0.004
R9477 S.n6019 S.n6018 0.004
R9478 S.n5701 S.n5700 0.004
R9479 S.n5254 S.n5253 0.004
R9480 S.n4920 S.n4919 0.004
R9481 S.n4477 S.n4476 0.004
R9482 S.n4121 S.n4120 0.004
R9483 S.n3677 S.n3676 0.004
R9484 S.n3237 S.n3236 0.004
R9485 S.n2865 S.n2864 0.004
R9486 S.n2473 S.n2472 0.004
R9487 S.n2028 S.n2027 0.004
R9488 S.n1617 S.n1616 0.004
R9489 S.n464 S.n463 0.004
R9490 S.n8440 S.n8439 0.004
R9491 S.n7778 S.n7777 0.004
R9492 S.n7521 S.n7520 0.004
R9493 S.n7225 S.n7224 0.004
R9494 S.n6791 S.n6790 0.004
R9495 S.n6479 S.n6478 0.004
R9496 S.n6049 S.n6048 0.004
R9497 S.n5724 S.n5723 0.004
R9498 S.n5284 S.n5283 0.004
R9499 S.n4943 S.n4942 0.004
R9500 S.n4507 S.n4506 0.004
R9501 S.n4144 S.n4143 0.004
R9502 S.n3707 S.n3706 0.004
R9503 S.n3260 S.n3259 0.004
R9504 S.n2895 S.n2894 0.004
R9505 S.n2496 S.n2495 0.004
R9506 S.n2058 S.n2057 0.004
R9507 S.n1640 S.n1639 0.004
R9508 S.n1241 S.n1240 0.004
R9509 S.n696 S.n695 0.004
R9510 S.n679 S.n678 0.004
R9511 S.n394 S.n393 0.004
R9512 S.n1154 S.n1153 0.004
R9513 S.n6251 S.n6250 0.004
R9514 S.n5665 S.n5664 0.004
R9515 S.n5193 S.n5192 0.004
R9516 S.n4884 S.n4883 0.004
R9517 S.n4416 S.n4415 0.004
R9518 S.n4085 S.n4084 0.004
R9519 S.n3616 S.n3615 0.004
R9520 S.n3201 S.n3200 0.004
R9521 S.n2804 S.n2803 0.004
R9522 S.n2437 S.n2436 0.004
R9523 S.n1967 S.n1966 0.004
R9524 S.n1581 S.n1580 0.004
R9525 S.n417 S.n416 0.004
R9526 S.n7003 S.n7002 0.004
R9527 S.n6443 S.n6442 0.004
R9528 S.n5988 S.n5987 0.004
R9529 S.n5688 S.n5687 0.004
R9530 S.n5223 S.n5222 0.004
R9531 S.n4907 S.n4906 0.004
R9532 S.n4446 S.n4445 0.004
R9533 S.n4108 S.n4107 0.004
R9534 S.n3646 S.n3645 0.004
R9535 S.n3224 S.n3223 0.004
R9536 S.n2834 S.n2833 0.004
R9537 S.n2460 S.n2459 0.004
R9538 S.n1997 S.n1996 0.004
R9539 S.n1604 S.n1603 0.004
R9540 S.n1182 S.n1181 0.004
R9541 S.n663 S.n662 0.004
R9542 S.n646 S.n645 0.004
R9543 S.n350 S.n349 0.004
R9544 S.n1095 S.n1094 0.004
R9545 S.n4709 S.n4708 0.004
R9546 S.n4049 S.n4048 0.004
R9547 S.n3555 S.n3554 0.004
R9548 S.n3165 S.n3164 0.004
R9549 S.n2743 S.n2742 0.004
R9550 S.n2401 S.n2400 0.004
R9551 S.n1906 S.n1905 0.004
R9552 S.n1545 S.n1544 0.004
R9553 S.n373 S.n372 0.004
R9554 S.n5496 S.n5495 0.004
R9555 S.n4871 S.n4870 0.004
R9556 S.n4385 S.n4384 0.004
R9557 S.n4072 S.n4071 0.004
R9558 S.n3585 S.n3584 0.004
R9559 S.n3188 S.n3187 0.004
R9560 S.n2773 S.n2772 0.004
R9561 S.n2424 S.n2423 0.004
R9562 S.n1939 S.n1938 0.004
R9563 S.n1568 S.n1567 0.004
R9564 S.n1123 S.n1122 0.004
R9565 S.n630 S.n629 0.004
R9566 S.n613 S.n612 0.004
R9567 S.n306 S.n305 0.004
R9568 S.n1036 S.n1035 0.004
R9569 S.n3097 S.n3096 0.004
R9570 S.n2365 S.n2364 0.004
R9571 S.n1845 S.n1844 0.004
R9572 S.n1509 S.n1508 0.004
R9573 S.n329 S.n328 0.004
R9574 S.n3919 S.n3918 0.004
R9575 S.n3152 S.n3151 0.004
R9576 S.n2712 S.n2711 0.004
R9577 S.n2388 S.n2387 0.004
R9578 S.n1875 S.n1874 0.004
R9579 S.n1532 S.n1531 0.004
R9580 S.n1064 S.n1063 0.004
R9581 S.n597 S.n596 0.004
R9582 S.n580 S.n579 0.004
R9583 S.n262 S.n261 0.004
R9584 S.n1443 S.n1442 0.004
R9585 S.n285 S.n284 0.004
R9586 S.n2272 S.n2271 0.004
R9587 S.n1496 S.n1495 0.004
R9588 S.n1005 S.n1004 0.004
R9589 S.n564 S.n563 0.004
R9590 S.n547 S.n546 0.004
R9591 S.n963 S.n962 0.004
R9592 S.n802 S.n801 0.004
R9593 S.n1805 S.n1804 0.004
R9594 S.n1794 S.n1793 0.004
R9595 S.n2312 S.n2311 0.004
R9596 S.n2300 S.n2299 0.004
R9597 S.n3440 S.n3439 0.004
R9598 S.n3428 S.n3427 0.004
R9599 S.n3959 S.n3958 0.004
R9600 S.n3947 S.n3946 0.004
R9601 S.n4754 S.n4753 0.004
R9602 S.n4742 S.n4741 0.004
R9603 S.n5536 S.n5535 0.004
R9604 S.n5524 S.n5523 0.004
R9605 S.n6296 S.n6295 0.004
R9606 S.n6284 S.n6283 0.004
R9607 S.n7043 S.n7042 0.004
R9608 S.n7031 S.n7030 0.004
R9609 S.n8054 S.n8053 0.004
R9610 S.n8042 S.n8041 0.004
R9611 S.n8766 S.n8765 0.004
R9612 S.n8754 S.n8753 0.004
R9613 S.n9170 S.n9169 0.004
R9614 S.n9158 S.n9157 0.004
R9615 S.n9847 S.n9846 0.004
R9616 S.n9835 S.n9834 0.004
R9617 S.n10505 S.n10504 0.004
R9618 S.n10493 S.n10492 0.004
R9619 S.n11133 S.n11132 0.004
R9620 S.n11121 S.n11120 0.004
R9621 S.n12061 S.n12060 0.004
R9622 S.n12340 S.n12339 0.004
R9623 S.n11865 S.n11864 0.004
R9624 S.n1821 S.n1820 0.004
R9625 S.n1777 S.n1776 0.004
R9626 S.n2329 S.n2328 0.004
R9627 S.n11848 S.n11847 0.004
R9628 S.n12355 S.n12354 0.004
R9629 S.n12078 S.n12077 0.004
R9630 S.n11158 S.n11157 0.004
R9631 S.n11150 S.n11149 0.004
R9632 S.n10530 S.n10529 0.004
R9633 S.n10522 S.n10521 0.004
R9634 S.n9872 S.n9871 0.004
R9635 S.n9864 S.n9863 0.004
R9636 S.n9195 S.n9194 0.004
R9637 S.n9187 S.n9186 0.004
R9638 S.n8791 S.n8790 0.004
R9639 S.n8783 S.n8782 0.004
R9640 S.n8079 S.n8078 0.004
R9641 S.n8071 S.n8070 0.004
R9642 S.n7068 S.n7067 0.004
R9643 S.n7060 S.n7059 0.004
R9644 S.n6321 S.n6320 0.004
R9645 S.n6313 S.n6312 0.004
R9646 S.n5561 S.n5560 0.004
R9647 S.n5553 S.n5552 0.004
R9648 S.n4779 S.n4778 0.004
R9649 S.n4771 S.n4770 0.004
R9650 S.n3984 S.n3983 0.004
R9651 S.n3976 S.n3975 0.004
R9652 S.n3465 S.n3464 0.004
R9653 S.n3457 S.n3456 0.004
R9654 S.n2337 S.n2336 0.004
R9655 S.n2664 S.n2663 0.004
R9656 S.n2628 S.n2627 0.004
R9657 S.n3488 S.n3487 0.004
R9658 S.n11833 S.n11832 0.004
R9659 S.n12370 S.n12369 0.004
R9660 S.n12094 S.n12093 0.004
R9661 S.n11412 S.n11411 0.004
R9662 S.n11181 S.n11180 0.004
R9663 S.n10796 S.n10795 0.004
R9664 S.n10553 S.n10552 0.004
R9665 S.n10146 S.n10145 0.004
R9666 S.n9895 S.n9894 0.004
R9667 S.n9470 S.n9469 0.004
R9668 S.n9218 S.n9217 0.004
R9669 S.n8603 S.n8602 0.004
R9670 S.n8814 S.n8813 0.004
R9671 S.n7907 S.n7906 0.004
R9672 S.n8102 S.n8101 0.004
R9673 S.n7354 S.n7353 0.004
R9674 S.n7091 S.n7090 0.004
R9675 S.n6608 S.n6607 0.004
R9676 S.n6344 S.n6343 0.004
R9677 S.n5853 S.n5852 0.004
R9678 S.n5584 S.n5583 0.004
R9679 S.n5072 S.n5071 0.004
R9680 S.n4802 S.n4801 0.004
R9681 S.n4273 S.n4272 0.004
R9682 S.n4007 S.n4006 0.004
R9683 S.n3389 S.n3388 0.004
R9684 S.n11820 S.n11819 0.004
R9685 S.n12389 S.n12388 0.004
R9686 S.n12111 S.n12110 0.004
R9687 S.n11431 S.n11430 0.004
R9688 S.n11198 S.n11197 0.004
R9689 S.n10815 S.n10814 0.004
R9690 S.n10570 S.n10569 0.004
R9691 S.n10165 S.n10164 0.004
R9692 S.n9912 S.n9911 0.004
R9693 S.n9489 S.n9488 0.004
R9694 S.n9235 S.n9234 0.004
R9695 S.n8622 S.n8621 0.004
R9696 S.n8831 S.n8830 0.004
R9697 S.n7926 S.n7925 0.004
R9698 S.n8119 S.n8118 0.004
R9699 S.n7373 S.n7372 0.004
R9700 S.n7108 S.n7107 0.004
R9701 S.n6627 S.n6626 0.004
R9702 S.n6361 S.n6360 0.004
R9703 S.n5872 S.n5871 0.004
R9704 S.n5601 S.n5600 0.004
R9705 S.n5091 S.n5090 0.004
R9706 S.n4819 S.n4818 0.004
R9707 S.n4313 S.n4312 0.004
R9708 S.n4322 S.n4321 0.004
R9709 S.n3407 S.n3406 0.004
R9710 S.n3505 S.n3504 0.004
R9711 S.n4337 S.n4336 0.004
R9712 S.n4292 S.n4291 0.004
R9713 S.n4832 S.n4831 0.004
R9714 S.n11803 S.n11802 0.004
R9715 S.n12402 S.n12401 0.004
R9716 S.n12124 S.n12123 0.004
R9717 S.n11444 S.n11443 0.004
R9718 S.n11211 S.n11210 0.004
R9719 S.n10828 S.n10827 0.004
R9720 S.n10583 S.n10582 0.004
R9721 S.n10178 S.n10177 0.004
R9722 S.n9925 S.n9924 0.004
R9723 S.n9502 S.n9501 0.004
R9724 S.n9248 S.n9247 0.004
R9725 S.n8635 S.n8634 0.004
R9726 S.n8844 S.n8843 0.004
R9727 S.n7939 S.n7938 0.004
R9728 S.n8132 S.n8131 0.004
R9729 S.n7386 S.n7385 0.004
R9730 S.n7121 S.n7120 0.004
R9731 S.n6640 S.n6639 0.004
R9732 S.n6374 S.n6373 0.004
R9733 S.n5885 S.n5884 0.004
R9734 S.n5614 S.n5613 0.004
R9735 S.n4840 S.n4839 0.004
R9736 S.n5143 S.n5142 0.004
R9737 S.n5107 S.n5106 0.004
R9738 S.n5629 S.n5628 0.004
R9739 S.n11788 S.n11787 0.004
R9740 S.n12418 S.n12417 0.004
R9741 S.n12139 S.n12138 0.004
R9742 S.n11460 S.n11459 0.004
R9743 S.n11226 S.n11225 0.004
R9744 S.n10844 S.n10843 0.004
R9745 S.n10598 S.n10597 0.004
R9746 S.n10194 S.n10193 0.004
R9747 S.n9940 S.n9939 0.004
R9748 S.n9518 S.n9517 0.004
R9749 S.n9263 S.n9262 0.004
R9750 S.n8651 S.n8650 0.004
R9751 S.n8859 S.n8858 0.004
R9752 S.n7955 S.n7954 0.004
R9753 S.n8147 S.n8146 0.004
R9754 S.n7402 S.n7401 0.004
R9755 S.n7136 S.n7135 0.004
R9756 S.n6656 S.n6655 0.004
R9757 S.n6389 S.n6388 0.004
R9758 S.n5637 S.n5636 0.004
R9759 S.n5940 S.n5939 0.004
R9760 S.n5904 S.n5903 0.004
R9761 S.n6404 S.n6403 0.004
R9762 S.n11773 S.n11772 0.004
R9763 S.n12434 S.n12433 0.004
R9764 S.n12154 S.n12153 0.004
R9765 S.n11476 S.n11475 0.004
R9766 S.n11241 S.n11240 0.004
R9767 S.n10860 S.n10859 0.004
R9768 S.n10613 S.n10612 0.004
R9769 S.n10210 S.n10209 0.004
R9770 S.n9955 S.n9954 0.004
R9771 S.n9534 S.n9533 0.004
R9772 S.n9278 S.n9277 0.004
R9773 S.n8667 S.n8666 0.004
R9774 S.n8874 S.n8873 0.004
R9775 S.n7971 S.n7970 0.004
R9776 S.n8162 S.n8161 0.004
R9777 S.n7418 S.n7417 0.004
R9778 S.n7151 S.n7150 0.004
R9779 S.n6412 S.n6411 0.004
R9780 S.n6711 S.n6710 0.004
R9781 S.n6675 S.n6674 0.004
R9782 S.n7166 S.n7165 0.004
R9783 S.n11758 S.n11757 0.004
R9784 S.n12450 S.n12449 0.004
R9785 S.n12169 S.n12168 0.004
R9786 S.n11492 S.n11491 0.004
R9787 S.n11256 S.n11255 0.004
R9788 S.n10876 S.n10875 0.004
R9789 S.n10628 S.n10627 0.004
R9790 S.n10226 S.n10225 0.004
R9791 S.n9970 S.n9969 0.004
R9792 S.n9550 S.n9549 0.004
R9793 S.n9293 S.n9292 0.004
R9794 S.n8683 S.n8682 0.004
R9795 S.n8889 S.n8888 0.004
R9796 S.n7987 S.n7986 0.004
R9797 S.n8177 S.n8176 0.004
R9798 S.n7174 S.n7173 0.004
R9799 S.n7473 S.n7472 0.004
R9800 S.n7437 S.n7436 0.004
R9801 S.n8192 S.n8191 0.004
R9802 S.n11743 S.n11742 0.004
R9803 S.n12466 S.n12465 0.004
R9804 S.n12184 S.n12183 0.004
R9805 S.n11508 S.n11507 0.004
R9806 S.n11271 S.n11270 0.004
R9807 S.n10892 S.n10891 0.004
R9808 S.n10643 S.n10642 0.004
R9809 S.n10242 S.n10241 0.004
R9810 S.n9985 S.n9984 0.004
R9811 S.n9566 S.n9565 0.004
R9812 S.n9308 S.n9307 0.004
R9813 S.n8699 S.n8698 0.004
R9814 S.n8904 S.n8903 0.004
R9815 S.n8003 S.n8002 0.004
R9816 S.n8209 S.n8208 0.004
R9817 S.n8021 S.n8020 0.004
R9818 S.n8919 S.n8918 0.004
R9819 S.n11728 S.n11727 0.004
R9820 S.n12482 S.n12481 0.004
R9821 S.n12199 S.n12198 0.004
R9822 S.n11524 S.n11523 0.004
R9823 S.n11286 S.n11285 0.004
R9824 S.n10908 S.n10907 0.004
R9825 S.n10658 S.n10657 0.004
R9826 S.n10258 S.n10257 0.004
R9827 S.n10000 S.n9999 0.004
R9828 S.n9582 S.n9581 0.004
R9829 S.n9323 S.n9322 0.004
R9830 S.n8715 S.n8714 0.004
R9831 S.n8936 S.n8935 0.004
R9832 S.n8733 S.n8732 0.004
R9833 S.n9338 S.n9337 0.004
R9834 S.n11713 S.n11712 0.004
R9835 S.n12498 S.n12497 0.004
R9836 S.n12214 S.n12213 0.004
R9837 S.n11540 S.n11539 0.004
R9838 S.n11301 S.n11300 0.004
R9839 S.n10924 S.n10923 0.004
R9840 S.n10673 S.n10672 0.004
R9841 S.n10274 S.n10273 0.004
R9842 S.n10015 S.n10014 0.004
R9843 S.n9346 S.n9345 0.004
R9844 S.n9637 S.n9636 0.004
R9845 S.n9601 S.n9600 0.004
R9846 S.n10030 S.n10029 0.004
R9847 S.n11698 S.n11697 0.004
R9848 S.n12514 S.n12513 0.004
R9849 S.n12229 S.n12228 0.004
R9850 S.n11556 S.n11555 0.004
R9851 S.n11316 S.n11315 0.004
R9852 S.n10940 S.n10939 0.004
R9853 S.n10688 S.n10687 0.004
R9854 S.n10038 S.n10037 0.004
R9855 S.n10329 S.n10328 0.004
R9856 S.n10293 S.n10292 0.004
R9857 S.n10703 S.n10702 0.004
R9858 S.n11683 S.n11682 0.004
R9859 S.n12530 S.n12529 0.004
R9860 S.n12244 S.n12243 0.004
R9861 S.n11572 S.n11571 0.004
R9862 S.n11331 S.n11330 0.004
R9863 S.n10711 S.n10710 0.004
R9864 S.n10995 S.n10994 0.004
R9865 S.n10959 S.n10958 0.004
R9866 S.n11346 S.n11345 0.004
R9867 S.n11668 S.n11667 0.004
R9868 S.n12546 S.n12545 0.004
R9869 S.n12259 S.n12258 0.004
R9870 S.n11354 S.n11353 0.004
R9871 S.n11630 S.n11629 0.004
R9872 S.n11589 S.n11588 0.004
R9873 S.n12579 S.n12578 0.004
R9874 S.n11655 S.n11654 0.004
R9875 S.n12566 S.n12565 0.004
R9876 S.t7 S.n177 0.004
R9877 S.n920 S.n919 0.004
R9878 S.n507 S.n506 0.004
R9879 S.n484 S.n483 0.004
R9880 S.n466 S.n465 0.004
R9881 S.n440 S.n439 0.004
R9882 S.n419 S.n418 0.004
R9883 S.n396 S.n395 0.004
R9884 S.n375 S.n374 0.004
R9885 S.n352 S.n351 0.004
R9886 S.n331 S.n330 0.004
R9887 S.n308 S.n307 0.004
R9888 S.n287 S.n286 0.004
R9889 S.n264 S.n263 0.004
R9890 S.t7 S.n190 0.004
R9891 S.n534 S.n519 0.004
R9892 S.n10725 S.n10724 0.004
R9893 S.n10384 S.n10383 0.004
R9894 S.n9724 S.n9723 0.004
R9895 S.n9052 S.n9051 0.004
R9896 S.n8357 S.n8356 0.004
R9897 S.n7650 S.n7649 0.004
R9898 S.n6920 S.n6919 0.004
R9899 S.n6178 S.n6177 0.004
R9900 S.n5413 S.n5412 0.004
R9901 S.n4636 S.n4635 0.004
R9902 S.n3836 S.n3835 0.004
R9903 S.n3024 S.n3023 0.004
R9904 S.n2188 S.n2187 0.004
R9905 S.n1353 S.n1352 0.004
R9906 S.n845 S.n844 0.004
R9907 S.n10725 S.n10723 0.004
R9908 S.n770 S.n758 0.004
R9909 S.n1743 S.n1742 0.004
R9910 S.n2594 S.n2582 0.004
R9911 S.n3358 S.n3346 0.004
R9912 S.n4242 S.n4230 0.004
R9913 S.n5041 S.n5029 0.004
R9914 S.n5822 S.n5810 0.004
R9915 S.n6577 S.n6565 0.004
R9916 S.n7323 S.n7311 0.004
R9917 S.n7876 S.n7864 0.004
R9918 S.n8572 S.n8560 0.004
R9919 S.n9439 S.n9427 0.004
R9920 S.n10115 S.n10103 0.004
R9921 S.n10765 S.n10753 0.004
R9922 S.n11382 S.n11370 0.004
R9923 S.n12285 S.n12283 0.004
R9924 S.n10056 S.n10055 0.004
R9925 S.n731 S.n722 0.004
R9926 S.n9363 S.n9361 0.004
R9927 S.n8477 S.n8476 0.004
R9928 S.n698 S.n689 0.004
R9929 S.n7764 S.n7762 0.004
R9930 S.n7192 S.n7191 0.004
R9931 S.n665 S.n656 0.004
R9932 S.n6429 S.n6427 0.004
R9933 S.n5655 S.n5654 0.004
R9934 S.n632 S.n623 0.004
R9935 S.n4857 S.n4855 0.004
R9936 S.n4039 S.n4038 0.004
R9937 S.n599 S.n590 0.004
R9938 S.n3138 S.n3136 0.004
R9939 S.n2355 S.n2354 0.004
R9940 S.n566 S.n557 0.004
R9941 S.n1482 S.n1480 0.004
R9942 S.n534 S.n533 0.004
R9943 S.n1335 S.n1334 0.004
R9944 S.n9680 S.n9679 0.004
R9945 S.n9008 S.n9007 0.004
R9946 S.n8313 S.n8312 0.004
R9947 S.n7606 S.n7605 0.004
R9948 S.n6876 S.n6875 0.004
R9949 S.n6134 S.n6133 0.004
R9950 S.n5369 S.n5368 0.004
R9951 S.n4592 S.n4591 0.004
R9952 S.n3792 S.n3791 0.004
R9953 S.n2980 S.n2979 0.004
R9954 S.n2144 S.n2143 0.004
R9955 S.n11363 S.n11358 0.004
R9956 S.n10392 S.n10390 0.004
R9957 S.n9732 S.n9730 0.004
R9958 S.n9060 S.n9058 0.004
R9959 S.n8365 S.n8363 0.004
R9960 S.n7658 S.n7656 0.004
R9961 S.n6928 S.n6926 0.004
R9962 S.n6186 S.n6184 0.004
R9963 S.n5421 S.n5419 0.004
R9964 S.n4644 S.n4642 0.004
R9965 S.n3844 S.n3842 0.004
R9966 S.n3032 S.n3030 0.004
R9967 S.n2196 S.n2194 0.004
R9968 S.n1361 S.n1359 0.004
R9969 S.n1702 S.n1701 0.004
R9970 S.n9816 S.n9815 0.004
R9971 S.n10056 S.n10040 0.004
R9972 S.n8449 S.n8448 0.004
R9973 S.n8477 S.n8461 0.004
R9974 S.n7012 S.n7011 0.004
R9975 S.n7192 S.n7176 0.004
R9976 S.n5505 S.n5504 0.004
R9977 S.n5655 S.n5639 0.004
R9978 S.n3928 S.n3927 0.004
R9979 S.n4039 S.n4023 0.004
R9980 S.n2281 S.n2280 0.004
R9981 S.n2355 S.n2339 0.004
R9982 S.n2695 S.n2681 0.004
R9983 S.n2696 S.n2695 0.004
R9984 S.n3537 S.n3536 0.004
R9985 S.n3536 S.n3522 0.004
R9986 S.n4368 S.n4354 0.004
R9987 S.n4369 S.n4368 0.004
R9988 S.n5174 S.n5160 0.004
R9989 S.n5175 S.n5174 0.004
R9990 S.n5971 S.n5957 0.004
R9991 S.n5972 S.n5971 0.004
R9992 S.n6742 S.n6728 0.004
R9993 S.n6743 S.n6742 0.004
R9994 S.n7504 S.n7490 0.004
R9995 S.n7505 S.n7504 0.004
R9996 S.n8240 S.n8226 0.004
R9997 S.n8241 S.n8240 0.004
R9998 S.n8967 S.n8953 0.004
R9999 S.n8968 S.n8967 0.004
R10000 S.n9668 S.n9654 0.004
R10001 S.n9669 S.n9668 0.004
R10002 S.n10360 S.n10346 0.004
R10003 S.n10361 S.n10360 0.004
R10004 S.n11024 S.n11010 0.004
R10005 S.n11025 S.n11024 0.004
R10006 S.n12274 S.n12272 0.004
R10007 S.n11635 S.n11634 0.004
R10008 S.n11644 S.n11643 0.004
R10009 S.t0 S.n11993 0.004
R10010 S.t244 S.n537 0.004
R10011 S.t7 S.n211 0.004
R10012 S.t7 S.n208 0.004
R10013 S.t7 S.n160 0.004
R10014 S.t225 S.n9366 0.004
R10015 S.t7 S.n235 0.004
R10016 S.t124 S.n10059 0.004
R10017 S.t7 S.n175 0.004
R10018 S.t144 S.n10728 0.004
R10019 S.t7 S.n189 0.004
R10020 S.t47 S.n11366 0.004
R10021 S.t106 S.n12288 0.004
R10022 S.t7 S.n199 0.004
R10023 S.t7 S.n148 0.004
R10024 S.t11 S.n7767 0.004
R10025 S.t7 S.n231 0.004
R10026 S.t40 S.n8480 0.004
R10027 S.t7 S.n136 0.004
R10028 S.t4 S.n6432 0.004
R10029 S.t7 S.n227 0.004
R10030 S.t102 S.n7195 0.004
R10031 S.t7 S.n123 0.004
R10032 S.t77 S.n4860 0.004
R10033 S.t7 S.n223 0.004
R10034 S.t25 S.n5658 0.004
R10035 S.t7 S.n110 0.004
R10036 S.t38 S.n3141 0.004
R10037 S.t7 S.n219 0.004
R10038 S.t94 S.n4042 0.004
R10039 S.t7 S.n97 0.004
R10040 S.t175 S.n1485 0.004
R10041 S.t7 S.n215 0.004
R10042 S.t187 S.n2358 0.004
R10043 S.t7 S.n84 0.004
R10044 S.t0 S.n11933 0.004
R10045 S.t0 S.n11937 0.004
R10046 S.t0 S.n11941 0.004
R10047 S.t0 S.n11945 0.004
R10048 S.t0 S.n11949 0.004
R10049 S.t0 S.n11953 0.004
R10050 S.t0 S.n11957 0.004
R10051 S.t0 S.n11961 0.004
R10052 S.t0 S.n11965 0.004
R10053 S.t0 S.n11969 0.004
R10054 S.t0 S.n11973 0.004
R10055 S.t0 S.n11977 0.004
R10056 S.t0 S.n11981 0.004
R10057 S.t0 S.n11985 0.004
R10058 S.t0 S.n11989 0.004
R10059 S.t0 S.n11928 0.004
R10060 S.t7 S.n206 0.004
R10061 S.t65 S.n11919 0.004
R10062 S.t7 S.n7 0.004
R10063 S.t7 S.n15 0.004
R10064 S.t7 S.n24 0.004
R10065 S.t7 S.n33 0.004
R10066 S.t7 S.n42 0.004
R10067 S.t7 S.n51 0.004
R10068 S.t7 S.n55 0.004
R10069 S.n822 S.n821 0.004
R10070 S.t7 S.n203 0.004
R10071 S.t7 S.n152 0.004
R10072 S.t7 S.n140 0.004
R10073 S.t7 S.n127 0.004
R10074 S.t7 S.n114 0.004
R10075 S.t7 S.n101 0.004
R10076 S.t7 S.n88 0.004
R10077 S.n12285 S.n12284 0.004
R10078 S.n10074 S.n10063 0.004
R10079 S.n9398 S.n9387 0.004
R10080 S.n8531 S.n8520 0.004
R10081 S.n7835 S.n7824 0.004
R10082 S.n7282 S.n7271 0.004
R10083 S.n6536 S.n6525 0.004
R10084 S.n5781 S.n5770 0.004
R10085 S.n5000 S.n4989 0.004
R10086 S.n4201 S.n4190 0.004
R10087 S.n3317 S.n3306 0.004
R10088 S.n2553 S.n2542 0.004
R10089 S.n11914 S.n11913 0.003
R10090 S.n12333 S.n12332 0.003
R10091 S.n12591 S.n12590 0.003
R10092 S.n953 S.n952 0.003
R10093 S.n926 S.n925 0.003
R10094 S.n1437 S.n1436 0.003
R10095 S.n11897 S.n11896 0.003
R10096 S.n12309 S.n12308 0.003
R10097 S.n12029 S.n12028 0.003
R10098 S.n11407 S.n11406 0.003
R10099 S.n11081 S.n11080 0.003
R10100 S.n10790 S.n10789 0.003
R10101 S.n10451 S.n10450 0.003
R10102 S.n10140 S.n10139 0.003
R10103 S.n9791 S.n9790 0.003
R10104 S.n9464 S.n9463 0.003
R10105 S.n9119 S.n9118 0.003
R10106 S.n8597 S.n8596 0.003
R10107 S.n8424 S.n8423 0.003
R10108 S.n7901 S.n7900 0.003
R10109 S.n7717 S.n7716 0.003
R10110 S.n7348 S.n7347 0.003
R10111 S.n6987 S.n6986 0.003
R10112 S.n6602 S.n6601 0.003
R10113 S.n6245 S.n6244 0.003
R10114 S.n5847 S.n5846 0.003
R10115 S.n5480 S.n5479 0.003
R10116 S.n5066 S.n5065 0.003
R10117 S.n4703 S.n4702 0.003
R10118 S.n4267 S.n4266 0.003
R10119 S.n3903 S.n3902 0.003
R10120 S.n3383 S.n3382 0.003
R10121 S.n3091 S.n3090 0.003
R10122 S.n2619 S.n2618 0.003
R10123 S.n2256 S.n2255 0.003
R10124 S.n1768 S.n1767 0.003
R10125 S.n793 S.n792 0.003
R10126 S.n490 S.n489 0.003
R10127 S.n1288 S.n1287 0.003
R10128 S.n9142 S.n9141 0.003
R10129 S.n8501 S.n8500 0.003
R10130 S.n8277 S.n8276 0.003
R10131 S.n7805 S.n7804 0.003
R10132 S.n7570 S.n7569 0.003
R10133 S.n7252 S.n7251 0.003
R10134 S.n6840 S.n6839 0.003
R10135 S.n6506 S.n6505 0.003
R10136 S.n6098 S.n6097 0.003
R10137 S.n5751 S.n5750 0.003
R10138 S.n5333 S.n5332 0.003
R10139 S.n4970 S.n4969 0.003
R10140 S.n4556 S.n4555 0.003
R10141 S.n4171 S.n4170 0.003
R10142 S.n3756 S.n3755 0.003
R10143 S.n3287 S.n3286 0.003
R10144 S.n2944 S.n2943 0.003
R10145 S.n2523 S.n2522 0.003
R10146 S.n2107 S.n2106 0.003
R10147 S.n1667 S.n1666 0.003
R10148 S.n513 S.n512 0.003
R10149 S.n9819 S.n9818 0.003
R10150 S.n9385 S.n9384 0.003
R10151 S.n9001 S.n9000 0.003
R10152 S.n8518 S.n8517 0.003
R10153 S.n8306 S.n8305 0.003
R10154 S.n7822 S.n7821 0.003
R10155 S.n7599 S.n7598 0.003
R10156 S.n7269 S.n7268 0.003
R10157 S.n6869 S.n6868 0.003
R10158 S.n6523 S.n6522 0.003
R10159 S.n6127 S.n6126 0.003
R10160 S.n5768 S.n5767 0.003
R10161 S.n5362 S.n5361 0.003
R10162 S.n4987 S.n4986 0.003
R10163 S.n4585 S.n4584 0.003
R10164 S.n4188 S.n4187 0.003
R10165 S.n3785 S.n3784 0.003
R10166 S.n3304 S.n3303 0.003
R10167 S.n2973 S.n2972 0.003
R10168 S.n2540 S.n2539 0.003
R10169 S.n2136 S.n2135 0.003
R10170 S.n1686 S.n1685 0.003
R10171 S.n1708 S.n1707 0.003
R10172 S.n1350 S.n1349 0.003
R10173 S.n814 S.n813 0.003
R10174 S.n843 S.n842 0.003
R10175 S.n2169 S.n2168 0.003
R10176 S.n3005 S.n3004 0.003
R10177 S.n3817 S.n3816 0.003
R10178 S.n4617 S.n4616 0.003
R10179 S.n5394 S.n5393 0.003
R10180 S.n6159 S.n6158 0.003
R10181 S.n6901 S.n6900 0.003
R10182 S.n7631 S.n7630 0.003
R10183 S.n8338 S.n8337 0.003
R10184 S.n9033 S.n9032 0.003
R10185 S.n9705 S.n9704 0.003
R10186 S.n10477 S.n10476 0.003
R10187 S.n10080 S.n10079 0.003
R10188 S.n9404 S.n9403 0.003
R10189 S.n8537 S.n8536 0.003
R10190 S.n7841 S.n7840 0.003
R10191 S.n7288 S.n7287 0.003
R10192 S.n6542 S.n6541 0.003
R10193 S.n5787 S.n5786 0.003
R10194 S.n5006 S.n5005 0.003
R10195 S.n4207 S.n4206 0.003
R10196 S.n3323 S.n3322 0.003
R10197 S.n2559 S.n2558 0.003
R10198 S.n1384 S.n1383 0.003
R10199 S.n757 S.n756 0.003
R10200 S.n876 S.n875 0.003
R10201 S.n11105 S.n11104 0.003
R10202 S.n10751 S.n10750 0.003
R10203 S.n10399 S.n10398 0.003
R10204 S.n10101 S.n10100 0.003
R10205 S.n9739 S.n9738 0.003
R10206 S.n9425 S.n9424 0.003
R10207 S.n9067 S.n9066 0.003
R10208 S.n8558 S.n8557 0.003
R10209 S.n8372 S.n8371 0.003
R10210 S.n7862 S.n7861 0.003
R10211 S.n7665 S.n7664 0.003
R10212 S.n7309 S.n7308 0.003
R10213 S.n6935 S.n6934 0.003
R10214 S.n6563 S.n6562 0.003
R10215 S.n6193 S.n6192 0.003
R10216 S.n5808 S.n5807 0.003
R10217 S.n5428 S.n5427 0.003
R10218 S.n5027 S.n5026 0.003
R10219 S.n4651 S.n4650 0.003
R10220 S.n4228 S.n4227 0.003
R10221 S.n3851 S.n3850 0.003
R10222 S.n3344 S.n3343 0.003
R10223 S.n3039 S.n3038 0.003
R10224 S.n2580 S.n2579 0.003
R10225 S.n2203 S.n2202 0.003
R10226 S.n1729 S.n1728 0.003
R10227 S.n1412 S.n1411 0.003
R10228 S.n776 S.n775 0.003
R10229 S.n1749 S.n1748 0.003
R10230 S.n2224 S.n2223 0.003
R10231 S.n2600 S.n2599 0.003
R10232 S.n3059 S.n3058 0.003
R10233 S.n3364 S.n3363 0.003
R10234 S.n3871 S.n3870 0.003
R10235 S.n4248 S.n4247 0.003
R10236 S.n4671 S.n4670 0.003
R10237 S.n5047 S.n5046 0.003
R10238 S.n5448 S.n5447 0.003
R10239 S.n5828 S.n5827 0.003
R10240 S.n6213 S.n6212 0.003
R10241 S.n6583 S.n6582 0.003
R10242 S.n6955 S.n6954 0.003
R10243 S.n7329 S.n7328 0.003
R10244 S.n7685 S.n7684 0.003
R10245 S.n7882 S.n7881 0.003
R10246 S.n8392 S.n8391 0.003
R10247 S.n8578 S.n8577 0.003
R10248 S.n9087 S.n9086 0.003
R10249 S.n9445 S.n9444 0.003
R10250 S.n9759 S.n9758 0.003
R10251 S.n10121 S.n10120 0.003
R10252 S.n10419 S.n10418 0.003
R10253 S.n10771 S.n10770 0.003
R10254 S.n11049 S.n11048 0.003
R10255 S.n11388 S.n11387 0.003
R10256 S.n12050 S.n12049 0.003
R10257 S.n905 S.n904 0.003
R10258 S.n1316 S.n1315 0.003
R10259 S.n737 S.n736 0.003
R10260 S.n720 S.n719 0.003
R10261 S.n446 S.n445 0.003
R10262 S.n1229 S.n1228 0.003
R10263 S.n7740 S.n7739 0.003
R10264 S.n7216 S.n7215 0.003
R10265 S.n6779 S.n6778 0.003
R10266 S.n6470 S.n6469 0.003
R10267 S.n6037 S.n6036 0.003
R10268 S.n5715 S.n5714 0.003
R10269 S.n5272 S.n5271 0.003
R10270 S.n4934 S.n4933 0.003
R10271 S.n4495 S.n4494 0.003
R10272 S.n4135 S.n4134 0.003
R10273 S.n3695 S.n3694 0.003
R10274 S.n3251 S.n3250 0.003
R10275 S.n2883 S.n2882 0.003
R10276 S.n2487 S.n2486 0.003
R10277 S.n2046 S.n2045 0.003
R10278 S.n1631 S.n1630 0.003
R10279 S.n461 S.n460 0.003
R10280 S.n8452 S.n8451 0.003
R10281 S.n7786 S.n7785 0.003
R10282 S.n7538 S.n7537 0.003
R10283 S.n7233 S.n7232 0.003
R10284 S.n6808 S.n6807 0.003
R10285 S.n6487 S.n6486 0.003
R10286 S.n6066 S.n6065 0.003
R10287 S.n5732 S.n5731 0.003
R10288 S.n5301 S.n5300 0.003
R10289 S.n4951 S.n4950 0.003
R10290 S.n4524 S.n4523 0.003
R10291 S.n4152 S.n4151 0.003
R10292 S.n3724 S.n3723 0.003
R10293 S.n3268 S.n3267 0.003
R10294 S.n2912 S.n2911 0.003
R10295 S.n2504 S.n2503 0.003
R10296 S.n2075 S.n2074 0.003
R10297 S.n1648 S.n1647 0.003
R10298 S.n1258 S.n1257 0.003
R10299 S.n704 S.n703 0.003
R10300 S.n687 S.n686 0.003
R10301 S.n402 S.n401 0.003
R10302 S.n1170 S.n1169 0.003
R10303 S.n6268 S.n6267 0.003
R10304 S.n5679 S.n5678 0.003
R10305 S.n5211 S.n5210 0.003
R10306 S.n4898 S.n4897 0.003
R10307 S.n4434 S.n4433 0.003
R10308 S.n4099 S.n4098 0.003
R10309 S.n3634 S.n3633 0.003
R10310 S.n3215 S.n3214 0.003
R10311 S.n2822 S.n2821 0.003
R10312 S.n2451 S.n2450 0.003
R10313 S.n1985 S.n1984 0.003
R10314 S.n1595 S.n1594 0.003
R10315 S.n425 S.n424 0.003
R10316 S.n7015 S.n7014 0.003
R10317 S.n6451 S.n6450 0.003
R10318 S.n6005 S.n6004 0.003
R10319 S.n5696 S.n5695 0.003
R10320 S.n5240 S.n5239 0.003
R10321 S.n4915 S.n4914 0.003
R10322 S.n4463 S.n4462 0.003
R10323 S.n4116 S.n4115 0.003
R10324 S.n3663 S.n3662 0.003
R10325 S.n3232 S.n3231 0.003
R10326 S.n2851 S.n2850 0.003
R10327 S.n2468 S.n2467 0.003
R10328 S.n2014 S.n2013 0.003
R10329 S.n1612 S.n1611 0.003
R10330 S.n1199 S.n1198 0.003
R10331 S.n671 S.n670 0.003
R10332 S.n654 S.n653 0.003
R10333 S.n358 S.n357 0.003
R10334 S.n1111 S.n1110 0.003
R10335 S.n4726 S.n4725 0.003
R10336 S.n4063 S.n4062 0.003
R10337 S.n3573 S.n3572 0.003
R10338 S.n3179 S.n3178 0.003
R10339 S.n2761 S.n2760 0.003
R10340 S.n2415 S.n2414 0.003
R10341 S.n1924 S.n1923 0.003
R10342 S.n1559 S.n1558 0.003
R10343 S.n381 S.n380 0.003
R10344 S.n5508 S.n5507 0.003
R10345 S.n4879 S.n4878 0.003
R10346 S.n4402 S.n4401 0.003
R10347 S.n4080 S.n4079 0.003
R10348 S.n3602 S.n3601 0.003
R10349 S.n3196 S.n3195 0.003
R10350 S.n2790 S.n2789 0.003
R10351 S.n2432 S.n2431 0.003
R10352 S.n1953 S.n1952 0.003
R10353 S.n1576 S.n1575 0.003
R10354 S.n1140 S.n1139 0.003
R10355 S.n638 S.n637 0.003
R10356 S.n621 S.n620 0.003
R10357 S.n314 S.n313 0.003
R10358 S.n1052 S.n1051 0.003
R10359 S.n3114 S.n3113 0.003
R10360 S.n2379 S.n2378 0.003
R10361 S.n1863 S.n1862 0.003
R10362 S.n1523 S.n1522 0.003
R10363 S.n337 S.n336 0.003
R10364 S.n3931 S.n3930 0.003
R10365 S.n3160 S.n3159 0.003
R10366 S.n2729 S.n2728 0.003
R10367 S.n2396 S.n2395 0.003
R10368 S.n1892 S.n1891 0.003
R10369 S.n1540 S.n1539 0.003
R10370 S.n1081 S.n1080 0.003
R10371 S.n605 S.n604 0.003
R10372 S.n588 S.n587 0.003
R10373 S.n270 S.n269 0.003
R10374 S.n1458 S.n1457 0.003
R10375 S.n293 S.n292 0.003
R10376 S.n2284 S.n2283 0.003
R10377 S.n1504 S.n1503 0.003
R10378 S.n1022 S.n1021 0.003
R10379 S.n572 S.n571 0.003
R10380 S.n555 S.n554 0.003
R10381 S.n959 S.n958 0.003
R10382 S.n808 S.n807 0.003
R10383 S.n1811 S.n1810 0.003
R10384 S.n1788 S.n1787 0.003
R10385 S.n2321 S.n2320 0.003
R10386 S.n2294 S.n2293 0.003
R10387 S.n3449 S.n3448 0.003
R10388 S.n3422 S.n3421 0.003
R10389 S.n3968 S.n3967 0.003
R10390 S.n3941 S.n3940 0.003
R10391 S.n4763 S.n4762 0.003
R10392 S.n4736 S.n4735 0.003
R10393 S.n5545 S.n5544 0.003
R10394 S.n5518 S.n5517 0.003
R10395 S.n6305 S.n6304 0.003
R10396 S.n6278 S.n6277 0.003
R10397 S.n7052 S.n7051 0.003
R10398 S.n7025 S.n7024 0.003
R10399 S.n8063 S.n8062 0.003
R10400 S.n8036 S.n8035 0.003
R10401 S.n8775 S.n8774 0.003
R10402 S.n8748 S.n8747 0.003
R10403 S.n9179 S.n9178 0.003
R10404 S.n9152 S.n9151 0.003
R10405 S.n9856 S.n9855 0.003
R10406 S.n9829 S.n9828 0.003
R10407 S.n10514 S.n10513 0.003
R10408 S.n10487 S.n10486 0.003
R10409 S.n11142 S.n11141 0.003
R10410 S.n11115 S.n11114 0.003
R10411 S.n12070 S.n12069 0.003
R10412 S.n12347 S.n12346 0.003
R10413 S.n11876 S.n11875 0.003
R10414 S.n1817 S.n1816 0.003
R10415 S.n1782 S.n1781 0.003
R10416 S.n2654 S.n2653 0.003
R10417 S.n11858 S.n11857 0.003
R10418 S.n12362 S.n12361 0.003
R10419 S.n12086 S.n12085 0.003
R10420 S.n11164 S.n11163 0.003
R10421 S.n11173 S.n11172 0.003
R10422 S.n10536 S.n10535 0.003
R10423 S.n10545 S.n10544 0.003
R10424 S.n9878 S.n9877 0.003
R10425 S.n9887 S.n9886 0.003
R10426 S.n9201 S.n9200 0.003
R10427 S.n9210 S.n9209 0.003
R10428 S.n8797 S.n8796 0.003
R10429 S.n8806 S.n8805 0.003
R10430 S.n8085 S.n8084 0.003
R10431 S.n8094 S.n8093 0.003
R10432 S.n7074 S.n7073 0.003
R10433 S.n7083 S.n7082 0.003
R10434 S.n6327 S.n6326 0.003
R10435 S.n6336 S.n6335 0.003
R10436 S.n5567 S.n5566 0.003
R10437 S.n5576 S.n5575 0.003
R10438 S.n4785 S.n4784 0.003
R10439 S.n4794 S.n4793 0.003
R10440 S.n3990 S.n3989 0.003
R10441 S.n3999 S.n3998 0.003
R10442 S.n3471 S.n3470 0.003
R10443 S.n3480 S.n3479 0.003
R10444 S.n2646 S.n2645 0.003
R10445 S.n2660 S.n2659 0.003
R10446 S.n2637 S.n2636 0.003
R10447 S.n3495 S.n3494 0.003
R10448 S.n11843 S.n11842 0.003
R10449 S.n12378 S.n12377 0.003
R10450 S.n12101 S.n12100 0.003
R10451 S.n11420 S.n11419 0.003
R10452 S.n11188 S.n11187 0.003
R10453 S.n10804 S.n10803 0.003
R10454 S.n10560 S.n10559 0.003
R10455 S.n10154 S.n10153 0.003
R10456 S.n9902 S.n9901 0.003
R10457 S.n9478 S.n9477 0.003
R10458 S.n9225 S.n9224 0.003
R10459 S.n8611 S.n8610 0.003
R10460 S.n8821 S.n8820 0.003
R10461 S.n7915 S.n7914 0.003
R10462 S.n8109 S.n8108 0.003
R10463 S.n7362 S.n7361 0.003
R10464 S.n7098 S.n7097 0.003
R10465 S.n6616 S.n6615 0.003
R10466 S.n6351 S.n6350 0.003
R10467 S.n5861 S.n5860 0.003
R10468 S.n5591 S.n5590 0.003
R10469 S.n5080 S.n5079 0.003
R10470 S.n4809 S.n4808 0.003
R10471 S.n4281 S.n4280 0.003
R10472 S.n4014 S.n4013 0.003
R10473 S.n3396 S.n3395 0.003
R10474 S.n11828 S.n11827 0.003
R10475 S.n12394 S.n12393 0.003
R10476 S.n12116 S.n12115 0.003
R10477 S.n11436 S.n11435 0.003
R10478 S.n11203 S.n11202 0.003
R10479 S.n10820 S.n10819 0.003
R10480 S.n10575 S.n10574 0.003
R10481 S.n10170 S.n10169 0.003
R10482 S.n9917 S.n9916 0.003
R10483 S.n9494 S.n9493 0.003
R10484 S.n9240 S.n9239 0.003
R10485 S.n8627 S.n8626 0.003
R10486 S.n8836 S.n8835 0.003
R10487 S.n7931 S.n7930 0.003
R10488 S.n8124 S.n8123 0.003
R10489 S.n7378 S.n7377 0.003
R10490 S.n7113 S.n7112 0.003
R10491 S.n6632 S.n6631 0.003
R10492 S.n6366 S.n6365 0.003
R10493 S.n5877 S.n5876 0.003
R10494 S.n5606 S.n5605 0.003
R10495 S.n5096 S.n5095 0.003
R10496 S.n4824 S.n4823 0.003
R10497 S.n4307 S.n4306 0.003
R10498 S.n4327 S.n4326 0.003
R10499 S.n3416 S.n3415 0.003
R10500 S.n3501 S.n3500 0.003
R10501 S.n4333 S.n4332 0.003
R10502 S.n4301 S.n4300 0.003
R10503 S.n5133 S.n5132 0.003
R10504 S.n11813 S.n11812 0.003
R10505 S.n12410 S.n12409 0.003
R10506 S.n12131 S.n12130 0.003
R10507 S.n11452 S.n11451 0.003
R10508 S.n11218 S.n11217 0.003
R10509 S.n10836 S.n10835 0.003
R10510 S.n10590 S.n10589 0.003
R10511 S.n10186 S.n10185 0.003
R10512 S.n9932 S.n9931 0.003
R10513 S.n9510 S.n9509 0.003
R10514 S.n9255 S.n9254 0.003
R10515 S.n8643 S.n8642 0.003
R10516 S.n8851 S.n8850 0.003
R10517 S.n7947 S.n7946 0.003
R10518 S.n8139 S.n8138 0.003
R10519 S.n7394 S.n7393 0.003
R10520 S.n7128 S.n7127 0.003
R10521 S.n6648 S.n6647 0.003
R10522 S.n6381 S.n6380 0.003
R10523 S.n5893 S.n5892 0.003
R10524 S.n5621 S.n5620 0.003
R10525 S.n5125 S.n5124 0.003
R10526 S.n5139 S.n5138 0.003
R10527 S.n5116 S.n5115 0.003
R10528 S.n5930 S.n5929 0.003
R10529 S.n11798 S.n11797 0.003
R10530 S.n12426 S.n12425 0.003
R10531 S.n12146 S.n12145 0.003
R10532 S.n11468 S.n11467 0.003
R10533 S.n11233 S.n11232 0.003
R10534 S.n10852 S.n10851 0.003
R10535 S.n10605 S.n10604 0.003
R10536 S.n10202 S.n10201 0.003
R10537 S.n9947 S.n9946 0.003
R10538 S.n9526 S.n9525 0.003
R10539 S.n9270 S.n9269 0.003
R10540 S.n8659 S.n8658 0.003
R10541 S.n8866 S.n8865 0.003
R10542 S.n7963 S.n7962 0.003
R10543 S.n8154 S.n8153 0.003
R10544 S.n7410 S.n7409 0.003
R10545 S.n7143 S.n7142 0.003
R10546 S.n6664 S.n6663 0.003
R10547 S.n6396 S.n6395 0.003
R10548 S.n5922 S.n5921 0.003
R10549 S.n5936 S.n5935 0.003
R10550 S.n5913 S.n5912 0.003
R10551 S.n6701 S.n6700 0.003
R10552 S.n11783 S.n11782 0.003
R10553 S.n12442 S.n12441 0.003
R10554 S.n12161 S.n12160 0.003
R10555 S.n11484 S.n11483 0.003
R10556 S.n11248 S.n11247 0.003
R10557 S.n10868 S.n10867 0.003
R10558 S.n10620 S.n10619 0.003
R10559 S.n10218 S.n10217 0.003
R10560 S.n9962 S.n9961 0.003
R10561 S.n9542 S.n9541 0.003
R10562 S.n9285 S.n9284 0.003
R10563 S.n8675 S.n8674 0.003
R10564 S.n8881 S.n8880 0.003
R10565 S.n7979 S.n7978 0.003
R10566 S.n8169 S.n8168 0.003
R10567 S.n7426 S.n7425 0.003
R10568 S.n7158 S.n7157 0.003
R10569 S.n6693 S.n6692 0.003
R10570 S.n6707 S.n6706 0.003
R10571 S.n6684 S.n6683 0.003
R10572 S.n7463 S.n7462 0.003
R10573 S.n11768 S.n11767 0.003
R10574 S.n12458 S.n12457 0.003
R10575 S.n12176 S.n12175 0.003
R10576 S.n11500 S.n11499 0.003
R10577 S.n11263 S.n11262 0.003
R10578 S.n10884 S.n10883 0.003
R10579 S.n10635 S.n10634 0.003
R10580 S.n10234 S.n10233 0.003
R10581 S.n9977 S.n9976 0.003
R10582 S.n9558 S.n9557 0.003
R10583 S.n9300 S.n9299 0.003
R10584 S.n8691 S.n8690 0.003
R10585 S.n8896 S.n8895 0.003
R10586 S.n7995 S.n7994 0.003
R10587 S.n8184 S.n8183 0.003
R10588 S.n7455 S.n7454 0.003
R10589 S.n7469 S.n7468 0.003
R10590 S.n7446 S.n7445 0.003
R10591 S.n8199 S.n8198 0.003
R10592 S.n11753 S.n11752 0.003
R10593 S.n12474 S.n12473 0.003
R10594 S.n12191 S.n12190 0.003
R10595 S.n11516 S.n11515 0.003
R10596 S.n11278 S.n11277 0.003
R10597 S.n10900 S.n10899 0.003
R10598 S.n10650 S.n10649 0.003
R10599 S.n10250 S.n10249 0.003
R10600 S.n9992 S.n9991 0.003
R10601 S.n9574 S.n9573 0.003
R10602 S.n9315 S.n9314 0.003
R10603 S.n8707 S.n8706 0.003
R10604 S.n8911 S.n8910 0.003
R10605 S.n8010 S.n8009 0.003
R10606 S.n8205 S.n8204 0.003
R10607 S.n8030 S.n8029 0.003
R10608 S.n8926 S.n8925 0.003
R10609 S.n11738 S.n11737 0.003
R10610 S.n12490 S.n12489 0.003
R10611 S.n12206 S.n12205 0.003
R10612 S.n11532 S.n11531 0.003
R10613 S.n11293 S.n11292 0.003
R10614 S.n10916 S.n10915 0.003
R10615 S.n10665 S.n10664 0.003
R10616 S.n10266 S.n10265 0.003
R10617 S.n10007 S.n10006 0.003
R10618 S.n9590 S.n9589 0.003
R10619 S.n9330 S.n9329 0.003
R10620 S.n8722 S.n8721 0.003
R10621 S.n8932 S.n8931 0.003
R10622 S.n8742 S.n8741 0.003
R10623 S.n9627 S.n9626 0.003
R10624 S.n11723 S.n11722 0.003
R10625 S.n12506 S.n12505 0.003
R10626 S.n12221 S.n12220 0.003
R10627 S.n11548 S.n11547 0.003
R10628 S.n11308 S.n11307 0.003
R10629 S.n10932 S.n10931 0.003
R10630 S.n10680 S.n10679 0.003
R10631 S.n10282 S.n10281 0.003
R10632 S.n10022 S.n10021 0.003
R10633 S.n9619 S.n9618 0.003
R10634 S.n9633 S.n9632 0.003
R10635 S.n9610 S.n9609 0.003
R10636 S.n10319 S.n10318 0.003
R10637 S.n11708 S.n11707 0.003
R10638 S.n12522 S.n12521 0.003
R10639 S.n12236 S.n12235 0.003
R10640 S.n11564 S.n11563 0.003
R10641 S.n11323 S.n11322 0.003
R10642 S.n10948 S.n10947 0.003
R10643 S.n10695 S.n10694 0.003
R10644 S.n10311 S.n10310 0.003
R10645 S.n10325 S.n10324 0.003
R10646 S.n10302 S.n10301 0.003
R10647 S.n10985 S.n10984 0.003
R10648 S.n11693 S.n11692 0.003
R10649 S.n12538 S.n12537 0.003
R10650 S.n12251 S.n12250 0.003
R10651 S.n11580 S.n11579 0.003
R10652 S.n11338 S.n11337 0.003
R10653 S.n10977 S.n10976 0.003
R10654 S.n10991 S.n10990 0.003
R10655 S.n10968 S.n10967 0.003
R10656 S.n11620 S.n11619 0.003
R10657 S.n11678 S.n11677 0.003
R10658 S.n12554 S.n12553 0.003
R10659 S.n12266 S.n12265 0.003
R10660 S.n11612 S.n11611 0.003
R10661 S.n11626 S.n11625 0.003
R10662 S.n11603 S.n11602 0.003
R10663 S.n12585 S.n12584 0.003
R10664 S.n11663 S.n11662 0.003
R10665 S.n12560 S.n12559 0.003
R10666 S.n1680 S.n1679 0.003
R10667 S.n11911 S.n11906 0.003
R10668 S.n12327 S.n12315 0.003
R10669 S.n950 S.n938 0.003
R10670 S.n920 S.n915 0.003
R10671 S.n1431 S.n1420 0.003
R10672 S.n11891 S.n11886 0.003
R10673 S.n12303 S.n12298 0.003
R10674 S.n12023 S.n12014 0.003
R10675 S.n11401 S.n11396 0.003
R10676 S.n11075 S.n11066 0.003
R10677 S.n10784 S.n10779 0.003
R10678 S.n10445 S.n10436 0.003
R10679 S.n10134 S.n10129 0.003
R10680 S.n9785 S.n9776 0.003
R10681 S.n9458 S.n9453 0.003
R10682 S.n9113 S.n9104 0.003
R10683 S.n8591 S.n8586 0.003
R10684 S.n8418 S.n8409 0.003
R10685 S.n7895 S.n7890 0.003
R10686 S.n7711 S.n7702 0.003
R10687 S.n7342 S.n7337 0.003
R10688 S.n6981 S.n6972 0.003
R10689 S.n6596 S.n6591 0.003
R10690 S.n6239 S.n6230 0.003
R10691 S.n5841 S.n5836 0.003
R10692 S.n5474 S.n5465 0.003
R10693 S.n5060 S.n5055 0.003
R10694 S.n4697 S.n4688 0.003
R10695 S.n4261 S.n4256 0.003
R10696 S.n3897 S.n3888 0.003
R10697 S.n3377 S.n3372 0.003
R10698 S.n3085 S.n3076 0.003
R10699 S.n2613 S.n2608 0.003
R10700 S.n2250 S.n2241 0.003
R10701 S.n1762 S.n1757 0.003
R10702 S.n787 S.n782 0.003
R10703 S.n484 S.n479 0.003
R10704 S.n1282 S.n1275 0.003
R10705 S.n9139 S.n9128 0.003
R10706 S.n8495 S.n8490 0.003
R10707 S.n8271 S.n8262 0.003
R10708 S.n7799 S.n7794 0.003
R10709 S.n7564 S.n7555 0.003
R10710 S.n7246 S.n7241 0.003
R10711 S.n6834 S.n6825 0.003
R10712 S.n6500 S.n6495 0.003
R10713 S.n6092 S.n6083 0.003
R10714 S.n5745 S.n5740 0.003
R10715 S.n5327 S.n5318 0.003
R10716 S.n4964 S.n4959 0.003
R10717 S.n4550 S.n4541 0.003
R10718 S.n4165 S.n4160 0.003
R10719 S.n3750 S.n3741 0.003
R10720 S.n3281 S.n3276 0.003
R10721 S.n2938 S.n2929 0.003
R10722 S.n2517 S.n2512 0.003
R10723 S.n2101 S.n2092 0.003
R10724 S.n1661 S.n1656 0.003
R10725 S.n507 S.n502 0.003
R10726 S.n9816 S.n9804 0.003
R10727 S.n9379 S.n9374 0.003
R10728 S.n8995 S.n8981 0.003
R10729 S.n8512 S.n8507 0.003
R10730 S.n8300 S.n8286 0.003
R10731 S.n7816 S.n7811 0.003
R10732 S.n7593 S.n7579 0.003
R10733 S.n7263 S.n7258 0.003
R10734 S.n6863 S.n6849 0.003
R10735 S.n6517 S.n6512 0.003
R10736 S.n6121 S.n6107 0.003
R10737 S.n5762 S.n5757 0.003
R10738 S.n5356 S.n5342 0.003
R10739 S.n4981 S.n4976 0.003
R10740 S.n4579 S.n4565 0.003
R10741 S.n4182 S.n4177 0.003
R10742 S.n3779 S.n3765 0.003
R10743 S.n3298 S.n3293 0.003
R10744 S.n2967 S.n2953 0.003
R10745 S.n2534 S.n2529 0.003
R10746 S.n2130 S.n2116 0.003
R10747 S.n1680 S.n1673 0.003
R10748 S.n1702 S.n1694 0.003
R10749 S.n1344 S.n1326 0.003
R10750 S.n822 S.n517 0.003
R10751 S.n837 S.n828 0.003
R10752 S.n2163 S.n2154 0.003
R10753 S.n2999 S.n2990 0.003
R10754 S.n3811 S.n3802 0.003
R10755 S.n4611 S.n4602 0.003
R10756 S.n5388 S.n5379 0.003
R10757 S.n6153 S.n6144 0.003
R10758 S.n6895 S.n6886 0.003
R10759 S.n7625 S.n7616 0.003
R10760 S.n8332 S.n8323 0.003
R10761 S.n9027 S.n9018 0.003
R10762 S.n9699 S.n9690 0.003
R10763 S.n10474 S.n10463 0.003
R10764 S.n10074 S.n10069 0.003
R10765 S.n9398 S.n9393 0.003
R10766 S.n8531 S.n8526 0.003
R10767 S.n7835 S.n7830 0.003
R10768 S.n7282 S.n7277 0.003
R10769 S.n6536 S.n6531 0.003
R10770 S.n5781 S.n5776 0.003
R10771 S.n5000 S.n4995 0.003
R10772 S.n4201 S.n4196 0.003
R10773 S.n3317 S.n3312 0.003
R10774 S.n2553 S.n2548 0.003
R10775 S.n1378 S.n1365 0.003
R10776 S.n751 S.n742 0.003
R10777 S.n870 S.n860 0.003
R10778 S.n11102 S.n11097 0.003
R10779 S.n10745 S.n10743 0.003
R10780 S.n10393 S.n10381 0.003
R10781 S.n10095 S.n10093 0.003
R10782 S.n9733 S.n9721 0.003
R10783 S.n9419 S.n9417 0.003
R10784 S.n9061 S.n9049 0.003
R10785 S.n8552 S.n8550 0.003
R10786 S.n8366 S.n8354 0.003
R10787 S.n7856 S.n7854 0.003
R10788 S.n7659 S.n7647 0.003
R10789 S.n7303 S.n7301 0.003
R10790 S.n6929 S.n6917 0.003
R10791 S.n6557 S.n6555 0.003
R10792 S.n6187 S.n6175 0.003
R10793 S.n5802 S.n5800 0.003
R10794 S.n5422 S.n5410 0.003
R10795 S.n5021 S.n5019 0.003
R10796 S.n4645 S.n4633 0.003
R10797 S.n4222 S.n4220 0.003
R10798 S.n3845 S.n3833 0.003
R10799 S.n3338 S.n3336 0.003
R10800 S.n3033 S.n3021 0.003
R10801 S.n2574 S.n2572 0.003
R10802 S.n2197 S.n2185 0.003
R10803 S.n1723 S.n1721 0.003
R10804 S.n1406 S.n1393 0.003
R10805 S.n770 S.n762 0.003
R10806 S.n1743 S.n1740 0.003
R10807 S.n2218 S.n2212 0.003
R10808 S.n2594 S.n2586 0.003
R10809 S.n3053 S.n3048 0.003
R10810 S.n3358 S.n3350 0.003
R10811 S.n3865 S.n3860 0.003
R10812 S.n4242 S.n4234 0.003
R10813 S.n4665 S.n4660 0.003
R10814 S.n5041 S.n5033 0.003
R10815 S.n5442 S.n5437 0.003
R10816 S.n5822 S.n5814 0.003
R10817 S.n6207 S.n6202 0.003
R10818 S.n6577 S.n6569 0.003
R10819 S.n6949 S.n6944 0.003
R10820 S.n7323 S.n7315 0.003
R10821 S.n7679 S.n7674 0.003
R10822 S.n7876 S.n7868 0.003
R10823 S.n8386 S.n8381 0.003
R10824 S.n8572 S.n8564 0.003
R10825 S.n9081 S.n9076 0.003
R10826 S.n9439 S.n9431 0.003
R10827 S.n9753 S.n9748 0.003
R10828 S.n10115 S.n10107 0.003
R10829 S.n10413 S.n10408 0.003
R10830 S.n10765 S.n10757 0.003
R10831 S.n11043 S.n11038 0.003
R10832 S.n11382 S.n11374 0.003
R10833 S.n12047 S.n12042 0.003
R10834 S.n899 S.n886 0.003
R10835 S.n1310 S.n1297 0.003
R10836 S.n731 S.n726 0.003
R10837 S.n714 S.n709 0.003
R10838 S.n440 S.n435 0.003
R10839 S.n1223 S.n1216 0.003
R10840 S.n7737 S.n7726 0.003
R10841 S.n7210 S.n7205 0.003
R10842 S.n6773 S.n6764 0.003
R10843 S.n6464 S.n6459 0.003
R10844 S.n6031 S.n6022 0.003
R10845 S.n5709 S.n5704 0.003
R10846 S.n5266 S.n5257 0.003
R10847 S.n4928 S.n4923 0.003
R10848 S.n4489 S.n4480 0.003
R10849 S.n4129 S.n4124 0.003
R10850 S.n3689 S.n3680 0.003
R10851 S.n3245 S.n3240 0.003
R10852 S.n2877 S.n2868 0.003
R10853 S.n2481 S.n2476 0.003
R10854 S.n2040 S.n2031 0.003
R10855 S.n1625 S.n1620 0.003
R10856 S.n466 S.n458 0.003
R10857 S.n8449 S.n8437 0.003
R10858 S.n7780 S.n7775 0.003
R10859 S.n7532 S.n7518 0.003
R10860 S.n7227 S.n7222 0.003
R10861 S.n6802 S.n6788 0.003
R10862 S.n6481 S.n6476 0.003
R10863 S.n6060 S.n6046 0.003
R10864 S.n5726 S.n5721 0.003
R10865 S.n5295 S.n5281 0.003
R10866 S.n4945 S.n4940 0.003
R10867 S.n4518 S.n4504 0.003
R10868 S.n4146 S.n4141 0.003
R10869 S.n3718 S.n3704 0.003
R10870 S.n3262 S.n3257 0.003
R10871 S.n2906 S.n2892 0.003
R10872 S.n2498 S.n2493 0.003
R10873 S.n2069 S.n2055 0.003
R10874 S.n1642 S.n1637 0.003
R10875 S.n1252 S.n1238 0.003
R10876 S.n698 S.n693 0.003
R10877 S.n681 S.n676 0.003
R10878 S.n396 S.n391 0.003
R10879 S.n1164 S.n1157 0.003
R10880 S.n6265 S.n6254 0.003
R10881 S.n5673 S.n5668 0.003
R10882 S.n5205 S.n5196 0.003
R10883 S.n4892 S.n4887 0.003
R10884 S.n4428 S.n4419 0.003
R10885 S.n4093 S.n4088 0.003
R10886 S.n3628 S.n3619 0.003
R10887 S.n3209 S.n3204 0.003
R10888 S.n2816 S.n2807 0.003
R10889 S.n2445 S.n2440 0.003
R10890 S.n1979 S.n1970 0.003
R10891 S.n1589 S.n1584 0.003
R10892 S.n419 S.n414 0.003
R10893 S.n7012 S.n7000 0.003
R10894 S.n6445 S.n6440 0.003
R10895 S.n5999 S.n5985 0.003
R10896 S.n5690 S.n5685 0.003
R10897 S.n5234 S.n5220 0.003
R10898 S.n4909 S.n4904 0.003
R10899 S.n4457 S.n4443 0.003
R10900 S.n4110 S.n4105 0.003
R10901 S.n3657 S.n3643 0.003
R10902 S.n3226 S.n3221 0.003
R10903 S.n2845 S.n2831 0.003
R10904 S.n2462 S.n2457 0.003
R10905 S.n2008 S.n1994 0.003
R10906 S.n1606 S.n1601 0.003
R10907 S.n1193 S.n1179 0.003
R10908 S.n665 S.n660 0.003
R10909 S.n648 S.n643 0.003
R10910 S.n352 S.n347 0.003
R10911 S.n1105 S.n1098 0.003
R10912 S.n4723 S.n4712 0.003
R10913 S.n4057 S.n4052 0.003
R10914 S.n3567 S.n3558 0.003
R10915 S.n3173 S.n3168 0.003
R10916 S.n2755 S.n2746 0.003
R10917 S.n2409 S.n2404 0.003
R10918 S.n1918 S.n1909 0.003
R10919 S.n1553 S.n1548 0.003
R10920 S.n375 S.n370 0.003
R10921 S.n5505 S.n5493 0.003
R10922 S.n4873 S.n4868 0.003
R10923 S.n4396 S.n4382 0.003
R10924 S.n4074 S.n4069 0.003
R10925 S.n3596 S.n3582 0.003
R10926 S.n3190 S.n3185 0.003
R10927 S.n2784 S.n2770 0.003
R10928 S.n2426 S.n2421 0.003
R10929 S.n1950 S.n1933 0.003
R10930 S.n1570 S.n1565 0.003
R10931 S.n1134 S.n1120 0.003
R10932 S.n632 S.n627 0.003
R10933 S.n615 S.n610 0.003
R10934 S.n308 S.n303 0.003
R10935 S.n1046 S.n1039 0.003
R10936 S.n3111 S.n3100 0.003
R10937 S.n2373 S.n2368 0.003
R10938 S.n1857 S.n1848 0.003
R10939 S.n1517 S.n1512 0.003
R10940 S.n331 S.n326 0.003
R10941 S.n3928 S.n3916 0.003
R10942 S.n3154 S.n3149 0.003
R10943 S.n2723 S.n2709 0.003
R10944 S.n2390 S.n2385 0.003
R10945 S.n1886 S.n1872 0.003
R10946 S.n1534 S.n1529 0.003
R10947 S.n1075 S.n1061 0.003
R10948 S.n599 S.n594 0.003
R10949 S.n582 S.n577 0.003
R10950 S.n264 S.n259 0.003
R10951 S.n1455 S.n1446 0.003
R10952 S.n287 S.n282 0.003
R10953 S.n2281 S.n2269 0.003
R10954 S.n1498 S.n1493 0.003
R10955 S.n1016 S.n1002 0.003
R10956 S.n566 S.n561 0.003
R10957 S.n549 S.n544 0.003
R10958 S.n805 S.n799 0.003
R10959 S.n1808 S.n1802 0.003
R10960 S.n1798 S.n1465 0.003
R10961 S.n2318 S.n2309 0.003
R10962 S.n2304 S.n2291 0.003
R10963 S.n3446 S.n3437 0.003
R10964 S.n3432 S.n3121 0.003
R10965 S.n3965 S.n3956 0.003
R10966 S.n3951 S.n3938 0.003
R10967 S.n4760 S.n4751 0.003
R10968 S.n4746 S.n4733 0.003
R10969 S.n5542 S.n5533 0.003
R10970 S.n5528 S.n5515 0.003
R10971 S.n6302 S.n6293 0.003
R10972 S.n6288 S.n6275 0.003
R10973 S.n7049 S.n7040 0.003
R10974 S.n7035 S.n7022 0.003
R10975 S.n8060 S.n8051 0.003
R10976 S.n8046 S.n7747 0.003
R10977 S.n8772 S.n8763 0.003
R10978 S.n8758 S.n8459 0.003
R10979 S.n9176 S.n9167 0.003
R10980 S.n9162 S.n9149 0.003
R10981 S.n9853 S.n9844 0.003
R10982 S.n9839 S.n9826 0.003
R10983 S.n10511 S.n10502 0.003
R10984 S.n10497 S.n10484 0.003
R10985 S.n11139 S.n11130 0.003
R10986 S.n11125 S.n11112 0.003
R10987 S.n12067 S.n12058 0.003
R10988 S.n12344 S.n12337 0.003
R10989 S.n11870 S.n11862 0.003
R10990 S.n1779 S.n1774 0.003
R10991 S.n2651 S.n2332 0.003
R10992 S.n11852 S.n11851 0.003
R10993 S.n12359 S.n12358 0.003
R10994 S.n12083 S.n12081 0.003
R10995 S.n11168 S.n11167 0.003
R10996 S.n11170 S.n11153 0.003
R10997 S.n10540 S.n10539 0.003
R10998 S.n10542 S.n10525 0.003
R10999 S.n9882 S.n9881 0.003
R11000 S.n9884 S.n9867 0.003
R11001 S.n9205 S.n9204 0.003
R11002 S.n9207 S.n9190 0.003
R11003 S.n8801 S.n8800 0.003
R11004 S.n8803 S.n8786 0.003
R11005 S.n8089 S.n8088 0.003
R11006 S.n8091 S.n8074 0.003
R11007 S.n7078 S.n7077 0.003
R11008 S.n7080 S.n7063 0.003
R11009 S.n6331 S.n6330 0.003
R11010 S.n6333 S.n6316 0.003
R11011 S.n5571 S.n5570 0.003
R11012 S.n5573 S.n5556 0.003
R11013 S.n4789 S.n4788 0.003
R11014 S.n4791 S.n4774 0.003
R11015 S.n3994 S.n3993 0.003
R11016 S.n3996 S.n3979 0.003
R11017 S.n3475 S.n3474 0.003
R11018 S.n3477 S.n3460 0.003
R11019 S.n2650 S.n2649 0.003
R11020 S.n2634 S.n2625 0.003
R11021 S.n3492 S.n3491 0.003
R11022 S.n11837 S.n11836 0.003
R11023 S.n12375 S.n12373 0.003
R11024 S.n12098 S.n12097 0.003
R11025 S.n11417 S.n11415 0.003
R11026 S.n11185 S.n11184 0.003
R11027 S.n10801 S.n10799 0.003
R11028 S.n10557 S.n10556 0.003
R11029 S.n10151 S.n10149 0.003
R11030 S.n9899 S.n9898 0.003
R11031 S.n9475 S.n9473 0.003
R11032 S.n9222 S.n9221 0.003
R11033 S.n8608 S.n8606 0.003
R11034 S.n8818 S.n8817 0.003
R11035 S.n7912 S.n7910 0.003
R11036 S.n8106 S.n8105 0.003
R11037 S.n7359 S.n7357 0.003
R11038 S.n7095 S.n7094 0.003
R11039 S.n6613 S.n6611 0.003
R11040 S.n6348 S.n6347 0.003
R11041 S.n5858 S.n5856 0.003
R11042 S.n5588 S.n5587 0.003
R11043 S.n5077 S.n5075 0.003
R11044 S.n4806 S.n4805 0.003
R11045 S.n4278 S.n4276 0.003
R11046 S.n4011 S.n4010 0.003
R11047 S.n3393 S.n3392 0.003
R11048 S.n11822 S.n11817 0.003
R11049 S.n12391 S.n12386 0.003
R11050 S.n12113 S.n12108 0.003
R11051 S.n11433 S.n11428 0.003
R11052 S.n11200 S.n11195 0.003
R11053 S.n10817 S.n10812 0.003
R11054 S.n10572 S.n10567 0.003
R11055 S.n10167 S.n10162 0.003
R11056 S.n9914 S.n9909 0.003
R11057 S.n9491 S.n9486 0.003
R11058 S.n9237 S.n9232 0.003
R11059 S.n8624 S.n8619 0.003
R11060 S.n8833 S.n8828 0.003
R11061 S.n7928 S.n7923 0.003
R11062 S.n8121 S.n8116 0.003
R11063 S.n7375 S.n7370 0.003
R11064 S.n7110 S.n7105 0.003
R11065 S.n6629 S.n6624 0.003
R11066 S.n6363 S.n6358 0.003
R11067 S.n5874 S.n5869 0.003
R11068 S.n5603 S.n5598 0.003
R11069 S.n5093 S.n5088 0.003
R11070 S.n4821 S.n4816 0.003
R11071 S.n4315 S.n4021 0.003
R11072 S.n4324 S.n4319 0.003
R11073 S.n3413 S.n3404 0.003
R11074 S.n4298 S.n4289 0.003
R11075 S.n5130 S.n4835 0.003
R11076 S.n11807 S.n11806 0.003
R11077 S.n12407 S.n12405 0.003
R11078 S.n12128 S.n12127 0.003
R11079 S.n11449 S.n11447 0.003
R11080 S.n11215 S.n11214 0.003
R11081 S.n10833 S.n10831 0.003
R11082 S.n10587 S.n10586 0.003
R11083 S.n10183 S.n10181 0.003
R11084 S.n9929 S.n9928 0.003
R11085 S.n9507 S.n9505 0.003
R11086 S.n9252 S.n9251 0.003
R11087 S.n8640 S.n8638 0.003
R11088 S.n8848 S.n8847 0.003
R11089 S.n7944 S.n7942 0.003
R11090 S.n8136 S.n8135 0.003
R11091 S.n7391 S.n7389 0.003
R11092 S.n7125 S.n7124 0.003
R11093 S.n6645 S.n6643 0.003
R11094 S.n6378 S.n6377 0.003
R11095 S.n5890 S.n5888 0.003
R11096 S.n5618 S.n5617 0.003
R11097 S.n5129 S.n5128 0.003
R11098 S.n5113 S.n5104 0.003
R11099 S.n5927 S.n5632 0.003
R11100 S.n11792 S.n11791 0.003
R11101 S.n12423 S.n12421 0.003
R11102 S.n12143 S.n12142 0.003
R11103 S.n11465 S.n11463 0.003
R11104 S.n11230 S.n11229 0.003
R11105 S.n10849 S.n10847 0.003
R11106 S.n10602 S.n10601 0.003
R11107 S.n10199 S.n10197 0.003
R11108 S.n9944 S.n9943 0.003
R11109 S.n9523 S.n9521 0.003
R11110 S.n9267 S.n9266 0.003
R11111 S.n8656 S.n8654 0.003
R11112 S.n8863 S.n8862 0.003
R11113 S.n7960 S.n7958 0.003
R11114 S.n8151 S.n8150 0.003
R11115 S.n7407 S.n7405 0.003
R11116 S.n7140 S.n7139 0.003
R11117 S.n6661 S.n6659 0.003
R11118 S.n6393 S.n6392 0.003
R11119 S.n5926 S.n5925 0.003
R11120 S.n5910 S.n5901 0.003
R11121 S.n6698 S.n6407 0.003
R11122 S.n11777 S.n11776 0.003
R11123 S.n12439 S.n12437 0.003
R11124 S.n12158 S.n12157 0.003
R11125 S.n11481 S.n11479 0.003
R11126 S.n11245 S.n11244 0.003
R11127 S.n10865 S.n10863 0.003
R11128 S.n10617 S.n10616 0.003
R11129 S.n10215 S.n10213 0.003
R11130 S.n9959 S.n9958 0.003
R11131 S.n9539 S.n9537 0.003
R11132 S.n9282 S.n9281 0.003
R11133 S.n8672 S.n8670 0.003
R11134 S.n8878 S.n8877 0.003
R11135 S.n7976 S.n7974 0.003
R11136 S.n8166 S.n8165 0.003
R11137 S.n7423 S.n7421 0.003
R11138 S.n7155 S.n7154 0.003
R11139 S.n6697 S.n6696 0.003
R11140 S.n6681 S.n6672 0.003
R11141 S.n7460 S.n7169 0.003
R11142 S.n11762 S.n11761 0.003
R11143 S.n12455 S.n12453 0.003
R11144 S.n12173 S.n12172 0.003
R11145 S.n11497 S.n11495 0.003
R11146 S.n11260 S.n11259 0.003
R11147 S.n10881 S.n10879 0.003
R11148 S.n10632 S.n10631 0.003
R11149 S.n10231 S.n10229 0.003
R11150 S.n9974 S.n9973 0.003
R11151 S.n9555 S.n9553 0.003
R11152 S.n9297 S.n9296 0.003
R11153 S.n8688 S.n8686 0.003
R11154 S.n8893 S.n8892 0.003
R11155 S.n7992 S.n7990 0.003
R11156 S.n8181 S.n8180 0.003
R11157 S.n7459 S.n7458 0.003
R11158 S.n7443 S.n7434 0.003
R11159 S.n8196 S.n8195 0.003
R11160 S.n11747 S.n11746 0.003
R11161 S.n12471 S.n12469 0.003
R11162 S.n12188 S.n12187 0.003
R11163 S.n11513 S.n11511 0.003
R11164 S.n11275 S.n11274 0.003
R11165 S.n10897 S.n10895 0.003
R11166 S.n10647 S.n10646 0.003
R11167 S.n10247 S.n10245 0.003
R11168 S.n9989 S.n9988 0.003
R11169 S.n9571 S.n9569 0.003
R11170 S.n9312 S.n9311 0.003
R11171 S.n8704 S.n8702 0.003
R11172 S.n8908 S.n8907 0.003
R11173 S.n8007 S.n8006 0.003
R11174 S.n8027 S.n8018 0.003
R11175 S.n8923 S.n8922 0.003
R11176 S.n11732 S.n11731 0.003
R11177 S.n12487 S.n12485 0.003
R11178 S.n12203 S.n12202 0.003
R11179 S.n11529 S.n11527 0.003
R11180 S.n11290 S.n11289 0.003
R11181 S.n10913 S.n10911 0.003
R11182 S.n10662 S.n10661 0.003
R11183 S.n10263 S.n10261 0.003
R11184 S.n10004 S.n10003 0.003
R11185 S.n9587 S.n9585 0.003
R11186 S.n9327 S.n9326 0.003
R11187 S.n8719 S.n8718 0.003
R11188 S.n8739 S.n8730 0.003
R11189 S.n9624 S.n9341 0.003
R11190 S.n11717 S.n11716 0.003
R11191 S.n12503 S.n12501 0.003
R11192 S.n12218 S.n12217 0.003
R11193 S.n11545 S.n11543 0.003
R11194 S.n11305 S.n11304 0.003
R11195 S.n10929 S.n10927 0.003
R11196 S.n10677 S.n10676 0.003
R11197 S.n10279 S.n10277 0.003
R11198 S.n10019 S.n10018 0.003
R11199 S.n9623 S.n9622 0.003
R11200 S.n9607 S.n9598 0.003
R11201 S.n10316 S.n10033 0.003
R11202 S.n11702 S.n11701 0.003
R11203 S.n12519 S.n12517 0.003
R11204 S.n12233 S.n12232 0.003
R11205 S.n11561 S.n11559 0.003
R11206 S.n11320 S.n11319 0.003
R11207 S.n10945 S.n10943 0.003
R11208 S.n10692 S.n10691 0.003
R11209 S.n10315 S.n10314 0.003
R11210 S.n10299 S.n10290 0.003
R11211 S.n10982 S.n10706 0.003
R11212 S.n11687 S.n11686 0.003
R11213 S.n12535 S.n12533 0.003
R11214 S.n12248 S.n12247 0.003
R11215 S.n11577 S.n11575 0.003
R11216 S.n11335 S.n11334 0.003
R11217 S.n10981 S.n10980 0.003
R11218 S.n10965 S.n10956 0.003
R11219 S.n11617 S.n11349 0.003
R11220 S.n11672 S.n11671 0.003
R11221 S.n12551 S.n12549 0.003
R11222 S.n12263 S.n12262 0.003
R11223 S.n11616 S.n11615 0.003
R11224 S.n11600 S.n11586 0.003
R11225 S.n12582 S.n12576 0.003
R11226 S.n11657 S.n11652 0.003
R11227 S.n12568 S.n12278 0.003
R11228 S.n980 S.n979 0.003
R11229 S.n2 S.n1 0.003
R11230 S.n10 S.n9 0.003
R11231 S.n18 S.n17 0.003
R11232 S.n27 S.n26 0.003
R11233 S.n36 S.n35 0.003
R11234 S.n45 S.n44 0.003
R11235 S.n59 S.n58 0.003
R11236 S.n11363 S.n11362 0.003
R11237 S.n945 S.n944 0.003
R11238 S.n835 S.n834 0.003
R11239 S.n11360 S.n11359 0.003
R11240 S.n10393 S.n10392 0.003
R11241 S.n9733 S.n9732 0.003
R11242 S.n9061 S.n9060 0.003
R11243 S.n8366 S.n8365 0.003
R11244 S.n7659 S.n7658 0.003
R11245 S.n6929 S.n6928 0.003
R11246 S.n6187 S.n6186 0.003
R11247 S.n5422 S.n5421 0.003
R11248 S.n4645 S.n4644 0.003
R11249 S.n3845 S.n3844 0.003
R11250 S.n3033 S.n3032 0.003
R11251 S.n2197 S.n2196 0.003
R11252 S.n1378 S.n1361 0.003
R11253 S.n12568 S.n12274 0.003
R11254 S.n11923 S.n11922 0.003
R11255 S.t0 S.n11925 0.003
R11256 S.n9363 S.n9362 0.003
R11257 S.n7764 S.n7763 0.003
R11258 S.n6429 S.n6428 0.003
R11259 S.n4857 S.n4856 0.003
R11260 S.n3138 S.n3137 0.003
R11261 S.n1482 S.n1481 0.003
R11262 S.n12038 S.n12037 0.003
R11263 S.n9379 S.n9370 0.003
R11264 S.n8512 S.n8503 0.003
R11265 S.n7816 S.n7807 0.003
R11266 S.n7263 S.n7254 0.003
R11267 S.n6517 S.n6508 0.003
R11268 S.n5762 S.n5753 0.003
R11269 S.n4981 S.n4972 0.003
R11270 S.n4182 S.n4173 0.003
R11271 S.n3298 S.n3289 0.003
R11272 S.n2534 S.n2525 0.003
R11273 S.n1680 S.n1669 0.003
R11274 S.n7780 S.n7771 0.003
R11275 S.n7227 S.n7218 0.003
R11276 S.n6481 S.n6472 0.003
R11277 S.n5726 S.n5717 0.003
R11278 S.n4945 S.n4936 0.003
R11279 S.n4146 S.n4137 0.003
R11280 S.n3262 S.n3253 0.003
R11281 S.n2498 S.n2489 0.003
R11282 S.n1642 S.n1633 0.003
R11283 S.n6445 S.n6436 0.003
R11284 S.n5690 S.n5681 0.003
R11285 S.n4909 S.n4900 0.003
R11286 S.n4110 S.n4101 0.003
R11287 S.n3226 S.n3217 0.003
R11288 S.n2462 S.n2453 0.003
R11289 S.n1606 S.n1597 0.003
R11290 S.n4873 S.n4864 0.003
R11291 S.n4074 S.n4065 0.003
R11292 S.n3190 S.n3181 0.003
R11293 S.n2426 S.n2417 0.003
R11294 S.n1570 S.n1561 0.003
R11295 S.n3154 S.n3145 0.003
R11296 S.n2390 S.n2381 0.003
R11297 S.n1534 S.n1525 0.003
R11298 S.n1498 S.n1489 0.003
R11299 S.n11911 S.n11902 0.003
R11300 S.n1449 S.n1448 0.003
R11301 S.n911 S.n910 0.003
R11302 S.n851 S.n850 0.003
R11303 S.n507 S.n499 0.002
R11304 S.n731 S.n723 0.002
R11305 S.n1310 S.n1289 0.002
R11306 S.n1680 S.n1670 0.002
R11307 S.n2130 S.n2113 0.002
R11308 S.n2534 S.n2526 0.002
R11309 S.n2967 S.n2950 0.002
R11310 S.n3298 S.n3290 0.002
R11311 S.n3779 S.n3762 0.002
R11312 S.n4182 S.n4174 0.002
R11313 S.n4579 S.n4562 0.002
R11314 S.n4981 S.n4973 0.002
R11315 S.n5356 S.n5339 0.002
R11316 S.n5762 S.n5754 0.002
R11317 S.n6121 S.n6104 0.002
R11318 S.n6517 S.n6509 0.002
R11319 S.n6863 S.n6846 0.002
R11320 S.n7263 S.n7255 0.002
R11321 S.n7593 S.n7576 0.002
R11322 S.n7816 S.n7808 0.002
R11323 S.n8300 S.n8283 0.002
R11324 S.n8512 S.n8504 0.002
R11325 S.n8995 S.n8978 0.002
R11326 S.n9379 S.n9371 0.002
R11327 S.n870 S.n857 0.002
R11328 S.n751 S.n739 0.002
R11329 S.n1378 S.n1362 0.002
R11330 S.n1723 S.n1709 0.002
R11331 S.n2197 S.n2170 0.002
R11332 S.n2574 S.n2560 0.002
R11333 S.n3033 S.n3006 0.002
R11334 S.n3338 S.n3324 0.002
R11335 S.n3845 S.n3818 0.002
R11336 S.n4222 S.n4208 0.002
R11337 S.n4645 S.n4618 0.002
R11338 S.n5021 S.n5007 0.002
R11339 S.n5422 S.n5395 0.002
R11340 S.n5802 S.n5788 0.002
R11341 S.n6187 S.n6160 0.002
R11342 S.n6557 S.n6543 0.002
R11343 S.n6929 S.n6902 0.002
R11344 S.n7303 S.n7289 0.002
R11345 S.n7659 S.n7632 0.002
R11346 S.n7856 S.n7842 0.002
R11347 S.n8366 S.n8339 0.002
R11348 S.n8552 S.n8538 0.002
R11349 S.n9061 S.n9034 0.002
R11350 S.n9419 S.n9405 0.002
R11351 S.n9733 S.n9706 0.002
R11352 S.n10095 S.n10081 0.002
R11353 S.n10393 S.n10366 0.002
R11354 S.n10745 S.n10731 0.002
R11355 S.n11382 S.n11371 0.002
R11356 S.n11043 S.n11035 0.002
R11357 S.n10765 S.n10754 0.002
R11358 S.n10413 S.n10405 0.002
R11359 S.n10115 S.n10104 0.002
R11360 S.n9753 S.n9745 0.002
R11361 S.n9439 S.n9428 0.002
R11362 S.n9081 S.n9073 0.002
R11363 S.n8572 S.n8561 0.002
R11364 S.n8386 S.n8378 0.002
R11365 S.n7876 S.n7865 0.002
R11366 S.n7679 S.n7671 0.002
R11367 S.n7323 S.n7312 0.002
R11368 S.n6949 S.n6941 0.002
R11369 S.n6577 S.n6566 0.002
R11370 S.n6207 S.n6199 0.002
R11371 S.n5822 S.n5811 0.002
R11372 S.n5442 S.n5434 0.002
R11373 S.n5041 S.n5030 0.002
R11374 S.n4665 S.n4657 0.002
R11375 S.n4242 S.n4231 0.002
R11376 S.n3865 S.n3857 0.002
R11377 S.n3358 S.n3347 0.002
R11378 S.n3053 S.n3045 0.002
R11379 S.n2594 S.n2583 0.002
R11380 S.n2218 S.n2209 0.002
R11381 S.n1743 S.n1730 0.002
R11382 S.n1406 S.n1390 0.002
R11383 S.n770 S.n759 0.002
R11384 S.n899 S.n877 0.002
R11385 S.n466 S.n455 0.002
R11386 S.n698 S.n690 0.002
R11387 S.n1252 S.n1230 0.002
R11388 S.n1642 S.n1634 0.002
R11389 S.n2069 S.n2052 0.002
R11390 S.n2498 S.n2490 0.002
R11391 S.n2906 S.n2889 0.002
R11392 S.n3262 S.n3254 0.002
R11393 S.n3718 S.n3701 0.002
R11394 S.n4146 S.n4138 0.002
R11395 S.n4518 S.n4501 0.002
R11396 S.n4945 S.n4937 0.002
R11397 S.n5295 S.n5278 0.002
R11398 S.n5726 S.n5718 0.002
R11399 S.n6060 S.n6043 0.002
R11400 S.n6481 S.n6473 0.002
R11401 S.n6802 S.n6785 0.002
R11402 S.n7227 S.n7219 0.002
R11403 S.n7532 S.n7515 0.002
R11404 S.n7780 S.n7772 0.002
R11405 S.n419 S.n411 0.002
R11406 S.n665 S.n657 0.002
R11407 S.n1193 S.n1171 0.002
R11408 S.n1606 S.n1598 0.002
R11409 S.n2008 S.n1991 0.002
R11410 S.n2462 S.n2454 0.002
R11411 S.n2845 S.n2828 0.002
R11412 S.n3226 S.n3218 0.002
R11413 S.n3657 S.n3640 0.002
R11414 S.n4110 S.n4102 0.002
R11415 S.n4457 S.n4440 0.002
R11416 S.n4909 S.n4901 0.002
R11417 S.n5234 S.n5217 0.002
R11418 S.n5690 S.n5682 0.002
R11419 S.n5999 S.n5982 0.002
R11420 S.n6445 S.n6437 0.002
R11421 S.n375 S.n367 0.002
R11422 S.n632 S.n624 0.002
R11423 S.n1134 S.n1112 0.002
R11424 S.n1570 S.n1562 0.002
R11425 S.n1950 S.n1930 0.002
R11426 S.n2426 S.n2418 0.002
R11427 S.n2784 S.n2767 0.002
R11428 S.n3190 S.n3182 0.002
R11429 S.n3596 S.n3579 0.002
R11430 S.n4074 S.n4066 0.002
R11431 S.n4396 S.n4379 0.002
R11432 S.n4873 S.n4865 0.002
R11433 S.n331 S.n323 0.002
R11434 S.n599 S.n591 0.002
R11435 S.n1075 S.n1053 0.002
R11436 S.n1534 S.n1526 0.002
R11437 S.n1886 S.n1869 0.002
R11438 S.n2390 S.n2382 0.002
R11439 S.n2723 S.n2706 0.002
R11440 S.n3154 S.n3146 0.002
R11441 S.n287 S.n279 0.002
R11442 S.n566 S.n558 0.002
R11443 S.n1016 S.n994 0.002
R11444 S.n1498 S.n1490 0.002
R11445 S.n11870 S.n11859 0.002
R11446 S.n12344 S.n12334 0.002
R11447 S.n12067 S.n12055 0.002
R11448 S.n11125 S.n11109 0.002
R11449 S.n11139 S.n11127 0.002
R11450 S.n10497 S.n10481 0.002
R11451 S.n10511 S.n10499 0.002
R11452 S.n9839 S.n9823 0.002
R11453 S.n9853 S.n9841 0.002
R11454 S.n9162 S.n9146 0.002
R11455 S.n9176 S.n9164 0.002
R11456 S.n8758 S.n8456 0.002
R11457 S.n8772 S.n8760 0.002
R11458 S.n8046 S.n7744 0.002
R11459 S.n8060 S.n8048 0.002
R11460 S.n7035 S.n7019 0.002
R11461 S.n7049 S.n7037 0.002
R11462 S.n6288 S.n6272 0.002
R11463 S.n6302 S.n6290 0.002
R11464 S.n5528 S.n5512 0.002
R11465 S.n5542 S.n5530 0.002
R11466 S.n4746 S.n4730 0.002
R11467 S.n4760 S.n4748 0.002
R11468 S.n3951 S.n3935 0.002
R11469 S.n3965 S.n3953 0.002
R11470 S.n3432 S.n3118 0.002
R11471 S.n3446 S.n3434 0.002
R11472 S.n2304 S.n2288 0.002
R11473 S.n2318 S.n2306 0.002
R11474 S.n1798 S.n1462 0.002
R11475 S.n1808 S.n1799 0.002
R11476 S.n11852 S.n11844 0.002
R11477 S.n12359 S.n12351 0.002
R11478 S.n12083 S.n12074 0.002
R11479 S.n11168 S.n11154 0.002
R11480 S.n11170 S.n11146 0.002
R11481 S.n10540 S.n10526 0.002
R11482 S.n10542 S.n10518 0.002
R11483 S.n9882 S.n9868 0.002
R11484 S.n9884 S.n9860 0.002
R11485 S.n9205 S.n9191 0.002
R11486 S.n9207 S.n9183 0.002
R11487 S.n8801 S.n8787 0.002
R11488 S.n8803 S.n8779 0.002
R11489 S.n8089 S.n8075 0.002
R11490 S.n8091 S.n8067 0.002
R11491 S.n7078 S.n7064 0.002
R11492 S.n7080 S.n7056 0.002
R11493 S.n6331 S.n6317 0.002
R11494 S.n6333 S.n6309 0.002
R11495 S.n5571 S.n5557 0.002
R11496 S.n5573 S.n5549 0.002
R11497 S.n4789 S.n4775 0.002
R11498 S.n4791 S.n4767 0.002
R11499 S.n3994 S.n3980 0.002
R11500 S.n3996 S.n3972 0.002
R11501 S.n3475 S.n3461 0.002
R11502 S.n3477 S.n3453 0.002
R11503 S.n2650 S.n2333 0.002
R11504 S.n2651 S.n2325 0.002
R11505 S.n1779 S.n1771 0.002
R11506 S.n11837 S.n11829 0.002
R11507 S.n12375 S.n12366 0.002
R11508 S.n12098 S.n12090 0.002
R11509 S.n11417 S.n11408 0.002
R11510 S.n11185 S.n11177 0.002
R11511 S.n10801 S.n10792 0.002
R11512 S.n10557 S.n10549 0.002
R11513 S.n10151 S.n10142 0.002
R11514 S.n9899 S.n9891 0.002
R11515 S.n9475 S.n9466 0.002
R11516 S.n9222 S.n9214 0.002
R11517 S.n8608 S.n8599 0.002
R11518 S.n8818 S.n8810 0.002
R11519 S.n7912 S.n7903 0.002
R11520 S.n8106 S.n8098 0.002
R11521 S.n7359 S.n7350 0.002
R11522 S.n7095 S.n7087 0.002
R11523 S.n6613 S.n6604 0.002
R11524 S.n6348 S.n6340 0.002
R11525 S.n5858 S.n5849 0.002
R11526 S.n5588 S.n5580 0.002
R11527 S.n5077 S.n5068 0.002
R11528 S.n4806 S.n4798 0.002
R11529 S.n4278 S.n4269 0.002
R11530 S.n4011 S.n4003 0.002
R11531 S.n3393 S.n3385 0.002
R11532 S.n3492 S.n3484 0.002
R11533 S.n2634 S.n2622 0.002
R11534 S.n11822 S.n11814 0.002
R11535 S.n12391 S.n12383 0.002
R11536 S.n12113 S.n12105 0.002
R11537 S.n11433 S.n11425 0.002
R11538 S.n11200 S.n11192 0.002
R11539 S.n10817 S.n10809 0.002
R11540 S.n10572 S.n10564 0.002
R11541 S.n10167 S.n10159 0.002
R11542 S.n9914 S.n9906 0.002
R11543 S.n9491 S.n9483 0.002
R11544 S.n9237 S.n9229 0.002
R11545 S.n8624 S.n8616 0.002
R11546 S.n8833 S.n8825 0.002
R11547 S.n7928 S.n7920 0.002
R11548 S.n8121 S.n8113 0.002
R11549 S.n7375 S.n7367 0.002
R11550 S.n7110 S.n7102 0.002
R11551 S.n6629 S.n6621 0.002
R11552 S.n6363 S.n6355 0.002
R11553 S.n5874 S.n5866 0.002
R11554 S.n5603 S.n5595 0.002
R11555 S.n5093 S.n5085 0.002
R11556 S.n4821 S.n4813 0.002
R11557 S.n4315 S.n4018 0.002
R11558 S.n4324 S.n4316 0.002
R11559 S.n3413 S.n3401 0.002
R11560 S.n11807 S.n11799 0.002
R11561 S.n12407 S.n12398 0.002
R11562 S.n12128 S.n12120 0.002
R11563 S.n11449 S.n11440 0.002
R11564 S.n11215 S.n11207 0.002
R11565 S.n10833 S.n10824 0.002
R11566 S.n10587 S.n10579 0.002
R11567 S.n10183 S.n10174 0.002
R11568 S.n9929 S.n9921 0.002
R11569 S.n9507 S.n9498 0.002
R11570 S.n9252 S.n9244 0.002
R11571 S.n8640 S.n8631 0.002
R11572 S.n8848 S.n8840 0.002
R11573 S.n7944 S.n7935 0.002
R11574 S.n8136 S.n8128 0.002
R11575 S.n7391 S.n7382 0.002
R11576 S.n7125 S.n7117 0.002
R11577 S.n6645 S.n6636 0.002
R11578 S.n6378 S.n6370 0.002
R11579 S.n5890 S.n5881 0.002
R11580 S.n5618 S.n5610 0.002
R11581 S.n5129 S.n4836 0.002
R11582 S.n5130 S.n4828 0.002
R11583 S.n4298 S.n4286 0.002
R11584 S.n11792 S.n11784 0.002
R11585 S.n12423 S.n12414 0.002
R11586 S.n12143 S.n12135 0.002
R11587 S.n11465 S.n11456 0.002
R11588 S.n11230 S.n11222 0.002
R11589 S.n10849 S.n10840 0.002
R11590 S.n10602 S.n10594 0.002
R11591 S.n10199 S.n10190 0.002
R11592 S.n9944 S.n9936 0.002
R11593 S.n9523 S.n9514 0.002
R11594 S.n9267 S.n9259 0.002
R11595 S.n8656 S.n8647 0.002
R11596 S.n8863 S.n8855 0.002
R11597 S.n7960 S.n7951 0.002
R11598 S.n8151 S.n8143 0.002
R11599 S.n7407 S.n7398 0.002
R11600 S.n7140 S.n7132 0.002
R11601 S.n6661 S.n6652 0.002
R11602 S.n6393 S.n6385 0.002
R11603 S.n5926 S.n5633 0.002
R11604 S.n5927 S.n5625 0.002
R11605 S.n5113 S.n5101 0.002
R11606 S.n11777 S.n11769 0.002
R11607 S.n12439 S.n12430 0.002
R11608 S.n12158 S.n12150 0.002
R11609 S.n11481 S.n11472 0.002
R11610 S.n11245 S.n11237 0.002
R11611 S.n10865 S.n10856 0.002
R11612 S.n10617 S.n10609 0.002
R11613 S.n10215 S.n10206 0.002
R11614 S.n9959 S.n9951 0.002
R11615 S.n9539 S.n9530 0.002
R11616 S.n9282 S.n9274 0.002
R11617 S.n8672 S.n8663 0.002
R11618 S.n8878 S.n8870 0.002
R11619 S.n7976 S.n7967 0.002
R11620 S.n8166 S.n8158 0.002
R11621 S.n7423 S.n7414 0.002
R11622 S.n7155 S.n7147 0.002
R11623 S.n6697 S.n6408 0.002
R11624 S.n6698 S.n6400 0.002
R11625 S.n5910 S.n5898 0.002
R11626 S.n11762 S.n11754 0.002
R11627 S.n12455 S.n12446 0.002
R11628 S.n12173 S.n12165 0.002
R11629 S.n11497 S.n11488 0.002
R11630 S.n11260 S.n11252 0.002
R11631 S.n10881 S.n10872 0.002
R11632 S.n10632 S.n10624 0.002
R11633 S.n10231 S.n10222 0.002
R11634 S.n9974 S.n9966 0.002
R11635 S.n9555 S.n9546 0.002
R11636 S.n9297 S.n9289 0.002
R11637 S.n8688 S.n8679 0.002
R11638 S.n8893 S.n8885 0.002
R11639 S.n7992 S.n7983 0.002
R11640 S.n8181 S.n8173 0.002
R11641 S.n7459 S.n7170 0.002
R11642 S.n7460 S.n7162 0.002
R11643 S.n6681 S.n6669 0.002
R11644 S.n11747 S.n11739 0.002
R11645 S.n12471 S.n12462 0.002
R11646 S.n12188 S.n12180 0.002
R11647 S.n11513 S.n11504 0.002
R11648 S.n11275 S.n11267 0.002
R11649 S.n10897 S.n10888 0.002
R11650 S.n10647 S.n10639 0.002
R11651 S.n10247 S.n10238 0.002
R11652 S.n9989 S.n9981 0.002
R11653 S.n9571 S.n9562 0.002
R11654 S.n9312 S.n9304 0.002
R11655 S.n8704 S.n8695 0.002
R11656 S.n8908 S.n8900 0.002
R11657 S.n8007 S.n7999 0.002
R11658 S.n8196 S.n8188 0.002
R11659 S.n7443 S.n7431 0.002
R11660 S.n11732 S.n11724 0.002
R11661 S.n12487 S.n12478 0.002
R11662 S.n12203 S.n12195 0.002
R11663 S.n11529 S.n11520 0.002
R11664 S.n11290 S.n11282 0.002
R11665 S.n10913 S.n10904 0.002
R11666 S.n10662 S.n10654 0.002
R11667 S.n10263 S.n10254 0.002
R11668 S.n10004 S.n9996 0.002
R11669 S.n9587 S.n9578 0.002
R11670 S.n9327 S.n9319 0.002
R11671 S.n8719 S.n8711 0.002
R11672 S.n8923 S.n8915 0.002
R11673 S.n8027 S.n8015 0.002
R11674 S.n11717 S.n11709 0.002
R11675 S.n12503 S.n12494 0.002
R11676 S.n12218 S.n12210 0.002
R11677 S.n11545 S.n11536 0.002
R11678 S.n11305 S.n11297 0.002
R11679 S.n10929 S.n10920 0.002
R11680 S.n10677 S.n10669 0.002
R11681 S.n10279 S.n10270 0.002
R11682 S.n10019 S.n10011 0.002
R11683 S.n9623 S.n9342 0.002
R11684 S.n9624 S.n9334 0.002
R11685 S.n8739 S.n8727 0.002
R11686 S.n11702 S.n11694 0.002
R11687 S.n12519 S.n12510 0.002
R11688 S.n12233 S.n12225 0.002
R11689 S.n11561 S.n11552 0.002
R11690 S.n11320 S.n11312 0.002
R11691 S.n10945 S.n10936 0.002
R11692 S.n10692 S.n10684 0.002
R11693 S.n10315 S.n10034 0.002
R11694 S.n10316 S.n10026 0.002
R11695 S.n9607 S.n9595 0.002
R11696 S.n11687 S.n11679 0.002
R11697 S.n12535 S.n12526 0.002
R11698 S.n12248 S.n12240 0.002
R11699 S.n11577 S.n11568 0.002
R11700 S.n11335 S.n11327 0.002
R11701 S.n10981 S.n10707 0.002
R11702 S.n10982 S.n10699 0.002
R11703 S.n10299 S.n10287 0.002
R11704 S.n11672 S.n11664 0.002
R11705 S.n12551 S.n12542 0.002
R11706 S.n12263 S.n12255 0.002
R11707 S.n11616 S.n11350 0.002
R11708 S.n11617 S.n11342 0.002
R11709 S.n10965 S.n10953 0.002
R11710 S.n12568 S.n12275 0.002
R11711 S.n11657 S.n11649 0.002
R11712 S.n11600 S.n11590 0.002
R11713 S.n12582 S.n12573 0.002
R11714 S.n12327 S.n12312 0.002
R11715 S.n11911 S.n11903 0.002
R11716 S.n950 S.n935 0.002
R11717 S.n9816 S.n9801 0.002
R11718 S.n11102 S.n11083 0.002
R11719 S.n8449 S.n8434 0.002
R11720 S.n7012 S.n6997 0.002
R11721 S.n5505 S.n5490 0.002
R11722 S.n3928 S.n3913 0.002
R11723 S.n2281 S.n2266 0.002
R11724 S.n12047 S.n12039 0.002
R11725 S.n2694 S.n2693 0.002
R11726 S.n3535 S.n3534 0.002
R11727 S.n4367 S.n4366 0.002
R11728 S.n5173 S.n5172 0.002
R11729 S.n5970 S.n5969 0.002
R11730 S.n6741 S.n6740 0.002
R11731 S.n7503 S.n7502 0.002
R11732 S.n8239 S.n8238 0.002
R11733 S.n8966 S.n8965 0.002
R11734 S.n9667 S.n9666 0.002
R11735 S.n10359 S.n10358 0.002
R11736 S.n11023 S.n11022 0.002
R11737 S.t7 S.n197 0.002
R11738 S.n1808 S.n1807 0.002
R11739 S.n934 S.n933 0.002
R11740 S.n11890 S.n11889 0.002
R11741 S.n10468 S.n10467 0.002
R11742 S.n9133 S.n9132 0.002
R11743 S.n7731 S.n7730 0.002
R11744 S.n6259 S.n6258 0.002
R11745 S.n4717 S.n4716 0.002
R11746 S.n3105 S.n3104 0.002
R11747 S.n1431 S.n1414 0.002
R11748 S.n1282 S.n1269 0.002
R11749 S.n2130 S.n2129 0.002
R11750 S.n2534 S.n2533 0.002
R11751 S.n2967 S.n2966 0.002
R11752 S.n3298 S.n3297 0.002
R11753 S.n3779 S.n3778 0.002
R11754 S.n4182 S.n4181 0.002
R11755 S.n4579 S.n4578 0.002
R11756 S.n4981 S.n4980 0.002
R11757 S.n5356 S.n5355 0.002
R11758 S.n5762 S.n5761 0.002
R11759 S.n6121 S.n6120 0.002
R11760 S.n6517 S.n6516 0.002
R11761 S.n6863 S.n6862 0.002
R11762 S.n7263 S.n7262 0.002
R11763 S.n7593 S.n7592 0.002
R11764 S.n7816 S.n7815 0.002
R11765 S.n8300 S.n8299 0.002
R11766 S.n8512 S.n8511 0.002
R11767 S.n8995 S.n8994 0.002
R11768 S.n9379 S.n9378 0.002
R11769 S.n1223 S.n1210 0.002
R11770 S.n1642 S.n1641 0.002
R11771 S.n2069 S.n2068 0.002
R11772 S.n2498 S.n2497 0.002
R11773 S.n2906 S.n2905 0.002
R11774 S.n3262 S.n3261 0.002
R11775 S.n3718 S.n3717 0.002
R11776 S.n4146 S.n4145 0.002
R11777 S.n4518 S.n4517 0.002
R11778 S.n4945 S.n4944 0.002
R11779 S.n5295 S.n5294 0.002
R11780 S.n5726 S.n5725 0.002
R11781 S.n6060 S.n6059 0.002
R11782 S.n6481 S.n6480 0.002
R11783 S.n6802 S.n6801 0.002
R11784 S.n7227 S.n7226 0.002
R11785 S.n7532 S.n7531 0.002
R11786 S.n7780 S.n7779 0.002
R11787 S.n1164 S.n1151 0.002
R11788 S.n1606 S.n1605 0.002
R11789 S.n2008 S.n2007 0.002
R11790 S.n2462 S.n2461 0.002
R11791 S.n2845 S.n2844 0.002
R11792 S.n3226 S.n3225 0.002
R11793 S.n3657 S.n3656 0.002
R11794 S.n4110 S.n4109 0.002
R11795 S.n4457 S.n4456 0.002
R11796 S.n4909 S.n4908 0.002
R11797 S.n5234 S.n5233 0.002
R11798 S.n5690 S.n5689 0.002
R11799 S.n5999 S.n5998 0.002
R11800 S.n6445 S.n6444 0.002
R11801 S.n1105 S.n1092 0.002
R11802 S.n1570 S.n1569 0.002
R11803 S.n1950 S.n1949 0.002
R11804 S.n2426 S.n2425 0.002
R11805 S.n2784 S.n2783 0.002
R11806 S.n3190 S.n3189 0.002
R11807 S.n3596 S.n3595 0.002
R11808 S.n4074 S.n4073 0.002
R11809 S.n4396 S.n4395 0.002
R11810 S.n4873 S.n4872 0.002
R11811 S.n1046 S.n1033 0.002
R11812 S.n1534 S.n1533 0.002
R11813 S.n1886 S.n1885 0.002
R11814 S.n2390 S.n2389 0.002
R11815 S.n2723 S.n2722 0.002
R11816 S.n3154 S.n3153 0.002
R11817 S.n1498 S.n1497 0.002
R11818 S.n2651 S.n2326 0.002
R11819 S.n3492 S.n3485 0.002
R11820 S.n3413 S.n3412 0.002
R11821 S.n4324 S.n4323 0.002
R11822 S.n4315 S.n4314 0.002
R11823 S.n4821 S.n4820 0.002
R11824 S.n5093 S.n5092 0.002
R11825 S.n5603 S.n5602 0.002
R11826 S.n5874 S.n5873 0.002
R11827 S.n6363 S.n6362 0.002
R11828 S.n6629 S.n6628 0.002
R11829 S.n7110 S.n7109 0.002
R11830 S.n7375 S.n7374 0.002
R11831 S.n8121 S.n8120 0.002
R11832 S.n7928 S.n7927 0.002
R11833 S.n8833 S.n8832 0.002
R11834 S.n8624 S.n8623 0.002
R11835 S.n9237 S.n9236 0.002
R11836 S.n9491 S.n9490 0.002
R11837 S.n9914 S.n9913 0.002
R11838 S.n10167 S.n10166 0.002
R11839 S.n10572 S.n10571 0.002
R11840 S.n10817 S.n10816 0.002
R11841 S.n11200 S.n11199 0.002
R11842 S.n11433 S.n11432 0.002
R11843 S.n12113 S.n12112 0.002
R11844 S.n12391 S.n12390 0.002
R11845 S.n11822 S.n11821 0.002
R11846 S.n5130 S.n4829 0.002
R11847 S.n5927 S.n5626 0.002
R11848 S.n6698 S.n6401 0.002
R11849 S.n7460 S.n7163 0.002
R11850 S.n8196 S.n8189 0.002
R11851 S.n8923 S.n8916 0.002
R11852 S.n9624 S.n9335 0.002
R11853 S.n10316 S.n10027 0.002
R11854 S.n10982 S.n10700 0.002
R11855 S.n11617 S.n11343 0.002
R11856 S.n12568 S.n12567 0.002
R11857 S.n11657 S.n11656 0.002
R11858 S.n12327 S.n12326 0.002
R11859 S.n11911 S.n11910 0.002
R11860 S.n9800 S.n9799 0.002
R11861 S.n8433 S.n8432 0.002
R11862 S.n6996 S.n6995 0.002
R11863 S.n5489 S.n5488 0.002
R11864 S.n3912 S.n3911 0.002
R11865 S.n2265 S.n2264 0.002
R11866 S.n78 S.n75 0.002
R11867 S.n12303 S.n12292 0.002
R11868 S.n12023 S.n12008 0.002
R11869 S.n11401 S.n11390 0.002
R11870 S.n11075 S.n11060 0.002
R11871 S.n10784 S.n10773 0.002
R11872 S.n10445 S.n10430 0.002
R11873 S.n10134 S.n10123 0.002
R11874 S.n9785 S.n9770 0.002
R11875 S.n9458 S.n9447 0.002
R11876 S.n9113 S.n9098 0.002
R11877 S.n8591 S.n8580 0.002
R11878 S.n8418 S.n8403 0.002
R11879 S.n7895 S.n7884 0.002
R11880 S.n7711 S.n7696 0.002
R11881 S.n7342 S.n7331 0.002
R11882 S.n6981 S.n6966 0.002
R11883 S.n6596 S.n6585 0.002
R11884 S.n6239 S.n6224 0.002
R11885 S.n5841 S.n5830 0.002
R11886 S.n5474 S.n5459 0.002
R11887 S.n5060 S.n5049 0.002
R11888 S.n4697 S.n4682 0.002
R11889 S.n4261 S.n4250 0.002
R11890 S.n3897 S.n3882 0.002
R11891 S.n3377 S.n3366 0.002
R11892 S.n3085 S.n3070 0.002
R11893 S.n2613 S.n2602 0.002
R11894 S.n2250 S.n2235 0.002
R11895 S.n1762 S.n1751 0.002
R11896 S.n787 S.n786 0.002
R11897 S.n8495 S.n8484 0.002
R11898 S.n8271 S.n8256 0.002
R11899 S.n7799 S.n7788 0.002
R11900 S.n7564 S.n7549 0.002
R11901 S.n7246 S.n7235 0.002
R11902 S.n6834 S.n6819 0.002
R11903 S.n6500 S.n6489 0.002
R11904 S.n6092 S.n6077 0.002
R11905 S.n5745 S.n5734 0.002
R11906 S.n5327 S.n5312 0.002
R11907 S.n4964 S.n4953 0.002
R11908 S.n4550 S.n4535 0.002
R11909 S.n4165 S.n4154 0.002
R11910 S.n3750 S.n3735 0.002
R11911 S.n3281 S.n3270 0.002
R11912 S.n2938 S.n2923 0.002
R11913 S.n2517 S.n2506 0.002
R11914 S.n2101 S.n2086 0.002
R11915 S.n1661 S.n1650 0.002
R11916 S.n1310 S.n1309 0.002
R11917 S.n731 S.n730 0.002
R11918 S.n714 S.n713 0.002
R11919 S.n7210 S.n7199 0.002
R11920 S.n6773 S.n6758 0.002
R11921 S.n6464 S.n6453 0.002
R11922 S.n6031 S.n6016 0.002
R11923 S.n5709 S.n5698 0.002
R11924 S.n5266 S.n5251 0.002
R11925 S.n4928 S.n4917 0.002
R11926 S.n4489 S.n4474 0.002
R11927 S.n4129 S.n4118 0.002
R11928 S.n3689 S.n3674 0.002
R11929 S.n3245 S.n3234 0.002
R11930 S.n2877 S.n2862 0.002
R11931 S.n2481 S.n2470 0.002
R11932 S.n2040 S.n2025 0.002
R11933 S.n1625 S.n1614 0.002
R11934 S.n1252 S.n1251 0.002
R11935 S.n698 S.n697 0.002
R11936 S.n681 S.n680 0.002
R11937 S.n5673 S.n5662 0.002
R11938 S.n5205 S.n5190 0.002
R11939 S.n4892 S.n4881 0.002
R11940 S.n4428 S.n4413 0.002
R11941 S.n4093 S.n4082 0.002
R11942 S.n3628 S.n3613 0.002
R11943 S.n3209 S.n3198 0.002
R11944 S.n2816 S.n2801 0.002
R11945 S.n2445 S.n2434 0.002
R11946 S.n1979 S.n1964 0.002
R11947 S.n1589 S.n1578 0.002
R11948 S.n1193 S.n1192 0.002
R11949 S.n665 S.n664 0.002
R11950 S.n648 S.n647 0.002
R11951 S.n4057 S.n4046 0.002
R11952 S.n3567 S.n3552 0.002
R11953 S.n3173 S.n3162 0.002
R11954 S.n2755 S.n2740 0.002
R11955 S.n2409 S.n2398 0.002
R11956 S.n1918 S.n1903 0.002
R11957 S.n1553 S.n1542 0.002
R11958 S.n1134 S.n1133 0.002
R11959 S.n632 S.n631 0.002
R11960 S.n615 S.n614 0.002
R11961 S.n2373 S.n2362 0.002
R11962 S.n1857 S.n1842 0.002
R11963 S.n1517 S.n1506 0.002
R11964 S.n1075 S.n1074 0.002
R11965 S.n599 S.n598 0.002
R11966 S.n582 S.n581 0.002
R11967 S.n1016 S.n1015 0.002
R11968 S.n566 S.n565 0.002
R11969 S.n549 S.n548 0.002
R11970 S.n11852 S.n11845 0.002
R11971 S.n12359 S.n12352 0.002
R11972 S.n12083 S.n12075 0.002
R11973 S.n11168 S.n11155 0.002
R11974 S.n11170 S.n11147 0.002
R11975 S.n10540 S.n10527 0.002
R11976 S.n10542 S.n10519 0.002
R11977 S.n9882 S.n9869 0.002
R11978 S.n9884 S.n9861 0.002
R11979 S.n9205 S.n9192 0.002
R11980 S.n9207 S.n9184 0.002
R11981 S.n8801 S.n8788 0.002
R11982 S.n8803 S.n8780 0.002
R11983 S.n8089 S.n8076 0.002
R11984 S.n8091 S.n8068 0.002
R11985 S.n7078 S.n7065 0.002
R11986 S.n7080 S.n7057 0.002
R11987 S.n6331 S.n6318 0.002
R11988 S.n6333 S.n6310 0.002
R11989 S.n5571 S.n5558 0.002
R11990 S.n5573 S.n5550 0.002
R11991 S.n4789 S.n4776 0.002
R11992 S.n4791 S.n4768 0.002
R11993 S.n3994 S.n3981 0.002
R11994 S.n3996 S.n3973 0.002
R11995 S.n3475 S.n3462 0.002
R11996 S.n3477 S.n3454 0.002
R11997 S.n2650 S.n2334 0.002
R11998 S.n1779 S.n1778 0.002
R11999 S.n11837 S.n11830 0.002
R12000 S.n12375 S.n12367 0.002
R12001 S.n12098 S.n12091 0.002
R12002 S.n11417 S.n11409 0.002
R12003 S.n11185 S.n11178 0.002
R12004 S.n10801 S.n10793 0.002
R12005 S.n10557 S.n10550 0.002
R12006 S.n10151 S.n10143 0.002
R12007 S.n9899 S.n9892 0.002
R12008 S.n9475 S.n9467 0.002
R12009 S.n9222 S.n9215 0.002
R12010 S.n8608 S.n8600 0.002
R12011 S.n8818 S.n8811 0.002
R12012 S.n7912 S.n7904 0.002
R12013 S.n8106 S.n8099 0.002
R12014 S.n7359 S.n7351 0.002
R12015 S.n7095 S.n7088 0.002
R12016 S.n6613 S.n6605 0.002
R12017 S.n6348 S.n6341 0.002
R12018 S.n5858 S.n5850 0.002
R12019 S.n5588 S.n5581 0.002
R12020 S.n5077 S.n5069 0.002
R12021 S.n4806 S.n4799 0.002
R12022 S.n4278 S.n4270 0.002
R12023 S.n4011 S.n4004 0.002
R12024 S.n3393 S.n3386 0.002
R12025 S.n2634 S.n2633 0.002
R12026 S.n11807 S.n11800 0.002
R12027 S.n12407 S.n12399 0.002
R12028 S.n12128 S.n12121 0.002
R12029 S.n11449 S.n11441 0.002
R12030 S.n11215 S.n11208 0.002
R12031 S.n10833 S.n10825 0.002
R12032 S.n10587 S.n10580 0.002
R12033 S.n10183 S.n10175 0.002
R12034 S.n9929 S.n9922 0.002
R12035 S.n9507 S.n9499 0.002
R12036 S.n9252 S.n9245 0.002
R12037 S.n8640 S.n8632 0.002
R12038 S.n8848 S.n8841 0.002
R12039 S.n7944 S.n7936 0.002
R12040 S.n8136 S.n8129 0.002
R12041 S.n7391 S.n7383 0.002
R12042 S.n7125 S.n7118 0.002
R12043 S.n6645 S.n6637 0.002
R12044 S.n6378 S.n6371 0.002
R12045 S.n5890 S.n5882 0.002
R12046 S.n5618 S.n5611 0.002
R12047 S.n5129 S.n4837 0.002
R12048 S.n4298 S.n4297 0.002
R12049 S.n11792 S.n11785 0.002
R12050 S.n12423 S.n12415 0.002
R12051 S.n12143 S.n12136 0.002
R12052 S.n11465 S.n11457 0.002
R12053 S.n11230 S.n11223 0.002
R12054 S.n10849 S.n10841 0.002
R12055 S.n10602 S.n10595 0.002
R12056 S.n10199 S.n10191 0.002
R12057 S.n9944 S.n9937 0.002
R12058 S.n9523 S.n9515 0.002
R12059 S.n9267 S.n9260 0.002
R12060 S.n8656 S.n8648 0.002
R12061 S.n8863 S.n8856 0.002
R12062 S.n7960 S.n7952 0.002
R12063 S.n8151 S.n8144 0.002
R12064 S.n7407 S.n7399 0.002
R12065 S.n7140 S.n7133 0.002
R12066 S.n6661 S.n6653 0.002
R12067 S.n6393 S.n6386 0.002
R12068 S.n5926 S.n5634 0.002
R12069 S.n5113 S.n5112 0.002
R12070 S.n11777 S.n11770 0.002
R12071 S.n12439 S.n12431 0.002
R12072 S.n12158 S.n12151 0.002
R12073 S.n11481 S.n11473 0.002
R12074 S.n11245 S.n11238 0.002
R12075 S.n10865 S.n10857 0.002
R12076 S.n10617 S.n10610 0.002
R12077 S.n10215 S.n10207 0.002
R12078 S.n9959 S.n9952 0.002
R12079 S.n9539 S.n9531 0.002
R12080 S.n9282 S.n9275 0.002
R12081 S.n8672 S.n8664 0.002
R12082 S.n8878 S.n8871 0.002
R12083 S.n7976 S.n7968 0.002
R12084 S.n8166 S.n8159 0.002
R12085 S.n7423 S.n7415 0.002
R12086 S.n7155 S.n7148 0.002
R12087 S.n6697 S.n6409 0.002
R12088 S.n5910 S.n5909 0.002
R12089 S.n11762 S.n11755 0.002
R12090 S.n12455 S.n12447 0.002
R12091 S.n12173 S.n12166 0.002
R12092 S.n11497 S.n11489 0.002
R12093 S.n11260 S.n11253 0.002
R12094 S.n10881 S.n10873 0.002
R12095 S.n10632 S.n10625 0.002
R12096 S.n10231 S.n10223 0.002
R12097 S.n9974 S.n9967 0.002
R12098 S.n9555 S.n9547 0.002
R12099 S.n9297 S.n9290 0.002
R12100 S.n8688 S.n8680 0.002
R12101 S.n8893 S.n8886 0.002
R12102 S.n7992 S.n7984 0.002
R12103 S.n8181 S.n8174 0.002
R12104 S.n7459 S.n7171 0.002
R12105 S.n6681 S.n6680 0.002
R12106 S.n11747 S.n11740 0.002
R12107 S.n12471 S.n12463 0.002
R12108 S.n12188 S.n12181 0.002
R12109 S.n11513 S.n11505 0.002
R12110 S.n11275 S.n11268 0.002
R12111 S.n10897 S.n10889 0.002
R12112 S.n10647 S.n10640 0.002
R12113 S.n10247 S.n10239 0.002
R12114 S.n9989 S.n9982 0.002
R12115 S.n9571 S.n9563 0.002
R12116 S.n9312 S.n9305 0.002
R12117 S.n8704 S.n8696 0.002
R12118 S.n8908 S.n8901 0.002
R12119 S.n8007 S.n8000 0.002
R12120 S.n7443 S.n7442 0.002
R12121 S.n11732 S.n11725 0.002
R12122 S.n12487 S.n12479 0.002
R12123 S.n12203 S.n12196 0.002
R12124 S.n11529 S.n11521 0.002
R12125 S.n11290 S.n11283 0.002
R12126 S.n10913 S.n10905 0.002
R12127 S.n10662 S.n10655 0.002
R12128 S.n10263 S.n10255 0.002
R12129 S.n10004 S.n9997 0.002
R12130 S.n9587 S.n9579 0.002
R12131 S.n9327 S.n9320 0.002
R12132 S.n8719 S.n8712 0.002
R12133 S.n8027 S.n8026 0.002
R12134 S.n11717 S.n11710 0.002
R12135 S.n12503 S.n12495 0.002
R12136 S.n12218 S.n12211 0.002
R12137 S.n11545 S.n11537 0.002
R12138 S.n11305 S.n11298 0.002
R12139 S.n10929 S.n10921 0.002
R12140 S.n10677 S.n10670 0.002
R12141 S.n10279 S.n10271 0.002
R12142 S.n10019 S.n10012 0.002
R12143 S.n9623 S.n9343 0.002
R12144 S.n8739 S.n8738 0.002
R12145 S.n11702 S.n11695 0.002
R12146 S.n12519 S.n12511 0.002
R12147 S.n12233 S.n12226 0.002
R12148 S.n11561 S.n11553 0.002
R12149 S.n11320 S.n11313 0.002
R12150 S.n10945 S.n10937 0.002
R12151 S.n10692 S.n10685 0.002
R12152 S.n10315 S.n10035 0.002
R12153 S.n9607 S.n9606 0.002
R12154 S.n11687 S.n11680 0.002
R12155 S.n12535 S.n12527 0.002
R12156 S.n12248 S.n12241 0.002
R12157 S.n11577 S.n11569 0.002
R12158 S.n11335 S.n11328 0.002
R12159 S.n10981 S.n10708 0.002
R12160 S.n10299 S.n10298 0.002
R12161 S.n11672 S.n11665 0.002
R12162 S.n12551 S.n12543 0.002
R12163 S.n12263 S.n12256 0.002
R12164 S.n11616 S.n11351 0.002
R12165 S.n10965 S.n10964 0.002
R12166 S.n12582 S.n12581 0.002
R12167 S.n870 S.n856 0.002
R12168 S.n899 S.n896 0.002
R12169 S.n11600 S.n11596 0.002
R12170 S.n11891 S.n11880 0.002
R12171 S.n9139 S.n9122 0.002
R12172 S.n7737 S.n7720 0.002
R12173 S.n6265 S.n6248 0.002
R12174 S.n4723 S.n4706 0.002
R12175 S.n3111 S.n3094 0.002
R12176 S.n1455 S.n1440 0.002
R12177 S.n82 S.n81 0.002
R12178 S.n12047 S.n12046 0.002
R12179 S.n11043 S.n11042 0.002
R12180 S.n10413 S.n10412 0.002
R12181 S.n9753 S.n9752 0.002
R12182 S.n9081 S.n9080 0.002
R12183 S.n8386 S.n8385 0.002
R12184 S.n7679 S.n7678 0.002
R12185 S.n6949 S.n6948 0.002
R12186 S.n6207 S.n6206 0.002
R12187 S.n5442 S.n5441 0.002
R12188 S.n4665 S.n4664 0.002
R12189 S.n3865 S.n3864 0.002
R12190 S.n3053 S.n3052 0.002
R12191 S.n2218 S.n2217 0.002
R12192 S.n2634 S.n2621 0.002
R12193 S.n4278 S.n4277 0.002
R12194 S.n5077 S.n5076 0.002
R12195 S.n5858 S.n5857 0.002
R12196 S.n6613 S.n6612 0.002
R12197 S.n7359 S.n7358 0.002
R12198 S.n7912 S.n7911 0.002
R12199 S.n8608 S.n8607 0.002
R12200 S.n9475 S.n9474 0.002
R12201 S.n10151 S.n10150 0.002
R12202 S.n10801 S.n10800 0.002
R12203 S.n11417 S.n11416 0.002
R12204 S.n12375 S.n12374 0.002
R12205 S.n4298 S.n4285 0.002
R12206 S.n5890 S.n5889 0.002
R12207 S.n6645 S.n6644 0.002
R12208 S.n7391 S.n7390 0.002
R12209 S.n7944 S.n7943 0.002
R12210 S.n8640 S.n8639 0.002
R12211 S.n9507 S.n9506 0.002
R12212 S.n10183 S.n10182 0.002
R12213 S.n10833 S.n10832 0.002
R12214 S.n11449 S.n11448 0.002
R12215 S.n12407 S.n12406 0.002
R12216 S.n5113 S.n5100 0.002
R12217 S.n6661 S.n6660 0.002
R12218 S.n7407 S.n7406 0.002
R12219 S.n7960 S.n7959 0.002
R12220 S.n8656 S.n8655 0.002
R12221 S.n9523 S.n9522 0.002
R12222 S.n10199 S.n10198 0.002
R12223 S.n10849 S.n10848 0.002
R12224 S.n11465 S.n11464 0.002
R12225 S.n12423 S.n12422 0.002
R12226 S.n5910 S.n5897 0.002
R12227 S.n7423 S.n7422 0.002
R12228 S.n7976 S.n7975 0.002
R12229 S.n8672 S.n8671 0.002
R12230 S.n9539 S.n9538 0.002
R12231 S.n10215 S.n10214 0.002
R12232 S.n10865 S.n10864 0.002
R12233 S.n11481 S.n11480 0.002
R12234 S.n12439 S.n12438 0.002
R12235 S.n6681 S.n6668 0.002
R12236 S.n7992 S.n7991 0.002
R12237 S.n8688 S.n8687 0.002
R12238 S.n9555 S.n9554 0.002
R12239 S.n10231 S.n10230 0.002
R12240 S.n10881 S.n10880 0.002
R12241 S.n11497 S.n11496 0.002
R12242 S.n12455 S.n12454 0.002
R12243 S.n7443 S.n7430 0.002
R12244 S.n8704 S.n8703 0.002
R12245 S.n9571 S.n9570 0.002
R12246 S.n10247 S.n10246 0.002
R12247 S.n10897 S.n10896 0.002
R12248 S.n11513 S.n11512 0.002
R12249 S.n12471 S.n12470 0.002
R12250 S.n8027 S.n8014 0.002
R12251 S.n9587 S.n9586 0.002
R12252 S.n10263 S.n10262 0.002
R12253 S.n10913 S.n10912 0.002
R12254 S.n11529 S.n11528 0.002
R12255 S.n12487 S.n12486 0.002
R12256 S.n8739 S.n8726 0.002
R12257 S.n10279 S.n10278 0.002
R12258 S.n10929 S.n10928 0.002
R12259 S.n11545 S.n11544 0.002
R12260 S.n12503 S.n12502 0.002
R12261 S.n9607 S.n9594 0.002
R12262 S.n10945 S.n10944 0.002
R12263 S.n11561 S.n11560 0.002
R12264 S.n12519 S.n12518 0.002
R12265 S.n10299 S.n10286 0.002
R12266 S.n11577 S.n11576 0.002
R12267 S.n12535 S.n12534 0.002
R12268 S.n10965 S.n10952 0.002
R12269 S.n12551 S.n12550 0.002
R12270 S.n3413 S.n3400 0.002
R12271 S.n5093 S.n5084 0.002
R12272 S.n5874 S.n5865 0.002
R12273 S.n6629 S.n6620 0.002
R12274 S.n7375 S.n7366 0.002
R12275 S.n7928 S.n7919 0.002
R12276 S.n8624 S.n8615 0.002
R12277 S.n9491 S.n9482 0.002
R12278 S.n10167 S.n10158 0.002
R12279 S.n10817 S.n10808 0.002
R12280 S.n11433 S.n11424 0.002
R12281 S.n12391 S.n12382 0.002
R12282 S.n10745 S.n10744 0.002
R12283 S.n10095 S.n10094 0.002
R12284 S.n9419 S.n9418 0.002
R12285 S.n8552 S.n8551 0.002
R12286 S.n7856 S.n7855 0.002
R12287 S.n7303 S.n7302 0.002
R12288 S.n6557 S.n6556 0.002
R12289 S.n5802 S.n5801 0.002
R12290 S.n5021 S.n5020 0.002
R12291 S.n4222 S.n4221 0.002
R12292 S.n3338 S.n3337 0.002
R12293 S.n2574 S.n2573 0.002
R12294 S.n1723 S.n1722 0.002
R12295 S.n751 S.n738 0.002
R12296 S.n805 S.n795 0.002
R12297 S.n2305 S.n2304 0.002
R12298 S.n3433 S.n3432 0.002
R12299 S.n3952 S.n3951 0.002
R12300 S.n4747 S.n4746 0.002
R12301 S.n5529 S.n5528 0.002
R12302 S.n6289 S.n6288 0.002
R12303 S.n7036 S.n7035 0.002
R12304 S.n8047 S.n8046 0.002
R12305 S.n8759 S.n8758 0.002
R12306 S.n9163 S.n9162 0.002
R12307 S.n9840 S.n9839 0.002
R12308 S.n10498 S.n10497 0.002
R12309 S.n11126 S.n11125 0.002
R12310 S.n1779 S.n1770 0.002
R12311 S.n3476 S.n3475 0.002
R12312 S.n3995 S.n3994 0.002
R12313 S.n4790 S.n4789 0.002
R12314 S.n5572 S.n5571 0.002
R12315 S.n6332 S.n6331 0.002
R12316 S.n7079 S.n7078 0.002
R12317 S.n8090 S.n8089 0.002
R12318 S.n8802 S.n8801 0.002
R12319 S.n9206 S.n9205 0.002
R12320 S.n9883 S.n9882 0.002
R12321 S.n10541 S.n10540 0.002
R12322 S.n11169 S.n11168 0.002
R12323 S.n11891 S.n11879 0.002
R12324 S.n12303 S.n12291 0.002
R12325 S.n12023 S.n11998 0.002
R12326 S.n11401 S.n11389 0.002
R12327 S.n11075 S.n11050 0.002
R12328 S.n10784 S.n10772 0.002
R12329 S.n10445 S.n10420 0.002
R12330 S.n10134 S.n10122 0.002
R12331 S.n9785 S.n9760 0.002
R12332 S.n9458 S.n9446 0.002
R12333 S.n9113 S.n9088 0.002
R12334 S.n8591 S.n8579 0.002
R12335 S.n8418 S.n8393 0.002
R12336 S.n7895 S.n7883 0.002
R12337 S.n7711 S.n7686 0.002
R12338 S.n7342 S.n7330 0.002
R12339 S.n6981 S.n6956 0.002
R12340 S.n6596 S.n6584 0.002
R12341 S.n6239 S.n6214 0.002
R12342 S.n5841 S.n5829 0.002
R12343 S.n5474 S.n5449 0.002
R12344 S.n5060 S.n5048 0.002
R12345 S.n4697 S.n4672 0.002
R12346 S.n4261 S.n4249 0.002
R12347 S.n3897 S.n3872 0.002
R12348 S.n3377 S.n3365 0.002
R12349 S.n3085 S.n3060 0.002
R12350 S.n2613 S.n2601 0.002
R12351 S.n2250 S.n2225 0.002
R12352 S.n1762 S.n1750 0.002
R12353 S.n1431 S.n1413 0.002
R12354 S.n787 S.n777 0.002
R12355 S.n920 S.n912 0.002
R12356 S.n10474 S.n10453 0.002
R12357 S.n10074 S.n10062 0.002
R12358 S.n9699 S.n9674 0.002
R12359 S.n9398 S.n9386 0.002
R12360 S.n9027 S.n9002 0.002
R12361 S.n8531 S.n8519 0.002
R12362 S.n8332 S.n8307 0.002
R12363 S.n7835 S.n7823 0.002
R12364 S.n7625 S.n7600 0.002
R12365 S.n7282 S.n7270 0.002
R12366 S.n6895 S.n6870 0.002
R12367 S.n6536 S.n6524 0.002
R12368 S.n6153 S.n6128 0.002
R12369 S.n5781 S.n5769 0.002
R12370 S.n5388 S.n5363 0.002
R12371 S.n5000 S.n4988 0.002
R12372 S.n4611 S.n4586 0.002
R12373 S.n4201 S.n4189 0.002
R12374 S.n3811 S.n3786 0.002
R12375 S.n3317 S.n3305 0.002
R12376 S.n2999 S.n2974 0.002
R12377 S.n2553 S.n2541 0.002
R12378 S.n2163 S.n2137 0.002
R12379 S.n1702 S.n1691 0.002
R12380 S.n1344 S.n1323 0.002
R12381 S.n837 S.n825 0.002
R12382 S.n822 S.n514 0.002
R12383 S.n9139 S.n9121 0.002
R12384 S.n8495 S.n8483 0.002
R12385 S.n8271 S.n8246 0.002
R12386 S.n7799 S.n7787 0.002
R12387 S.n7564 S.n7539 0.002
R12388 S.n7246 S.n7234 0.002
R12389 S.n6834 S.n6809 0.002
R12390 S.n6500 S.n6488 0.002
R12391 S.n6092 S.n6067 0.002
R12392 S.n5745 S.n5733 0.002
R12393 S.n5327 S.n5302 0.002
R12394 S.n4964 S.n4952 0.002
R12395 S.n4550 S.n4525 0.002
R12396 S.n4165 S.n4153 0.002
R12397 S.n3750 S.n3725 0.002
R12398 S.n3281 S.n3269 0.002
R12399 S.n2938 S.n2913 0.002
R12400 S.n2517 S.n2505 0.002
R12401 S.n2101 S.n2076 0.002
R12402 S.n1661 S.n1649 0.002
R12403 S.n1282 S.n1259 0.002
R12404 S.n714 S.n705 0.002
R12405 S.n484 S.n476 0.002
R12406 S.n7737 S.n7719 0.002
R12407 S.n7210 S.n7198 0.002
R12408 S.n6773 S.n6748 0.002
R12409 S.n6464 S.n6452 0.002
R12410 S.n6031 S.n6006 0.002
R12411 S.n5709 S.n5697 0.002
R12412 S.n5266 S.n5241 0.002
R12413 S.n4928 S.n4916 0.002
R12414 S.n4489 S.n4464 0.002
R12415 S.n4129 S.n4117 0.002
R12416 S.n3689 S.n3664 0.002
R12417 S.n3245 S.n3233 0.002
R12418 S.n2877 S.n2852 0.002
R12419 S.n2481 S.n2469 0.002
R12420 S.n2040 S.n2015 0.002
R12421 S.n1625 S.n1613 0.002
R12422 S.n1223 S.n1200 0.002
R12423 S.n681 S.n672 0.002
R12424 S.n440 S.n432 0.002
R12425 S.n6265 S.n6247 0.002
R12426 S.n5673 S.n5661 0.002
R12427 S.n5205 S.n5180 0.002
R12428 S.n4892 S.n4880 0.002
R12429 S.n4428 S.n4403 0.002
R12430 S.n4093 S.n4081 0.002
R12431 S.n3628 S.n3603 0.002
R12432 S.n3209 S.n3197 0.002
R12433 S.n2816 S.n2791 0.002
R12434 S.n2445 S.n2433 0.002
R12435 S.n1979 S.n1954 0.002
R12436 S.n1589 S.n1577 0.002
R12437 S.n1164 S.n1141 0.002
R12438 S.n648 S.n639 0.002
R12439 S.n396 S.n388 0.002
R12440 S.n4723 S.n4705 0.002
R12441 S.n4057 S.n4045 0.002
R12442 S.n3567 S.n3542 0.002
R12443 S.n3173 S.n3161 0.002
R12444 S.n2755 S.n2730 0.002
R12445 S.n2409 S.n2397 0.002
R12446 S.n1918 S.n1893 0.002
R12447 S.n1553 S.n1541 0.002
R12448 S.n1105 S.n1082 0.002
R12449 S.n615 S.n606 0.002
R12450 S.n352 S.n344 0.002
R12451 S.n3111 S.n3093 0.002
R12452 S.n2373 S.n2361 0.002
R12453 S.n1857 S.n1832 0.002
R12454 S.n1517 S.n1505 0.002
R12455 S.n1046 S.n1023 0.002
R12456 S.n582 S.n573 0.002
R12457 S.n308 S.n300 0.002
R12458 S.n1455 S.n1439 0.002
R12459 S.n549 S.n540 0.002
R12460 S.n264 S.n256 0.002
R12461 S.n11995 S.n11994 0.002
R12462 S.n883 S.n882 0.002
R12463 S.n1322 S.n1321 0.001
R12464 S.n1277 S.n1276 0.001
R12465 S.n1218 S.n1217 0.001
R12466 S.n1159 S.n1158 0.001
R12467 S.n1100 S.n1099 0.001
R12468 S.n1041 S.n1040 0.001
R12469 S.n83 S.n82 0.001
R12470 S.t7 S.n83 0.001
R12471 S.n11034 S.n11033 0.001
R12472 S.n10404 S.n10403 0.001
R12473 S.n9744 S.n9743 0.001
R12474 S.n9072 S.n9071 0.001
R12475 S.n8377 S.n8376 0.001
R12476 S.n7670 S.n7669 0.001
R12477 S.n6940 S.n6939 0.001
R12478 S.n6198 S.n6197 0.001
R12479 S.n5433 S.n5432 0.001
R12480 S.n4656 S.n4655 0.001
R12481 S.n3856 S.n3855 0.001
R12482 S.n3044 S.n3043 0.001
R12483 S.n2208 S.n2207 0.001
R12484 S.n1389 S.n1388 0.001
R12485 S.n11994 S.t0 0.001
R12486 S.t7 S.n57 0.001
R12487 S.t7 S.n3 0.001
R12488 S.t7 S.n169 0.001
R12489 S.t7 S.n180 0.001
R12490 S.t7 S.n11 0.001
R12491 S.t7 S.n20 0.001
R12492 S.t7 S.n29 0.001
R12493 S.t7 S.n38 0.001
R12494 S.t7 S.n47 0.001
R12495 S.n11633 S.n11632 0.001
R12496 S.n2163 S.n2148 0.001
R12497 S.n9815 S.n9814 0.001
R12498 S.n8448 S.n8447 0.001
R12499 S.n7011 S.n7010 0.001
R12500 S.n5504 S.n5503 0.001
R12501 S.n3927 S.n3926 0.001
R12502 S.n2280 S.n2279 0.001
R12503 S.n12608 S.n12607 0.001
R12504 S.n1428 S.n1427 0.001
R12505 S.n1759 S.n1758 0.001
R12506 S.n2247 S.n2246 0.001
R12507 S.n2610 S.n2609 0.001
R12508 S.n3082 S.n3081 0.001
R12509 S.n3374 S.n3373 0.001
R12510 S.n3894 S.n3893 0.001
R12511 S.n4258 S.n4257 0.001
R12512 S.n4694 S.n4693 0.001
R12513 S.n5057 S.n5056 0.001
R12514 S.n5471 S.n5470 0.001
R12515 S.n5838 S.n5837 0.001
R12516 S.n6236 S.n6235 0.001
R12517 S.n6593 S.n6592 0.001
R12518 S.n6978 S.n6977 0.001
R12519 S.n7339 S.n7338 0.001
R12520 S.n7708 S.n7707 0.001
R12521 S.n7892 S.n7891 0.001
R12522 S.n8415 S.n8414 0.001
R12523 S.n8588 S.n8587 0.001
R12524 S.n9110 S.n9109 0.001
R12525 S.n9455 S.n9454 0.001
R12526 S.n9782 S.n9781 0.001
R12527 S.n10131 S.n10130 0.001
R12528 S.n10442 S.n10441 0.001
R12529 S.n10781 S.n10780 0.001
R12530 S.n11072 S.n11071 0.001
R12531 S.n11398 S.n11397 0.001
R12532 S.n12020 S.n12019 0.001
R12533 S.n12300 S.n12299 0.001
R12534 S.n779 S.n778 0.001
R12535 S.n1690 S.n1689 0.001
R12536 S.n2160 S.n2159 0.001
R12537 S.n2550 S.n2549 0.001
R12538 S.n2996 S.n2995 0.001
R12539 S.n3314 S.n3313 0.001
R12540 S.n3808 S.n3807 0.001
R12541 S.n4198 S.n4197 0.001
R12542 S.n4608 S.n4607 0.001
R12543 S.n4997 S.n4996 0.001
R12544 S.n5385 S.n5384 0.001
R12545 S.n5778 S.n5777 0.001
R12546 S.n6150 S.n6149 0.001
R12547 S.n6533 S.n6532 0.001
R12548 S.n6892 S.n6891 0.001
R12549 S.n7279 S.n7278 0.001
R12550 S.n7622 S.n7621 0.001
R12551 S.n7832 S.n7831 0.001
R12552 S.n8329 S.n8328 0.001
R12553 S.n8528 S.n8527 0.001
R12554 S.n9024 S.n9023 0.001
R12555 S.n9395 S.n9394 0.001
R12556 S.n9696 S.n9695 0.001
R12557 S.n10071 S.n10070 0.001
R12558 S.n1658 S.n1657 0.001
R12559 S.n2098 S.n2097 0.001
R12560 S.n2514 S.n2513 0.001
R12561 S.n2935 S.n2934 0.001
R12562 S.n3278 S.n3277 0.001
R12563 S.n3747 S.n3746 0.001
R12564 S.n4162 S.n4161 0.001
R12565 S.n4547 S.n4546 0.001
R12566 S.n4961 S.n4960 0.001
R12567 S.n5324 S.n5323 0.001
R12568 S.n5742 S.n5741 0.001
R12569 S.n6089 S.n6088 0.001
R12570 S.n6497 S.n6496 0.001
R12571 S.n6831 S.n6830 0.001
R12572 S.n7243 S.n7242 0.001
R12573 S.n7561 S.n7560 0.001
R12574 S.n7796 S.n7795 0.001
R12575 S.n8268 S.n8267 0.001
R12576 S.n8492 S.n8491 0.001
R12577 S.n1622 S.n1621 0.001
R12578 S.n2037 S.n2036 0.001
R12579 S.n2478 S.n2477 0.001
R12580 S.n2874 S.n2873 0.001
R12581 S.n3242 S.n3241 0.001
R12582 S.n3686 S.n3685 0.001
R12583 S.n4126 S.n4125 0.001
R12584 S.n4486 S.n4485 0.001
R12585 S.n4925 S.n4924 0.001
R12586 S.n5263 S.n5262 0.001
R12587 S.n5706 S.n5705 0.001
R12588 S.n6028 S.n6027 0.001
R12589 S.n6461 S.n6460 0.001
R12590 S.n6770 S.n6769 0.001
R12591 S.n7207 S.n7206 0.001
R12592 S.n1586 S.n1585 0.001
R12593 S.n1976 S.n1975 0.001
R12594 S.n2442 S.n2441 0.001
R12595 S.n2813 S.n2812 0.001
R12596 S.n3206 S.n3205 0.001
R12597 S.n3625 S.n3624 0.001
R12598 S.n4090 S.n4089 0.001
R12599 S.n4425 S.n4424 0.001
R12600 S.n4889 S.n4888 0.001
R12601 S.n5202 S.n5201 0.001
R12602 S.n5670 S.n5669 0.001
R12603 S.n1550 S.n1549 0.001
R12604 S.n1915 S.n1914 0.001
R12605 S.n2406 S.n2405 0.001
R12606 S.n2752 S.n2751 0.001
R12607 S.n3170 S.n3169 0.001
R12608 S.n3564 S.n3563 0.001
R12609 S.n4054 S.n4053 0.001
R12610 S.n1514 S.n1513 0.001
R12611 S.n1854 S.n1853 0.001
R12612 S.n2370 S.n2369 0.001
R12613 S.n8977 S.n8976 0.001
R12614 S.n8282 S.n8281 0.001
R12615 S.n7575 S.n7574 0.001
R12616 S.n6845 S.n6844 0.001
R12617 S.n6103 S.n6102 0.001
R12618 S.n5338 S.n5337 0.001
R12619 S.n4561 S.n4560 0.001
R12620 S.n3761 S.n3760 0.001
R12621 S.n2949 S.n2948 0.001
R12622 S.n2112 S.n2111 0.001
R12623 S.n1294 S.n1293 0.001
R12624 S.n7514 S.n7513 0.001
R12625 S.n6784 S.n6783 0.001
R12626 S.n6042 S.n6041 0.001
R12627 S.n5277 S.n5276 0.001
R12628 S.n4500 S.n4499 0.001
R12629 S.n3700 S.n3699 0.001
R12630 S.n2888 S.n2887 0.001
R12631 S.n2051 S.n2050 0.001
R12632 S.n1235 S.n1234 0.001
R12633 S.n5981 S.n5980 0.001
R12634 S.n5216 S.n5215 0.001
R12635 S.n4439 S.n4438 0.001
R12636 S.n3639 S.n3638 0.001
R12637 S.n2827 S.n2826 0.001
R12638 S.n1990 S.n1989 0.001
R12639 S.n1176 S.n1175 0.001
R12640 S.n4378 S.n4377 0.001
R12641 S.n3578 S.n3577 0.001
R12642 S.n2766 S.n2765 0.001
R12643 S.n1929 S.n1928 0.001
R12644 S.n1117 S.n1116 0.001
R12645 S.n2705 S.n2704 0.001
R12646 S.n1868 S.n1867 0.001
R12647 S.n1058 S.n1057 0.001
R12648 S.n999 S.n998 0.001
R12649 S.n805 S.n796 0.001
R12650 S.n530 S.n529 0.001
R12651 S.n1477 S.n1476 0.001
R12652 S.n2351 S.n2350 0.001
R12653 S.n3133 S.n3132 0.001
R12654 S.n4035 S.n4034 0.001
R12655 S.n4852 S.n4851 0.001
R12656 S.n5651 S.n5650 0.001
R12657 S.n6424 S.n6423 0.001
R12658 S.n7188 S.n7187 0.001
R12659 S.n7759 S.n7758 0.001
R12660 S.n8473 S.n8472 0.001
R12661 S.n9358 S.n9357 0.001
R12662 S.n10052 S.n10051 0.001
R12663 S.n10720 S.n10719 0.001
R12664 S.n79 S.n78 0.001
R12665 S.n9699 S.n9684 0.001
R12666 S.n9027 S.n9012 0.001
R12667 S.n8332 S.n8317 0.001
R12668 S.n7625 S.n7610 0.001
R12669 S.n6895 S.n6880 0.001
R12670 S.n6153 S.n6138 0.001
R12671 S.n5388 S.n5373 0.001
R12672 S.n4611 S.n4596 0.001
R12673 S.n3811 S.n3796 0.001
R12674 S.n2999 S.n2984 0.001
R12675 S.n237 S.t7 0.001
R12676 S.t7 S.n193 0.001
R12677 S.t7 S.n155 0.001
R12678 S.t7 S.n143 0.001
R12679 S.t7 S.n131 0.001
R12680 S.t7 S.n118 0.001
R12681 S.t7 S.n105 0.001
R12682 S.t7 S.n92 0.001
R12683 S.n9364 S.n9363 0.001
R12684 S.n10726 S.n10725 0.001
R12685 S.n11364 S.n11363 0.001
R12686 S.n12286 S.n12285 0.001
R12687 S.n10057 S.n10056 0.001
R12688 S.n7765 S.n7764 0.001
R12689 S.n8478 S.n8477 0.001
R12690 S.n6430 S.n6429 0.001
R12691 S.n7193 S.n7192 0.001
R12692 S.n4858 S.n4857 0.001
R12693 S.n5656 S.n5655 0.001
R12694 S.n3139 S.n3138 0.001
R12695 S.n4040 S.n4039 0.001
R12696 S.n1483 S.n1482 0.001
R12697 S.n2356 S.n2355 0.001
R12698 S.n535 S.n534 0.001
R12699 S.n11923 S.n11920 0.001
R12700 S.n78 S.n77 0.001
R12701 S.n10474 S.n10455 0.001
R12702 S.n11870 S.n11869 0.001
R12703 S.n12344 S.n12343 0.001
R12704 S.n12067 S.n12066 0.001
R12705 S.n11125 S.n11124 0.001
R12706 S.n11139 S.n11138 0.001
R12707 S.n10497 S.n10496 0.001
R12708 S.n10511 S.n10510 0.001
R12709 S.n9839 S.n9838 0.001
R12710 S.n9853 S.n9852 0.001
R12711 S.n9162 S.n9161 0.001
R12712 S.n9176 S.n9175 0.001
R12713 S.n8758 S.n8757 0.001
R12714 S.n8772 S.n8771 0.001
R12715 S.n8046 S.n8045 0.001
R12716 S.n8060 S.n8059 0.001
R12717 S.n7035 S.n7034 0.001
R12718 S.n7049 S.n7048 0.001
R12719 S.n6288 S.n6287 0.001
R12720 S.n6302 S.n6301 0.001
R12721 S.n5528 S.n5527 0.001
R12722 S.n5542 S.n5541 0.001
R12723 S.n4746 S.n4745 0.001
R12724 S.n4760 S.n4759 0.001
R12725 S.n3951 S.n3950 0.001
R12726 S.n3965 S.n3964 0.001
R12727 S.n3432 S.n3431 0.001
R12728 S.n3446 S.n3445 0.001
R12729 S.n2304 S.n2303 0.001
R12730 S.n2318 S.n2317 0.001
R12731 S.n1798 S.n1797 0.001
R12732 S.n528 S.n527 0.001
R12733 S.n1475 S.n1474 0.001
R12734 S.n2349 S.n2348 0.001
R12735 S.n3131 S.n3130 0.001
R12736 S.n4033 S.n4032 0.001
R12737 S.n4850 S.n4849 0.001
R12738 S.n5649 S.n5648 0.001
R12739 S.n6422 S.n6421 0.001
R12740 S.n7186 S.n7185 0.001
R12741 S.n7757 S.n7756 0.001
R12742 S.n8471 S.n8470 0.001
R12743 S.n9356 S.n9355 0.001
R12744 S.n10050 S.n10049 0.001
R12745 S.n10718 S.n10717 0.001
R12746 S.n11920 S.t65 0.001
R12747 S.t244 S.n535 0.001
R12748 S.t225 S.n9364 0.001
R12749 S.t124 S.n10057 0.001
R12750 S.t144 S.n10726 0.001
R12751 S.t47 S.n11364 0.001
R12752 S.t106 S.n12286 0.001
R12753 S.t11 S.n7765 0.001
R12754 S.t40 S.n8478 0.001
R12755 S.t4 S.n6430 0.001
R12756 S.t102 S.n7193 0.001
R12757 S.t77 S.n4858 0.001
R12758 S.t25 S.n5656 0.001
R12759 S.t38 S.n3139 0.001
R12760 S.t94 S.n4040 0.001
R12761 S.t175 S.n1483 0.001
R12762 S.t187 S.n2356 0.001
R12763 S.n1827 S.n1826 0.001
R12764 S.n529 S.n528 0.001
R12765 S.n1476 S.n1475 0.001
R12766 S.n2350 S.n2349 0.001
R12767 S.n3132 S.n3131 0.001
R12768 S.n4034 S.n4033 0.001
R12769 S.n4851 S.n4850 0.001
R12770 S.n5650 S.n5649 0.001
R12771 S.n6423 S.n6422 0.001
R12772 S.n7187 S.n7186 0.001
R12773 S.n7758 S.n7757 0.001
R12774 S.n8472 S.n8471 0.001
R12775 S.n9357 S.n9356 0.001
R12776 S.n10051 S.n10050 0.001
R12777 S.n10719 S.n10718 0.001
R12778 S.n12311 S.n12310 0.001
R12779 S.n823 S.n822 0.001
R12780 S.n714 S.n706 0.001
R12781 S.n681 S.n673 0.001
R12782 S.n648 S.n640 0.001
R12783 S.n615 S.n607 0.001
R12784 S.n582 S.n574 0.001
R12785 S.n549 S.n541 0.001
R12786 S.n973 S.n972 0.001
R12787 S.n986 S.n985 0.001
R12788 S.n2671 S.n2670 0.001
R12789 S.n3513 S.n3512 0.001
R12790 S.n4344 S.n4343 0.001
R12791 S.n5150 S.n5149 0.001
R12792 S.n5947 S.n5946 0.001
R12793 S.n6718 S.n6717 0.001
R12794 S.n7480 S.n7479 0.001
R12795 S.n8216 S.n8215 0.001
R12796 S.n8943 S.n8942 0.001
R12797 S.n9644 S.n9643 0.001
R12798 S.n10336 S.n10335 0.001
R12799 S.n11000 S.n10999 0.001
R12800 S.n865 S.n864 0.001
R12801 S.n78 S.n68 0.001
R12802 S.n78 S.n74 0.001
R12803 S.n78 S.n73 0.001
R12804 S.n78 S.n72 0.001
R12805 S.n78 S.n71 0.001
R12806 S.n78 S.n70 0.001
R12807 S.n78 S.n69 0.001
R12808 S.n11906 S.n11905 0.001
R12809 S.n12315 S.n12314 0.001
R12810 S.n938 S.n937 0.001
R12811 S.n915 S.n914 0.001
R12812 S.n1420 S.n1419 0.001
R12813 S.n11886 S.n11885 0.001
R12814 S.n12298 S.n12297 0.001
R12815 S.n12014 S.n12013 0.001
R12816 S.n11396 S.n11395 0.001
R12817 S.n11066 S.n11065 0.001
R12818 S.n10779 S.n10778 0.001
R12819 S.n10436 S.n10435 0.001
R12820 S.n10129 S.n10128 0.001
R12821 S.n9776 S.n9775 0.001
R12822 S.n9453 S.n9452 0.001
R12823 S.n9104 S.n9103 0.001
R12824 S.n8586 S.n8585 0.001
R12825 S.n8409 S.n8408 0.001
R12826 S.n7890 S.n7889 0.001
R12827 S.n7702 S.n7701 0.001
R12828 S.n7337 S.n7336 0.001
R12829 S.n6972 S.n6971 0.001
R12830 S.n6591 S.n6590 0.001
R12831 S.n6230 S.n6229 0.001
R12832 S.n5836 S.n5835 0.001
R12833 S.n5465 S.n5464 0.001
R12834 S.n5055 S.n5054 0.001
R12835 S.n4688 S.n4687 0.001
R12836 S.n4256 S.n4255 0.001
R12837 S.n3888 S.n3887 0.001
R12838 S.n3372 S.n3371 0.001
R12839 S.n3076 S.n3075 0.001
R12840 S.n2608 S.n2607 0.001
R12841 S.n2241 S.n2240 0.001
R12842 S.n1757 S.n1756 0.001
R12843 S.n782 S.n781 0.001
R12844 S.n479 S.n478 0.001
R12845 S.n1275 S.n1274 0.001
R12846 S.n9128 S.n9127 0.001
R12847 S.n8490 S.n8489 0.001
R12848 S.n8262 S.n8261 0.001
R12849 S.n7794 S.n7793 0.001
R12850 S.n7555 S.n7554 0.001
R12851 S.n7241 S.n7240 0.001
R12852 S.n6825 S.n6824 0.001
R12853 S.n6495 S.n6494 0.001
R12854 S.n6083 S.n6082 0.001
R12855 S.n5740 S.n5739 0.001
R12856 S.n5318 S.n5317 0.001
R12857 S.n4959 S.n4958 0.001
R12858 S.n4541 S.n4540 0.001
R12859 S.n4160 S.n4159 0.001
R12860 S.n3741 S.n3740 0.001
R12861 S.n3276 S.n3275 0.001
R12862 S.n2929 S.n2928 0.001
R12863 S.n2512 S.n2511 0.001
R12864 S.n2092 S.n2091 0.001
R12865 S.n1656 S.n1655 0.001
R12866 S.n502 S.n501 0.001
R12867 S.n9804 S.n9803 0.001
R12868 S.n9374 S.n9373 0.001
R12869 S.n8981 S.n8980 0.001
R12870 S.n8507 S.n8506 0.001
R12871 S.n8286 S.n8285 0.001
R12872 S.n7811 S.n7810 0.001
R12873 S.n7579 S.n7578 0.001
R12874 S.n7258 S.n7257 0.001
R12875 S.n6849 S.n6848 0.001
R12876 S.n6512 S.n6511 0.001
R12877 S.n6107 S.n6106 0.001
R12878 S.n5757 S.n5756 0.001
R12879 S.n5342 S.n5341 0.001
R12880 S.n4976 S.n4975 0.001
R12881 S.n4565 S.n4564 0.001
R12882 S.n4177 S.n4176 0.001
R12883 S.n3765 S.n3764 0.001
R12884 S.n3293 S.n3292 0.001
R12885 S.n2953 S.n2952 0.001
R12886 S.n2529 S.n2528 0.001
R12887 S.n2116 S.n2115 0.001
R12888 S.n1673 S.n1672 0.001
R12889 S.n1694 S.n1693 0.001
R12890 S.n1326 S.n1325 0.001
R12891 S.n517 S.n516 0.001
R12892 S.n828 S.n827 0.001
R12893 S.n2154 S.n2153 0.001
R12894 S.n2990 S.n2989 0.001
R12895 S.n3802 S.n3801 0.001
R12896 S.n4602 S.n4601 0.001
R12897 S.n5379 S.n5378 0.001
R12898 S.n6144 S.n6143 0.001
R12899 S.n6886 S.n6885 0.001
R12900 S.n7616 S.n7615 0.001
R12901 S.n8323 S.n8322 0.001
R12902 S.n9018 S.n9017 0.001
R12903 S.n9690 S.n9689 0.001
R12904 S.n10463 S.n10462 0.001
R12905 S.n10069 S.n10068 0.001
R12906 S.n9393 S.n9392 0.001
R12907 S.n8526 S.n8525 0.001
R12908 S.n7830 S.n7829 0.001
R12909 S.n7277 S.n7276 0.001
R12910 S.n6531 S.n6530 0.001
R12911 S.n5776 S.n5775 0.001
R12912 S.n4995 S.n4994 0.001
R12913 S.n4196 S.n4195 0.001
R12914 S.n3312 S.n3311 0.001
R12915 S.n2548 S.n2547 0.001
R12916 S.n1365 S.n1364 0.001
R12917 S.n742 S.n741 0.001
R12918 S.n860 S.n859 0.001
R12919 S.n11097 S.n11096 0.001
R12920 S.n10743 S.n10742 0.001
R12921 S.n10381 S.n10380 0.001
R12922 S.n10093 S.n10092 0.001
R12923 S.n9721 S.n9720 0.001
R12924 S.n9417 S.n9416 0.001
R12925 S.n9049 S.n9048 0.001
R12926 S.n8550 S.n8549 0.001
R12927 S.n8354 S.n8353 0.001
R12928 S.n7854 S.n7853 0.001
R12929 S.n7647 S.n7646 0.001
R12930 S.n7301 S.n7300 0.001
R12931 S.n6917 S.n6916 0.001
R12932 S.n6555 S.n6554 0.001
R12933 S.n6175 S.n6174 0.001
R12934 S.n5800 S.n5799 0.001
R12935 S.n5410 S.n5409 0.001
R12936 S.n5019 S.n5018 0.001
R12937 S.n4633 S.n4632 0.001
R12938 S.n4220 S.n4219 0.001
R12939 S.n3833 S.n3832 0.001
R12940 S.n3336 S.n3335 0.001
R12941 S.n3021 S.n3020 0.001
R12942 S.n2572 S.n2571 0.001
R12943 S.n2185 S.n2184 0.001
R12944 S.n1721 S.n1720 0.001
R12945 S.n1393 S.n1392 0.001
R12946 S.n762 S.n761 0.001
R12947 S.n1740 S.n1739 0.001
R12948 S.n2212 S.n2211 0.001
R12949 S.n2586 S.n2585 0.001
R12950 S.n3048 S.n3047 0.001
R12951 S.n3350 S.n3349 0.001
R12952 S.n3860 S.n3859 0.001
R12953 S.n4234 S.n4233 0.001
R12954 S.n4660 S.n4659 0.001
R12955 S.n5033 S.n5032 0.001
R12956 S.n5437 S.n5436 0.001
R12957 S.n5814 S.n5813 0.001
R12958 S.n6202 S.n6201 0.001
R12959 S.n6569 S.n6568 0.001
R12960 S.n6944 S.n6943 0.001
R12961 S.n7315 S.n7314 0.001
R12962 S.n7674 S.n7673 0.001
R12963 S.n7868 S.n7867 0.001
R12964 S.n8381 S.n8380 0.001
R12965 S.n8564 S.n8563 0.001
R12966 S.n9076 S.n9075 0.001
R12967 S.n9431 S.n9430 0.001
R12968 S.n9748 S.n9747 0.001
R12969 S.n10107 S.n10106 0.001
R12970 S.n10408 S.n10407 0.001
R12971 S.n10757 S.n10756 0.001
R12972 S.n11038 S.n11037 0.001
R12973 S.n11374 S.n11373 0.001
R12974 S.n12042 S.n12041 0.001
R12975 S.n886 S.n885 0.001
R12976 S.n1297 S.n1296 0.001
R12977 S.n726 S.n725 0.001
R12978 S.n709 S.n708 0.001
R12979 S.n435 S.n434 0.001
R12980 S.n1216 S.n1215 0.001
R12981 S.n7726 S.n7725 0.001
R12982 S.n7205 S.n7204 0.001
R12983 S.n6764 S.n6763 0.001
R12984 S.n6459 S.n6458 0.001
R12985 S.n6022 S.n6021 0.001
R12986 S.n5704 S.n5703 0.001
R12987 S.n5257 S.n5256 0.001
R12988 S.n4923 S.n4922 0.001
R12989 S.n4480 S.n4479 0.001
R12990 S.n4124 S.n4123 0.001
R12991 S.n3680 S.n3679 0.001
R12992 S.n3240 S.n3239 0.001
R12993 S.n2868 S.n2867 0.001
R12994 S.n2476 S.n2475 0.001
R12995 S.n2031 S.n2030 0.001
R12996 S.n1620 S.n1619 0.001
R12997 S.n458 S.n457 0.001
R12998 S.n8437 S.n8436 0.001
R12999 S.n7775 S.n7774 0.001
R13000 S.n7518 S.n7517 0.001
R13001 S.n7222 S.n7221 0.001
R13002 S.n6788 S.n6787 0.001
R13003 S.n6476 S.n6475 0.001
R13004 S.n6046 S.n6045 0.001
R13005 S.n5721 S.n5720 0.001
R13006 S.n5281 S.n5280 0.001
R13007 S.n4940 S.n4939 0.001
R13008 S.n4504 S.n4503 0.001
R13009 S.n4141 S.n4140 0.001
R13010 S.n3704 S.n3703 0.001
R13011 S.n3257 S.n3256 0.001
R13012 S.n2892 S.n2891 0.001
R13013 S.n2493 S.n2492 0.001
R13014 S.n2055 S.n2054 0.001
R13015 S.n1637 S.n1636 0.001
R13016 S.n1238 S.n1237 0.001
R13017 S.n693 S.n692 0.001
R13018 S.n676 S.n675 0.001
R13019 S.n391 S.n390 0.001
R13020 S.n1157 S.n1156 0.001
R13021 S.n6254 S.n6253 0.001
R13022 S.n5668 S.n5667 0.001
R13023 S.n5196 S.n5195 0.001
R13024 S.n4887 S.n4886 0.001
R13025 S.n4419 S.n4418 0.001
R13026 S.n4088 S.n4087 0.001
R13027 S.n3619 S.n3618 0.001
R13028 S.n3204 S.n3203 0.001
R13029 S.n2807 S.n2806 0.001
R13030 S.n2440 S.n2439 0.001
R13031 S.n1970 S.n1969 0.001
R13032 S.n1584 S.n1583 0.001
R13033 S.n414 S.n413 0.001
R13034 S.n7000 S.n6999 0.001
R13035 S.n6440 S.n6439 0.001
R13036 S.n5985 S.n5984 0.001
R13037 S.n5685 S.n5684 0.001
R13038 S.n5220 S.n5219 0.001
R13039 S.n4904 S.n4903 0.001
R13040 S.n4443 S.n4442 0.001
R13041 S.n4105 S.n4104 0.001
R13042 S.n3643 S.n3642 0.001
R13043 S.n3221 S.n3220 0.001
R13044 S.n2831 S.n2830 0.001
R13045 S.n2457 S.n2456 0.001
R13046 S.n1994 S.n1993 0.001
R13047 S.n1601 S.n1600 0.001
R13048 S.n1179 S.n1178 0.001
R13049 S.n660 S.n659 0.001
R13050 S.n643 S.n642 0.001
R13051 S.n347 S.n346 0.001
R13052 S.n1098 S.n1097 0.001
R13053 S.n4712 S.n4711 0.001
R13054 S.n4052 S.n4051 0.001
R13055 S.n3558 S.n3557 0.001
R13056 S.n3168 S.n3167 0.001
R13057 S.n2746 S.n2745 0.001
R13058 S.n2404 S.n2403 0.001
R13059 S.n1909 S.n1908 0.001
R13060 S.n1548 S.n1547 0.001
R13061 S.n370 S.n369 0.001
R13062 S.n5493 S.n5492 0.001
R13063 S.n4868 S.n4867 0.001
R13064 S.n4382 S.n4381 0.001
R13065 S.n4069 S.n4068 0.001
R13066 S.n3582 S.n3581 0.001
R13067 S.n3185 S.n3184 0.001
R13068 S.n2770 S.n2769 0.001
R13069 S.n2421 S.n2420 0.001
R13070 S.n1933 S.n1932 0.001
R13071 S.n1565 S.n1564 0.001
R13072 S.n1120 S.n1119 0.001
R13073 S.n627 S.n626 0.001
R13074 S.n610 S.n609 0.001
R13075 S.n303 S.n302 0.001
R13076 S.n1039 S.n1038 0.001
R13077 S.n3100 S.n3099 0.001
R13078 S.n2368 S.n2367 0.001
R13079 S.n1848 S.n1847 0.001
R13080 S.n1512 S.n1511 0.001
R13081 S.n326 S.n325 0.001
R13082 S.n3916 S.n3915 0.001
R13083 S.n3149 S.n3148 0.001
R13084 S.n2709 S.n2708 0.001
R13085 S.n2385 S.n2384 0.001
R13086 S.n1872 S.n1871 0.001
R13087 S.n1529 S.n1528 0.001
R13088 S.n1061 S.n1060 0.001
R13089 S.n594 S.n593 0.001
R13090 S.n577 S.n576 0.001
R13091 S.n259 S.n258 0.001
R13092 S.n1446 S.n1445 0.001
R13093 S.n282 S.n281 0.001
R13094 S.n2269 S.n2268 0.001
R13095 S.n1493 S.n1492 0.001
R13096 S.n1002 S.n1001 0.001
R13097 S.n561 S.n560 0.001
R13098 S.n544 S.n543 0.001
R13099 S.n799 S.n798 0.001
R13100 S.n1802 S.n1801 0.001
R13101 S.n1465 S.n1464 0.001
R13102 S.n2309 S.n2308 0.001
R13103 S.n2291 S.n2290 0.001
R13104 S.n3437 S.n3436 0.001
R13105 S.n3121 S.n3120 0.001
R13106 S.n3956 S.n3955 0.001
R13107 S.n3938 S.n3937 0.001
R13108 S.n4751 S.n4750 0.001
R13109 S.n4733 S.n4732 0.001
R13110 S.n5533 S.n5532 0.001
R13111 S.n5515 S.n5514 0.001
R13112 S.n6293 S.n6292 0.001
R13113 S.n6275 S.n6274 0.001
R13114 S.n7040 S.n7039 0.001
R13115 S.n7022 S.n7021 0.001
R13116 S.n8051 S.n8050 0.001
R13117 S.n7747 S.n7746 0.001
R13118 S.n8763 S.n8762 0.001
R13119 S.n8459 S.n8458 0.001
R13120 S.n9167 S.n9166 0.001
R13121 S.n9149 S.n9148 0.001
R13122 S.n9844 S.n9843 0.001
R13123 S.n9826 S.n9825 0.001
R13124 S.n10502 S.n10501 0.001
R13125 S.n10484 S.n10483 0.001
R13126 S.n11130 S.n11129 0.001
R13127 S.n11112 S.n11111 0.001
R13128 S.n12058 S.n12057 0.001
R13129 S.n12337 S.n12336 0.001
R13130 S.n11862 S.n11861 0.001
R13131 S.n1774 S.n1773 0.001
R13132 S.n2332 S.n2331 0.001
R13133 S.n11851 S.n11850 0.001
R13134 S.n12358 S.n12357 0.001
R13135 S.n12081 S.n12080 0.001
R13136 S.n11167 S.n11166 0.001
R13137 S.n11153 S.n11152 0.001
R13138 S.n10539 S.n10538 0.001
R13139 S.n10525 S.n10524 0.001
R13140 S.n9881 S.n9880 0.001
R13141 S.n9867 S.n9866 0.001
R13142 S.n9204 S.n9203 0.001
R13143 S.n9190 S.n9189 0.001
R13144 S.n8800 S.n8799 0.001
R13145 S.n8786 S.n8785 0.001
R13146 S.n8088 S.n8087 0.001
R13147 S.n8074 S.n8073 0.001
R13148 S.n7077 S.n7076 0.001
R13149 S.n7063 S.n7062 0.001
R13150 S.n6330 S.n6329 0.001
R13151 S.n6316 S.n6315 0.001
R13152 S.n5570 S.n5569 0.001
R13153 S.n5556 S.n5555 0.001
R13154 S.n4788 S.n4787 0.001
R13155 S.n4774 S.n4773 0.001
R13156 S.n3993 S.n3992 0.001
R13157 S.n3979 S.n3978 0.001
R13158 S.n3474 S.n3473 0.001
R13159 S.n3460 S.n3459 0.001
R13160 S.n2649 S.n2648 0.001
R13161 S.n2625 S.n2624 0.001
R13162 S.n3491 S.n3490 0.001
R13163 S.n11836 S.n11835 0.001
R13164 S.n12373 S.n12372 0.001
R13165 S.n12097 S.n12096 0.001
R13166 S.n11415 S.n11414 0.001
R13167 S.n11184 S.n11183 0.001
R13168 S.n10799 S.n10798 0.001
R13169 S.n10556 S.n10555 0.001
R13170 S.n10149 S.n10148 0.001
R13171 S.n9898 S.n9897 0.001
R13172 S.n9473 S.n9472 0.001
R13173 S.n9221 S.n9220 0.001
R13174 S.n8606 S.n8605 0.001
R13175 S.n8817 S.n8816 0.001
R13176 S.n7910 S.n7909 0.001
R13177 S.n8105 S.n8104 0.001
R13178 S.n7357 S.n7356 0.001
R13179 S.n7094 S.n7093 0.001
R13180 S.n6611 S.n6610 0.001
R13181 S.n6347 S.n6346 0.001
R13182 S.n5856 S.n5855 0.001
R13183 S.n5587 S.n5586 0.001
R13184 S.n5075 S.n5074 0.001
R13185 S.n4805 S.n4804 0.001
R13186 S.n4276 S.n4275 0.001
R13187 S.n4010 S.n4009 0.001
R13188 S.n3392 S.n3391 0.001
R13189 S.n11817 S.n11816 0.001
R13190 S.n12386 S.n12385 0.001
R13191 S.n12108 S.n12107 0.001
R13192 S.n11428 S.n11427 0.001
R13193 S.n11195 S.n11194 0.001
R13194 S.n10812 S.n10811 0.001
R13195 S.n10567 S.n10566 0.001
R13196 S.n10162 S.n10161 0.001
R13197 S.n9909 S.n9908 0.001
R13198 S.n9486 S.n9485 0.001
R13199 S.n9232 S.n9231 0.001
R13200 S.n8619 S.n8618 0.001
R13201 S.n8828 S.n8827 0.001
R13202 S.n7923 S.n7922 0.001
R13203 S.n8116 S.n8115 0.001
R13204 S.n7370 S.n7369 0.001
R13205 S.n7105 S.n7104 0.001
R13206 S.n6624 S.n6623 0.001
R13207 S.n6358 S.n6357 0.001
R13208 S.n5869 S.n5868 0.001
R13209 S.n5598 S.n5597 0.001
R13210 S.n5088 S.n5087 0.001
R13211 S.n4816 S.n4815 0.001
R13212 S.n4021 S.n4020 0.001
R13213 S.n4319 S.n4318 0.001
R13214 S.n3404 S.n3403 0.001
R13215 S.n4289 S.n4288 0.001
R13216 S.n4835 S.n4834 0.001
R13217 S.n11806 S.n11805 0.001
R13218 S.n12405 S.n12404 0.001
R13219 S.n12127 S.n12126 0.001
R13220 S.n11447 S.n11446 0.001
R13221 S.n11214 S.n11213 0.001
R13222 S.n10831 S.n10830 0.001
R13223 S.n10586 S.n10585 0.001
R13224 S.n10181 S.n10180 0.001
R13225 S.n9928 S.n9927 0.001
R13226 S.n9505 S.n9504 0.001
R13227 S.n9251 S.n9250 0.001
R13228 S.n8638 S.n8637 0.001
R13229 S.n8847 S.n8846 0.001
R13230 S.n7942 S.n7941 0.001
R13231 S.n8135 S.n8134 0.001
R13232 S.n7389 S.n7388 0.001
R13233 S.n7124 S.n7123 0.001
R13234 S.n6643 S.n6642 0.001
R13235 S.n6377 S.n6376 0.001
R13236 S.n5888 S.n5887 0.001
R13237 S.n5617 S.n5616 0.001
R13238 S.n5128 S.n5127 0.001
R13239 S.n5104 S.n5103 0.001
R13240 S.n5632 S.n5631 0.001
R13241 S.n11791 S.n11790 0.001
R13242 S.n12421 S.n12420 0.001
R13243 S.n12142 S.n12141 0.001
R13244 S.n11463 S.n11462 0.001
R13245 S.n11229 S.n11228 0.001
R13246 S.n10847 S.n10846 0.001
R13247 S.n10601 S.n10600 0.001
R13248 S.n10197 S.n10196 0.001
R13249 S.n9943 S.n9942 0.001
R13250 S.n9521 S.n9520 0.001
R13251 S.n9266 S.n9265 0.001
R13252 S.n8654 S.n8653 0.001
R13253 S.n8862 S.n8861 0.001
R13254 S.n7958 S.n7957 0.001
R13255 S.n8150 S.n8149 0.001
R13256 S.n7405 S.n7404 0.001
R13257 S.n7139 S.n7138 0.001
R13258 S.n6659 S.n6658 0.001
R13259 S.n6392 S.n6391 0.001
R13260 S.n5925 S.n5924 0.001
R13261 S.n5901 S.n5900 0.001
R13262 S.n6407 S.n6406 0.001
R13263 S.n11776 S.n11775 0.001
R13264 S.n12437 S.n12436 0.001
R13265 S.n12157 S.n12156 0.001
R13266 S.n11479 S.n11478 0.001
R13267 S.n11244 S.n11243 0.001
R13268 S.n10863 S.n10862 0.001
R13269 S.n10616 S.n10615 0.001
R13270 S.n10213 S.n10212 0.001
R13271 S.n9958 S.n9957 0.001
R13272 S.n9537 S.n9536 0.001
R13273 S.n9281 S.n9280 0.001
R13274 S.n8670 S.n8669 0.001
R13275 S.n8877 S.n8876 0.001
R13276 S.n7974 S.n7973 0.001
R13277 S.n8165 S.n8164 0.001
R13278 S.n7421 S.n7420 0.001
R13279 S.n7154 S.n7153 0.001
R13280 S.n6696 S.n6695 0.001
R13281 S.n6672 S.n6671 0.001
R13282 S.n7169 S.n7168 0.001
R13283 S.n11761 S.n11760 0.001
R13284 S.n12453 S.n12452 0.001
R13285 S.n12172 S.n12171 0.001
R13286 S.n11495 S.n11494 0.001
R13287 S.n11259 S.n11258 0.001
R13288 S.n10879 S.n10878 0.001
R13289 S.n10631 S.n10630 0.001
R13290 S.n10229 S.n10228 0.001
R13291 S.n9973 S.n9972 0.001
R13292 S.n9553 S.n9552 0.001
R13293 S.n9296 S.n9295 0.001
R13294 S.n8686 S.n8685 0.001
R13295 S.n8892 S.n8891 0.001
R13296 S.n7990 S.n7989 0.001
R13297 S.n8180 S.n8179 0.001
R13298 S.n7458 S.n7457 0.001
R13299 S.n7434 S.n7433 0.001
R13300 S.n8195 S.n8194 0.001
R13301 S.n11746 S.n11745 0.001
R13302 S.n12469 S.n12468 0.001
R13303 S.n12187 S.n12186 0.001
R13304 S.n11511 S.n11510 0.001
R13305 S.n11274 S.n11273 0.001
R13306 S.n10895 S.n10894 0.001
R13307 S.n10646 S.n10645 0.001
R13308 S.n10245 S.n10244 0.001
R13309 S.n9988 S.n9987 0.001
R13310 S.n9569 S.n9568 0.001
R13311 S.n9311 S.n9310 0.001
R13312 S.n8702 S.n8701 0.001
R13313 S.n8907 S.n8906 0.001
R13314 S.n8006 S.n8005 0.001
R13315 S.n8018 S.n8017 0.001
R13316 S.n8922 S.n8921 0.001
R13317 S.n11731 S.n11730 0.001
R13318 S.n12485 S.n12484 0.001
R13319 S.n12202 S.n12201 0.001
R13320 S.n11527 S.n11526 0.001
R13321 S.n11289 S.n11288 0.001
R13322 S.n10911 S.n10910 0.001
R13323 S.n10661 S.n10660 0.001
R13324 S.n10261 S.n10260 0.001
R13325 S.n10003 S.n10002 0.001
R13326 S.n9585 S.n9584 0.001
R13327 S.n9326 S.n9325 0.001
R13328 S.n8718 S.n8717 0.001
R13329 S.n8730 S.n8729 0.001
R13330 S.n9341 S.n9340 0.001
R13331 S.n11716 S.n11715 0.001
R13332 S.n12501 S.n12500 0.001
R13333 S.n12217 S.n12216 0.001
R13334 S.n11543 S.n11542 0.001
R13335 S.n11304 S.n11303 0.001
R13336 S.n10927 S.n10926 0.001
R13337 S.n10676 S.n10675 0.001
R13338 S.n10277 S.n10276 0.001
R13339 S.n10018 S.n10017 0.001
R13340 S.n9622 S.n9621 0.001
R13341 S.n9598 S.n9597 0.001
R13342 S.n10033 S.n10032 0.001
R13343 S.n11701 S.n11700 0.001
R13344 S.n12517 S.n12516 0.001
R13345 S.n12232 S.n12231 0.001
R13346 S.n11559 S.n11558 0.001
R13347 S.n11319 S.n11318 0.001
R13348 S.n10943 S.n10942 0.001
R13349 S.n10691 S.n10690 0.001
R13350 S.n10314 S.n10313 0.001
R13351 S.n10290 S.n10289 0.001
R13352 S.n10706 S.n10705 0.001
R13353 S.n11686 S.n11685 0.001
R13354 S.n12533 S.n12532 0.001
R13355 S.n12247 S.n12246 0.001
R13356 S.n11575 S.n11574 0.001
R13357 S.n11334 S.n11333 0.001
R13358 S.n10980 S.n10979 0.001
R13359 S.n10956 S.n10955 0.001
R13360 S.n11349 S.n11348 0.001
R13361 S.n11671 S.n11670 0.001
R13362 S.n12549 S.n12548 0.001
R13363 S.n12262 S.n12261 0.001
R13364 S.n11615 S.n11614 0.001
R13365 S.n11586 S.n11585 0.001
R13366 S.n12576 S.n12575 0.001
R13367 S.n11652 S.n11651 0.001
R13368 S.n12278 S.n12277 0.001
R13369 S.n78 S.n76 0.001
R13370 S.n10722 S.n10721 0.001
R13371 S.n10054 S.n10053 0.001
R13372 S.n9360 S.n9359 0.001
R13373 S.n8475 S.n8474 0.001
R13374 S.n7761 S.n7760 0.001
R13375 S.n7190 S.n7189 0.001
R13376 S.n6426 S.n6425 0.001
R13377 S.n5653 S.n5652 0.001
R13378 S.n4854 S.n4853 0.001
R13379 S.n4037 S.n4036 0.001
R13380 S.n3135 S.n3134 0.001
R13381 S.n2353 S.n2352 0.001
R13382 S.n1479 S.n1478 0.001
R13383 S.n532 S.n531 0.001
R13384 S.t65 S.n11914 0.001
R13385 S.t65 S.n11917 0.001
R13386 S.t106 S.n12333 0.001
R13387 S.t106 S.n12330 0.001
R13388 S.n12330 S.n12327 0.001
R13389 S.n12591 S.t157 0.001
R13390 S.n12611 S.n12593 0.001
R13391 S.t159 S.n953 0.001
R13392 S.t159 S.n956 0.001
R13393 S.t159 S.n926 0.001
R13394 S.t159 S.n923 0.001
R13395 S.n923 S.n920 0.001
R13396 S.t72 S.n1437 0.001
R13397 S.t72 S.n1434 0.001
R13398 S.n1434 S.n1431 0.001
R13399 S.t65 S.n11897 0.001
R13400 S.t65 S.n11894 0.001
R13401 S.n11894 S.n11891 0.001
R13402 S.t106 S.n12309 0.001
R13403 S.t106 S.n12306 0.001
R13404 S.n12306 S.n12303 0.001
R13405 S.t157 S.n12029 0.001
R13406 S.t157 S.n12026 0.001
R13407 S.n12026 S.n12023 0.001
R13408 S.t47 S.n11407 0.001
R13409 S.t47 S.n11404 0.001
R13410 S.n11404 S.n11401 0.001
R13411 S.t115 S.n11081 0.001
R13412 S.t115 S.n11078 0.001
R13413 S.n11078 S.n11075 0.001
R13414 S.t144 S.n10790 0.001
R13415 S.t144 S.n10787 0.001
R13416 S.n10787 S.n10784 0.001
R13417 S.t35 S.n10451 0.001
R13418 S.t35 S.n10448 0.001
R13419 S.n10448 S.n10445 0.001
R13420 S.t124 S.n10140 0.001
R13421 S.t124 S.n10137 0.001
R13422 S.n10137 S.n10134 0.001
R13423 S.t61 S.n9791 0.001
R13424 S.t61 S.n9788 0.001
R13425 S.n9788 S.n9785 0.001
R13426 S.t225 S.n9464 0.001
R13427 S.t225 S.n9461 0.001
R13428 S.n9461 S.n9458 0.001
R13429 S.t31 S.n9119 0.001
R13430 S.t31 S.n9116 0.001
R13431 S.n9116 S.n9113 0.001
R13432 S.t40 S.n8597 0.001
R13433 S.t40 S.n8594 0.001
R13434 S.n8594 S.n8591 0.001
R13435 S.t300 S.n8424 0.001
R13436 S.t300 S.n8421 0.001
R13437 S.n8421 S.n8418 0.001
R13438 S.t11 S.n7901 0.001
R13439 S.t11 S.n7898 0.001
R13440 S.n7898 S.n7895 0.001
R13441 S.t27 S.n7717 0.001
R13442 S.t27 S.n7714 0.001
R13443 S.n7714 S.n7711 0.001
R13444 S.t102 S.n7348 0.001
R13445 S.t102 S.n7345 0.001
R13446 S.n7345 S.n7342 0.001
R13447 S.t130 S.n6987 0.001
R13448 S.t130 S.n6984 0.001
R13449 S.n6984 S.n6981 0.001
R13450 S.t4 S.n6602 0.001
R13451 S.t4 S.n6599 0.001
R13452 S.n6599 S.n6596 0.001
R13453 S.t69 S.n6245 0.001
R13454 S.t69 S.n6242 0.001
R13455 S.n6242 S.n6239 0.001
R13456 S.t25 S.n5847 0.001
R13457 S.t25 S.n5844 0.001
R13458 S.n5844 S.n5841 0.001
R13459 S.t109 S.n5480 0.001
R13460 S.t109 S.n5477 0.001
R13461 S.n5477 S.n5474 0.001
R13462 S.t77 S.n5066 0.001
R13463 S.t77 S.n5063 0.001
R13464 S.n5063 S.n5060 0.001
R13465 S.t33 S.n4703 0.001
R13466 S.t33 S.n4700 0.001
R13467 S.n4700 S.n4697 0.001
R13468 S.t94 S.n4267 0.001
R13469 S.t94 S.n4264 0.001
R13470 S.n4264 S.n4261 0.001
R13471 S.t53 S.n3903 0.001
R13472 S.t53 S.n3900 0.001
R13473 S.n3900 S.n3897 0.001
R13474 S.t38 S.n3383 0.001
R13475 S.t38 S.n3380 0.001
R13476 S.n3380 S.n3377 0.001
R13477 S.t84 S.n3091 0.001
R13478 S.t84 S.n3088 0.001
R13479 S.n3088 S.n3085 0.001
R13480 S.t187 S.n2619 0.001
R13481 S.t187 S.n2616 0.001
R13482 S.n2616 S.n2613 0.001
R13483 S.t259 S.n2256 0.001
R13484 S.t259 S.n2253 0.001
R13485 S.n2253 S.n2250 0.001
R13486 S.t175 S.n1768 0.001
R13487 S.t175 S.n1765 0.001
R13488 S.n1765 S.n1762 0.001
R13489 S.t244 S.n793 0.001
R13490 S.t244 S.n790 0.001
R13491 S.n790 S.n787 0.001
R13492 S.t159 S.n490 0.001
R13493 S.t159 S.n487 0.001
R13494 S.n487 S.n484 0.001
R13495 S.t72 S.n1288 0.001
R13496 S.t72 S.n1285 0.001
R13497 S.n1285 S.n1282 0.001
R13498 S.t31 S.n9142 0.001
R13499 S.t31 S.n9145 0.001
R13500 S.t40 S.n8501 0.001
R13501 S.t40 S.n8498 0.001
R13502 S.n8498 S.n8495 0.001
R13503 S.t300 S.n8277 0.001
R13504 S.t300 S.n8274 0.001
R13505 S.n8274 S.n8271 0.001
R13506 S.t11 S.n7805 0.001
R13507 S.t11 S.n7802 0.001
R13508 S.n7802 S.n7799 0.001
R13509 S.t27 S.n7570 0.001
R13510 S.t27 S.n7567 0.001
R13511 S.n7567 S.n7564 0.001
R13512 S.t102 S.n7252 0.001
R13513 S.t102 S.n7249 0.001
R13514 S.n7249 S.n7246 0.001
R13515 S.t130 S.n6840 0.001
R13516 S.t130 S.n6837 0.001
R13517 S.n6837 S.n6834 0.001
R13518 S.t4 S.n6506 0.001
R13519 S.t4 S.n6503 0.001
R13520 S.n6503 S.n6500 0.001
R13521 S.t69 S.n6098 0.001
R13522 S.t69 S.n6095 0.001
R13523 S.n6095 S.n6092 0.001
R13524 S.t25 S.n5751 0.001
R13525 S.t25 S.n5748 0.001
R13526 S.n5748 S.n5745 0.001
R13527 S.t109 S.n5333 0.001
R13528 S.t109 S.n5330 0.001
R13529 S.n5330 S.n5327 0.001
R13530 S.t77 S.n4970 0.001
R13531 S.t77 S.n4967 0.001
R13532 S.n4967 S.n4964 0.001
R13533 S.t33 S.n4556 0.001
R13534 S.t33 S.n4553 0.001
R13535 S.n4553 S.n4550 0.001
R13536 S.t94 S.n4171 0.001
R13537 S.t94 S.n4168 0.001
R13538 S.n4168 S.n4165 0.001
R13539 S.t53 S.n3756 0.001
R13540 S.t53 S.n3753 0.001
R13541 S.n3753 S.n3750 0.001
R13542 S.t38 S.n3287 0.001
R13543 S.t38 S.n3284 0.001
R13544 S.n3284 S.n3281 0.001
R13545 S.t84 S.n2944 0.001
R13546 S.t84 S.n2941 0.001
R13547 S.n2941 S.n2938 0.001
R13548 S.t187 S.n2523 0.001
R13549 S.t187 S.n2520 0.001
R13550 S.n2520 S.n2517 0.001
R13551 S.t259 S.n2107 0.001
R13552 S.t259 S.n2104 0.001
R13553 S.n2104 S.n2101 0.001
R13554 S.t175 S.n1667 0.001
R13555 S.t175 S.n1664 0.001
R13556 S.n1664 S.n1661 0.001
R13557 S.t159 S.n513 0.001
R13558 S.t159 S.n510 0.001
R13559 S.n510 S.n507 0.001
R13560 S.t61 S.n9819 0.001
R13561 S.t61 S.n9822 0.001
R13562 S.t225 S.n9385 0.001
R13563 S.t225 S.n9382 0.001
R13564 S.n9382 S.n9379 0.001
R13565 S.t31 S.n9001 0.001
R13566 S.t31 S.n8998 0.001
R13567 S.n8998 S.n8995 0.001
R13568 S.t40 S.n8518 0.001
R13569 S.t40 S.n8515 0.001
R13570 S.n8515 S.n8512 0.001
R13571 S.t300 S.n8306 0.001
R13572 S.t300 S.n8303 0.001
R13573 S.n8303 S.n8300 0.001
R13574 S.t11 S.n7822 0.001
R13575 S.t11 S.n7819 0.001
R13576 S.n7819 S.n7816 0.001
R13577 S.t27 S.n7599 0.001
R13578 S.t27 S.n7596 0.001
R13579 S.n7596 S.n7593 0.001
R13580 S.t102 S.n7269 0.001
R13581 S.t102 S.n7266 0.001
R13582 S.n7266 S.n7263 0.001
R13583 S.t130 S.n6869 0.001
R13584 S.t130 S.n6866 0.001
R13585 S.n6866 S.n6863 0.001
R13586 S.t4 S.n6523 0.001
R13587 S.t4 S.n6520 0.001
R13588 S.n6520 S.n6517 0.001
R13589 S.t69 S.n6127 0.001
R13590 S.t69 S.n6124 0.001
R13591 S.n6124 S.n6121 0.001
R13592 S.t25 S.n5768 0.001
R13593 S.t25 S.n5765 0.001
R13594 S.n5765 S.n5762 0.001
R13595 S.t109 S.n5362 0.001
R13596 S.t109 S.n5359 0.001
R13597 S.n5359 S.n5356 0.001
R13598 S.t77 S.n4987 0.001
R13599 S.t77 S.n4984 0.001
R13600 S.n4984 S.n4981 0.001
R13601 S.t33 S.n4585 0.001
R13602 S.t33 S.n4582 0.001
R13603 S.n4582 S.n4579 0.001
R13604 S.t94 S.n4188 0.001
R13605 S.t94 S.n4185 0.001
R13606 S.n4185 S.n4182 0.001
R13607 S.t53 S.n3785 0.001
R13608 S.t53 S.n3782 0.001
R13609 S.n3782 S.n3779 0.001
R13610 S.t38 S.n3304 0.001
R13611 S.t38 S.n3301 0.001
R13612 S.n3301 S.n3298 0.001
R13613 S.t84 S.n2973 0.001
R13614 S.t84 S.n2970 0.001
R13615 S.n2970 S.n2967 0.001
R13616 S.t187 S.n2540 0.001
R13617 S.t187 S.n2537 0.001
R13618 S.n2537 S.n2534 0.001
R13619 S.t259 S.n2136 0.001
R13620 S.t259 S.n2133 0.001
R13621 S.n2133 S.n2130 0.001
R13622 S.t175 S.n1686 0.001
R13623 S.t175 S.n1683 0.001
R13624 S.n1683 S.n1680 0.001
R13625 S.t175 S.n1708 0.001
R13626 S.t175 S.n1705 0.001
R13627 S.n1705 S.n1702 0.001
R13628 S.t72 S.n1350 0.001
R13629 S.t72 S.n1347 0.001
R13630 S.n1347 S.n1344 0.001
R13631 S.n814 S.t244 0.001
R13632 S.n822 S.n817 0.001
R13633 S.t159 S.n843 0.001
R13634 S.t159 S.n840 0.001
R13635 S.n840 S.n837 0.001
R13636 S.t259 S.n2169 0.001
R13637 S.t259 S.n2166 0.001
R13638 S.n2166 S.n2163 0.001
R13639 S.t84 S.n3005 0.001
R13640 S.t84 S.n3002 0.001
R13641 S.n3002 S.n2999 0.001
R13642 S.t53 S.n3817 0.001
R13643 S.t53 S.n3814 0.001
R13644 S.n3814 S.n3811 0.001
R13645 S.t33 S.n4617 0.001
R13646 S.t33 S.n4614 0.001
R13647 S.n4614 S.n4611 0.001
R13648 S.t109 S.n5394 0.001
R13649 S.t109 S.n5391 0.001
R13650 S.n5391 S.n5388 0.001
R13651 S.t69 S.n6159 0.001
R13652 S.t69 S.n6156 0.001
R13653 S.n6156 S.n6153 0.001
R13654 S.t130 S.n6901 0.001
R13655 S.t130 S.n6898 0.001
R13656 S.n6898 S.n6895 0.001
R13657 S.t27 S.n7631 0.001
R13658 S.t27 S.n7628 0.001
R13659 S.n7628 S.n7625 0.001
R13660 S.t300 S.n8338 0.001
R13661 S.t300 S.n8335 0.001
R13662 S.n8335 S.n8332 0.001
R13663 S.t31 S.n9033 0.001
R13664 S.t31 S.n9030 0.001
R13665 S.n9030 S.n9027 0.001
R13666 S.t61 S.n9705 0.001
R13667 S.t61 S.n9702 0.001
R13668 S.n9702 S.n9699 0.001
R13669 S.t35 S.n10477 0.001
R13670 S.t35 S.n10480 0.001
R13671 S.t124 S.n10080 0.001
R13672 S.t124 S.n10077 0.001
R13673 S.n10077 S.n10074 0.001
R13674 S.t225 S.n9404 0.001
R13675 S.t225 S.n9401 0.001
R13676 S.n9401 S.n9398 0.001
R13677 S.t40 S.n8537 0.001
R13678 S.t40 S.n8534 0.001
R13679 S.n8534 S.n8531 0.001
R13680 S.t11 S.n7841 0.001
R13681 S.t11 S.n7838 0.001
R13682 S.n7838 S.n7835 0.001
R13683 S.t102 S.n7288 0.001
R13684 S.t102 S.n7285 0.001
R13685 S.n7285 S.n7282 0.001
R13686 S.t4 S.n6542 0.001
R13687 S.t4 S.n6539 0.001
R13688 S.n6539 S.n6536 0.001
R13689 S.t25 S.n5787 0.001
R13690 S.t25 S.n5784 0.001
R13691 S.n5784 S.n5781 0.001
R13692 S.t77 S.n5006 0.001
R13693 S.t77 S.n5003 0.001
R13694 S.n5003 S.n5000 0.001
R13695 S.t94 S.n4207 0.001
R13696 S.t94 S.n4204 0.001
R13697 S.n4204 S.n4201 0.001
R13698 S.t38 S.n3323 0.001
R13699 S.t38 S.n3320 0.001
R13700 S.n3320 S.n3317 0.001
R13701 S.t187 S.n2559 0.001
R13702 S.t187 S.n2556 0.001
R13703 S.n2556 S.n2553 0.001
R13704 S.t72 S.n1384 0.001
R13705 S.t72 S.n1381 0.001
R13706 S.n1381 S.n1378 0.001
R13707 S.t244 S.n757 0.001
R13708 S.t244 S.n754 0.001
R13709 S.n754 S.n751 0.001
R13710 S.t159 S.n876 0.001
R13711 S.t159 S.n873 0.001
R13712 S.n873 S.n870 0.001
R13713 S.t115 S.n11105 0.001
R13714 S.t115 S.n11108 0.001
R13715 S.t144 S.n10751 0.001
R13716 S.t144 S.n10748 0.001
R13717 S.n10748 S.n10745 0.001
R13718 S.t35 S.n10399 0.001
R13719 S.t35 S.n10396 0.001
R13720 S.n10396 S.n10393 0.001
R13721 S.t124 S.n10101 0.001
R13722 S.t124 S.n10098 0.001
R13723 S.n10098 S.n10095 0.001
R13724 S.t61 S.n9739 0.001
R13725 S.t61 S.n9736 0.001
R13726 S.n9736 S.n9733 0.001
R13727 S.t225 S.n9425 0.001
R13728 S.t225 S.n9422 0.001
R13729 S.n9422 S.n9419 0.001
R13730 S.t31 S.n9067 0.001
R13731 S.t31 S.n9064 0.001
R13732 S.n9064 S.n9061 0.001
R13733 S.t40 S.n8558 0.001
R13734 S.t40 S.n8555 0.001
R13735 S.n8555 S.n8552 0.001
R13736 S.t300 S.n8372 0.001
R13737 S.t300 S.n8369 0.001
R13738 S.n8369 S.n8366 0.001
R13739 S.t11 S.n7862 0.001
R13740 S.t11 S.n7859 0.001
R13741 S.n7859 S.n7856 0.001
R13742 S.t27 S.n7665 0.001
R13743 S.t27 S.n7662 0.001
R13744 S.n7662 S.n7659 0.001
R13745 S.t102 S.n7309 0.001
R13746 S.t102 S.n7306 0.001
R13747 S.n7306 S.n7303 0.001
R13748 S.t130 S.n6935 0.001
R13749 S.t130 S.n6932 0.001
R13750 S.n6932 S.n6929 0.001
R13751 S.t4 S.n6563 0.001
R13752 S.t4 S.n6560 0.001
R13753 S.n6560 S.n6557 0.001
R13754 S.t69 S.n6193 0.001
R13755 S.t69 S.n6190 0.001
R13756 S.n6190 S.n6187 0.001
R13757 S.t25 S.n5808 0.001
R13758 S.t25 S.n5805 0.001
R13759 S.n5805 S.n5802 0.001
R13760 S.t109 S.n5428 0.001
R13761 S.t109 S.n5425 0.001
R13762 S.n5425 S.n5422 0.001
R13763 S.t77 S.n5027 0.001
R13764 S.t77 S.n5024 0.001
R13765 S.n5024 S.n5021 0.001
R13766 S.t33 S.n4651 0.001
R13767 S.t33 S.n4648 0.001
R13768 S.n4648 S.n4645 0.001
R13769 S.t94 S.n4228 0.001
R13770 S.t94 S.n4225 0.001
R13771 S.n4225 S.n4222 0.001
R13772 S.t53 S.n3851 0.001
R13773 S.t53 S.n3848 0.001
R13774 S.n3848 S.n3845 0.001
R13775 S.t38 S.n3344 0.001
R13776 S.t38 S.n3341 0.001
R13777 S.n3341 S.n3338 0.001
R13778 S.t84 S.n3039 0.001
R13779 S.t84 S.n3036 0.001
R13780 S.n3036 S.n3033 0.001
R13781 S.t187 S.n2580 0.001
R13782 S.t187 S.n2577 0.001
R13783 S.n2577 S.n2574 0.001
R13784 S.t259 S.n2203 0.001
R13785 S.t259 S.n2200 0.001
R13786 S.n2200 S.n2197 0.001
R13787 S.t175 S.n1729 0.001
R13788 S.t175 S.n1726 0.001
R13789 S.n1726 S.n1723 0.001
R13790 S.t72 S.n1412 0.001
R13791 S.t72 S.n1409 0.001
R13792 S.n1409 S.n1406 0.001
R13793 S.t244 S.n776 0.001
R13794 S.t244 S.n773 0.001
R13795 S.n773 S.n770 0.001
R13796 S.t175 S.n1749 0.001
R13797 S.t175 S.n1746 0.001
R13798 S.n1746 S.n1743 0.001
R13799 S.t259 S.n2224 0.001
R13800 S.t259 S.n2221 0.001
R13801 S.n2221 S.n2218 0.001
R13802 S.t187 S.n2600 0.001
R13803 S.t187 S.n2597 0.001
R13804 S.n2597 S.n2594 0.001
R13805 S.t84 S.n3059 0.001
R13806 S.t84 S.n3056 0.001
R13807 S.n3056 S.n3053 0.001
R13808 S.t38 S.n3364 0.001
R13809 S.t38 S.n3361 0.001
R13810 S.n3361 S.n3358 0.001
R13811 S.t53 S.n3871 0.001
R13812 S.t53 S.n3868 0.001
R13813 S.n3868 S.n3865 0.001
R13814 S.t94 S.n4248 0.001
R13815 S.t94 S.n4245 0.001
R13816 S.n4245 S.n4242 0.001
R13817 S.t33 S.n4671 0.001
R13818 S.t33 S.n4668 0.001
R13819 S.n4668 S.n4665 0.001
R13820 S.t77 S.n5047 0.001
R13821 S.t77 S.n5044 0.001
R13822 S.n5044 S.n5041 0.001
R13823 S.t109 S.n5448 0.001
R13824 S.t109 S.n5445 0.001
R13825 S.n5445 S.n5442 0.001
R13826 S.t25 S.n5828 0.001
R13827 S.t25 S.n5825 0.001
R13828 S.n5825 S.n5822 0.001
R13829 S.t69 S.n6213 0.001
R13830 S.t69 S.n6210 0.001
R13831 S.n6210 S.n6207 0.001
R13832 S.t4 S.n6583 0.001
R13833 S.t4 S.n6580 0.001
R13834 S.n6580 S.n6577 0.001
R13835 S.t130 S.n6955 0.001
R13836 S.t130 S.n6952 0.001
R13837 S.n6952 S.n6949 0.001
R13838 S.t102 S.n7329 0.001
R13839 S.t102 S.n7326 0.001
R13840 S.n7326 S.n7323 0.001
R13841 S.t27 S.n7685 0.001
R13842 S.t27 S.n7682 0.001
R13843 S.n7682 S.n7679 0.001
R13844 S.t11 S.n7882 0.001
R13845 S.t11 S.n7879 0.001
R13846 S.n7879 S.n7876 0.001
R13847 S.t300 S.n8392 0.001
R13848 S.t300 S.n8389 0.001
R13849 S.n8389 S.n8386 0.001
R13850 S.t40 S.n8578 0.001
R13851 S.t40 S.n8575 0.001
R13852 S.n8575 S.n8572 0.001
R13853 S.t31 S.n9087 0.001
R13854 S.t31 S.n9084 0.001
R13855 S.n9084 S.n9081 0.001
R13856 S.t225 S.n9445 0.001
R13857 S.t225 S.n9442 0.001
R13858 S.n9442 S.n9439 0.001
R13859 S.t61 S.n9759 0.001
R13860 S.t61 S.n9756 0.001
R13861 S.n9756 S.n9753 0.001
R13862 S.t124 S.n10121 0.001
R13863 S.t124 S.n10118 0.001
R13864 S.n10118 S.n10115 0.001
R13865 S.t35 S.n10419 0.001
R13866 S.t35 S.n10416 0.001
R13867 S.n10416 S.n10413 0.001
R13868 S.t144 S.n10771 0.001
R13869 S.t144 S.n10768 0.001
R13870 S.n10768 S.n10765 0.001
R13871 S.t115 S.n11049 0.001
R13872 S.t115 S.n11046 0.001
R13873 S.n11046 S.n11043 0.001
R13874 S.t47 S.n11388 0.001
R13875 S.t47 S.n11385 0.001
R13876 S.n11385 S.n11382 0.001
R13877 S.t157 S.n12050 0.001
R13878 S.t157 S.n12053 0.001
R13879 S.t159 S.n905 0.001
R13880 S.t159 S.n902 0.001
R13881 S.n902 S.n899 0.001
R13882 S.t72 S.n1316 0.001
R13883 S.t72 S.n1313 0.001
R13884 S.n1313 S.n1310 0.001
R13885 S.t244 S.n737 0.001
R13886 S.t244 S.n734 0.001
R13887 S.n734 S.n731 0.001
R13888 S.t244 S.n720 0.001
R13889 S.t244 S.n717 0.001
R13890 S.n717 S.n714 0.001
R13891 S.t159 S.n446 0.001
R13892 S.t159 S.n443 0.001
R13893 S.n443 S.n440 0.001
R13894 S.t72 S.n1229 0.001
R13895 S.t72 S.n1226 0.001
R13896 S.n1226 S.n1223 0.001
R13897 S.t27 S.n7740 0.001
R13898 S.t27 S.n7743 0.001
R13899 S.t102 S.n7216 0.001
R13900 S.t102 S.n7213 0.001
R13901 S.n7213 S.n7210 0.001
R13902 S.t130 S.n6779 0.001
R13903 S.t130 S.n6776 0.001
R13904 S.n6776 S.n6773 0.001
R13905 S.t4 S.n6470 0.001
R13906 S.t4 S.n6467 0.001
R13907 S.n6467 S.n6464 0.001
R13908 S.t69 S.n6037 0.001
R13909 S.t69 S.n6034 0.001
R13910 S.n6034 S.n6031 0.001
R13911 S.t25 S.n5715 0.001
R13912 S.t25 S.n5712 0.001
R13913 S.n5712 S.n5709 0.001
R13914 S.t109 S.n5272 0.001
R13915 S.t109 S.n5269 0.001
R13916 S.n5269 S.n5266 0.001
R13917 S.t77 S.n4934 0.001
R13918 S.t77 S.n4931 0.001
R13919 S.n4931 S.n4928 0.001
R13920 S.t33 S.n4495 0.001
R13921 S.t33 S.n4492 0.001
R13922 S.n4492 S.n4489 0.001
R13923 S.t94 S.n4135 0.001
R13924 S.t94 S.n4132 0.001
R13925 S.n4132 S.n4129 0.001
R13926 S.t53 S.n3695 0.001
R13927 S.t53 S.n3692 0.001
R13928 S.n3692 S.n3689 0.001
R13929 S.t38 S.n3251 0.001
R13930 S.t38 S.n3248 0.001
R13931 S.n3248 S.n3245 0.001
R13932 S.t84 S.n2883 0.001
R13933 S.t84 S.n2880 0.001
R13934 S.n2880 S.n2877 0.001
R13935 S.t187 S.n2487 0.001
R13936 S.t187 S.n2484 0.001
R13937 S.n2484 S.n2481 0.001
R13938 S.t259 S.n2046 0.001
R13939 S.t259 S.n2043 0.001
R13940 S.n2043 S.n2040 0.001
R13941 S.t175 S.n1631 0.001
R13942 S.t175 S.n1628 0.001
R13943 S.n1628 S.n1625 0.001
R13944 S.t159 S.n469 0.001
R13945 S.n469 S.n466 0.001
R13946 S.t300 S.n8452 0.001
R13947 S.t300 S.n8455 0.001
R13948 S.t11 S.n7786 0.001
R13949 S.t11 S.n7783 0.001
R13950 S.n7783 S.n7780 0.001
R13951 S.t27 S.n7538 0.001
R13952 S.t27 S.n7535 0.001
R13953 S.n7535 S.n7532 0.001
R13954 S.t102 S.n7233 0.001
R13955 S.t102 S.n7230 0.001
R13956 S.n7230 S.n7227 0.001
R13957 S.t130 S.n6808 0.001
R13958 S.t130 S.n6805 0.001
R13959 S.n6805 S.n6802 0.001
R13960 S.t4 S.n6487 0.001
R13961 S.t4 S.n6484 0.001
R13962 S.n6484 S.n6481 0.001
R13963 S.t69 S.n6066 0.001
R13964 S.t69 S.n6063 0.001
R13965 S.n6063 S.n6060 0.001
R13966 S.t25 S.n5732 0.001
R13967 S.t25 S.n5729 0.001
R13968 S.n5729 S.n5726 0.001
R13969 S.t109 S.n5301 0.001
R13970 S.t109 S.n5298 0.001
R13971 S.n5298 S.n5295 0.001
R13972 S.t77 S.n4951 0.001
R13973 S.t77 S.n4948 0.001
R13974 S.n4948 S.n4945 0.001
R13975 S.t33 S.n4524 0.001
R13976 S.t33 S.n4521 0.001
R13977 S.n4521 S.n4518 0.001
R13978 S.t94 S.n4152 0.001
R13979 S.t94 S.n4149 0.001
R13980 S.n4149 S.n4146 0.001
R13981 S.t53 S.n3724 0.001
R13982 S.t53 S.n3721 0.001
R13983 S.n3721 S.n3718 0.001
R13984 S.t38 S.n3268 0.001
R13985 S.t38 S.n3265 0.001
R13986 S.n3265 S.n3262 0.001
R13987 S.t84 S.n2912 0.001
R13988 S.t84 S.n2909 0.001
R13989 S.n2909 S.n2906 0.001
R13990 S.t187 S.n2504 0.001
R13991 S.t187 S.n2501 0.001
R13992 S.n2501 S.n2498 0.001
R13993 S.t259 S.n2075 0.001
R13994 S.t259 S.n2072 0.001
R13995 S.n2072 S.n2069 0.001
R13996 S.t175 S.n1648 0.001
R13997 S.t175 S.n1645 0.001
R13998 S.n1645 S.n1642 0.001
R13999 S.t72 S.n1258 0.001
R14000 S.t72 S.n1255 0.001
R14001 S.n1255 S.n1252 0.001
R14002 S.t244 S.n704 0.001
R14003 S.t244 S.n701 0.001
R14004 S.n701 S.n698 0.001
R14005 S.t244 S.n687 0.001
R14006 S.t244 S.n684 0.001
R14007 S.n684 S.n681 0.001
R14008 S.t159 S.n402 0.001
R14009 S.t159 S.n399 0.001
R14010 S.n399 S.n396 0.001
R14011 S.t72 S.n1170 0.001
R14012 S.t72 S.n1167 0.001
R14013 S.n1167 S.n1164 0.001
R14014 S.t69 S.n6268 0.001
R14015 S.t69 S.n6271 0.001
R14016 S.t25 S.n5679 0.001
R14017 S.t25 S.n5676 0.001
R14018 S.n5676 S.n5673 0.001
R14019 S.t109 S.n5211 0.001
R14020 S.t109 S.n5208 0.001
R14021 S.n5208 S.n5205 0.001
R14022 S.t77 S.n4898 0.001
R14023 S.t77 S.n4895 0.001
R14024 S.n4895 S.n4892 0.001
R14025 S.t33 S.n4434 0.001
R14026 S.t33 S.n4431 0.001
R14027 S.n4431 S.n4428 0.001
R14028 S.t94 S.n4099 0.001
R14029 S.t94 S.n4096 0.001
R14030 S.n4096 S.n4093 0.001
R14031 S.t53 S.n3634 0.001
R14032 S.t53 S.n3631 0.001
R14033 S.n3631 S.n3628 0.001
R14034 S.t38 S.n3215 0.001
R14035 S.t38 S.n3212 0.001
R14036 S.n3212 S.n3209 0.001
R14037 S.t84 S.n2822 0.001
R14038 S.t84 S.n2819 0.001
R14039 S.n2819 S.n2816 0.001
R14040 S.t187 S.n2451 0.001
R14041 S.t187 S.n2448 0.001
R14042 S.n2448 S.n2445 0.001
R14043 S.t259 S.n1985 0.001
R14044 S.t259 S.n1982 0.001
R14045 S.n1982 S.n1979 0.001
R14046 S.t175 S.n1595 0.001
R14047 S.t175 S.n1592 0.001
R14048 S.n1592 S.n1589 0.001
R14049 S.t159 S.n425 0.001
R14050 S.t159 S.n422 0.001
R14051 S.n422 S.n419 0.001
R14052 S.t130 S.n7015 0.001
R14053 S.t130 S.n7018 0.001
R14054 S.t4 S.n6451 0.001
R14055 S.t4 S.n6448 0.001
R14056 S.n6448 S.n6445 0.001
R14057 S.t69 S.n6005 0.001
R14058 S.t69 S.n6002 0.001
R14059 S.n6002 S.n5999 0.001
R14060 S.t25 S.n5696 0.001
R14061 S.t25 S.n5693 0.001
R14062 S.n5693 S.n5690 0.001
R14063 S.t109 S.n5240 0.001
R14064 S.t109 S.n5237 0.001
R14065 S.n5237 S.n5234 0.001
R14066 S.t77 S.n4915 0.001
R14067 S.t77 S.n4912 0.001
R14068 S.n4912 S.n4909 0.001
R14069 S.t33 S.n4463 0.001
R14070 S.t33 S.n4460 0.001
R14071 S.n4460 S.n4457 0.001
R14072 S.t94 S.n4116 0.001
R14073 S.t94 S.n4113 0.001
R14074 S.n4113 S.n4110 0.001
R14075 S.t53 S.n3663 0.001
R14076 S.t53 S.n3660 0.001
R14077 S.n3660 S.n3657 0.001
R14078 S.t38 S.n3232 0.001
R14079 S.t38 S.n3229 0.001
R14080 S.n3229 S.n3226 0.001
R14081 S.t84 S.n2851 0.001
R14082 S.t84 S.n2848 0.001
R14083 S.n2848 S.n2845 0.001
R14084 S.t187 S.n2468 0.001
R14085 S.t187 S.n2465 0.001
R14086 S.n2465 S.n2462 0.001
R14087 S.t259 S.n2014 0.001
R14088 S.t259 S.n2011 0.001
R14089 S.n2011 S.n2008 0.001
R14090 S.t175 S.n1612 0.001
R14091 S.t175 S.n1609 0.001
R14092 S.n1609 S.n1606 0.001
R14093 S.t72 S.n1199 0.001
R14094 S.t72 S.n1196 0.001
R14095 S.n1196 S.n1193 0.001
R14096 S.t244 S.n671 0.001
R14097 S.t244 S.n668 0.001
R14098 S.n668 S.n665 0.001
R14099 S.t244 S.n654 0.001
R14100 S.t244 S.n651 0.001
R14101 S.n651 S.n648 0.001
R14102 S.t159 S.n358 0.001
R14103 S.t159 S.n355 0.001
R14104 S.n355 S.n352 0.001
R14105 S.t72 S.n1111 0.001
R14106 S.t72 S.n1108 0.001
R14107 S.n1108 S.n1105 0.001
R14108 S.t33 S.n4726 0.001
R14109 S.t33 S.n4729 0.001
R14110 S.t94 S.n4063 0.001
R14111 S.t94 S.n4060 0.001
R14112 S.n4060 S.n4057 0.001
R14113 S.t53 S.n3573 0.001
R14114 S.t53 S.n3570 0.001
R14115 S.n3570 S.n3567 0.001
R14116 S.t38 S.n3179 0.001
R14117 S.t38 S.n3176 0.001
R14118 S.n3176 S.n3173 0.001
R14119 S.t84 S.n2761 0.001
R14120 S.t84 S.n2758 0.001
R14121 S.n2758 S.n2755 0.001
R14122 S.t187 S.n2415 0.001
R14123 S.t187 S.n2412 0.001
R14124 S.n2412 S.n2409 0.001
R14125 S.t259 S.n1924 0.001
R14126 S.t259 S.n1921 0.001
R14127 S.n1921 S.n1918 0.001
R14128 S.t175 S.n1559 0.001
R14129 S.t175 S.n1556 0.001
R14130 S.n1556 S.n1553 0.001
R14131 S.t159 S.n381 0.001
R14132 S.t159 S.n378 0.001
R14133 S.n378 S.n375 0.001
R14134 S.t109 S.n5508 0.001
R14135 S.t109 S.n5511 0.001
R14136 S.t77 S.n4879 0.001
R14137 S.t77 S.n4876 0.001
R14138 S.n4876 S.n4873 0.001
R14139 S.t33 S.n4402 0.001
R14140 S.t33 S.n4399 0.001
R14141 S.n4399 S.n4396 0.001
R14142 S.t94 S.n4080 0.001
R14143 S.t94 S.n4077 0.001
R14144 S.n4077 S.n4074 0.001
R14145 S.t53 S.n3602 0.001
R14146 S.t53 S.n3599 0.001
R14147 S.n3599 S.n3596 0.001
R14148 S.t38 S.n3196 0.001
R14149 S.t38 S.n3193 0.001
R14150 S.n3193 S.n3190 0.001
R14151 S.t84 S.n2790 0.001
R14152 S.t84 S.n2787 0.001
R14153 S.n2787 S.n2784 0.001
R14154 S.t187 S.n2432 0.001
R14155 S.t187 S.n2429 0.001
R14156 S.n2429 S.n2426 0.001
R14157 S.t259 S.n1953 0.001
R14158 S.n1950 S.n1936 0.001
R14159 S.t175 S.n1576 0.001
R14160 S.t175 S.n1573 0.001
R14161 S.n1573 S.n1570 0.001
R14162 S.t72 S.n1140 0.001
R14163 S.t72 S.n1137 0.001
R14164 S.n1137 S.n1134 0.001
R14165 S.t244 S.n638 0.001
R14166 S.t244 S.n635 0.001
R14167 S.n635 S.n632 0.001
R14168 S.t244 S.n621 0.001
R14169 S.t244 S.n618 0.001
R14170 S.n618 S.n615 0.001
R14171 S.t159 S.n314 0.001
R14172 S.t159 S.n311 0.001
R14173 S.n311 S.n308 0.001
R14174 S.t72 S.n1052 0.001
R14175 S.t72 S.n1049 0.001
R14176 S.n1049 S.n1046 0.001
R14177 S.t84 S.n3114 0.001
R14178 S.t84 S.n3117 0.001
R14179 S.t187 S.n2379 0.001
R14180 S.t187 S.n2376 0.001
R14181 S.n2376 S.n2373 0.001
R14182 S.t259 S.n1863 0.001
R14183 S.t259 S.n1860 0.001
R14184 S.n1860 S.n1857 0.001
R14185 S.t175 S.n1523 0.001
R14186 S.t175 S.n1520 0.001
R14187 S.n1520 S.n1517 0.001
R14188 S.t159 S.n337 0.001
R14189 S.t159 S.n334 0.001
R14190 S.n334 S.n331 0.001
R14191 S.t53 S.n3931 0.001
R14192 S.t53 S.n3934 0.001
R14193 S.t38 S.n3160 0.001
R14194 S.t38 S.n3157 0.001
R14195 S.n3157 S.n3154 0.001
R14196 S.t84 S.n2729 0.001
R14197 S.t84 S.n2726 0.001
R14198 S.n2726 S.n2723 0.001
R14199 S.t187 S.n2396 0.001
R14200 S.t187 S.n2393 0.001
R14201 S.n2393 S.n2390 0.001
R14202 S.t259 S.n1892 0.001
R14203 S.t259 S.n1889 0.001
R14204 S.n1889 S.n1886 0.001
R14205 S.t175 S.n1540 0.001
R14206 S.t175 S.n1537 0.001
R14207 S.n1537 S.n1534 0.001
R14208 S.t72 S.n1081 0.001
R14209 S.t72 S.n1078 0.001
R14210 S.n1078 S.n1075 0.001
R14211 S.t244 S.n605 0.001
R14212 S.t244 S.n602 0.001
R14213 S.n602 S.n599 0.001
R14214 S.t244 S.n588 0.001
R14215 S.t244 S.n585 0.001
R14216 S.n585 S.n582 0.001
R14217 S.t159 S.n270 0.001
R14218 S.t159 S.n267 0.001
R14219 S.n267 S.n264 0.001
R14220 S.t72 S.n1458 0.001
R14221 S.t72 S.n1461 0.001
R14222 S.t159 S.n293 0.001
R14223 S.t159 S.n290 0.001
R14224 S.n290 S.n287 0.001
R14225 S.t259 S.n2284 0.001
R14226 S.t259 S.n2287 0.001
R14227 S.t175 S.n1504 0.001
R14228 S.t175 S.n1501 0.001
R14229 S.n1501 S.n1498 0.001
R14230 S.t72 S.n1022 0.001
R14231 S.t72 S.n1019 0.001
R14232 S.n1019 S.n1016 0.001
R14233 S.t244 S.n572 0.001
R14234 S.t244 S.n569 0.001
R14235 S.n569 S.n566 0.001
R14236 S.t244 S.n555 0.001
R14237 S.t244 S.n552 0.001
R14238 S.n552 S.n549 0.001
R14239 S.n959 S.t159 0.001
R14240 S.n980 S.n961 0.001
R14241 S.t244 S.n808 0.001
R14242 S.t244 S.n811 0.001
R14243 S.t72 S.n1811 0.001
R14244 S.t72 S.n1814 0.001
R14245 S.n1788 S.t175 0.001
R14246 S.n1798 S.n1791 0.001
R14247 S.t259 S.n2321 0.001
R14248 S.t259 S.n2324 0.001
R14249 S.n2304 S.n2297 0.001
R14250 S.t84 S.n3449 0.001
R14251 S.t84 S.n3452 0.001
R14252 S.n3422 S.t38 0.001
R14253 S.n3432 S.n3425 0.001
R14254 S.t53 S.n3968 0.001
R14255 S.t53 S.n3971 0.001
R14256 S.n3951 S.n3944 0.001
R14257 S.t33 S.n4763 0.001
R14258 S.t33 S.n4766 0.001
R14259 S.n4746 S.n4739 0.001
R14260 S.t109 S.n5545 0.001
R14261 S.t109 S.n5548 0.001
R14262 S.n5528 S.n5521 0.001
R14263 S.t69 S.n6305 0.001
R14264 S.t69 S.n6308 0.001
R14265 S.n6288 S.n6281 0.001
R14266 S.t130 S.n7052 0.001
R14267 S.t130 S.n7055 0.001
R14268 S.n7035 S.n7028 0.001
R14269 S.t27 S.n8063 0.001
R14270 S.t27 S.n8066 0.001
R14271 S.n8036 S.t11 0.001
R14272 S.n8046 S.n8039 0.001
R14273 S.t300 S.n8775 0.001
R14274 S.t300 S.n8778 0.001
R14275 S.n8748 S.t40 0.001
R14276 S.n8758 S.n8751 0.001
R14277 S.t31 S.n9179 0.001
R14278 S.t31 S.n9182 0.001
R14279 S.n9162 S.n9155 0.001
R14280 S.t61 S.n9856 0.001
R14281 S.t61 S.n9859 0.001
R14282 S.n9839 S.n9832 0.001
R14283 S.t35 S.n10514 0.001
R14284 S.t35 S.n10517 0.001
R14285 S.n10497 S.n10490 0.001
R14286 S.t115 S.n11142 0.001
R14287 S.t115 S.n11145 0.001
R14288 S.n11125 S.n11118 0.001
R14289 S.t157 S.n12070 0.001
R14290 S.t157 S.n12073 0.001
R14291 S.t106 S.n12347 0.001
R14292 S.t106 S.n12350 0.001
R14293 S.t65 S.n11876 0.001
R14294 S.t65 S.n11873 0.001
R14295 S.n11873 S.n11870 0.001
R14296 S.n11869 S.n11868 0.001
R14297 S.n12343 S.n12342 0.001
R14298 S.n12066 S.n12065 0.001
R14299 S.n11124 S.n11123 0.001
R14300 S.n11138 S.n11137 0.001
R14301 S.n10496 S.n10495 0.001
R14302 S.n10510 S.n10509 0.001
R14303 S.n9838 S.n9837 0.001
R14304 S.n9852 S.n9851 0.001
R14305 S.n9161 S.n9160 0.001
R14306 S.n9175 S.n9174 0.001
R14307 S.n8757 S.n8756 0.001
R14308 S.n8771 S.n8770 0.001
R14309 S.n8045 S.n8044 0.001
R14310 S.n8059 S.n8058 0.001
R14311 S.n7034 S.n7033 0.001
R14312 S.n7048 S.n7047 0.001
R14313 S.n6287 S.n6286 0.001
R14314 S.n6301 S.n6300 0.001
R14315 S.n5527 S.n5526 0.001
R14316 S.n5541 S.n5540 0.001
R14317 S.n4745 S.n4744 0.001
R14318 S.n4759 S.n4758 0.001
R14319 S.n3950 S.n3949 0.001
R14320 S.n3964 S.n3963 0.001
R14321 S.n3431 S.n3430 0.001
R14322 S.n3445 S.n3444 0.001
R14323 S.n2303 S.n2302 0.001
R14324 S.n2317 S.n2316 0.001
R14325 S.n1797 S.n1796 0.001
R14326 S.n1817 S.t72 0.001
R14327 S.n1826 S.n1819 0.001
R14328 S.t175 S.n1782 0.001
R14329 S.t175 S.n1785 0.001
R14330 S.t259 S.n2654 0.001
R14331 S.t259 S.n2657 0.001
R14332 S.t65 S.n11858 0.001
R14333 S.t65 S.n11855 0.001
R14334 S.n11855 S.n11852 0.001
R14335 S.t106 S.n12362 0.001
R14336 S.t106 S.n12365 0.001
R14337 S.t157 S.n12086 0.001
R14338 S.t157 S.n12089 0.001
R14339 S.n11168 S.n11161 0.001
R14340 S.t115 S.n11173 0.001
R14341 S.t115 S.n11176 0.001
R14342 S.n10540 S.n10533 0.001
R14343 S.t35 S.n10545 0.001
R14344 S.t35 S.n10548 0.001
R14345 S.n9882 S.n9875 0.001
R14346 S.t61 S.n9887 0.001
R14347 S.t61 S.n9890 0.001
R14348 S.n9205 S.n9198 0.001
R14349 S.t31 S.n9210 0.001
R14350 S.t31 S.n9213 0.001
R14351 S.n8801 S.n8794 0.001
R14352 S.t300 S.n8806 0.001
R14353 S.t300 S.n8809 0.001
R14354 S.n8089 S.n8082 0.001
R14355 S.t27 S.n8094 0.001
R14356 S.t27 S.n8097 0.001
R14357 S.n7078 S.n7071 0.001
R14358 S.t130 S.n7083 0.001
R14359 S.t130 S.n7086 0.001
R14360 S.n6331 S.n6324 0.001
R14361 S.t69 S.n6336 0.001
R14362 S.t69 S.n6339 0.001
R14363 S.n5571 S.n5564 0.001
R14364 S.t109 S.n5576 0.001
R14365 S.t109 S.n5579 0.001
R14366 S.n4789 S.n4782 0.001
R14367 S.t33 S.n4794 0.001
R14368 S.t33 S.n4797 0.001
R14369 S.n3994 S.n3987 0.001
R14370 S.t53 S.n3999 0.001
R14371 S.t53 S.n4002 0.001
R14372 S.n3475 S.n3468 0.001
R14373 S.t84 S.n3480 0.001
R14374 S.t84 S.n3483 0.001
R14375 S.n2643 S.t187 0.001
R14376 S.n2650 S.n2643 0.001
R14377 S.n2660 S.t259 0.001
R14378 S.n2696 S.n2662 0.001
R14379 S.t187 S.n2637 0.001
R14380 S.t187 S.n2640 0.001
R14381 S.t84 S.n3495 0.001
R14382 S.t84 S.n3498 0.001
R14383 S.t65 S.n11843 0.001
R14384 S.t65 S.n11840 0.001
R14385 S.n11840 S.n11837 0.001
R14386 S.t106 S.n12378 0.001
R14387 S.t106 S.n12381 0.001
R14388 S.t157 S.n12101 0.001
R14389 S.t157 S.n12104 0.001
R14390 S.t47 S.n11420 0.001
R14391 S.t47 S.n11423 0.001
R14392 S.t115 S.n11188 0.001
R14393 S.t115 S.n11191 0.001
R14394 S.t144 S.n10804 0.001
R14395 S.t144 S.n10807 0.001
R14396 S.t35 S.n10560 0.001
R14397 S.t35 S.n10563 0.001
R14398 S.t124 S.n10154 0.001
R14399 S.t124 S.n10157 0.001
R14400 S.t61 S.n9902 0.001
R14401 S.t61 S.n9905 0.001
R14402 S.t225 S.n9478 0.001
R14403 S.t225 S.n9481 0.001
R14404 S.t31 S.n9225 0.001
R14405 S.t31 S.n9228 0.001
R14406 S.t40 S.n8611 0.001
R14407 S.t40 S.n8614 0.001
R14408 S.t300 S.n8821 0.001
R14409 S.t300 S.n8824 0.001
R14410 S.t11 S.n7915 0.001
R14411 S.t11 S.n7918 0.001
R14412 S.t27 S.n8109 0.001
R14413 S.t27 S.n8112 0.001
R14414 S.t102 S.n7362 0.001
R14415 S.t102 S.n7365 0.001
R14416 S.t130 S.n7098 0.001
R14417 S.t130 S.n7101 0.001
R14418 S.t4 S.n6616 0.001
R14419 S.t4 S.n6619 0.001
R14420 S.t69 S.n6351 0.001
R14421 S.t69 S.n6354 0.001
R14422 S.t25 S.n5861 0.001
R14423 S.t25 S.n5864 0.001
R14424 S.t109 S.n5591 0.001
R14425 S.t109 S.n5594 0.001
R14426 S.t77 S.n5080 0.001
R14427 S.t77 S.n5083 0.001
R14428 S.t33 S.n4809 0.001
R14429 S.t33 S.n4812 0.001
R14430 S.t94 S.n4281 0.001
R14431 S.t94 S.n4284 0.001
R14432 S.t53 S.n4014 0.001
R14433 S.t53 S.n4017 0.001
R14434 S.t38 S.n3396 0.001
R14435 S.t38 S.n3399 0.001
R14436 S.t65 S.n11828 0.001
R14437 S.t65 S.n11825 0.001
R14438 S.n11825 S.n11822 0.001
R14439 S.t106 S.n12394 0.001
R14440 S.t106 S.n12397 0.001
R14441 S.t157 S.n12116 0.001
R14442 S.t157 S.n12119 0.001
R14443 S.t47 S.n11436 0.001
R14444 S.t47 S.n11439 0.001
R14445 S.t115 S.n11203 0.001
R14446 S.t115 S.n11206 0.001
R14447 S.t144 S.n10820 0.001
R14448 S.t144 S.n10823 0.001
R14449 S.t35 S.n10575 0.001
R14450 S.t35 S.n10578 0.001
R14451 S.t124 S.n10170 0.001
R14452 S.t124 S.n10173 0.001
R14453 S.t61 S.n9917 0.001
R14454 S.t61 S.n9920 0.001
R14455 S.t225 S.n9494 0.001
R14456 S.t225 S.n9497 0.001
R14457 S.t31 S.n9240 0.001
R14458 S.t31 S.n9243 0.001
R14459 S.t40 S.n8627 0.001
R14460 S.t40 S.n8630 0.001
R14461 S.t300 S.n8836 0.001
R14462 S.t300 S.n8839 0.001
R14463 S.t11 S.n7931 0.001
R14464 S.t11 S.n7934 0.001
R14465 S.t27 S.n8124 0.001
R14466 S.t27 S.n8127 0.001
R14467 S.t102 S.n7378 0.001
R14468 S.t102 S.n7381 0.001
R14469 S.t130 S.n7113 0.001
R14470 S.t130 S.n7116 0.001
R14471 S.t4 S.n6632 0.001
R14472 S.t4 S.n6635 0.001
R14473 S.t69 S.n6366 0.001
R14474 S.t69 S.n6369 0.001
R14475 S.t25 S.n5877 0.001
R14476 S.t25 S.n5880 0.001
R14477 S.t109 S.n5606 0.001
R14478 S.t109 S.n5609 0.001
R14479 S.t77 S.n5096 0.001
R14480 S.t77 S.n5099 0.001
R14481 S.t33 S.n4824 0.001
R14482 S.t33 S.n4827 0.001
R14483 S.n4307 S.t94 0.001
R14484 S.n4315 S.n4310 0.001
R14485 S.t53 S.n4327 0.001
R14486 S.t53 S.n4330 0.001
R14487 S.t38 S.n3416 0.001
R14488 S.t38 S.n3419 0.001
R14489 S.n3501 S.t84 0.001
R14490 S.n3537 S.n3503 0.001
R14491 S.n4333 S.t53 0.001
R14492 S.n4369 S.n4335 0.001
R14493 S.t94 S.n4301 0.001
R14494 S.t94 S.n4304 0.001
R14495 S.t33 S.n5133 0.001
R14496 S.t33 S.n5136 0.001
R14497 S.t65 S.n11813 0.001
R14498 S.t65 S.n11810 0.001
R14499 S.n11810 S.n11807 0.001
R14500 S.t106 S.n12410 0.001
R14501 S.t106 S.n12413 0.001
R14502 S.t157 S.n12131 0.001
R14503 S.t157 S.n12134 0.001
R14504 S.t47 S.n11452 0.001
R14505 S.t47 S.n11455 0.001
R14506 S.t115 S.n11218 0.001
R14507 S.t115 S.n11221 0.001
R14508 S.t144 S.n10836 0.001
R14509 S.t144 S.n10839 0.001
R14510 S.t35 S.n10590 0.001
R14511 S.t35 S.n10593 0.001
R14512 S.t124 S.n10186 0.001
R14513 S.t124 S.n10189 0.001
R14514 S.t61 S.n9932 0.001
R14515 S.t61 S.n9935 0.001
R14516 S.t225 S.n9510 0.001
R14517 S.t225 S.n9513 0.001
R14518 S.t31 S.n9255 0.001
R14519 S.t31 S.n9258 0.001
R14520 S.t40 S.n8643 0.001
R14521 S.t40 S.n8646 0.001
R14522 S.t300 S.n8851 0.001
R14523 S.t300 S.n8854 0.001
R14524 S.t11 S.n7947 0.001
R14525 S.t11 S.n7950 0.001
R14526 S.t27 S.n8139 0.001
R14527 S.t27 S.n8142 0.001
R14528 S.t102 S.n7394 0.001
R14529 S.t102 S.n7397 0.001
R14530 S.t130 S.n7128 0.001
R14531 S.t130 S.n7131 0.001
R14532 S.t4 S.n6648 0.001
R14533 S.t4 S.n6651 0.001
R14534 S.t69 S.n6381 0.001
R14535 S.t69 S.n6384 0.001
R14536 S.t25 S.n5893 0.001
R14537 S.t25 S.n5896 0.001
R14538 S.t109 S.n5621 0.001
R14539 S.t109 S.n5624 0.001
R14540 S.n5122 S.t77 0.001
R14541 S.n5129 S.n5122 0.001
R14542 S.n5139 S.t33 0.001
R14543 S.n5175 S.n5141 0.001
R14544 S.t77 S.n5116 0.001
R14545 S.t77 S.n5119 0.001
R14546 S.t109 S.n5930 0.001
R14547 S.t109 S.n5933 0.001
R14548 S.t65 S.n11798 0.001
R14549 S.t65 S.n11795 0.001
R14550 S.n11795 S.n11792 0.001
R14551 S.t106 S.n12426 0.001
R14552 S.t106 S.n12429 0.001
R14553 S.t157 S.n12146 0.001
R14554 S.t157 S.n12149 0.001
R14555 S.t47 S.n11468 0.001
R14556 S.t47 S.n11471 0.001
R14557 S.t115 S.n11233 0.001
R14558 S.t115 S.n11236 0.001
R14559 S.t144 S.n10852 0.001
R14560 S.t144 S.n10855 0.001
R14561 S.t35 S.n10605 0.001
R14562 S.t35 S.n10608 0.001
R14563 S.t124 S.n10202 0.001
R14564 S.t124 S.n10205 0.001
R14565 S.t61 S.n9947 0.001
R14566 S.t61 S.n9950 0.001
R14567 S.t225 S.n9526 0.001
R14568 S.t225 S.n9529 0.001
R14569 S.t31 S.n9270 0.001
R14570 S.t31 S.n9273 0.001
R14571 S.t40 S.n8659 0.001
R14572 S.t40 S.n8662 0.001
R14573 S.t300 S.n8866 0.001
R14574 S.t300 S.n8869 0.001
R14575 S.t11 S.n7963 0.001
R14576 S.t11 S.n7966 0.001
R14577 S.t27 S.n8154 0.001
R14578 S.t27 S.n8157 0.001
R14579 S.t102 S.n7410 0.001
R14580 S.t102 S.n7413 0.001
R14581 S.t130 S.n7143 0.001
R14582 S.t130 S.n7146 0.001
R14583 S.t4 S.n6664 0.001
R14584 S.t4 S.n6667 0.001
R14585 S.t69 S.n6396 0.001
R14586 S.t69 S.n6399 0.001
R14587 S.n5919 S.t25 0.001
R14588 S.n5926 S.n5919 0.001
R14589 S.n5936 S.t109 0.001
R14590 S.n5972 S.n5938 0.001
R14591 S.t25 S.n5913 0.001
R14592 S.t25 S.n5916 0.001
R14593 S.t69 S.n6701 0.001
R14594 S.t69 S.n6704 0.001
R14595 S.t65 S.n11783 0.001
R14596 S.t65 S.n11780 0.001
R14597 S.n11780 S.n11777 0.001
R14598 S.t106 S.n12442 0.001
R14599 S.t106 S.n12445 0.001
R14600 S.t157 S.n12161 0.001
R14601 S.t157 S.n12164 0.001
R14602 S.t47 S.n11484 0.001
R14603 S.t47 S.n11487 0.001
R14604 S.t115 S.n11248 0.001
R14605 S.t115 S.n11251 0.001
R14606 S.t144 S.n10868 0.001
R14607 S.t144 S.n10871 0.001
R14608 S.t35 S.n10620 0.001
R14609 S.t35 S.n10623 0.001
R14610 S.t124 S.n10218 0.001
R14611 S.t124 S.n10221 0.001
R14612 S.t61 S.n9962 0.001
R14613 S.t61 S.n9965 0.001
R14614 S.t225 S.n9542 0.001
R14615 S.t225 S.n9545 0.001
R14616 S.t31 S.n9285 0.001
R14617 S.t31 S.n9288 0.001
R14618 S.t40 S.n8675 0.001
R14619 S.t40 S.n8678 0.001
R14620 S.t300 S.n8881 0.001
R14621 S.t300 S.n8884 0.001
R14622 S.t11 S.n7979 0.001
R14623 S.t11 S.n7982 0.001
R14624 S.t27 S.n8169 0.001
R14625 S.t27 S.n8172 0.001
R14626 S.t102 S.n7426 0.001
R14627 S.t102 S.n7429 0.001
R14628 S.t130 S.n7158 0.001
R14629 S.t130 S.n7161 0.001
R14630 S.n6690 S.t4 0.001
R14631 S.n6697 S.n6690 0.001
R14632 S.n6707 S.t69 0.001
R14633 S.n6743 S.n6709 0.001
R14634 S.t4 S.n6684 0.001
R14635 S.t4 S.n6687 0.001
R14636 S.t130 S.n7463 0.001
R14637 S.t130 S.n7466 0.001
R14638 S.t65 S.n11768 0.001
R14639 S.t65 S.n11765 0.001
R14640 S.n11765 S.n11762 0.001
R14641 S.t106 S.n12458 0.001
R14642 S.t106 S.n12461 0.001
R14643 S.t157 S.n12176 0.001
R14644 S.t157 S.n12179 0.001
R14645 S.t47 S.n11500 0.001
R14646 S.t47 S.n11503 0.001
R14647 S.t115 S.n11263 0.001
R14648 S.t115 S.n11266 0.001
R14649 S.t144 S.n10884 0.001
R14650 S.t144 S.n10887 0.001
R14651 S.t35 S.n10635 0.001
R14652 S.t35 S.n10638 0.001
R14653 S.t124 S.n10234 0.001
R14654 S.t124 S.n10237 0.001
R14655 S.t61 S.n9977 0.001
R14656 S.t61 S.n9980 0.001
R14657 S.t225 S.n9558 0.001
R14658 S.t225 S.n9561 0.001
R14659 S.t31 S.n9300 0.001
R14660 S.t31 S.n9303 0.001
R14661 S.t40 S.n8691 0.001
R14662 S.t40 S.n8694 0.001
R14663 S.t300 S.n8896 0.001
R14664 S.t300 S.n8899 0.001
R14665 S.t11 S.n7995 0.001
R14666 S.t11 S.n7998 0.001
R14667 S.t27 S.n8184 0.001
R14668 S.t27 S.n8187 0.001
R14669 S.n7452 S.t102 0.001
R14670 S.n7459 S.n7452 0.001
R14671 S.n7469 S.t130 0.001
R14672 S.n7505 S.n7471 0.001
R14673 S.t102 S.n7446 0.001
R14674 S.t102 S.n7449 0.001
R14675 S.t27 S.n8199 0.001
R14676 S.t27 S.n8202 0.001
R14677 S.t65 S.n11753 0.001
R14678 S.t65 S.n11750 0.001
R14679 S.n11750 S.n11747 0.001
R14680 S.t106 S.n12474 0.001
R14681 S.t106 S.n12477 0.001
R14682 S.t157 S.n12191 0.001
R14683 S.t157 S.n12194 0.001
R14684 S.t47 S.n11516 0.001
R14685 S.t47 S.n11519 0.001
R14686 S.t115 S.n11278 0.001
R14687 S.t115 S.n11281 0.001
R14688 S.t144 S.n10900 0.001
R14689 S.t144 S.n10903 0.001
R14690 S.t35 S.n10650 0.001
R14691 S.t35 S.n10653 0.001
R14692 S.t124 S.n10250 0.001
R14693 S.t124 S.n10253 0.001
R14694 S.t61 S.n9992 0.001
R14695 S.t61 S.n9995 0.001
R14696 S.t225 S.n9574 0.001
R14697 S.t225 S.n9577 0.001
R14698 S.t31 S.n9315 0.001
R14699 S.t31 S.n9318 0.001
R14700 S.t40 S.n8707 0.001
R14701 S.t40 S.n8710 0.001
R14702 S.t300 S.n8911 0.001
R14703 S.t300 S.n8914 0.001
R14704 S.t11 S.n8010 0.001
R14705 S.t11 S.n8013 0.001
R14706 S.n8205 S.t27 0.001
R14707 S.n8241 S.n8207 0.001
R14708 S.t11 S.n8030 0.001
R14709 S.t11 S.n8033 0.001
R14710 S.t300 S.n8926 0.001
R14711 S.t300 S.n8929 0.001
R14712 S.t65 S.n11738 0.001
R14713 S.t65 S.n11735 0.001
R14714 S.n11735 S.n11732 0.001
R14715 S.t106 S.n12490 0.001
R14716 S.t106 S.n12493 0.001
R14717 S.t157 S.n12206 0.001
R14718 S.t157 S.n12209 0.001
R14719 S.t47 S.n11532 0.001
R14720 S.t47 S.n11535 0.001
R14721 S.t115 S.n11293 0.001
R14722 S.t115 S.n11296 0.001
R14723 S.t144 S.n10916 0.001
R14724 S.t144 S.n10919 0.001
R14725 S.t35 S.n10665 0.001
R14726 S.t35 S.n10668 0.001
R14727 S.t124 S.n10266 0.001
R14728 S.t124 S.n10269 0.001
R14729 S.t61 S.n10007 0.001
R14730 S.t61 S.n10010 0.001
R14731 S.t225 S.n9590 0.001
R14732 S.t225 S.n9593 0.001
R14733 S.t31 S.n9330 0.001
R14734 S.t31 S.n9333 0.001
R14735 S.t40 S.n8722 0.001
R14736 S.t40 S.n8725 0.001
R14737 S.n8932 S.t300 0.001
R14738 S.n8968 S.n8934 0.001
R14739 S.t40 S.n8742 0.001
R14740 S.t40 S.n8745 0.001
R14741 S.t31 S.n9627 0.001
R14742 S.t31 S.n9630 0.001
R14743 S.t65 S.n11723 0.001
R14744 S.t65 S.n11720 0.001
R14745 S.n11720 S.n11717 0.001
R14746 S.t106 S.n12506 0.001
R14747 S.t106 S.n12509 0.001
R14748 S.t157 S.n12221 0.001
R14749 S.t157 S.n12224 0.001
R14750 S.t47 S.n11548 0.001
R14751 S.t47 S.n11551 0.001
R14752 S.t115 S.n11308 0.001
R14753 S.t115 S.n11311 0.001
R14754 S.t144 S.n10932 0.001
R14755 S.t144 S.n10935 0.001
R14756 S.t35 S.n10680 0.001
R14757 S.t35 S.n10683 0.001
R14758 S.t124 S.n10282 0.001
R14759 S.t124 S.n10285 0.001
R14760 S.t61 S.n10022 0.001
R14761 S.t61 S.n10025 0.001
R14762 S.n9616 S.t225 0.001
R14763 S.n9623 S.n9616 0.001
R14764 S.n9633 S.t31 0.001
R14765 S.n9669 S.n9635 0.001
R14766 S.t225 S.n9610 0.001
R14767 S.t225 S.n9613 0.001
R14768 S.t61 S.n10319 0.001
R14769 S.t61 S.n10322 0.001
R14770 S.t65 S.n11708 0.001
R14771 S.t65 S.n11705 0.001
R14772 S.n11705 S.n11702 0.001
R14773 S.t106 S.n12522 0.001
R14774 S.t106 S.n12525 0.001
R14775 S.t157 S.n12236 0.001
R14776 S.t157 S.n12239 0.001
R14777 S.t47 S.n11564 0.001
R14778 S.t47 S.n11567 0.001
R14779 S.t115 S.n11323 0.001
R14780 S.t115 S.n11326 0.001
R14781 S.t144 S.n10948 0.001
R14782 S.t144 S.n10951 0.001
R14783 S.t35 S.n10695 0.001
R14784 S.t35 S.n10698 0.001
R14785 S.n10308 S.t124 0.001
R14786 S.n10315 S.n10308 0.001
R14787 S.n10325 S.t61 0.001
R14788 S.n10361 S.n10327 0.001
R14789 S.t124 S.n10302 0.001
R14790 S.t124 S.n10305 0.001
R14791 S.t35 S.n10985 0.001
R14792 S.t35 S.n10988 0.001
R14793 S.t65 S.n11693 0.001
R14794 S.t65 S.n11690 0.001
R14795 S.n11690 S.n11687 0.001
R14796 S.t106 S.n12538 0.001
R14797 S.t106 S.n12541 0.001
R14798 S.t157 S.n12251 0.001
R14799 S.t157 S.n12254 0.001
R14800 S.t47 S.n11580 0.001
R14801 S.t47 S.n11583 0.001
R14802 S.t115 S.n11338 0.001
R14803 S.t115 S.n11341 0.001
R14804 S.n10974 S.t144 0.001
R14805 S.n10981 S.n10974 0.001
R14806 S.n10991 S.t35 0.001
R14807 S.n11025 S.n10993 0.001
R14808 S.t144 S.n10968 0.001
R14809 S.t144 S.n10971 0.001
R14810 S.t115 S.n11620 0.001
R14811 S.t115 S.n11623 0.001
R14812 S.t65 S.n11678 0.001
R14813 S.t65 S.n11675 0.001
R14814 S.n11675 S.n11672 0.001
R14815 S.t106 S.n12554 0.001
R14816 S.t106 S.n12557 0.001
R14817 S.t157 S.n12266 0.001
R14818 S.t157 S.n12269 0.001
R14819 S.n11609 S.t47 0.001
R14820 S.n11616 S.n11609 0.001
R14821 S.n11626 S.t115 0.001
R14822 S.n11644 S.n11628 0.001
R14823 S.t47 S.n11603 0.001
R14824 S.t47 S.n11606 0.001
R14825 S.t157 S.n12585 0.001
R14826 S.t157 S.n12588 0.001
R14827 S.t65 S.n11663 0.001
R14828 S.t65 S.n11660 0.001
R14829 S.n11660 S.n11657 0.001
R14830 S.n12560 S.t106 0.001
R14831 S.n12568 S.n12563 0.001
R14832 S.n63 S.n62 0.001
R14833 S.n67 S.n66 0.001
R14834 S.n977 S.n976 0.001
R14835 S.n990 S.n989 0.001
R14836 S.n2675 S.n2674 0.001
R14837 S.n3516 S.n3508 0.001
R14838 S.n4348 S.n4347 0.001
R14839 S.n5154 S.n5153 0.001
R14840 S.n5951 S.n5950 0.001
R14841 S.n6722 S.n6721 0.001
R14842 S.n7484 S.n7483 0.001
R14843 S.n8220 S.n8219 0.001
R14844 S.n8947 S.n8946 0.001
R14845 S.n9648 S.n9647 0.001
R14846 S.n10340 S.n10339 0.001
R14847 S.n11004 S.n11003 0.001
R14848 S.n11638 S.n11637 0.001
R14849 S.n11914 S.n11911 0.001
R14850 S.n12611 S.n12591 0.001
R14851 S.n12050 S.n12047 0.001
R14852 S.n11105 S.n11102 0.001
R14853 S.n822 S.n814 0.001
R14854 S.n10477 S.n10474 0.001
R14855 S.n9819 S.n9816 0.001
R14856 S.n9142 S.n9139 0.001
R14857 S.n8452 S.n8449 0.001
R14858 S.n466 S.n461 0.001
R14859 S.n7740 S.n7737 0.001
R14860 S.n7015 S.n7012 0.001
R14861 S.n6268 S.n6265 0.001
R14862 S.n5508 S.n5505 0.001
R14863 S.n1953 S.n1950 0.001
R14864 S.n4726 S.n4723 0.001
R14865 S.n3931 S.n3928 0.001
R14866 S.n3114 S.n3111 0.001
R14867 S.n2284 S.n2281 0.001
R14868 S.n1458 S.n1455 0.001
R14869 S.n953 S.n950 0.001
R14870 S.n980 S.n959 0.001
R14871 S.n12347 S.n12344 0.001
R14872 S.n12070 S.n12067 0.001
R14873 S.n11125 S.n11115 0.001
R14874 S.n11142 S.n11139 0.001
R14875 S.n10497 S.n10487 0.001
R14876 S.n10514 S.n10511 0.001
R14877 S.n9839 S.n9829 0.001
R14878 S.n9856 S.n9853 0.001
R14879 S.n9162 S.n9152 0.001
R14880 S.n9179 S.n9176 0.001
R14881 S.n8758 S.n8748 0.001
R14882 S.n8775 S.n8772 0.001
R14883 S.n8046 S.n8036 0.001
R14884 S.n8063 S.n8060 0.001
R14885 S.n7035 S.n7025 0.001
R14886 S.n7052 S.n7049 0.001
R14887 S.n6288 S.n6278 0.001
R14888 S.n6305 S.n6302 0.001
R14889 S.n5528 S.n5518 0.001
R14890 S.n5545 S.n5542 0.001
R14891 S.n4746 S.n4736 0.001
R14892 S.n4763 S.n4760 0.001
R14893 S.n3951 S.n3941 0.001
R14894 S.n3968 S.n3965 0.001
R14895 S.n3432 S.n3422 0.001
R14896 S.n3449 S.n3446 0.001
R14897 S.n2304 S.n2294 0.001
R14898 S.n2321 S.n2318 0.001
R14899 S.n1798 S.n1788 0.001
R14900 S.n1811 S.n1808 0.001
R14901 S.n808 S.n805 0.001
R14902 S.n1826 S.n1817 0.001
R14903 S.n12362 S.n12359 0.001
R14904 S.n12086 S.n12083 0.001
R14905 S.n11168 S.n11164 0.001
R14906 S.n11173 S.n11170 0.001
R14907 S.n10540 S.n10536 0.001
R14908 S.n10545 S.n10542 0.001
R14909 S.n9882 S.n9878 0.001
R14910 S.n9887 S.n9884 0.001
R14911 S.n9205 S.n9201 0.001
R14912 S.n9210 S.n9207 0.001
R14913 S.n8801 S.n8797 0.001
R14914 S.n8806 S.n8803 0.001
R14915 S.n8089 S.n8085 0.001
R14916 S.n8094 S.n8091 0.001
R14917 S.n7078 S.n7074 0.001
R14918 S.n7083 S.n7080 0.001
R14919 S.n6331 S.n6327 0.001
R14920 S.n6336 S.n6333 0.001
R14921 S.n5571 S.n5567 0.001
R14922 S.n5576 S.n5573 0.001
R14923 S.n4789 S.n4785 0.001
R14924 S.n4794 S.n4791 0.001
R14925 S.n3994 S.n3990 0.001
R14926 S.n3999 S.n3996 0.001
R14927 S.n3475 S.n3471 0.001
R14928 S.n3480 S.n3477 0.001
R14929 S.n2650 S.n2646 0.001
R14930 S.n2654 S.n2651 0.001
R14931 S.n1782 S.n1779 0.001
R14932 S.n2696 S.n2660 0.001
R14933 S.n2637 S.n2634 0.001
R14934 S.n3495 S.n3492 0.001
R14935 S.n3396 S.n3393 0.001
R14936 S.n4014 S.n4011 0.001
R14937 S.n4281 S.n4278 0.001
R14938 S.n4809 S.n4806 0.001
R14939 S.n5080 S.n5077 0.001
R14940 S.n5591 S.n5588 0.001
R14941 S.n5861 S.n5858 0.001
R14942 S.n6351 S.n6348 0.001
R14943 S.n6616 S.n6613 0.001
R14944 S.n7098 S.n7095 0.001
R14945 S.n7362 S.n7359 0.001
R14946 S.n8109 S.n8106 0.001
R14947 S.n7915 S.n7912 0.001
R14948 S.n8821 S.n8818 0.001
R14949 S.n8611 S.n8608 0.001
R14950 S.n9225 S.n9222 0.001
R14951 S.n9478 S.n9475 0.001
R14952 S.n9902 S.n9899 0.001
R14953 S.n10154 S.n10151 0.001
R14954 S.n10560 S.n10557 0.001
R14955 S.n10804 S.n10801 0.001
R14956 S.n11188 S.n11185 0.001
R14957 S.n11420 S.n11417 0.001
R14958 S.n12101 S.n12098 0.001
R14959 S.n12378 S.n12375 0.001
R14960 S.n3537 S.n3501 0.001
R14961 S.n3416 S.n3413 0.001
R14962 S.n4327 S.n4324 0.001
R14963 S.n4315 S.n4307 0.001
R14964 S.n4824 S.n4821 0.001
R14965 S.n5096 S.n5093 0.001
R14966 S.n5606 S.n5603 0.001
R14967 S.n5877 S.n5874 0.001
R14968 S.n6366 S.n6363 0.001
R14969 S.n6632 S.n6629 0.001
R14970 S.n7113 S.n7110 0.001
R14971 S.n7378 S.n7375 0.001
R14972 S.n8124 S.n8121 0.001
R14973 S.n7931 S.n7928 0.001
R14974 S.n8836 S.n8833 0.001
R14975 S.n8627 S.n8624 0.001
R14976 S.n9240 S.n9237 0.001
R14977 S.n9494 S.n9491 0.001
R14978 S.n9917 S.n9914 0.001
R14979 S.n10170 S.n10167 0.001
R14980 S.n10575 S.n10572 0.001
R14981 S.n10820 S.n10817 0.001
R14982 S.n11203 S.n11200 0.001
R14983 S.n11436 S.n11433 0.001
R14984 S.n12116 S.n12113 0.001
R14985 S.n12394 S.n12391 0.001
R14986 S.n4369 S.n4333 0.001
R14987 S.n4301 S.n4298 0.001
R14988 S.n5133 S.n5130 0.001
R14989 S.n5129 S.n5125 0.001
R14990 S.n5621 S.n5618 0.001
R14991 S.n5893 S.n5890 0.001
R14992 S.n6381 S.n6378 0.001
R14993 S.n6648 S.n6645 0.001
R14994 S.n7128 S.n7125 0.001
R14995 S.n7394 S.n7391 0.001
R14996 S.n8139 S.n8136 0.001
R14997 S.n7947 S.n7944 0.001
R14998 S.n8851 S.n8848 0.001
R14999 S.n8643 S.n8640 0.001
R15000 S.n9255 S.n9252 0.001
R15001 S.n9510 S.n9507 0.001
R15002 S.n9932 S.n9929 0.001
R15003 S.n10186 S.n10183 0.001
R15004 S.n10590 S.n10587 0.001
R15005 S.n10836 S.n10833 0.001
R15006 S.n11218 S.n11215 0.001
R15007 S.n11452 S.n11449 0.001
R15008 S.n12131 S.n12128 0.001
R15009 S.n12410 S.n12407 0.001
R15010 S.n5175 S.n5139 0.001
R15011 S.n5116 S.n5113 0.001
R15012 S.n5930 S.n5927 0.001
R15013 S.n5926 S.n5922 0.001
R15014 S.n6396 S.n6393 0.001
R15015 S.n6664 S.n6661 0.001
R15016 S.n7143 S.n7140 0.001
R15017 S.n7410 S.n7407 0.001
R15018 S.n8154 S.n8151 0.001
R15019 S.n7963 S.n7960 0.001
R15020 S.n8866 S.n8863 0.001
R15021 S.n8659 S.n8656 0.001
R15022 S.n9270 S.n9267 0.001
R15023 S.n9526 S.n9523 0.001
R15024 S.n9947 S.n9944 0.001
R15025 S.n10202 S.n10199 0.001
R15026 S.n10605 S.n10602 0.001
R15027 S.n10852 S.n10849 0.001
R15028 S.n11233 S.n11230 0.001
R15029 S.n11468 S.n11465 0.001
R15030 S.n12146 S.n12143 0.001
R15031 S.n12426 S.n12423 0.001
R15032 S.n5972 S.n5936 0.001
R15033 S.n5913 S.n5910 0.001
R15034 S.n6701 S.n6698 0.001
R15035 S.n6697 S.n6693 0.001
R15036 S.n7158 S.n7155 0.001
R15037 S.n7426 S.n7423 0.001
R15038 S.n8169 S.n8166 0.001
R15039 S.n7979 S.n7976 0.001
R15040 S.n8881 S.n8878 0.001
R15041 S.n8675 S.n8672 0.001
R15042 S.n9285 S.n9282 0.001
R15043 S.n9542 S.n9539 0.001
R15044 S.n9962 S.n9959 0.001
R15045 S.n10218 S.n10215 0.001
R15046 S.n10620 S.n10617 0.001
R15047 S.n10868 S.n10865 0.001
R15048 S.n11248 S.n11245 0.001
R15049 S.n11484 S.n11481 0.001
R15050 S.n12161 S.n12158 0.001
R15051 S.n12442 S.n12439 0.001
R15052 S.n6743 S.n6707 0.001
R15053 S.n6684 S.n6681 0.001
R15054 S.n7463 S.n7460 0.001
R15055 S.n7459 S.n7455 0.001
R15056 S.n8184 S.n8181 0.001
R15057 S.n7995 S.n7992 0.001
R15058 S.n8896 S.n8893 0.001
R15059 S.n8691 S.n8688 0.001
R15060 S.n9300 S.n9297 0.001
R15061 S.n9558 S.n9555 0.001
R15062 S.n9977 S.n9974 0.001
R15063 S.n10234 S.n10231 0.001
R15064 S.n10635 S.n10632 0.001
R15065 S.n10884 S.n10881 0.001
R15066 S.n11263 S.n11260 0.001
R15067 S.n11500 S.n11497 0.001
R15068 S.n12176 S.n12173 0.001
R15069 S.n12458 S.n12455 0.001
R15070 S.n7505 S.n7469 0.001
R15071 S.n7446 S.n7443 0.001
R15072 S.n8199 S.n8196 0.001
R15073 S.n8010 S.n8007 0.001
R15074 S.n8911 S.n8908 0.001
R15075 S.n8707 S.n8704 0.001
R15076 S.n9315 S.n9312 0.001
R15077 S.n9574 S.n9571 0.001
R15078 S.n9992 S.n9989 0.001
R15079 S.n10250 S.n10247 0.001
R15080 S.n10650 S.n10647 0.001
R15081 S.n10900 S.n10897 0.001
R15082 S.n11278 S.n11275 0.001
R15083 S.n11516 S.n11513 0.001
R15084 S.n12191 S.n12188 0.001
R15085 S.n12474 S.n12471 0.001
R15086 S.n8241 S.n8205 0.001
R15087 S.n8030 S.n8027 0.001
R15088 S.n8926 S.n8923 0.001
R15089 S.n8722 S.n8719 0.001
R15090 S.n9330 S.n9327 0.001
R15091 S.n9590 S.n9587 0.001
R15092 S.n10007 S.n10004 0.001
R15093 S.n10266 S.n10263 0.001
R15094 S.n10665 S.n10662 0.001
R15095 S.n10916 S.n10913 0.001
R15096 S.n11293 S.n11290 0.001
R15097 S.n11532 S.n11529 0.001
R15098 S.n12206 S.n12203 0.001
R15099 S.n12490 S.n12487 0.001
R15100 S.n8968 S.n8932 0.001
R15101 S.n8742 S.n8739 0.001
R15102 S.n9627 S.n9624 0.001
R15103 S.n9623 S.n9619 0.001
R15104 S.n10022 S.n10019 0.001
R15105 S.n10282 S.n10279 0.001
R15106 S.n10680 S.n10677 0.001
R15107 S.n10932 S.n10929 0.001
R15108 S.n11308 S.n11305 0.001
R15109 S.n11548 S.n11545 0.001
R15110 S.n12221 S.n12218 0.001
R15111 S.n12506 S.n12503 0.001
R15112 S.n9669 S.n9633 0.001
R15113 S.n9610 S.n9607 0.001
R15114 S.n10319 S.n10316 0.001
R15115 S.n10315 S.n10311 0.001
R15116 S.n10695 S.n10692 0.001
R15117 S.n10948 S.n10945 0.001
R15118 S.n11323 S.n11320 0.001
R15119 S.n11564 S.n11561 0.001
R15120 S.n12236 S.n12233 0.001
R15121 S.n12522 S.n12519 0.001
R15122 S.n10361 S.n10325 0.001
R15123 S.n10302 S.n10299 0.001
R15124 S.n10985 S.n10982 0.001
R15125 S.n10981 S.n10977 0.001
R15126 S.n11338 S.n11335 0.001
R15127 S.n11580 S.n11577 0.001
R15128 S.n12251 S.n12248 0.001
R15129 S.n12538 S.n12535 0.001
R15130 S.n11025 S.n10991 0.001
R15131 S.n10968 S.n10965 0.001
R15132 S.n11620 S.n11617 0.001
R15133 S.n11616 S.n11612 0.001
R15134 S.n12266 S.n12263 0.001
R15135 S.n12554 S.n12551 0.001
R15136 S.n11644 S.n11626 0.001
R15137 S.n11603 S.n11600 0.001
R15138 S.n12585 S.n12582 0.001
R15139 S.n12568 S.n12560 0.001
C0 S D 4782.53fF
C1 G D 2242.34fF
C2 DNW S 5943.07fF
C3 DNW G 9.27fF
C4 S G 3017.69fF
C5 DNW D 518.88fF
C6 D VSUBS -62.04fF
C7 G VSUBS -303.14fF
C8 S VSUBS 385.63fF $ **FLOATING
C9 DNW VSUBS 11261.70fF $ **FLOATING
C10 S.n0 VSUBS 0.96fF $ **FLOATING
C11 S.n1 VSUBS 0.34fF $ **FLOATING
C12 S.n2 VSUBS 0.33fF $ **FLOATING
C13 S.n3 VSUBS 2.64fF $ **FLOATING
C14 S.n4 VSUBS 8.97fF $ **FLOATING
C15 S.n5 VSUBS 8.97fF $ **FLOATING
C16 S.n6 VSUBS 5.39fF $ **FLOATING
C17 S.n7 VSUBS 2.17fF $ **FLOATING
C18 S.n8 VSUBS 0.96fF $ **FLOATING
C19 S.n9 VSUBS 0.34fF $ **FLOATING
C20 S.n10 VSUBS 0.33fF $ **FLOATING
C21 S.n11 VSUBS 2.64fF $ **FLOATING
C22 S.n12 VSUBS 8.97fF $ **FLOATING
C23 S.n13 VSUBS 8.97fF $ **FLOATING
C24 S.n14 VSUBS 5.39fF $ **FLOATING
C25 S.n15 VSUBS 2.17fF $ **FLOATING
C26 S.n16 VSUBS 0.96fF $ **FLOATING
C27 S.n17 VSUBS 0.34fF $ **FLOATING
C28 S.n18 VSUBS 0.33fF $ **FLOATING
C29 S.n19 VSUBS 9.37fF $ **FLOATING
C30 S.n20 VSUBS 2.64fF $ **FLOATING
C31 S.n21 VSUBS 8.97fF $ **FLOATING
C32 S.n22 VSUBS 8.97fF $ **FLOATING
C33 S.n23 VSUBS 5.39fF $ **FLOATING
C34 S.n24 VSUBS 2.17fF $ **FLOATING
C35 S.n25 VSUBS 0.96fF $ **FLOATING
C36 S.n26 VSUBS 0.34fF $ **FLOATING
C37 S.n27 VSUBS 0.33fF $ **FLOATING
C38 S.n28 VSUBS 9.37fF $ **FLOATING
C39 S.n29 VSUBS 2.64fF $ **FLOATING
C40 S.n30 VSUBS 8.97fF $ **FLOATING
C41 S.n31 VSUBS 8.97fF $ **FLOATING
C42 S.n32 VSUBS 5.39fF $ **FLOATING
C43 S.n33 VSUBS 2.17fF $ **FLOATING
C44 S.n34 VSUBS 0.96fF $ **FLOATING
C45 S.n35 VSUBS 0.34fF $ **FLOATING
C46 S.n36 VSUBS 0.33fF $ **FLOATING
C47 S.n37 VSUBS 9.37fF $ **FLOATING
C48 S.n38 VSUBS 2.64fF $ **FLOATING
C49 S.n39 VSUBS 8.97fF $ **FLOATING
C50 S.n40 VSUBS 8.97fF $ **FLOATING
C51 S.n41 VSUBS 5.39fF $ **FLOATING
C52 S.n42 VSUBS 2.17fF $ **FLOATING
C53 S.n43 VSUBS 0.96fF $ **FLOATING
C54 S.n44 VSUBS 0.34fF $ **FLOATING
C55 S.n45 VSUBS 0.33fF $ **FLOATING
C56 S.n46 VSUBS 9.37fF $ **FLOATING
C57 S.n47 VSUBS 2.64fF $ **FLOATING
C58 S.n48 VSUBS 8.97fF $ **FLOATING
C59 S.n49 VSUBS 8.97fF $ **FLOATING
C60 S.n50 VSUBS 5.39fF $ **FLOATING
C61 S.n51 VSUBS 2.17fF $ **FLOATING
C62 S.n52 VSUBS 13.61fF $ **FLOATING
C63 S.n53 VSUBS 13.61fF $ **FLOATING
C64 S.n54 VSUBS 5.33fF $ **FLOATING
C65 S.n55 VSUBS 2.04fF $ **FLOATING
C66 S.n56 VSUBS 16.41fF $ **FLOATING
C67 S.n57 VSUBS 2.64fF $ **FLOATING
C68 S.n58 VSUBS 0.34fF $ **FLOATING
C69 S.n59 VSUBS 0.30fF $ **FLOATING
C70 S.n60 VSUBS 0.96fF $ **FLOATING
C71 S.t991 VSUBS 0.02fF
C72 S.n61 VSUBS 1.31fF $ **FLOATING
C73 S.n62 VSUBS 54.09fF $ **FLOATING
C74 S.n63 VSUBS 2.22fF $ **FLOATING
C75 S.n64 VSUBS 0.35fF $ **FLOATING
C76 S.n65 VSUBS 0.62fF $ **FLOATING
C77 S.n66 VSUBS 0.53fF $ **FLOATING
C78 S.n67 VSUBS 3.67fF $ **FLOATING
C79 S.n68 VSUBS 4.25fF $ **FLOATING
C80 S.n69 VSUBS 4.22fF $ **FLOATING
C81 S.n70 VSUBS 4.22fF $ **FLOATING
C82 S.n71 VSUBS 4.22fF $ **FLOATING
C83 S.n72 VSUBS 4.22fF $ **FLOATING
C84 S.n73 VSUBS 4.22fF $ **FLOATING
C85 S.n74 VSUBS 4.22fF $ **FLOATING
C86 S.n75 VSUBS 4.70fF $ **FLOATING
C87 S.n76 VSUBS 4.30fF $ **FLOATING
C88 S.n77 VSUBS 4.28fF $ **FLOATING
C89 S.n78 VSUBS 130.14fF $ **FLOATING
C90 S.n79 VSUBS 2.19fF $ **FLOATING
C91 S.n80 VSUBS 12.90fF $ **FLOATING
C92 S.n81 VSUBS 1.89fF $ **FLOATING
C93 S.n82 VSUBS 9.41fF $ **FLOATING
C94 S.n83 VSUBS 0.25fF $ **FLOATING
C95 S.t172 VSUBS 0.02fF
C96 S.n84 VSUBS 0.44fF $ **FLOATING
C97 S.n85 VSUBS 8.97fF $ **FLOATING
C98 S.n86 VSUBS 8.97fF $ **FLOATING
C99 S.n87 VSUBS 5.46fF $ **FLOATING
C100 S.n88 VSUBS 1.96fF $ **FLOATING
C101 S.t1874 VSUBS 0.02fF
C102 S.n89 VSUBS 0.89fF $ **FLOATING
C103 S.t46 VSUBS 0.02fF
C104 S.n90 VSUBS 0.89fF $ **FLOATING
C105 S.n91 VSUBS 9.43fF $ **FLOATING
C106 S.n92 VSUBS 3.28fF $ **FLOATING
C107 S.n93 VSUBS 0.38fF $ **FLOATING
C108 S.n94 VSUBS 0.31fF $ **FLOATING
C109 S.n95 VSUBS 1.00fF $ **FLOATING
C110 S.n96 VSUBS 0.02fF $ **FLOATING
C111 S.t2550 VSUBS 0.02fF
C112 S.n97 VSUBS 0.37fF $ **FLOATING
C113 S.n98 VSUBS 8.97fF $ **FLOATING
C114 S.n99 VSUBS 8.97fF $ **FLOATING
C115 S.n100 VSUBS 5.46fF $ **FLOATING
C116 S.n101 VSUBS 1.96fF $ **FLOATING
C117 S.t2263 VSUBS 0.02fF
C118 S.n102 VSUBS 0.89fF $ **FLOATING
C119 S.t610 VSUBS 0.02fF
C120 S.n103 VSUBS 0.89fF $ **FLOATING
C121 S.n104 VSUBS 9.43fF $ **FLOATING
C122 S.n105 VSUBS 3.28fF $ **FLOATING
C123 S.n106 VSUBS 0.38fF $ **FLOATING
C124 S.n107 VSUBS 0.31fF $ **FLOATING
C125 S.n108 VSUBS 1.00fF $ **FLOATING
C126 S.n109 VSUBS 0.02fF $ **FLOATING
C127 S.t561 VSUBS 0.02fF
C128 S.n110 VSUBS 0.37fF $ **FLOATING
C129 S.n111 VSUBS 8.97fF $ **FLOATING
C130 S.n112 VSUBS 8.97fF $ **FLOATING
C131 S.n113 VSUBS 5.46fF $ **FLOATING
C132 S.n114 VSUBS 1.96fF $ **FLOATING
C133 S.t1321 VSUBS 0.02fF
C134 S.n115 VSUBS 0.89fF $ **FLOATING
C135 S.t2187 VSUBS 0.02fF
C136 S.n116 VSUBS 0.89fF $ **FLOATING
C137 S.n117 VSUBS 9.43fF $ **FLOATING
C138 S.n118 VSUBS 3.28fF $ **FLOATING
C139 S.n119 VSUBS 0.38fF $ **FLOATING
C140 S.n120 VSUBS 0.31fF $ **FLOATING
C141 S.n121 VSUBS 1.00fF $ **FLOATING
C142 S.n122 VSUBS 0.02fF $ **FLOATING
C143 S.t2136 VSUBS 0.02fF
C144 S.n123 VSUBS 0.37fF $ **FLOATING
C145 S.n124 VSUBS 8.97fF $ **FLOATING
C146 S.n125 VSUBS 8.97fF $ **FLOATING
C147 S.n126 VSUBS 5.46fF $ **FLOATING
C148 S.n127 VSUBS 1.96fF $ **FLOATING
C149 S.t1847 VSUBS 0.02fF
C150 S.n128 VSUBS 0.89fF $ **FLOATING
C151 S.t1366 VSUBS 0.02fF
C152 S.n129 VSUBS 0.89fF $ **FLOATING
C153 S.n130 VSUBS 9.43fF $ **FLOATING
C154 S.n131 VSUBS 3.28fF $ **FLOATING
C155 S.n132 VSUBS 0.38fF $ **FLOATING
C156 S.n133 VSUBS 0.31fF $ **FLOATING
C157 S.n134 VSUBS 1.00fF $ **FLOATING
C158 S.n135 VSUBS 0.02fF $ **FLOATING
C159 S.t121 VSUBS 0.02fF
C160 S.n136 VSUBS 0.37fF $ **FLOATING
C161 S.n137 VSUBS 8.97fF $ **FLOATING
C162 S.n138 VSUBS 8.97fF $ **FLOATING
C163 S.n139 VSUBS 5.46fF $ **FLOATING
C164 S.n140 VSUBS 1.96fF $ **FLOATING
C165 S.t891 VSUBS 0.02fF
C166 S.n141 VSUBS 0.89fF $ **FLOATING
C167 S.t1760 VSUBS 0.02fF
C168 S.n142 VSUBS 0.89fF $ **FLOATING
C169 S.n143 VSUBS 3.28fF $ **FLOATING
C170 S.n144 VSUBS 0.38fF $ **FLOATING
C171 S.n145 VSUBS 0.31fF $ **FLOATING
C172 S.n146 VSUBS 1.00fF $ **FLOATING
C173 S.n147 VSUBS 0.02fF $ **FLOATING
C174 S.t1702 VSUBS 0.02fF
C175 S.n148 VSUBS 0.37fF $ **FLOATING
C176 S.n149 VSUBS 8.97fF $ **FLOATING
C177 S.n150 VSUBS 8.97fF $ **FLOATING
C178 S.n151 VSUBS 5.46fF $ **FLOATING
C179 S.n152 VSUBS 1.96fF $ **FLOATING
C180 S.t8 VSUBS 0.02fF
C181 S.n153 VSUBS 0.89fF $ **FLOATING
C182 S.t805 VSUBS 0.02fF
C183 S.n154 VSUBS 0.89fF $ **FLOATING
C184 S.n155 VSUBS 3.28fF $ **FLOATING
C185 S.n156 VSUBS 0.38fF $ **FLOATING
C186 S.n157 VSUBS 0.31fF $ **FLOATING
C187 S.n158 VSUBS 1.00fF $ **FLOATING
C188 S.n159 VSUBS 0.02fF $ **FLOATING
C189 S.t746 VSUBS 0.02fF
C190 S.n160 VSUBS 0.37fF $ **FLOATING
C191 S.n161 VSUBS 0.31fF $ **FLOATING
C192 S.n162 VSUBS 8.97fF $ **FLOATING
C193 S.n163 VSUBS 8.97fF $ **FLOATING
C194 S.n164 VSUBS 5.22fF $ **FLOATING
C195 S.n165 VSUBS 1.00fF $ **FLOATING
C196 S.n166 VSUBS 0.35fF $ **FLOATING
C197 S.t2160 VSUBS 0.02fF
C198 S.n167 VSUBS 0.89fF $ **FLOATING
C199 S.t506 VSUBS 0.02fF
C200 S.n168 VSUBS 0.89fF $ **FLOATING
C201 S.n169 VSUBS 3.39fF $ **FLOATING
C202 S.n170 VSUBS 0.27fF $ **FLOATING
C203 S.n171 VSUBS 1.05fF $ **FLOATING
C204 S.n172 VSUBS 1.15fF $ **FLOATING
C205 S.n173 VSUBS 0.42fF $ **FLOATING
C206 S.n174 VSUBS 0.02fF $ **FLOATING
C207 S.t1967 VSUBS 0.02fF
C208 S.n175 VSUBS 0.37fF $ **FLOATING
C209 S.n176 VSUBS 0.37fF $ **FLOATING
C210 S.n177 VSUBS 0.83fF $ **FLOATING
C211 S.t427 VSUBS 0.02fF
C212 S.n178 VSUBS 0.89fF $ **FLOATING
C213 S.t1292 VSUBS 0.02fF
C214 S.n179 VSUBS 0.89fF $ **FLOATING
C215 S.n180 VSUBS 2.64fF $ **FLOATING
C216 S.n181 VSUBS 8.97fF $ **FLOATING
C217 S.n182 VSUBS 8.97fF $ **FLOATING
C218 S.n183 VSUBS 5.76fF $ **FLOATING
C219 S.n184 VSUBS 1.77fF $ **FLOATING
C220 S.n185 VSUBS 1.13fF $ **FLOATING
C221 S.n186 VSUBS 0.00fF $ **FLOATING
C222 S.n187 VSUBS 0.39fF $ **FLOATING
C223 S.n188 VSUBS 0.02fF $ **FLOATING
C224 S.t227 VSUBS 0.02fF
C225 S.n189 VSUBS 0.37fF $ **FLOATING
C226 S.n190 VSUBS 1.62fF $ **FLOATING
C227 S.t1223 VSUBS 0.02fF
C228 S.n191 VSUBS 0.89fF $ **FLOATING
C229 S.t2081 VSUBS 0.02fF
C230 S.n192 VSUBS 0.89fF $ **FLOATING
C231 S.n193 VSUBS 2.64fF $ **FLOATING
C232 S.n194 VSUBS 8.97fF $ **FLOATING
C233 S.n195 VSUBS 8.97fF $ **FLOATING
C234 S.n196 VSUBS 5.53fF $ **FLOATING
C235 S.n197 VSUBS 1.51fF $ **FLOATING
C236 S.n198 VSUBS 0.02fF $ **FLOATING
C237 S.t1015 VSUBS 0.02fF
C238 S.n199 VSUBS 0.37fF $ **FLOATING
C239 S.n200 VSUBS 20.80fF $ **FLOATING
C240 S.n201 VSUBS 20.80fF $ **FLOATING
C241 S.n202 VSUBS 5.79fF $ **FLOATING
C242 S.n203 VSUBS 1.96fF $ **FLOATING
C243 S.t1585 VSUBS 0.02fF
C244 S.n204 VSUBS 0.89fF $ **FLOATING
C245 S.t353 VSUBS 0.02fF
C246 S.n205 VSUBS 0.89fF $ **FLOATING
C247 S.n206 VSUBS 1.62fF $ **FLOATING
C248 S.n207 VSUBS 0.02fF $ **FLOATING
C249 S.t1266 VSUBS 0.02fF
C250 S.n208 VSUBS 0.37fF $ **FLOATING
C251 S.t1829 VSUBS 0.02fF
C252 S.n209 VSUBS 0.89fF $ **FLOATING
C253 S.n210 VSUBS 0.02fF $ **FLOATING
C254 S.t1773 VSUBS 0.02fF
C255 S.n211 VSUBS 0.37fF $ **FLOATING
C256 S.t956 VSUBS 0.02fF
C257 S.n212 VSUBS 0.89fF $ **FLOATING
C258 S.t1007 VSUBS 0.02fF
C259 S.n213 VSUBS 0.89fF $ **FLOATING
C260 S.n214 VSUBS 0.02fF $ **FLOATING
C261 S.t950 VSUBS 0.02fF
C262 S.n215 VSUBS 0.37fF $ **FLOATING
C263 S.t119 VSUBS 0.02fF
C264 S.n216 VSUBS 0.89fF $ **FLOATING
C265 S.t1400 VSUBS 0.02fF
C266 S.n217 VSUBS 0.89fF $ **FLOATING
C267 S.n218 VSUBS 0.02fF $ **FLOATING
C268 S.t1348 VSUBS 0.02fF
C269 S.n219 VSUBS 0.37fF $ **FLOATING
C270 S.t533 VSUBS 0.02fF
C271 S.n220 VSUBS 0.89fF $ **FLOATING
C272 S.t453 VSUBS 0.02fF
C273 S.n221 VSUBS 0.89fF $ **FLOATING
C274 S.n222 VSUBS 0.02fF $ **FLOATING
C275 S.t405 VSUBS 0.02fF
C276 S.n223 VSUBS 0.37fF $ **FLOATING
C277 S.t2229 VSUBS 0.02fF
C278 S.n224 VSUBS 0.89fF $ **FLOATING
C279 S.t976 VSUBS 0.02fF
C280 S.n225 VSUBS 0.89fF $ **FLOATING
C281 S.n226 VSUBS 0.02fF $ **FLOATING
C282 S.t924 VSUBS 0.02fF
C283 S.n227 VSUBS 0.37fF $ **FLOATING
C284 S.t76 VSUBS 0.02fF
C285 S.n228 VSUBS 0.89fF $ **FLOATING
C286 S.t2541 VSUBS 0.02fF
C287 S.n229 VSUBS 0.89fF $ **FLOATING
C288 S.n230 VSUBS 0.02fF $ **FLOATING
C289 S.t2491 VSUBS 0.02fF
C290 S.n231 VSUBS 0.37fF $ **FLOATING
C291 S.t1671 VSUBS 0.02fF
C292 S.n232 VSUBS 0.89fF $ **FLOATING
C293 S.t2238 VSUBS 0.02fF
C294 S.n233 VSUBS 0.89fF $ **FLOATING
C295 S.n234 VSUBS 0.02fF $ **FLOATING
C296 S.t1184 VSUBS 0.02fF
C297 S.n235 VSUBS 0.37fF $ **FLOATING
C298 S.t1372 VSUBS 0.02fF
C299 S.n236 VSUBS 0.89fF $ **FLOATING
C300 S.t7 VSUBS 172.40fF
C301 S.n237 VSUBS 3.28fF $ **FLOATING
C302 S.n238 VSUBS 9.43fF $ **FLOATING
C303 S.n239 VSUBS 9.37fF $ **FLOATING
C304 S.n240 VSUBS 9.43fF $ **FLOATING
C305 S.n241 VSUBS 9.37fF $ **FLOATING
C306 S.n242 VSUBS 9.37fF $ **FLOATING
C307 S.n243 VSUBS 9.37fF $ **FLOATING
C308 S.n244 VSUBS 9.43fF $ **FLOATING
C309 S.n245 VSUBS 12.50fF $ **FLOATING
C310 S.n246 VSUBS 1.18fF $ **FLOATING
C311 S.n247 VSUBS 0.38fF $ **FLOATING
C312 S.n248 VSUBS 1.21fF $ **FLOATING
C313 S.n249 VSUBS 0.37fF $ **FLOATING
C314 S.n250 VSUBS 0.65fF $ **FLOATING
C315 S.n251 VSUBS 0.44fF $ **FLOATING
C316 S.n252 VSUBS 1.62fF $ **FLOATING
C317 S.n253 VSUBS 0.50fF $ **FLOATING
C318 S.n254 VSUBS 0.46fF $ **FLOATING
C319 S.n255 VSUBS 0.45fF $ **FLOATING
C320 S.n256 VSUBS 1.84fF $ **FLOATING
C321 S.n257 VSUBS 0.12fF $ **FLOATING
C322 S.t2320 VSUBS 0.02fF
C323 S.n258 VSUBS 0.14fF $ **FLOATING
C324 S.t616 VSUBS 0.02fF
C325 S.n260 VSUBS 0.24fF $ **FLOATING
C326 S.n261 VSUBS 0.36fF $ **FLOATING
C327 S.n262 VSUBS 0.61fF $ **FLOATING
C328 S.n263 VSUBS 2.49fF $ **FLOATING
C329 S.n264 VSUBS 2.02fF $ **FLOATING
C330 S.t903 VSUBS 0.02fF
C331 S.n265 VSUBS 0.24fF $ **FLOATING
C332 S.n266 VSUBS 0.91fF $ **FLOATING
C333 S.n267 VSUBS 0.05fF $ **FLOATING
C334 S.t665 VSUBS 0.02fF
C335 S.n268 VSUBS 0.12fF $ **FLOATING
C336 S.n269 VSUBS 0.14fF $ **FLOATING
C337 S.n271 VSUBS 0.18fF $ **FLOATING
C338 S.n272 VSUBS 0.10fF $ **FLOATING
C339 S.n273 VSUBS 0.94fF $ **FLOATING
C340 S.n274 VSUBS 0.46fF $ **FLOATING
C341 S.n275 VSUBS 0.77fF $ **FLOATING
C342 S.n276 VSUBS 0.21fF $ **FLOATING
C343 S.n277 VSUBS 0.36fF $ **FLOATING
C344 S.n278 VSUBS 0.53fF $ **FLOATING
C345 S.n279 VSUBS 1.62fF $ **FLOATING
C346 S.n280 VSUBS 0.12fF $ **FLOATING
C347 S.t702 VSUBS 0.02fF
C348 S.n281 VSUBS 0.14fF $ **FLOATING
C349 S.t1526 VSUBS 0.02fF
C350 S.n283 VSUBS 0.24fF $ **FLOATING
C351 S.n284 VSUBS 0.36fF $ **FLOATING
C352 S.n285 VSUBS 0.61fF $ **FLOATING
C353 S.n286 VSUBS 2.48fF $ **FLOATING
C354 S.n287 VSUBS 1.96fF $ **FLOATING
C355 S.t1820 VSUBS 0.02fF
C356 S.n288 VSUBS 0.24fF $ **FLOATING
C357 S.n289 VSUBS 0.91fF $ **FLOATING
C358 S.n290 VSUBS 0.05fF $ **FLOATING
C359 S.t1570 VSUBS 0.02fF
C360 S.n291 VSUBS 0.12fF $ **FLOATING
C361 S.n292 VSUBS 0.14fF $ **FLOATING
C362 S.n294 VSUBS 0.65fF $ **FLOATING
C363 S.n295 VSUBS 0.44fF $ **FLOATING
C364 S.n296 VSUBS 1.62fF $ **FLOATING
C365 S.n297 VSUBS 0.50fF $ **FLOATING
C366 S.n298 VSUBS 0.46fF $ **FLOATING
C367 S.n299 VSUBS 0.45fF $ **FLOATING
C368 S.n300 VSUBS 1.84fF $ **FLOATING
C369 S.n301 VSUBS 0.12fF $ **FLOATING
C370 S.t340 VSUBS 0.02fF
C371 S.n302 VSUBS 0.14fF $ **FLOATING
C372 S.t1155 VSUBS 0.02fF
C373 S.n304 VSUBS 0.24fF $ **FLOATING
C374 S.n305 VSUBS 0.36fF $ **FLOATING
C375 S.n306 VSUBS 0.61fF $ **FLOATING
C376 S.n307 VSUBS 2.49fF $ **FLOATING
C377 S.n308 VSUBS 2.02fF $ **FLOATING
C378 S.t1426 VSUBS 0.02fF
C379 S.n309 VSUBS 0.24fF $ **FLOATING
C380 S.n310 VSUBS 0.91fF $ **FLOATING
C381 S.n311 VSUBS 0.05fF $ **FLOATING
C382 S.t2361 VSUBS 0.02fF
C383 S.n312 VSUBS 0.12fF $ **FLOATING
C384 S.n313 VSUBS 0.14fF $ **FLOATING
C385 S.n315 VSUBS 0.18fF $ **FLOATING
C386 S.n316 VSUBS 0.10fF $ **FLOATING
C387 S.n317 VSUBS 0.94fF $ **FLOATING
C388 S.n318 VSUBS 0.46fF $ **FLOATING
C389 S.n319 VSUBS 0.77fF $ **FLOATING
C390 S.n320 VSUBS 0.21fF $ **FLOATING
C391 S.n321 VSUBS 0.36fF $ **FLOATING
C392 S.n322 VSUBS 0.53fF $ **FLOATING
C393 S.n323 VSUBS 1.62fF $ **FLOATING
C394 S.n324 VSUBS 0.12fF $ **FLOATING
C395 S.t1126 VSUBS 0.02fF
C396 S.n325 VSUBS 0.14fF $ **FLOATING
C397 S.t1939 VSUBS 0.02fF
C398 S.n327 VSUBS 0.24fF $ **FLOATING
C399 S.n328 VSUBS 0.36fF $ **FLOATING
C400 S.n329 VSUBS 0.61fF $ **FLOATING
C401 S.n330 VSUBS 2.48fF $ **FLOATING
C402 S.n331 VSUBS 1.96fF $ **FLOATING
C403 S.t2216 VSUBS 0.02fF
C404 S.n332 VSUBS 0.24fF $ **FLOATING
C405 S.n333 VSUBS 0.91fF $ **FLOATING
C406 S.n334 VSUBS 0.05fF $ **FLOATING
C407 S.t1988 VSUBS 0.02fF
C408 S.n335 VSUBS 0.12fF $ **FLOATING
C409 S.n336 VSUBS 0.14fF $ **FLOATING
C410 S.n338 VSUBS 0.65fF $ **FLOATING
C411 S.n339 VSUBS 0.44fF $ **FLOATING
C412 S.n340 VSUBS 1.62fF $ **FLOATING
C413 S.n341 VSUBS 0.50fF $ **FLOATING
C414 S.n342 VSUBS 0.46fF $ **FLOATING
C415 S.n343 VSUBS 0.45fF $ **FLOATING
C416 S.n344 VSUBS 1.84fF $ **FLOATING
C417 S.n345 VSUBS 0.12fF $ **FLOATING
C418 S.t1906 VSUBS 0.02fF
C419 S.n346 VSUBS 0.14fF $ **FLOATING
C420 S.t195 VSUBS 0.02fF
C421 S.n348 VSUBS 0.24fF $ **FLOATING
C422 S.n349 VSUBS 0.36fF $ **FLOATING
C423 S.n350 VSUBS 0.61fF $ **FLOATING
C424 S.n351 VSUBS 2.49fF $ **FLOATING
C425 S.n352 VSUBS 2.02fF $ **FLOATING
C426 S.t481 VSUBS 0.02fF
C427 S.n353 VSUBS 0.24fF $ **FLOATING
C428 S.n354 VSUBS 0.91fF $ **FLOATING
C429 S.n355 VSUBS 0.05fF $ **FLOATING
C430 S.t256 VSUBS 0.02fF
C431 S.n356 VSUBS 0.12fF $ **FLOATING
C432 S.n357 VSUBS 0.14fF $ **FLOATING
C433 S.n359 VSUBS 0.18fF $ **FLOATING
C434 S.n360 VSUBS 0.10fF $ **FLOATING
C435 S.n361 VSUBS 0.94fF $ **FLOATING
C436 S.n362 VSUBS 0.46fF $ **FLOATING
C437 S.n363 VSUBS 0.77fF $ **FLOATING
C438 S.n364 VSUBS 0.21fF $ **FLOATING
C439 S.n365 VSUBS 0.36fF $ **FLOATING
C440 S.n366 VSUBS 0.53fF $ **FLOATING
C441 S.n367 VSUBS 1.62fF $ **FLOATING
C442 S.n368 VSUBS 0.12fF $ **FLOATING
C443 S.t160 VSUBS 0.02fF
C444 S.n369 VSUBS 0.14fF $ **FLOATING
C445 S.t982 VSUBS 0.02fF
C446 S.n371 VSUBS 0.24fF $ **FLOATING
C447 S.n372 VSUBS 0.36fF $ **FLOATING
C448 S.n373 VSUBS 0.61fF $ **FLOATING
C449 S.n374 VSUBS 2.48fF $ **FLOATING
C450 S.n375 VSUBS 1.96fF $ **FLOATING
C451 S.t1270 VSUBS 0.02fF
C452 S.n376 VSUBS 0.24fF $ **FLOATING
C453 S.n377 VSUBS 0.91fF $ **FLOATING
C454 S.n378 VSUBS 0.05fF $ **FLOATING
C455 S.t1038 VSUBS 0.02fF
C456 S.n379 VSUBS 0.12fF $ **FLOATING
C457 S.n380 VSUBS 0.14fF $ **FLOATING
C458 S.n382 VSUBS 0.65fF $ **FLOATING
C459 S.n383 VSUBS 0.44fF $ **FLOATING
C460 S.n384 VSUBS 1.62fF $ **FLOATING
C461 S.n385 VSUBS 0.50fF $ **FLOATING
C462 S.n386 VSUBS 0.46fF $ **FLOATING
C463 S.n387 VSUBS 0.45fF $ **FLOATING
C464 S.n388 VSUBS 1.84fF $ **FLOATING
C465 S.n389 VSUBS 0.12fF $ **FLOATING
C466 S.t1082 VSUBS 0.02fF
C467 S.n390 VSUBS 0.14fF $ **FLOATING
C468 S.t1896 VSUBS 0.02fF
C469 S.n392 VSUBS 0.24fF $ **FLOATING
C470 S.n393 VSUBS 0.36fF $ **FLOATING
C471 S.n394 VSUBS 0.61fF $ **FLOATING
C472 S.n395 VSUBS 2.49fF $ **FLOATING
C473 S.n396 VSUBS 2.02fF $ **FLOATING
C474 S.t2178 VSUBS 0.02fF
C475 S.n397 VSUBS 0.24fF $ **FLOATING
C476 S.n398 VSUBS 0.91fF $ **FLOATING
C477 S.n399 VSUBS 0.05fF $ **FLOATING
C478 S.t1950 VSUBS 0.02fF
C479 S.n400 VSUBS 0.12fF $ **FLOATING
C480 S.n401 VSUBS 0.14fF $ **FLOATING
C481 S.n403 VSUBS 0.18fF $ **FLOATING
C482 S.n404 VSUBS 0.10fF $ **FLOATING
C483 S.n405 VSUBS 0.94fF $ **FLOATING
C484 S.n406 VSUBS 0.46fF $ **FLOATING
C485 S.n407 VSUBS 0.77fF $ **FLOATING
C486 S.n408 VSUBS 0.21fF $ **FLOATING
C487 S.n409 VSUBS 0.36fF $ **FLOATING
C488 S.n410 VSUBS 0.53fF $ **FLOATING
C489 S.n411 VSUBS 1.62fF $ **FLOATING
C490 S.n412 VSUBS 0.12fF $ **FLOATING
C491 S.t678 VSUBS 0.02fF
C492 S.n413 VSUBS 0.14fF $ **FLOATING
C493 S.t1498 VSUBS 0.02fF
C494 S.n415 VSUBS 0.24fF $ **FLOATING
C495 S.n416 VSUBS 0.36fF $ **FLOATING
C496 S.n417 VSUBS 0.61fF $ **FLOATING
C497 S.n418 VSUBS 2.48fF $ **FLOATING
C498 S.n419 VSUBS 1.96fF $ **FLOATING
C499 S.t1789 VSUBS 0.02fF
C500 S.n420 VSUBS 0.24fF $ **FLOATING
C501 S.n421 VSUBS 0.91fF $ **FLOATING
C502 S.n422 VSUBS 0.05fF $ **FLOATING
C503 S.t1549 VSUBS 0.02fF
C504 S.n423 VSUBS 0.12fF $ **FLOATING
C505 S.n424 VSUBS 0.14fF $ **FLOATING
C506 S.n426 VSUBS 0.65fF $ **FLOATING
C507 S.n427 VSUBS 0.44fF $ **FLOATING
C508 S.n428 VSUBS 1.62fF $ **FLOATING
C509 S.n429 VSUBS 0.50fF $ **FLOATING
C510 S.n430 VSUBS 0.46fF $ **FLOATING
C511 S.n431 VSUBS 0.45fF $ **FLOATING
C512 S.n432 VSUBS 1.84fF $ **FLOATING
C513 S.n433 VSUBS 0.12fF $ **FLOATING
C514 S.t1468 VSUBS 0.02fF
C515 S.n434 VSUBS 0.14fF $ **FLOATING
C516 S.t2284 VSUBS 0.02fF
C517 S.n436 VSUBS 0.24fF $ **FLOATING
C518 S.n437 VSUBS 0.36fF $ **FLOATING
C519 S.n438 VSUBS 0.61fF $ **FLOATING
C520 S.n439 VSUBS 2.49fF $ **FLOATING
C521 S.n440 VSUBS 2.02fF $ **FLOATING
C522 S.t2571 VSUBS 0.02fF
C523 S.n441 VSUBS 0.24fF $ **FLOATING
C524 S.n442 VSUBS 0.91fF $ **FLOATING
C525 S.n443 VSUBS 0.05fF $ **FLOATING
C526 S.t2335 VSUBS 0.02fF
C527 S.n444 VSUBS 0.12fF $ **FLOATING
C528 S.n445 VSUBS 0.14fF $ **FLOATING
C529 S.n447 VSUBS 0.18fF $ **FLOATING
C530 S.n448 VSUBS 0.10fF $ **FLOATING
C531 S.n449 VSUBS 0.94fF $ **FLOATING
C532 S.n450 VSUBS 0.46fF $ **FLOATING
C533 S.n451 VSUBS 0.77fF $ **FLOATING
C534 S.n452 VSUBS 0.21fF $ **FLOATING
C535 S.n453 VSUBS 0.36fF $ **FLOATING
C536 S.n454 VSUBS 0.53fF $ **FLOATING
C537 S.n455 VSUBS 1.62fF $ **FLOATING
C538 S.n456 VSUBS 0.12fF $ **FLOATING
C539 S.t2256 VSUBS 0.02fF
C540 S.n457 VSUBS 0.14fF $ **FLOATING
C541 S.t600 VSUBS 0.02fF
C542 S.n459 VSUBS 0.12fF $ **FLOATING
C543 S.n460 VSUBS 0.14fF $ **FLOATING
C544 S.t556 VSUBS 0.02fF
C545 S.n462 VSUBS 0.24fF $ **FLOATING
C546 S.n463 VSUBS 0.36fF $ **FLOATING
C547 S.n464 VSUBS 0.61fF $ **FLOATING
C548 S.n465 VSUBS 2.48fF $ **FLOATING
C549 S.n466 VSUBS 1.96fF $ **FLOATING
C550 S.t837 VSUBS 0.02fF
C551 S.n467 VSUBS 0.24fF $ **FLOATING
C552 S.n468 VSUBS 0.91fF $ **FLOATING
C553 S.n469 VSUBS 0.05fF $ **FLOATING
C554 S.n470 VSUBS 0.65fF $ **FLOATING
C555 S.n471 VSUBS 0.44fF $ **FLOATING
C556 S.n472 VSUBS 1.62fF $ **FLOATING
C557 S.n473 VSUBS 0.50fF $ **FLOATING
C558 S.n474 VSUBS 0.46fF $ **FLOATING
C559 S.n475 VSUBS 0.45fF $ **FLOATING
C560 S.n476 VSUBS 1.84fF $ **FLOATING
C561 S.n477 VSUBS 0.12fF $ **FLOATING
C562 S.t525 VSUBS 0.02fF
C563 S.n478 VSUBS 0.14fF $ **FLOATING
C564 S.t1344 VSUBS 0.02fF
C565 S.n480 VSUBS 0.24fF $ **FLOATING
C566 S.n481 VSUBS 0.36fF $ **FLOATING
C567 S.n482 VSUBS 0.61fF $ **FLOATING
C568 S.n483 VSUBS 2.49fF $ **FLOATING
C569 S.n484 VSUBS 2.02fF $ **FLOATING
C570 S.t1619 VSUBS 0.02fF
C571 S.n485 VSUBS 0.24fF $ **FLOATING
C572 S.n486 VSUBS 0.91fF $ **FLOATING
C573 S.n487 VSUBS 0.05fF $ **FLOATING
C574 S.t1392 VSUBS 0.02fF
C575 S.n488 VSUBS 0.12fF $ **FLOATING
C576 S.n489 VSUBS 0.14fF $ **FLOATING
C577 S.n491 VSUBS 0.18fF $ **FLOATING
C578 S.n492 VSUBS 0.10fF $ **FLOATING
C579 S.n493 VSUBS 0.94fF $ **FLOATING
C580 S.n494 VSUBS 0.46fF $ **FLOATING
C581 S.n495 VSUBS 0.77fF $ **FLOATING
C582 S.n496 VSUBS 0.21fF $ **FLOATING
C583 S.n497 VSUBS 0.36fF $ **FLOATING
C584 S.n498 VSUBS 0.53fF $ **FLOATING
C585 S.n499 VSUBS 1.62fF $ **FLOATING
C586 S.n500 VSUBS 0.12fF $ **FLOATING
C587 S.t1397 VSUBS 0.02fF
C588 S.n501 VSUBS 0.14fF $ **FLOATING
C589 S.t1212 VSUBS 0.02fF
C590 S.n503 VSUBS 0.24fF $ **FLOATING
C591 S.n504 VSUBS 0.36fF $ **FLOATING
C592 S.n505 VSUBS 0.61fF $ **FLOATING
C593 S.n506 VSUBS 2.48fF $ **FLOATING
C594 S.n507 VSUBS 1.96fF $ **FLOATING
C595 S.t2045 VSUBS 0.02fF
C596 S.n508 VSUBS 0.24fF $ **FLOATING
C597 S.n509 VSUBS 0.91fF $ **FLOATING
C598 S.n510 VSUBS 0.05fF $ **FLOATING
C599 S.t2299 VSUBS 0.02fF
C600 S.n511 VSUBS 0.12fF $ **FLOATING
C601 S.n512 VSUBS 0.14fF $ **FLOATING
C602 S.n514 VSUBS 1.89fF $ **FLOATING
C603 S.n515 VSUBS 0.12fF $ **FLOATING
C604 S.t2211 VSUBS 0.02fF
C605 S.n516 VSUBS 0.14fF $ **FLOATING
C606 S.t421 VSUBS 0.02fF
C607 S.n518 VSUBS 1.22fF $ **FLOATING
C608 S.n519 VSUBS 2.29fF $ **FLOATING
C609 S.n520 VSUBS 0.61fF $ **FLOATING
C610 S.n521 VSUBS 0.35fF $ **FLOATING
C611 S.n522 VSUBS 0.63fF $ **FLOATING
C612 S.n523 VSUBS 1.15fF $ **FLOATING
C613 S.n524 VSUBS 3.00fF $ **FLOATING
C614 S.n525 VSUBS 0.59fF $ **FLOATING
C615 S.n526 VSUBS 0.01fF $ **FLOATING
C616 S.n527 VSUBS 0.97fF $ **FLOATING
C617 S.t185 VSUBS 21.42fF
C618 S.n528 VSUBS 20.29fF $ **FLOATING
C619 S.n530 VSUBS 0.38fF $ **FLOATING
C620 S.n531 VSUBS 0.23fF $ **FLOATING
C621 S.n532 VSUBS 2.89fF $ **FLOATING
C622 S.n533 VSUBS 2.46fF $ **FLOATING
C623 S.n534 VSUBS 4.30fF $ **FLOATING
C624 S.n535 VSUBS 0.25fF $ **FLOATING
C625 S.n536 VSUBS 0.01fF $ **FLOATING
C626 S.t2126 VSUBS 0.02fF
C627 S.n537 VSUBS 0.26fF $ **FLOATING
C628 S.t693 VSUBS 0.02fF
C629 S.n538 VSUBS 0.95fF $ **FLOATING
C630 S.n539 VSUBS 0.71fF $ **FLOATING
C631 S.n540 VSUBS 1.89fF $ **FLOATING
C632 S.n541 VSUBS 1.78fF $ **FLOATING
C633 S.n542 VSUBS 0.12fF $ **FLOATING
C634 S.t395 VSUBS 0.02fF
C635 S.n543 VSUBS 0.14fF $ **FLOATING
C636 S.t1216 VSUBS 0.02fF
C637 S.n545 VSUBS 0.24fF $ **FLOATING
C638 S.n546 VSUBS 0.36fF $ **FLOATING
C639 S.n547 VSUBS 0.61fF $ **FLOATING
C640 S.n548 VSUBS 2.74fF $ **FLOATING
C641 S.n549 VSUBS 2.05fF $ **FLOATING
C642 S.t1485 VSUBS 0.02fF
C643 S.n550 VSUBS 0.24fF $ **FLOATING
C644 S.n551 VSUBS 0.91fF $ **FLOATING
C645 S.n552 VSUBS 0.05fF $ **FLOATING
C646 S.t1261 VSUBS 0.02fF
C647 S.n553 VSUBS 0.12fF $ **FLOATING
C648 S.n554 VSUBS 0.14fF $ **FLOATING
C649 S.n556 VSUBS 1.24fF $ **FLOATING
C650 S.n557 VSUBS 1.28fF $ **FLOATING
C651 S.n558 VSUBS 1.88fF $ **FLOATING
C652 S.n559 VSUBS 0.12fF $ **FLOATING
C653 S.t1299 VSUBS 0.02fF
C654 S.n560 VSUBS 0.14fF $ **FLOATING
C655 S.t1994 VSUBS 0.02fF
C656 S.n562 VSUBS 0.24fF $ **FLOATING
C657 S.n563 VSUBS 0.36fF $ **FLOATING
C658 S.n564 VSUBS 0.61fF $ **FLOATING
C659 S.n565 VSUBS 2.75fF $ **FLOATING
C660 S.n566 VSUBS 2.17fF $ **FLOATING
C661 S.t2266 VSUBS 0.02fF
C662 S.n567 VSUBS 0.24fF $ **FLOATING
C663 S.n568 VSUBS 0.91fF $ **FLOATING
C664 S.n569 VSUBS 0.05fF $ **FLOATING
C665 S.t2049 VSUBS 0.02fF
C666 S.n570 VSUBS 0.12fF $ **FLOATING
C667 S.n571 VSUBS 0.14fF $ **FLOATING
C668 S.n573 VSUBS 1.89fF $ **FLOATING
C669 S.n574 VSUBS 1.79fF $ **FLOATING
C670 S.n575 VSUBS 0.12fF $ **FLOATING
C671 S.t2089 VSUBS 0.02fF
C672 S.n576 VSUBS 0.14fF $ **FLOATING
C673 S.t386 VSUBS 0.02fF
C674 S.n578 VSUBS 0.24fF $ **FLOATING
C675 S.n579 VSUBS 0.36fF $ **FLOATING
C676 S.n580 VSUBS 0.61fF $ **FLOATING
C677 S.n581 VSUBS 2.73fF $ **FLOATING
C678 S.n582 VSUBS 2.05fF $ **FLOATING
C679 S.t657 VSUBS 0.02fF
C680 S.n583 VSUBS 0.24fF $ **FLOATING
C681 S.n584 VSUBS 0.91fF $ **FLOATING
C682 S.n585 VSUBS 0.05fF $ **FLOATING
C683 S.t435 VSUBS 0.02fF
C684 S.n586 VSUBS 0.12fF $ **FLOATING
C685 S.n587 VSUBS 0.14fF $ **FLOATING
C686 S.n589 VSUBS 1.24fF $ **FLOATING
C687 S.n590 VSUBS 1.28fF $ **FLOATING
C688 S.n591 VSUBS 1.88fF $ **FLOATING
C689 S.n592 VSUBS 0.12fF $ **FLOATING
C690 S.t1689 VSUBS 0.02fF
C691 S.n593 VSUBS 0.14fF $ **FLOATING
C692 S.t2507 VSUBS 0.02fF
C693 S.n595 VSUBS 0.24fF $ **FLOATING
C694 S.n596 VSUBS 0.36fF $ **FLOATING
C695 S.n597 VSUBS 0.61fF $ **FLOATING
C696 S.n598 VSUBS 2.75fF $ **FLOATING
C697 S.n599 VSUBS 2.17fF $ **FLOATING
C698 S.t287 VSUBS 0.02fF
C699 S.n600 VSUBS 0.24fF $ **FLOATING
C700 S.n601 VSUBS 0.91fF $ **FLOATING
C701 S.n602 VSUBS 0.05fF $ **FLOATING
C702 S.t2558 VSUBS 0.02fF
C703 S.n603 VSUBS 0.12fF $ **FLOATING
C704 S.n604 VSUBS 0.14fF $ **FLOATING
C705 S.n606 VSUBS 1.89fF $ **FLOATING
C706 S.n607 VSUBS 1.79fF $ **FLOATING
C707 S.n608 VSUBS 0.12fF $ **FLOATING
C708 S.t2477 VSUBS 0.02fF
C709 S.n609 VSUBS 0.14fF $ **FLOATING
C710 S.t767 VSUBS 0.02fF
C711 S.n611 VSUBS 0.24fF $ **FLOATING
C712 S.n612 VSUBS 0.36fF $ **FLOATING
C713 S.n613 VSUBS 0.61fF $ **FLOATING
C714 S.n614 VSUBS 2.73fF $ **FLOATING
C715 S.n615 VSUBS 2.05fF $ **FLOATING
C716 S.t1070 VSUBS 0.02fF
C717 S.n616 VSUBS 0.24fF $ **FLOATING
C718 S.n617 VSUBS 0.91fF $ **FLOATING
C719 S.n618 VSUBS 0.05fF $ **FLOATING
C720 S.t824 VSUBS 0.02fF
C721 S.n619 VSUBS 0.12fF $ **FLOATING
C722 S.n620 VSUBS 0.14fF $ **FLOATING
C723 S.n622 VSUBS 1.24fF $ **FLOATING
C724 S.n623 VSUBS 1.28fF $ **FLOATING
C725 S.n624 VSUBS 1.88fF $ **FLOATING
C726 S.n625 VSUBS 0.12fF $ **FLOATING
C727 S.t733 VSUBS 0.02fF
C728 S.n626 VSUBS 0.14fF $ **FLOATING
C729 S.t1553 VSUBS 0.02fF
C730 S.n628 VSUBS 0.24fF $ **FLOATING
C731 S.n629 VSUBS 0.36fF $ **FLOATING
C732 S.n630 VSUBS 0.61fF $ **FLOATING
C733 S.n631 VSUBS 2.75fF $ **FLOATING
C734 S.n632 VSUBS 2.17fF $ **FLOATING
C735 S.t1853 VSUBS 0.02fF
C736 S.n633 VSUBS 0.24fF $ **FLOATING
C737 S.n634 VSUBS 0.91fF $ **FLOATING
C738 S.n635 VSUBS 0.05fF $ **FLOATING
C739 S.t1606 VSUBS 0.02fF
C740 S.n636 VSUBS 0.12fF $ **FLOATING
C741 S.n637 VSUBS 0.14fF $ **FLOATING
C742 S.n639 VSUBS 1.89fF $ **FLOATING
C743 S.n640 VSUBS 1.79fF $ **FLOATING
C744 S.n641 VSUBS 0.12fF $ **FLOATING
C745 S.t1650 VSUBS 0.02fF
C746 S.n642 VSUBS 0.14fF $ **FLOATING
C747 S.t2340 VSUBS 0.02fF
C748 S.n644 VSUBS 0.24fF $ **FLOATING
C749 S.n645 VSUBS 0.36fF $ **FLOATING
C750 S.n646 VSUBS 0.61fF $ **FLOATING
C751 S.n647 VSUBS 2.73fF $ **FLOATING
C752 S.n648 VSUBS 2.05fF $ **FLOATING
C753 S.t88 VSUBS 0.02fF
C754 S.n649 VSUBS 0.24fF $ **FLOATING
C755 S.n650 VSUBS 0.91fF $ **FLOATING
C756 S.n651 VSUBS 0.05fF $ **FLOATING
C757 S.t2392 VSUBS 0.02fF
C758 S.n652 VSUBS 0.12fF $ **FLOATING
C759 S.n653 VSUBS 0.14fF $ **FLOATING
C760 S.n655 VSUBS 1.24fF $ **FLOATING
C761 S.n656 VSUBS 1.28fF $ **FLOATING
C762 S.n657 VSUBS 1.88fF $ **FLOATING
C763 S.n658 VSUBS 0.12fF $ **FLOATING
C764 S.t1274 VSUBS 0.02fF
C765 S.n659 VSUBS 0.14fF $ **FLOATING
C766 S.t2088 VSUBS 0.02fF
C767 S.n661 VSUBS 0.24fF $ **FLOATING
C768 S.n662 VSUBS 0.36fF $ **FLOATING
C769 S.n663 VSUBS 0.61fF $ **FLOATING
C770 S.n664 VSUBS 2.75fF $ **FLOATING
C771 S.n665 VSUBS 2.17fF $ **FLOATING
C772 S.t2362 VSUBS 0.02fF
C773 S.n666 VSUBS 0.24fF $ **FLOATING
C774 S.n667 VSUBS 0.91fF $ **FLOATING
C775 S.n668 VSUBS 0.05fF $ **FLOATING
C776 S.t780 VSUBS 0.02fF
C777 S.n669 VSUBS 0.12fF $ **FLOATING
C778 S.n670 VSUBS 0.14fF $ **FLOATING
C779 S.n672 VSUBS 1.89fF $ **FLOATING
C780 S.n673 VSUBS 1.79fF $ **FLOATING
C781 S.n674 VSUBS 0.12fF $ **FLOATING
C782 S.t2062 VSUBS 0.02fF
C783 S.n675 VSUBS 0.14fF $ **FLOATING
C784 S.t362 VSUBS 0.02fF
C785 S.n677 VSUBS 0.24fF $ **FLOATING
C786 S.n678 VSUBS 0.36fF $ **FLOATING
C787 S.n679 VSUBS 0.61fF $ **FLOATING
C788 S.n680 VSUBS 2.73fF $ **FLOATING
C789 S.n681 VSUBS 2.05fF $ **FLOATING
C790 S.t631 VSUBS 0.02fF
C791 S.n682 VSUBS 0.24fF $ **FLOATING
C792 S.n683 VSUBS 0.91fF $ **FLOATING
C793 S.n684 VSUBS 0.05fF $ **FLOATING
C794 S.t408 VSUBS 0.02fF
C795 S.n685 VSUBS 0.12fF $ **FLOATING
C796 S.n686 VSUBS 0.14fF $ **FLOATING
C797 S.n688 VSUBS 1.24fF $ **FLOATING
C798 S.n689 VSUBS 1.28fF $ **FLOATING
C799 S.n690 VSUBS 1.88fF $ **FLOATING
C800 S.n691 VSUBS 0.12fF $ **FLOATING
C801 S.t327 VSUBS 0.02fF
C802 S.n692 VSUBS 0.14fF $ **FLOATING
C803 S.t1147 VSUBS 0.02fF
C804 S.n694 VSUBS 0.24fF $ **FLOATING
C805 S.n695 VSUBS 0.36fF $ **FLOATING
C806 S.n696 VSUBS 0.61fF $ **FLOATING
C807 S.n697 VSUBS 2.75fF $ **FLOATING
C808 S.n698 VSUBS 2.17fF $ **FLOATING
C809 S.t1420 VSUBS 0.02fF
C810 S.n699 VSUBS 0.24fF $ **FLOATING
C811 S.n700 VSUBS 0.91fF $ **FLOATING
C812 S.n701 VSUBS 0.05fF $ **FLOATING
C813 S.t1200 VSUBS 0.02fF
C814 S.n702 VSUBS 0.12fF $ **FLOATING
C815 S.n703 VSUBS 0.14fF $ **FLOATING
C816 S.n705 VSUBS 1.89fF $ **FLOATING
C817 S.n706 VSUBS 1.79fF $ **FLOATING
C818 S.n707 VSUBS 0.12fF $ **FLOATING
C819 S.t1116 VSUBS 0.02fF
C820 S.n708 VSUBS 0.14fF $ **FLOATING
C821 S.t1929 VSUBS 0.02fF
C822 S.n710 VSUBS 0.24fF $ **FLOATING
C823 S.n711 VSUBS 0.36fF $ **FLOATING
C824 S.n712 VSUBS 0.61fF $ **FLOATING
C825 S.n713 VSUBS 2.73fF $ **FLOATING
C826 S.n714 VSUBS 2.05fF $ **FLOATING
C827 S.t2209 VSUBS 0.02fF
C828 S.n715 VSUBS 0.24fF $ **FLOATING
C829 S.n716 VSUBS 0.91fF $ **FLOATING
C830 S.n717 VSUBS 0.05fF $ **FLOATING
C831 S.t1980 VSUBS 0.02fF
C832 S.n718 VSUBS 0.12fF $ **FLOATING
C833 S.n719 VSUBS 0.14fF $ **FLOATING
C834 S.n721 VSUBS 1.24fF $ **FLOATING
C835 S.n722 VSUBS 1.28fF $ **FLOATING
C836 S.n723 VSUBS 1.88fF $ **FLOATING
C837 S.n724 VSUBS 0.12fF $ **FLOATING
C838 S.t2021 VSUBS 0.02fF
C839 S.n725 VSUBS 0.14fF $ **FLOATING
C840 S.t186 VSUBS 0.02fF
C841 S.n727 VSUBS 0.24fF $ **FLOATING
C842 S.n728 VSUBS 0.36fF $ **FLOATING
C843 S.n729 VSUBS 0.61fF $ **FLOATING
C844 S.n730 VSUBS 2.75fF $ **FLOATING
C845 S.n731 VSUBS 2.17fF $ **FLOATING
C846 S.t476 VSUBS 0.02fF
C847 S.n732 VSUBS 0.24fF $ **FLOATING
C848 S.n733 VSUBS 0.91fF $ **FLOATING
C849 S.n734 VSUBS 0.05fF $ **FLOATING
C850 S.t245 VSUBS 0.02fF
C851 S.n735 VSUBS 0.12fF $ **FLOATING
C852 S.n736 VSUBS 0.14fF $ **FLOATING
C853 S.n738 VSUBS 2.61fF $ **FLOATING
C854 S.n739 VSUBS 1.88fF $ **FLOATING
C855 S.n740 VSUBS 0.12fF $ **FLOATING
C856 S.t477 VSUBS 0.02fF
C857 S.n741 VSUBS 0.14fF $ **FLOATING
C858 S.t285 VSUBS 0.02fF
C859 S.n743 VSUBS 0.24fF $ **FLOATING
C860 S.n744 VSUBS 0.36fF $ **FLOATING
C861 S.n745 VSUBS 0.61fF $ **FLOATING
C862 S.n746 VSUBS 0.90fF $ **FLOATING
C863 S.n747 VSUBS 0.77fF $ **FLOATING
C864 S.n748 VSUBS 0.97fF $ **FLOATING
C865 S.n749 VSUBS 0.09fF $ **FLOATING
C866 S.n750 VSUBS 0.33fF $ **FLOATING
C867 S.n751 VSUBS 2.15fF $ **FLOATING
C868 S.t1127 VSUBS 0.02fF
C869 S.n752 VSUBS 0.24fF $ **FLOATING
C870 S.n753 VSUBS 0.91fF $ **FLOATING
C871 S.n754 VSUBS 0.05fF $ **FLOATING
C872 S.t1346 VSUBS 0.02fF
C873 S.n755 VSUBS 0.12fF $ **FLOATING
C874 S.n756 VSUBS 0.14fF $ **FLOATING
C875 S.n758 VSUBS 2.30fF $ **FLOATING
C876 S.n759 VSUBS 1.88fF $ **FLOATING
C877 S.n760 VSUBS 0.12fF $ **FLOATING
C878 S.t1264 VSUBS 0.02fF
C879 S.n761 VSUBS 0.14fF $ **FLOATING
C880 S.t1066 VSUBS 0.02fF
C881 S.n763 VSUBS 0.24fF $ **FLOATING
C882 S.n764 VSUBS 0.36fF $ **FLOATING
C883 S.n765 VSUBS 0.61fF $ **FLOATING
C884 S.n766 VSUBS 0.77fF $ **FLOATING
C885 S.n767 VSUBS 0.48fF $ **FLOATING
C886 S.n768 VSUBS 0.09fF $ **FLOATING
C887 S.n769 VSUBS 0.33fF $ **FLOATING
C888 S.n770 VSUBS 2.02fF $ **FLOATING
C889 S.t1910 VSUBS 0.02fF
C890 S.n771 VSUBS 0.24fF $ **FLOATING
C891 S.n772 VSUBS 0.91fF $ **FLOATING
C892 S.n773 VSUBS 0.05fF $ **FLOATING
C893 S.t2132 VSUBS 0.02fF
C894 S.n774 VSUBS 0.12fF $ **FLOATING
C895 S.n775 VSUBS 0.14fF $ **FLOATING
C896 S.n777 VSUBS 1.89fF $ **FLOATING
C897 S.n778 VSUBS 1.16fF $ **FLOATING
C898 S.n779 VSUBS 0.22fF $ **FLOATING
C899 S.n780 VSUBS 0.12fF $ **FLOATING
C900 S.t2053 VSUBS 0.02fF
C901 S.n781 VSUBS 0.14fF $ **FLOATING
C902 S.t1852 VSUBS 0.02fF
C903 S.n783 VSUBS 0.24fF $ **FLOATING
C904 S.n784 VSUBS 0.36fF $ **FLOATING
C905 S.n785 VSUBS 0.61fF $ **FLOATING
C906 S.n786 VSUBS 2.73fF $ **FLOATING
C907 S.n787 VSUBS 1.88fF $ **FLOATING
C908 S.t165 VSUBS 0.02fF
C909 S.n788 VSUBS 0.24fF $ **FLOATING
C910 S.n789 VSUBS 0.91fF $ **FLOATING
C911 S.n790 VSUBS 0.05fF $ **FLOATING
C912 S.t398 VSUBS 0.02fF
C913 S.n791 VSUBS 0.12fF $ **FLOATING
C914 S.n792 VSUBS 0.14fF $ **FLOATING
C915 S.n794 VSUBS 20.78fF $ **FLOATING
C916 S.n795 VSUBS 2.72fF $ **FLOATING
C917 S.n796 VSUBS 1.96fF $ **FLOATING
C918 S.n797 VSUBS 0.12fF $ **FLOATING
C919 S.t1383 VSUBS 0.02fF
C920 S.n798 VSUBS 0.14fF $ **FLOATING
C921 S.t989 VSUBS 0.02fF
C922 S.n800 VSUBS 0.24fF $ **FLOATING
C923 S.n801 VSUBS 0.36fF $ **FLOATING
C924 S.n802 VSUBS 0.61fF $ **FLOATING
C925 S.n803 VSUBS 1.56fF $ **FLOATING
C926 S.n804 VSUBS 0.28fF $ **FLOATING
C927 S.n805 VSUBS 2.10fF $ **FLOATING
C928 S.t1189 VSUBS 0.02fF
C929 S.n806 VSUBS 0.12fF $ **FLOATING
C930 S.n807 VSUBS 0.14fF $ **FLOATING
C931 S.t2377 VSUBS 0.02fF
C932 S.n809 VSUBS 0.24fF $ **FLOATING
C933 S.n810 VSUBS 0.91fF $ **FLOATING
C934 S.n811 VSUBS 0.05fF $ **FLOATING
C935 S.t244 VSUBS 48.27fF
C936 S.t557 VSUBS 0.02fF
C937 S.n812 VSUBS 0.12fF $ **FLOATING
C938 S.n813 VSUBS 0.14fF $ **FLOATING
C939 S.t341 VSUBS 0.02fF
C940 S.n815 VSUBS 0.24fF $ **FLOATING
C941 S.n816 VSUBS 0.91fF $ **FLOATING
C942 S.n817 VSUBS 0.05fF $ **FLOATING
C943 S.t2014 VSUBS 0.02fF
C944 S.n818 VSUBS 0.24fF $ **FLOATING
C945 S.n819 VSUBS 0.36fF $ **FLOATING
C946 S.n820 VSUBS 0.61fF $ **FLOATING
C947 S.n821 VSUBS 2.24fF $ **FLOATING
C948 S.n822 VSUBS 2.69fF $ **FLOATING
C949 S.n823 VSUBS 2.65fF $ **FLOATING
C950 S.n824 VSUBS 2.36fF $ **FLOATING
C951 S.n825 VSUBS 1.86fF $ **FLOATING
C952 S.n826 VSUBS 0.12fF $ **FLOATING
C953 S.t2185 VSUBS 0.02fF
C954 S.n827 VSUBS 0.14fF $ **FLOATING
C955 S.t1989 VSUBS 0.02fF
C956 S.n829 VSUBS 0.24fF $ **FLOATING
C957 S.n830 VSUBS 0.36fF $ **FLOATING
C958 S.n831 VSUBS 0.61fF $ **FLOATING
C959 S.n832 VSUBS 0.40fF $ **FLOATING
C960 S.n833 VSUBS 0.67fF $ **FLOATING
C961 S.n834 VSUBS 0.55fF $ **FLOATING
C962 S.n835 VSUBS 0.33fF $ **FLOATING
C963 S.n836 VSUBS 1.07fF $ **FLOATING
C964 S.n837 VSUBS 2.13fF $ **FLOATING
C965 S.t313 VSUBS 0.02fF
C966 S.n838 VSUBS 0.24fF $ **FLOATING
C967 S.n839 VSUBS 0.91fF $ **FLOATING
C968 S.n840 VSUBS 0.05fF $ **FLOATING
C969 S.t530 VSUBS 0.02fF
C970 S.n841 VSUBS 0.12fF $ **FLOATING
C971 S.n842 VSUBS 0.14fF $ **FLOATING
C972 S.n844 VSUBS 0.03fF $ **FLOATING
C973 S.n845 VSUBS 0.03fF $ **FLOATING
C974 S.n846 VSUBS 0.10fF $ **FLOATING
C975 S.n847 VSUBS 0.36fF $ **FLOATING
C976 S.n848 VSUBS 0.38fF $ **FLOATING
C977 S.n849 VSUBS 0.11fF $ **FLOATING
C978 S.n850 VSUBS 0.12fF $ **FLOATING
C979 S.n851 VSUBS 0.03fF $ **FLOATING
C980 S.n852 VSUBS 0.07fF $ **FLOATING
C981 S.n853 VSUBS 1.40fF $ **FLOATING
C982 S.n854 VSUBS 0.04fF $ **FLOATING
C983 S.n855 VSUBS 0.49fF $ **FLOATING
C984 S.n856 VSUBS 0.38fF $ **FLOATING
C985 S.n857 VSUBS 1.62fF $ **FLOATING
C986 S.n858 VSUBS 0.12fF $ **FLOATING
C987 S.t450 VSUBS 0.02fF
C988 S.n859 VSUBS 0.14fF $ **FLOATING
C989 S.t257 VSUBS 0.02fF
C990 S.n861 VSUBS 0.24fF $ **FLOATING
C991 S.n862 VSUBS 0.36fF $ **FLOATING
C992 S.n863 VSUBS 0.61fF $ **FLOATING
C993 S.n864 VSUBS 0.35fF $ **FLOATING
C994 S.n865 VSUBS 0.54fF $ **FLOATING
C995 S.n866 VSUBS 0.38fF $ **FLOATING
C996 S.n867 VSUBS 0.18fF $ **FLOATING
C997 S.n868 VSUBS 0.25fF $ **FLOATING
C998 S.n869 VSUBS 0.09fF $ **FLOATING
C999 S.n870 VSUBS 1.96fF $ **FLOATING
C1000 S.t1101 VSUBS 0.02fF
C1001 S.n871 VSUBS 0.24fF $ **FLOATING
C1002 S.n872 VSUBS 0.91fF $ **FLOATING
C1003 S.n873 VSUBS 0.05fF $ **FLOATING
C1004 S.t1317 VSUBS 0.02fF
C1005 S.n874 VSUBS 0.12fF $ **FLOATING
C1006 S.n875 VSUBS 0.14fF $ **FLOATING
C1007 S.n877 VSUBS 1.50fF $ **FLOATING
C1008 S.n878 VSUBS 0.25fF $ **FLOATING
C1009 S.n879 VSUBS 0.09fF $ **FLOATING
C1010 S.n880 VSUBS 0.78fF $ **FLOATING
C1011 S.n881 VSUBS 0.21fF $ **FLOATING
C1012 S.n882 VSUBS 1.73fF $ **FLOATING
C1013 S.n883 VSUBS 0.44fF $ **FLOATING
C1014 S.n884 VSUBS 0.12fF $ **FLOATING
C1015 S.t1240 VSUBS 0.02fF
C1016 S.n885 VSUBS 0.14fF $ **FLOATING
C1017 S.t1044 VSUBS 0.02fF
C1018 S.n887 VSUBS 0.24fF $ **FLOATING
C1019 S.n888 VSUBS 0.36fF $ **FLOATING
C1020 S.n889 VSUBS 0.61fF $ **FLOATING
C1021 S.n890 VSUBS 0.83fF $ **FLOATING
C1022 S.n891 VSUBS 0.32fF $ **FLOATING
C1023 S.n892 VSUBS 0.29fF $ **FLOATING
C1024 S.n893 VSUBS 0.25fF $ **FLOATING
C1025 S.n894 VSUBS 0.22fF $ **FLOATING
C1026 S.n895 VSUBS 0.60fF $ **FLOATING
C1027 S.n896 VSUBS 0.28fF $ **FLOATING
C1028 S.n897 VSUBS 0.14fF $ **FLOATING
C1029 S.n898 VSUBS 1.74fF $ **FLOATING
C1030 S.n899 VSUBS 1.93fF $ **FLOATING
C1031 S.t1883 VSUBS 0.02fF
C1032 S.n900 VSUBS 0.24fF $ **FLOATING
C1033 S.n901 VSUBS 0.91fF $ **FLOATING
C1034 S.n902 VSUBS 0.05fF $ **FLOATING
C1035 S.t2105 VSUBS 0.02fF
C1036 S.n903 VSUBS 0.12fF $ **FLOATING
C1037 S.n904 VSUBS 0.14fF $ **FLOATING
C1038 S.n906 VSUBS 0.19fF $ **FLOATING
C1039 S.n907 VSUBS 0.10fF $ **FLOATING
C1040 S.n908 VSUBS 0.68fF $ **FLOATING
C1041 S.n909 VSUBS 0.28fF $ **FLOATING
C1042 S.n910 VSUBS 1.74fF $ **FLOATING
C1043 S.n911 VSUBS 0.21fF $ **FLOATING
C1044 S.n912 VSUBS 1.84fF $ **FLOATING
C1045 S.n913 VSUBS 0.12fF $ **FLOATING
C1046 S.t2025 VSUBS 0.02fF
C1047 S.n914 VSUBS 0.14fF $ **FLOATING
C1048 S.t1823 VSUBS 0.02fF
C1049 S.n916 VSUBS 0.24fF $ **FLOATING
C1050 S.n917 VSUBS 0.36fF $ **FLOATING
C1051 S.n918 VSUBS 0.61fF $ **FLOATING
C1052 S.n919 VSUBS 2.49fF $ **FLOATING
C1053 S.n920 VSUBS 1.86fF $ **FLOATING
C1054 S.t127 VSUBS 0.02fF
C1055 S.n921 VSUBS 0.24fF $ **FLOATING
C1056 S.n922 VSUBS 0.91fF $ **FLOATING
C1057 S.n923 VSUBS 0.05fF $ **FLOATING
C1058 S.t375 VSUBS 0.02fF
C1059 S.n924 VSUBS 0.12fF $ **FLOATING
C1060 S.n925 VSUBS 0.14fF $ **FLOATING
C1061 S.n927 VSUBS 0.06fF $ **FLOATING
C1062 S.n928 VSUBS 0.20fF $ **FLOATING
C1063 S.n929 VSUBS 0.09fF $ **FLOATING
C1064 S.n930 VSUBS 0.21fF $ **FLOATING
C1065 S.n931 VSUBS 0.10fF $ **FLOATING
C1066 S.n932 VSUBS 0.30fF $ **FLOATING
C1067 S.n933 VSUBS 1.01fF $ **FLOATING
C1068 S.n934 VSUBS 0.45fF $ **FLOATING
C1069 S.n935 VSUBS 2.07fF $ **FLOATING
C1070 S.n936 VSUBS 0.12fF $ **FLOATING
C1071 S.t1534 VSUBS 0.02fF
C1072 S.n937 VSUBS 0.14fF $ **FLOATING
C1073 S.t2350 VSUBS 0.02fF
C1074 S.n939 VSUBS 0.24fF $ **FLOATING
C1075 S.n940 VSUBS 0.36fF $ **FLOATING
C1076 S.n941 VSUBS 0.61fF $ **FLOATING
C1077 S.n942 VSUBS 0.43fF $ **FLOATING
C1078 S.n943 VSUBS 0.96fF $ **FLOATING
C1079 S.n944 VSUBS 0.39fF $ **FLOATING
C1080 S.n945 VSUBS 0.44fF $ **FLOATING
C1081 S.n946 VSUBS 0.25fF $ **FLOATING
C1082 S.n947 VSUBS 0.79fF $ **FLOATING
C1083 S.n948 VSUBS 0.18fF $ **FLOATING
C1084 S.n949 VSUBS 0.09fF $ **FLOATING
C1085 S.n950 VSUBS 1.81fF $ **FLOATING
C1086 S.t2402 VSUBS 0.02fF
C1087 S.n951 VSUBS 0.12fF $ **FLOATING
C1088 S.n952 VSUBS 0.14fF $ **FLOATING
C1089 S.t93 VSUBS 0.02fF
C1090 S.n954 VSUBS 0.24fF $ **FLOATING
C1091 S.n955 VSUBS 0.91fF $ **FLOATING
C1092 S.n956 VSUBS 0.05fF $ **FLOATING
C1093 S.t159 VSUBS 47.89fF
C1094 S.t234 VSUBS 0.02fF
C1095 S.n957 VSUBS 0.01fF $ **FLOATING
C1096 S.n958 VSUBS 0.26fF $ **FLOATING
C1097 S.t1000 VSUBS 0.02fF
C1098 S.n960 VSUBS 1.19fF $ **FLOATING
C1099 S.n961 VSUBS 0.05fF $ **FLOATING
C1100 S.t698 VSUBS 0.02fF
C1101 S.n962 VSUBS 0.64fF $ **FLOATING
C1102 S.n963 VSUBS 0.61fF $ **FLOATING
C1103 S.n964 VSUBS 8.97fF $ **FLOATING
C1104 S.n965 VSUBS 20.37fF $ **FLOATING
C1105 S.n966 VSUBS 8.97fF $ **FLOATING
C1106 S.n967 VSUBS 20.37fF $ **FLOATING
C1107 S.n968 VSUBS 0.60fF $ **FLOATING
C1108 S.n969 VSUBS 0.22fF $ **FLOATING
C1109 S.n970 VSUBS 0.88fF $ **FLOATING
C1110 S.n971 VSUBS 0.88fF $ **FLOATING
C1111 S.n972 VSUBS 3.39fF $ **FLOATING
C1112 S.n973 VSUBS 0.29fF $ **FLOATING
C1113 S.t87 VSUBS 21.42fF
C1114 S.n974 VSUBS 21.71fF $ **FLOATING
C1115 S.n975 VSUBS 0.21fF $ **FLOATING
C1116 S.n976 VSUBS 1.42fF $ **FLOATING
C1117 S.n977 VSUBS 4.25fF $ **FLOATING
C1118 S.n978 VSUBS 1.14fF $ **FLOATING
C1119 S.n979 VSUBS 1.80fF $ **FLOATING
C1120 S.n980 VSUBS 4.23fF $ **FLOATING
C1121 S.n981 VSUBS 0.24fF $ **FLOATING
C1122 S.n982 VSUBS 0.60fF $ **FLOATING
C1123 S.n983 VSUBS 0.22fF $ **FLOATING
C1124 S.n984 VSUBS 0.59fF $ **FLOATING
C1125 S.n985 VSUBS 3.39fF $ **FLOATING
C1126 S.n986 VSUBS 0.29fF $ **FLOATING
C1127 S.t51 VSUBS 21.42fF
C1128 S.n987 VSUBS 21.71fF $ **FLOATING
C1129 S.n988 VSUBS 0.77fF $ **FLOATING
C1130 S.n989 VSUBS 0.28fF $ **FLOATING
C1131 S.n990 VSUBS 4.00fF $ **FLOATING
C1132 S.n991 VSUBS 1.50fF $ **FLOATING
C1133 S.n992 VSUBS 1.30fF $ **FLOATING
C1134 S.n993 VSUBS 0.28fF $ **FLOATING
C1135 S.n994 VSUBS 1.88fF $ **FLOATING
C1136 S.n995 VSUBS 0.25fF $ **FLOATING
C1137 S.n996 VSUBS 0.09fF $ **FLOATING
C1138 S.n997 VSUBS 0.21fF $ **FLOATING
C1139 S.n998 VSUBS 0.79fF $ **FLOATING
C1140 S.n999 VSUBS 0.44fF $ **FLOATING
C1141 S.n1000 VSUBS 0.12fF $ **FLOATING
C1142 S.t1755 VSUBS 0.02fF
C1143 S.n1001 VSUBS 0.14fF $ **FLOATING
C1144 S.t2565 VSUBS 0.02fF
C1145 S.n1003 VSUBS 0.24fF $ **FLOATING
C1146 S.n1004 VSUBS 0.36fF $ **FLOATING
C1147 S.n1005 VSUBS 0.61fF $ **FLOATING
C1148 S.n1006 VSUBS 0.02fF $ **FLOATING
C1149 S.n1007 VSUBS 0.01fF $ **FLOATING
C1150 S.n1008 VSUBS 0.02fF $ **FLOATING
C1151 S.n1009 VSUBS 0.08fF $ **FLOATING
C1152 S.n1010 VSUBS 0.06fF $ **FLOATING
C1153 S.n1011 VSUBS 0.03fF $ **FLOATING
C1154 S.n1012 VSUBS 0.04fF $ **FLOATING
C1155 S.n1013 VSUBS 1.00fF $ **FLOATING
C1156 S.n1014 VSUBS 0.36fF $ **FLOATING
C1157 S.n1015 VSUBS 1.85fF $ **FLOATING
C1158 S.n1016 VSUBS 1.98fF $ **FLOATING
C1159 S.t346 VSUBS 0.02fF
C1160 S.n1017 VSUBS 0.24fF $ **FLOATING
C1161 S.n1018 VSUBS 0.91fF $ **FLOATING
C1162 S.n1019 VSUBS 0.05fF $ **FLOATING
C1163 S.t73 VSUBS 0.02fF
C1164 S.n1020 VSUBS 0.12fF $ **FLOATING
C1165 S.n1021 VSUBS 0.14fF $ **FLOATING
C1166 S.n1023 VSUBS 1.89fF $ **FLOATING
C1167 S.n1024 VSUBS 0.06fF $ **FLOATING
C1168 S.n1025 VSUBS 0.03fF $ **FLOATING
C1169 S.n1026 VSUBS 0.04fF $ **FLOATING
C1170 S.n1027 VSUBS 0.99fF $ **FLOATING
C1171 S.n1028 VSUBS 0.02fF $ **FLOATING
C1172 S.n1029 VSUBS 0.01fF $ **FLOATING
C1173 S.n1030 VSUBS 0.02fF $ **FLOATING
C1174 S.n1031 VSUBS 0.08fF $ **FLOATING
C1175 S.n1032 VSUBS 0.36fF $ **FLOATING
C1176 S.n1033 VSUBS 1.86fF $ **FLOATING
C1177 S.t960 VSUBS 0.02fF
C1178 S.n1034 VSUBS 0.24fF $ **FLOATING
C1179 S.n1035 VSUBS 0.36fF $ **FLOATING
C1180 S.n1036 VSUBS 0.61fF $ **FLOATING
C1181 S.n1037 VSUBS 0.12fF $ **FLOATING
C1182 S.t135 VSUBS 0.02fF
C1183 S.n1038 VSUBS 0.14fF $ **FLOATING
C1184 S.n1040 VSUBS 0.95fF $ **FLOATING
C1185 S.n1041 VSUBS 0.59fF $ **FLOATING
C1186 S.n1042 VSUBS 0.25fF $ **FLOATING
C1187 S.n1043 VSUBS 0.70fF $ **FLOATING
C1188 S.n1044 VSUBS 0.23fF $ **FLOATING
C1189 S.n1045 VSUBS 0.09fF $ **FLOATING
C1190 S.n1046 VSUBS 1.88fF $ **FLOATING
C1191 S.t1251 VSUBS 0.02fF
C1192 S.n1047 VSUBS 0.24fF $ **FLOATING
C1193 S.n1048 VSUBS 0.91fF $ **FLOATING
C1194 S.n1049 VSUBS 0.05fF $ **FLOATING
C1195 S.t1018 VSUBS 0.02fF
C1196 S.n1050 VSUBS 0.12fF $ **FLOATING
C1197 S.n1051 VSUBS 0.14fF $ **FLOATING
C1198 S.n1053 VSUBS 1.88fF $ **FLOATING
C1199 S.n1054 VSUBS 0.25fF $ **FLOATING
C1200 S.n1055 VSUBS 0.09fF $ **FLOATING
C1201 S.n1056 VSUBS 0.21fF $ **FLOATING
C1202 S.n1057 VSUBS 0.79fF $ **FLOATING
C1203 S.n1058 VSUBS 0.44fF $ **FLOATING
C1204 S.n1059 VSUBS 0.12fF $ **FLOATING
C1205 S.t2273 VSUBS 0.02fF
C1206 S.n1060 VSUBS 0.14fF $ **FLOATING
C1207 S.t571 VSUBS 0.02fF
C1208 S.n1062 VSUBS 0.24fF $ **FLOATING
C1209 S.n1063 VSUBS 0.36fF $ **FLOATING
C1210 S.n1064 VSUBS 0.61fF $ **FLOATING
C1211 S.n1065 VSUBS 0.02fF $ **FLOATING
C1212 S.n1066 VSUBS 0.01fF $ **FLOATING
C1213 S.n1067 VSUBS 0.02fF $ **FLOATING
C1214 S.n1068 VSUBS 0.08fF $ **FLOATING
C1215 S.n1069 VSUBS 0.06fF $ **FLOATING
C1216 S.n1070 VSUBS 0.03fF $ **FLOATING
C1217 S.n1071 VSUBS 0.04fF $ **FLOATING
C1218 S.n1072 VSUBS 1.00fF $ **FLOATING
C1219 S.n1073 VSUBS 0.36fF $ **FLOATING
C1220 S.n1074 VSUBS 1.85fF $ **FLOATING
C1221 S.n1075 VSUBS 1.98fF $ **FLOATING
C1222 S.t855 VSUBS 0.02fF
C1223 S.n1076 VSUBS 0.24fF $ **FLOATING
C1224 S.n1077 VSUBS 0.91fF $ **FLOATING
C1225 S.n1078 VSUBS 0.05fF $ **FLOATING
C1226 S.t1798 VSUBS 0.02fF
C1227 S.n1079 VSUBS 0.12fF $ **FLOATING
C1228 S.n1080 VSUBS 0.14fF $ **FLOATING
C1229 S.n1082 VSUBS 1.89fF $ **FLOATING
C1230 S.n1083 VSUBS 0.06fF $ **FLOATING
C1231 S.n1084 VSUBS 0.03fF $ **FLOATING
C1232 S.n1085 VSUBS 0.04fF $ **FLOATING
C1233 S.n1086 VSUBS 0.99fF $ **FLOATING
C1234 S.n1087 VSUBS 0.02fF $ **FLOATING
C1235 S.n1088 VSUBS 0.01fF $ **FLOATING
C1236 S.n1089 VSUBS 0.02fF $ **FLOATING
C1237 S.n1090 VSUBS 0.08fF $ **FLOATING
C1238 S.n1091 VSUBS 0.36fF $ **FLOATING
C1239 S.n1092 VSUBS 1.86fF $ **FLOATING
C1240 S.t1358 VSUBS 0.02fF
C1241 S.n1093 VSUBS 0.24fF $ **FLOATING
C1242 S.n1094 VSUBS 0.36fF $ **FLOATING
C1243 S.n1095 VSUBS 0.61fF $ **FLOATING
C1244 S.n1096 VSUBS 0.12fF $ **FLOATING
C1245 S.t543 VSUBS 0.02fF
C1246 S.n1097 VSUBS 0.14fF $ **FLOATING
C1247 S.n1099 VSUBS 0.95fF $ **FLOATING
C1248 S.n1100 VSUBS 0.59fF $ **FLOATING
C1249 S.n1101 VSUBS 0.25fF $ **FLOATING
C1250 S.n1102 VSUBS 0.70fF $ **FLOATING
C1251 S.n1103 VSUBS 0.23fF $ **FLOATING
C1252 S.n1104 VSUBS 0.09fF $ **FLOATING
C1253 S.n1105 VSUBS 1.88fF $ **FLOATING
C1254 S.t1638 VSUBS 0.02fF
C1255 S.n1106 VSUBS 0.24fF $ **FLOATING
C1256 S.n1107 VSUBS 0.91fF $ **FLOATING
C1257 S.n1108 VSUBS 0.05fF $ **FLOATING
C1258 S.t1409 VSUBS 0.02fF
C1259 S.n1109 VSUBS 0.12fF $ **FLOATING
C1260 S.n1110 VSUBS 0.14fF $ **FLOATING
C1261 S.n1112 VSUBS 1.88fF $ **FLOATING
C1262 S.n1113 VSUBS 0.25fF $ **FLOATING
C1263 S.n1114 VSUBS 0.09fF $ **FLOATING
C1264 S.n1115 VSUBS 0.21fF $ **FLOATING
C1265 S.n1116 VSUBS 0.79fF $ **FLOATING
C1266 S.n1117 VSUBS 0.44fF $ **FLOATING
C1267 S.n1118 VSUBS 0.12fF $ **FLOATING
C1268 S.t1332 VSUBS 0.02fF
C1269 S.n1119 VSUBS 0.14fF $ **FLOATING
C1270 S.t2145 VSUBS 0.02fF
C1271 S.n1121 VSUBS 0.24fF $ **FLOATING
C1272 S.n1122 VSUBS 0.36fF $ **FLOATING
C1273 S.n1123 VSUBS 0.61fF $ **FLOATING
C1274 S.n1124 VSUBS 0.02fF $ **FLOATING
C1275 S.n1125 VSUBS 0.01fF $ **FLOATING
C1276 S.n1126 VSUBS 0.02fF $ **FLOATING
C1277 S.n1127 VSUBS 0.08fF $ **FLOATING
C1278 S.n1128 VSUBS 0.06fF $ **FLOATING
C1279 S.n1129 VSUBS 0.03fF $ **FLOATING
C1280 S.n1130 VSUBS 0.04fF $ **FLOATING
C1281 S.n1131 VSUBS 1.00fF $ **FLOATING
C1282 S.n1132 VSUBS 0.36fF $ **FLOATING
C1283 S.n1133 VSUBS 1.85fF $ **FLOATING
C1284 S.n1134 VSUBS 1.98fF $ **FLOATING
C1285 S.t2422 VSUBS 0.02fF
C1286 S.n1135 VSUBS 0.24fF $ **FLOATING
C1287 S.n1136 VSUBS 0.91fF $ **FLOATING
C1288 S.n1137 VSUBS 0.05fF $ **FLOATING
C1289 S.t2199 VSUBS 0.02fF
C1290 S.n1138 VSUBS 0.12fF $ **FLOATING
C1291 S.n1139 VSUBS 0.14fF $ **FLOATING
C1292 S.n1141 VSUBS 1.89fF $ **FLOATING
C1293 S.n1142 VSUBS 0.06fF $ **FLOATING
C1294 S.n1143 VSUBS 0.03fF $ **FLOATING
C1295 S.n1144 VSUBS 0.04fF $ **FLOATING
C1296 S.n1145 VSUBS 0.99fF $ **FLOATING
C1297 S.n1146 VSUBS 0.02fF $ **FLOATING
C1298 S.n1147 VSUBS 0.01fF $ **FLOATING
C1299 S.n1148 VSUBS 0.02fF $ **FLOATING
C1300 S.n1149 VSUBS 0.08fF $ **FLOATING
C1301 S.n1150 VSUBS 0.36fF $ **FLOATING
C1302 S.n1151 VSUBS 1.86fF $ **FLOATING
C1303 S.t412 VSUBS 0.02fF
C1304 S.n1152 VSUBS 0.24fF $ **FLOATING
C1305 S.n1153 VSUBS 0.36fF $ **FLOATING
C1306 S.n1154 VSUBS 0.61fF $ **FLOATING
C1307 S.n1155 VSUBS 0.12fF $ **FLOATING
C1308 S.t2116 VSUBS 0.02fF
C1309 S.n1156 VSUBS 0.14fF $ **FLOATING
C1310 S.n1158 VSUBS 0.95fF $ **FLOATING
C1311 S.n1159 VSUBS 0.59fF $ **FLOATING
C1312 S.n1160 VSUBS 0.25fF $ **FLOATING
C1313 S.n1161 VSUBS 0.70fF $ **FLOATING
C1314 S.n1162 VSUBS 0.23fF $ **FLOATING
C1315 S.n1163 VSUBS 0.09fF $ **FLOATING
C1316 S.n1164 VSUBS 1.88fF $ **FLOATING
C1317 S.t684 VSUBS 0.02fF
C1318 S.n1165 VSUBS 0.24fF $ **FLOATING
C1319 S.n1166 VSUBS 0.91fF $ **FLOATING
C1320 S.n1167 VSUBS 0.05fF $ **FLOATING
C1321 S.t465 VSUBS 0.02fF
C1322 S.n1168 VSUBS 0.12fF $ **FLOATING
C1323 S.n1169 VSUBS 0.14fF $ **FLOATING
C1324 S.n1171 VSUBS 1.88fF $ **FLOATING
C1325 S.n1172 VSUBS 0.25fF $ **FLOATING
C1326 S.n1173 VSUBS 0.09fF $ **FLOATING
C1327 S.n1174 VSUBS 0.21fF $ **FLOATING
C1328 S.n1175 VSUBS 0.79fF $ **FLOATING
C1329 S.n1176 VSUBS 0.44fF $ **FLOATING
C1330 S.n1177 VSUBS 0.12fF $ **FLOATING
C1331 S.t509 VSUBS 0.02fF
C1332 S.n1178 VSUBS 0.14fF $ **FLOATING
C1333 S.t1323 VSUBS 0.02fF
C1334 S.n1180 VSUBS 0.24fF $ **FLOATING
C1335 S.n1181 VSUBS 0.36fF $ **FLOATING
C1336 S.n1182 VSUBS 0.61fF $ **FLOATING
C1337 S.n1183 VSUBS 0.02fF $ **FLOATING
C1338 S.n1184 VSUBS 0.01fF $ **FLOATING
C1339 S.n1185 VSUBS 0.02fF $ **FLOATING
C1340 S.n1186 VSUBS 0.08fF $ **FLOATING
C1341 S.n1187 VSUBS 0.06fF $ **FLOATING
C1342 S.n1188 VSUBS 0.03fF $ **FLOATING
C1343 S.n1189 VSUBS 0.04fF $ **FLOATING
C1344 S.n1190 VSUBS 1.00fF $ **FLOATING
C1345 S.n1191 VSUBS 0.36fF $ **FLOATING
C1346 S.n1192 VSUBS 1.85fF $ **FLOATING
C1347 S.n1193 VSUBS 1.98fF $ **FLOATING
C1348 S.t1593 VSUBS 0.02fF
C1349 S.n1194 VSUBS 0.24fF $ **FLOATING
C1350 S.n1195 VSUBS 0.91fF $ **FLOATING
C1351 S.n1196 VSUBS 0.05fF $ **FLOATING
C1352 S.t1375 VSUBS 0.02fF
C1353 S.n1197 VSUBS 0.12fF $ **FLOATING
C1354 S.n1198 VSUBS 0.14fF $ **FLOATING
C1355 S.n1200 VSUBS 1.89fF $ **FLOATING
C1356 S.n1201 VSUBS 0.06fF $ **FLOATING
C1357 S.n1202 VSUBS 0.03fF $ **FLOATING
C1358 S.n1203 VSUBS 0.04fF $ **FLOATING
C1359 S.n1204 VSUBS 0.99fF $ **FLOATING
C1360 S.n1205 VSUBS 0.02fF $ **FLOATING
C1361 S.n1206 VSUBS 0.01fF $ **FLOATING
C1362 S.n1207 VSUBS 0.02fF $ **FLOATING
C1363 S.n1208 VSUBS 0.08fF $ **FLOATING
C1364 S.n1209 VSUBS 0.36fF $ **FLOATING
C1365 S.n1210 VSUBS 1.86fF $ **FLOATING
C1366 S.t933 VSUBS 0.02fF
C1367 S.n1211 VSUBS 0.24fF $ **FLOATING
C1368 S.n1212 VSUBS 0.36fF $ **FLOATING
C1369 S.n1213 VSUBS 0.61fF $ **FLOATING
C1370 S.n1214 VSUBS 0.12fF $ **FLOATING
C1371 S.t90 VSUBS 0.02fF
C1372 S.n1215 VSUBS 0.14fF $ **FLOATING
C1373 S.n1217 VSUBS 0.95fF $ **FLOATING
C1374 S.n1218 VSUBS 0.59fF $ **FLOATING
C1375 S.n1219 VSUBS 0.25fF $ **FLOATING
C1376 S.n1220 VSUBS 0.70fF $ **FLOATING
C1377 S.n1221 VSUBS 0.23fF $ **FLOATING
C1378 S.n1222 VSUBS 0.09fF $ **FLOATING
C1379 S.n1223 VSUBS 1.88fF $ **FLOATING
C1380 S.t1230 VSUBS 0.02fF
C1381 S.n1224 VSUBS 0.24fF $ **FLOATING
C1382 S.n1225 VSUBS 0.91fF $ **FLOATING
C1383 S.n1226 VSUBS 0.05fF $ **FLOATING
C1384 S.t987 VSUBS 0.02fF
C1385 S.n1227 VSUBS 0.12fF $ **FLOATING
C1386 S.n1228 VSUBS 0.14fF $ **FLOATING
C1387 S.n1230 VSUBS 1.88fF $ **FLOATING
C1388 S.n1231 VSUBS 0.25fF $ **FLOATING
C1389 S.n1232 VSUBS 0.09fF $ **FLOATING
C1390 S.n1233 VSUBS 0.21fF $ **FLOATING
C1391 S.n1234 VSUBS 0.79fF $ **FLOATING
C1392 S.n1235 VSUBS 0.44fF $ **FLOATING
C1393 S.n1236 VSUBS 0.12fF $ **FLOATING
C1394 S.t900 VSUBS 0.02fF
C1395 S.n1237 VSUBS 0.14fF $ **FLOATING
C1396 S.t1711 VSUBS 0.02fF
C1397 S.n1239 VSUBS 0.24fF $ **FLOATING
C1398 S.n1240 VSUBS 0.36fF $ **FLOATING
C1399 S.n1241 VSUBS 0.61fF $ **FLOATING
C1400 S.n1242 VSUBS 0.02fF $ **FLOATING
C1401 S.n1243 VSUBS 0.01fF $ **FLOATING
C1402 S.n1244 VSUBS 0.02fF $ **FLOATING
C1403 S.n1245 VSUBS 0.08fF $ **FLOATING
C1404 S.n1246 VSUBS 0.06fF $ **FLOATING
C1405 S.n1247 VSUBS 0.03fF $ **FLOATING
C1406 S.n1248 VSUBS 0.04fF $ **FLOATING
C1407 S.n1249 VSUBS 1.00fF $ **FLOATING
C1408 S.n1250 VSUBS 0.36fF $ **FLOATING
C1409 S.n1251 VSUBS 1.85fF $ **FLOATING
C1410 S.n1252 VSUBS 1.98fF $ **FLOATING
C1411 S.t2008 VSUBS 0.02fF
C1412 S.n1253 VSUBS 0.24fF $ **FLOATING
C1413 S.n1254 VSUBS 0.91fF $ **FLOATING
C1414 S.n1255 VSUBS 0.05fF $ **FLOATING
C1415 S.t1769 VSUBS 0.02fF
C1416 S.n1256 VSUBS 0.12fF $ **FLOATING
C1417 S.n1257 VSUBS 0.14fF $ **FLOATING
C1418 S.n1259 VSUBS 1.89fF $ **FLOATING
C1419 S.n1260 VSUBS 0.06fF $ **FLOATING
C1420 S.n1261 VSUBS 0.03fF $ **FLOATING
C1421 S.n1262 VSUBS 0.04fF $ **FLOATING
C1422 S.n1263 VSUBS 0.99fF $ **FLOATING
C1423 S.n1264 VSUBS 0.02fF $ **FLOATING
C1424 S.n1265 VSUBS 0.01fF $ **FLOATING
C1425 S.n1266 VSUBS 0.02fF $ **FLOATING
C1426 S.n1267 VSUBS 0.08fF $ **FLOATING
C1427 S.n1268 VSUBS 0.36fF $ **FLOATING
C1428 S.n1269 VSUBS 1.86fF $ **FLOATING
C1429 S.t2498 VSUBS 0.02fF
C1430 S.n1270 VSUBS 0.24fF $ **FLOATING
C1431 S.n1271 VSUBS 0.36fF $ **FLOATING
C1432 S.n1272 VSUBS 0.61fF $ **FLOATING
C1433 S.n1273 VSUBS 0.12fF $ **FLOATING
C1434 S.t1680 VSUBS 0.02fF
C1435 S.n1274 VSUBS 0.14fF $ **FLOATING
C1436 S.n1276 VSUBS 0.95fF $ **FLOATING
C1437 S.n1277 VSUBS 0.59fF $ **FLOATING
C1438 S.n1278 VSUBS 0.25fF $ **FLOATING
C1439 S.n1279 VSUBS 0.70fF $ **FLOATING
C1440 S.n1280 VSUBS 0.23fF $ **FLOATING
C1441 S.n1281 VSUBS 0.09fF $ **FLOATING
C1442 S.n1282 VSUBS 1.88fF $ **FLOATING
C1443 S.t280 VSUBS 0.02fF
C1444 S.n1283 VSUBS 0.24fF $ **FLOATING
C1445 S.n1284 VSUBS 0.91fF $ **FLOATING
C1446 S.n1285 VSUBS 0.05fF $ **FLOATING
C1447 S.t2547 VSUBS 0.02fF
C1448 S.n1286 VSUBS 0.12fF $ **FLOATING
C1449 S.n1287 VSUBS 0.14fF $ **FLOATING
C1450 S.n1289 VSUBS 1.88fF $ **FLOATING
C1451 S.n1290 VSUBS 0.25fF $ **FLOATING
C1452 S.n1291 VSUBS 0.09fF $ **FLOATING
C1453 S.n1292 VSUBS 0.21fF $ **FLOATING
C1454 S.n1293 VSUBS 0.79fF $ **FLOATING
C1455 S.n1294 VSUBS 0.44fF $ **FLOATING
C1456 S.n1295 VSUBS 0.12fF $ **FLOATING
C1457 S.t2466 VSUBS 0.02fF
C1458 S.n1296 VSUBS 0.14fF $ **FLOATING
C1459 S.t754 VSUBS 0.02fF
C1460 S.n1298 VSUBS 0.24fF $ **FLOATING
C1461 S.n1299 VSUBS 0.36fF $ **FLOATING
C1462 S.n1300 VSUBS 0.61fF $ **FLOATING
C1463 S.n1301 VSUBS 0.02fF $ **FLOATING
C1464 S.n1302 VSUBS 0.01fF $ **FLOATING
C1465 S.n1303 VSUBS 0.02fF $ **FLOATING
C1466 S.n1304 VSUBS 0.08fF $ **FLOATING
C1467 S.n1305 VSUBS 0.03fF $ **FLOATING
C1468 S.n1306 VSUBS 0.04fF $ **FLOATING
C1469 S.n1307 VSUBS 1.02fF $ **FLOATING
C1470 S.n1308 VSUBS 0.36fF $ **FLOATING
C1471 S.n1309 VSUBS 1.85fF $ **FLOATING
C1472 S.n1310 VSUBS 1.98fF $ **FLOATING
C1473 S.t1060 VSUBS 0.02fF
C1474 S.n1311 VSUBS 0.24fF $ **FLOATING
C1475 S.n1312 VSUBS 0.91fF $ **FLOATING
C1476 S.n1313 VSUBS 0.05fF $ **FLOATING
C1477 S.t813 VSUBS 0.02fF
C1478 S.n1314 VSUBS 0.12fF $ **FLOATING
C1479 S.n1315 VSUBS 0.14fF $ **FLOATING
C1480 S.n1317 VSUBS 0.25fF $ **FLOATING
C1481 S.n1318 VSUBS 0.70fF $ **FLOATING
C1482 S.n1319 VSUBS 0.23fF $ **FLOATING
C1483 S.n1320 VSUBS 0.09fF $ **FLOATING
C1484 S.n1321 VSUBS 0.95fF $ **FLOATING
C1485 S.n1322 VSUBS 0.59fF $ **FLOATING
C1486 S.n1323 VSUBS 1.89fF $ **FLOATING
C1487 S.n1324 VSUBS 0.12fF $ **FLOATING
C1488 S.t2235 VSUBS 0.02fF
C1489 S.n1325 VSUBS 0.14fF $ **FLOATING
C1490 S.t2039 VSUBS 0.02fF
C1491 S.n1327 VSUBS 0.24fF $ **FLOATING
C1492 S.n1328 VSUBS 0.36fF $ **FLOATING
C1493 S.n1329 VSUBS 0.61fF $ **FLOATING
C1494 S.n1330 VSUBS 0.18fF $ **FLOATING
C1495 S.n1331 VSUBS 0.21fF $ **FLOATING
C1496 S.n1332 VSUBS 0.47fF $ **FLOATING
C1497 S.n1333 VSUBS 0.33fF $ **FLOATING
C1498 S.n1334 VSUBS 0.01fF $ **FLOATING
C1499 S.n1335 VSUBS 0.01fF $ **FLOATING
C1500 S.n1336 VSUBS 0.01fF $ **FLOATING
C1501 S.n1337 VSUBS 0.07fF $ **FLOATING
C1502 S.n1338 VSUBS 0.07fF $ **FLOATING
C1503 S.n1339 VSUBS 0.04fF $ **FLOATING
C1504 S.n1340 VSUBS 0.05fF $ **FLOATING
C1505 S.n1341 VSUBS 0.41fF $ **FLOATING
C1506 S.n1342 VSUBS 0.58fF $ **FLOATING
C1507 S.n1343 VSUBS 0.19fF $ **FLOATING
C1508 S.n1344 VSUBS 1.97fF $ **FLOATING
C1509 S.t366 VSUBS 0.02fF
C1510 S.n1345 VSUBS 0.24fF $ **FLOATING
C1511 S.n1346 VSUBS 0.91fF $ **FLOATING
C1512 S.n1347 VSUBS 0.05fF $ **FLOATING
C1513 S.t1728 VSUBS 0.02fF
C1514 S.n1348 VSUBS 0.12fF $ **FLOATING
C1515 S.n1349 VSUBS 0.14fF $ **FLOATING
C1516 S.n1351 VSUBS 0.04fF $ **FLOATING
C1517 S.n1352 VSUBS 0.03fF $ **FLOATING
C1518 S.n1353 VSUBS 0.03fF $ **FLOATING
C1519 S.n1354 VSUBS 0.10fF $ **FLOATING
C1520 S.n1355 VSUBS 0.36fF $ **FLOATING
C1521 S.n1356 VSUBS 0.38fF $ **FLOATING
C1522 S.n1357 VSUBS 0.11fF $ **FLOATING
C1523 S.n1358 VSUBS 0.12fF $ **FLOATING
C1524 S.n1359 VSUBS 0.07fF $ **FLOATING
C1525 S.n1360 VSUBS 0.12fF $ **FLOATING
C1526 S.n1361 VSUBS 0.18fF $ **FLOATING
C1527 S.n1362 VSUBS 1.88fF $ **FLOATING
C1528 S.n1363 VSUBS 0.12fF $ **FLOATING
C1529 S.t504 VSUBS 0.02fF
C1530 S.n1364 VSUBS 0.14fF $ **FLOATING
C1531 S.t308 VSUBS 0.02fF
C1532 S.n1366 VSUBS 0.24fF $ **FLOATING
C1533 S.n1367 VSUBS 0.36fF $ **FLOATING
C1534 S.n1368 VSUBS 0.61fF $ **FLOATING
C1535 S.n1369 VSUBS 0.42fF $ **FLOATING
C1536 S.n1370 VSUBS 0.21fF $ **FLOATING
C1537 S.n1371 VSUBS 0.16fF $ **FLOATING
C1538 S.n1372 VSUBS 0.28fF $ **FLOATING
C1539 S.n1373 VSUBS 0.21fF $ **FLOATING
C1540 S.n1374 VSUBS 0.79fF $ **FLOATING
C1541 S.n1375 VSUBS 0.31fF $ **FLOATING
C1542 S.n1376 VSUBS 0.22fF $ **FLOATING
C1543 S.n1377 VSUBS 0.38fF $ **FLOATING
C1544 S.n1378 VSUBS 3.61fF $ **FLOATING
C1545 S.t1154 VSUBS 0.02fF
C1546 S.n1379 VSUBS 0.24fF $ **FLOATING
C1547 S.n1380 VSUBS 0.91fF $ **FLOATING
C1548 S.n1381 VSUBS 0.05fF $ **FLOATING
C1549 S.t1369 VSUBS 0.02fF
C1550 S.n1382 VSUBS 0.12fF $ **FLOATING
C1551 S.n1383 VSUBS 0.14fF $ **FLOATING
C1552 S.n1385 VSUBS 0.25fF $ **FLOATING
C1553 S.n1386 VSUBS 0.09fF $ **FLOATING
C1554 S.n1387 VSUBS 0.21fF $ **FLOATING
C1555 S.n1388 VSUBS 1.28fF $ **FLOATING
C1556 S.n1389 VSUBS 0.53fF $ **FLOATING
C1557 S.n1390 VSUBS 1.88fF $ **FLOATING
C1558 S.n1391 VSUBS 0.12fF $ **FLOATING
C1559 S.t1287 VSUBS 0.02fF
C1560 S.n1392 VSUBS 0.14fF $ **FLOATING
C1561 S.t1092 VSUBS 0.02fF
C1562 S.n1394 VSUBS 0.24fF $ **FLOATING
C1563 S.n1395 VSUBS 0.36fF $ **FLOATING
C1564 S.n1396 VSUBS 0.61fF $ **FLOATING
C1565 S.n1397 VSUBS 0.42fF $ **FLOATING
C1566 S.n1398 VSUBS 0.21fF $ **FLOATING
C1567 S.n1399 VSUBS 0.16fF $ **FLOATING
C1568 S.n1400 VSUBS 0.28fF $ **FLOATING
C1569 S.n1401 VSUBS 0.21fF $ **FLOATING
C1570 S.n1402 VSUBS 0.30fF $ **FLOATING
C1571 S.n1403 VSUBS 0.36fF $ **FLOATING
C1572 S.n1404 VSUBS 0.22fF $ **FLOATING
C1573 S.n1405 VSUBS 0.38fF $ **FLOATING
C1574 S.n1406 VSUBS 2.42fF $ **FLOATING
C1575 S.t1935 VSUBS 0.02fF
C1576 S.n1407 VSUBS 0.24fF $ **FLOATING
C1577 S.n1408 VSUBS 0.91fF $ **FLOATING
C1578 S.n1409 VSUBS 0.05fF $ **FLOATING
C1579 S.t2156 VSUBS 0.02fF
C1580 S.n1410 VSUBS 0.12fF $ **FLOATING
C1581 S.n1411 VSUBS 0.14fF $ **FLOATING
C1582 S.n1413 VSUBS 1.89fF $ **FLOATING
C1583 S.n1414 VSUBS 2.67fF $ **FLOATING
C1584 S.t1876 VSUBS 0.02fF
C1585 S.n1415 VSUBS 0.24fF $ **FLOATING
C1586 S.n1416 VSUBS 0.36fF $ **FLOATING
C1587 S.n1417 VSUBS 0.61fF $ **FLOATING
C1588 S.n1418 VSUBS 0.12fF $ **FLOATING
C1589 S.t2075 VSUBS 0.02fF
C1590 S.n1419 VSUBS 0.14fF $ **FLOATING
C1591 S.n1421 VSUBS 0.70fF $ **FLOATING
C1592 S.n1422 VSUBS 0.23fF $ **FLOATING
C1593 S.n1423 VSUBS 0.25fF $ **FLOATING
C1594 S.n1424 VSUBS 0.09fF $ **FLOATING
C1595 S.n1425 VSUBS 0.23fF $ **FLOATING
C1596 S.n1426 VSUBS 0.70fF $ **FLOATING
C1597 S.n1427 VSUBS 1.16fF $ **FLOATING
C1598 S.n1428 VSUBS 0.22fF $ **FLOATING
C1599 S.n1429 VSUBS 0.25fF $ **FLOATING
C1600 S.n1430 VSUBS 0.09fF $ **FLOATING
C1601 S.n1431 VSUBS 1.88fF $ **FLOATING
C1602 S.t194 VSUBS 0.02fF
C1603 S.n1432 VSUBS 0.24fF $ **FLOATING
C1604 S.n1433 VSUBS 0.91fF $ **FLOATING
C1605 S.n1434 VSUBS 0.05fF $ **FLOATING
C1606 S.t422 VSUBS 0.02fF
C1607 S.n1435 VSUBS 0.12fF $ **FLOATING
C1608 S.n1436 VSUBS 0.14fF $ **FLOATING
C1609 S.n1438 VSUBS 20.78fF $ **FLOATING
C1610 S.n1439 VSUBS 1.72fF $ **FLOATING
C1611 S.n1440 VSUBS 3.06fF $ **FLOATING
C1612 S.t1783 VSUBS 0.02fF
C1613 S.n1441 VSUBS 0.24fF $ **FLOATING
C1614 S.n1442 VSUBS 0.36fF $ **FLOATING
C1615 S.n1443 VSUBS 0.61fF $ **FLOATING
C1616 S.n1444 VSUBS 0.12fF $ **FLOATING
C1617 S.t968 VSUBS 0.02fF
C1618 S.n1445 VSUBS 0.14fF $ **FLOATING
C1619 S.n1447 VSUBS 0.28fF $ **FLOATING
C1620 S.n1448 VSUBS 0.74fF $ **FLOATING
C1621 S.n1449 VSUBS 0.60fF $ **FLOATING
C1622 S.n1450 VSUBS 0.21fF $ **FLOATING
C1623 S.n1451 VSUBS 0.20fF $ **FLOATING
C1624 S.n1452 VSUBS 0.06fF $ **FLOATING
C1625 S.n1453 VSUBS 0.09fF $ **FLOATING
C1626 S.n1454 VSUBS 0.10fF $ **FLOATING
C1627 S.n1455 VSUBS 1.99fF $ **FLOATING
C1628 S.t1838 VSUBS 0.02fF
C1629 S.n1456 VSUBS 0.12fF $ **FLOATING
C1630 S.n1457 VSUBS 0.14fF $ **FLOATING
C1631 S.t2073 VSUBS 0.02fF
C1632 S.n1459 VSUBS 0.24fF $ **FLOATING
C1633 S.n1460 VSUBS 0.91fF $ **FLOATING
C1634 S.n1461 VSUBS 0.05fF $ **FLOATING
C1635 S.n1462 VSUBS 1.88fF $ **FLOATING
C1636 S.n1463 VSUBS 0.12fF $ **FLOATING
C1637 S.t370 VSUBS 0.02fF
C1638 S.n1464 VSUBS 0.14fF $ **FLOATING
C1639 S.t2356 VSUBS 0.02fF
C1640 S.n1466 VSUBS 1.22fF $ **FLOATING
C1641 S.n1467 VSUBS 0.61fF $ **FLOATING
C1642 S.n1468 VSUBS 0.35fF $ **FLOATING
C1643 S.n1469 VSUBS 0.63fF $ **FLOATING
C1644 S.n1470 VSUBS 1.15fF $ **FLOATING
C1645 S.n1471 VSUBS 3.00fF $ **FLOATING
C1646 S.n1472 VSUBS 0.59fF $ **FLOATING
C1647 S.n1473 VSUBS 0.01fF $ **FLOATING
C1648 S.n1474 VSUBS 0.97fF $ **FLOATING
C1649 S.t97 VSUBS 21.42fF
C1650 S.n1475 VSUBS 20.29fF $ **FLOATING
C1651 S.n1477 VSUBS 0.38fF $ **FLOATING
C1652 S.n1478 VSUBS 0.23fF $ **FLOATING
C1653 S.n1479 VSUBS 2.90fF $ **FLOATING
C1654 S.n1480 VSUBS 2.46fF $ **FLOATING
C1655 S.n1481 VSUBS 1.96fF $ **FLOATING
C1656 S.n1482 VSUBS 3.94fF $ **FLOATING
C1657 S.n1483 VSUBS 0.25fF $ **FLOATING
C1658 S.n1484 VSUBS 0.01fF $ **FLOATING
C1659 S.t1542 VSUBS 0.02fF
C1660 S.n1485 VSUBS 0.26fF $ **FLOATING
C1661 S.t108 VSUBS 0.02fF
C1662 S.n1486 VSUBS 0.95fF $ **FLOATING
C1663 S.n1487 VSUBS 0.71fF $ **FLOATING
C1664 S.n1488 VSUBS 0.78fF $ **FLOATING
C1665 S.n1489 VSUBS 1.93fF $ **FLOATING
C1666 S.n1490 VSUBS 1.88fF $ **FLOATING
C1667 S.n1491 VSUBS 0.12fF $ **FLOATING
C1668 S.t2330 VSUBS 0.02fF
C1669 S.n1492 VSUBS 0.14fF $ **FLOATING
C1670 S.t623 VSUBS 0.02fF
C1671 S.n1494 VSUBS 0.24fF $ **FLOATING
C1672 S.n1495 VSUBS 0.36fF $ **FLOATING
C1673 S.n1496 VSUBS 0.61fF $ **FLOATING
C1674 S.n1497 VSUBS 1.52fF $ **FLOATING
C1675 S.n1498 VSUBS 2.99fF $ **FLOATING
C1676 S.t913 VSUBS 0.02fF
C1677 S.n1499 VSUBS 0.24fF $ **FLOATING
C1678 S.n1500 VSUBS 0.91fF $ **FLOATING
C1679 S.n1501 VSUBS 0.05fF $ **FLOATING
C1680 S.t674 VSUBS 0.02fF
C1681 S.n1502 VSUBS 0.12fF $ **FLOATING
C1682 S.n1503 VSUBS 0.14fF $ **FLOATING
C1683 S.n1505 VSUBS 1.89fF $ **FLOATING
C1684 S.n1506 VSUBS 1.88fF $ **FLOATING
C1685 S.t1416 VSUBS 0.02fF
C1686 S.n1507 VSUBS 0.24fF $ **FLOATING
C1687 S.n1508 VSUBS 0.36fF $ **FLOATING
C1688 S.n1509 VSUBS 0.61fF $ **FLOATING
C1689 S.n1510 VSUBS 0.12fF $ **FLOATING
C1690 S.t716 VSUBS 0.02fF
C1691 S.n1511 VSUBS 0.14fF $ **FLOATING
C1692 S.n1513 VSUBS 1.16fF $ **FLOATING
C1693 S.n1514 VSUBS 0.22fF $ **FLOATING
C1694 S.n1515 VSUBS 0.25fF $ **FLOATING
C1695 S.n1516 VSUBS 0.09fF $ **FLOATING
C1696 S.n1517 VSUBS 1.88fF $ **FLOATING
C1697 S.t1697 VSUBS 0.02fF
C1698 S.n1518 VSUBS 0.24fF $ **FLOATING
C1699 S.n1519 VSUBS 0.91fF $ **FLOATING
C1700 S.n1520 VSUBS 0.05fF $ **FLOATING
C1701 S.t1464 VSUBS 0.02fF
C1702 S.n1521 VSUBS 0.12fF $ **FLOATING
C1703 S.n1522 VSUBS 0.14fF $ **FLOATING
C1704 S.n1524 VSUBS 0.78fF $ **FLOATING
C1705 S.n1525 VSUBS 1.94fF $ **FLOATING
C1706 S.n1526 VSUBS 1.88fF $ **FLOATING
C1707 S.n1527 VSUBS 0.12fF $ **FLOATING
C1708 S.t1507 VSUBS 0.02fF
C1709 S.n1528 VSUBS 0.14fF $ **FLOATING
C1710 S.t2322 VSUBS 0.02fF
C1711 S.n1530 VSUBS 0.24fF $ **FLOATING
C1712 S.n1531 VSUBS 0.36fF $ **FLOATING
C1713 S.n1532 VSUBS 0.61fF $ **FLOATING
C1714 S.n1533 VSUBS 1.84fF $ **FLOATING
C1715 S.n1534 VSUBS 2.99fF $ **FLOATING
C1716 S.t52 VSUBS 0.02fF
C1717 S.n1535 VSUBS 0.24fF $ **FLOATING
C1718 S.n1536 VSUBS 0.91fF $ **FLOATING
C1719 S.n1537 VSUBS 0.05fF $ **FLOATING
C1720 S.t2373 VSUBS 0.02fF
C1721 S.n1538 VSUBS 0.12fF $ **FLOATING
C1722 S.n1539 VSUBS 0.14fF $ **FLOATING
C1723 S.n1541 VSUBS 1.89fF $ **FLOATING
C1724 S.n1542 VSUBS 1.88fF $ **FLOATING
C1725 S.t1946 VSUBS 0.02fF
C1726 S.n1543 VSUBS 0.24fF $ **FLOATING
C1727 S.n1544 VSUBS 0.36fF $ **FLOATING
C1728 S.n1545 VSUBS 0.61fF $ **FLOATING
C1729 S.n1546 VSUBS 0.12fF $ **FLOATING
C1730 S.t1139 VSUBS 0.02fF
C1731 S.n1547 VSUBS 0.14fF $ **FLOATING
C1732 S.n1549 VSUBS 1.16fF $ **FLOATING
C1733 S.n1550 VSUBS 0.22fF $ **FLOATING
C1734 S.n1551 VSUBS 0.25fF $ **FLOATING
C1735 S.n1552 VSUBS 0.09fF $ **FLOATING
C1736 S.n1553 VSUBS 1.88fF $ **FLOATING
C1737 S.t2224 VSUBS 0.02fF
C1738 S.n1554 VSUBS 0.24fF $ **FLOATING
C1739 S.n1555 VSUBS 0.91fF $ **FLOATING
C1740 S.n1556 VSUBS 0.05fF $ **FLOATING
C1741 S.t1999 VSUBS 0.02fF
C1742 S.n1557 VSUBS 0.12fF $ **FLOATING
C1743 S.n1558 VSUBS 0.14fF $ **FLOATING
C1744 S.n1560 VSUBS 0.78fF $ **FLOATING
C1745 S.n1561 VSUBS 1.94fF $ **FLOATING
C1746 S.n1562 VSUBS 1.88fF $ **FLOATING
C1747 S.n1563 VSUBS 0.12fF $ **FLOATING
C1748 S.t1920 VSUBS 0.02fF
C1749 S.n1564 VSUBS 0.14fF $ **FLOATING
C1750 S.t202 VSUBS 0.02fF
C1751 S.n1566 VSUBS 0.24fF $ **FLOATING
C1752 S.n1567 VSUBS 0.36fF $ **FLOATING
C1753 S.n1568 VSUBS 0.61fF $ **FLOATING
C1754 S.n1569 VSUBS 1.84fF $ **FLOATING
C1755 S.n1570 VSUBS 2.99fF $ **FLOATING
C1756 S.t492 VSUBS 0.02fF
C1757 S.n1571 VSUBS 0.24fF $ **FLOATING
C1758 S.n1572 VSUBS 0.91fF $ **FLOATING
C1759 S.n1573 VSUBS 0.05fF $ **FLOATING
C1760 S.t269 VSUBS 0.02fF
C1761 S.n1574 VSUBS 0.12fF $ **FLOATING
C1762 S.n1575 VSUBS 0.14fF $ **FLOATING
C1763 S.n1577 VSUBS 1.89fF $ **FLOATING
C1764 S.n1578 VSUBS 1.88fF $ **FLOATING
C1765 S.t994 VSUBS 0.02fF
C1766 S.n1579 VSUBS 0.24fF $ **FLOATING
C1767 S.n1580 VSUBS 0.36fF $ **FLOATING
C1768 S.n1581 VSUBS 0.61fF $ **FLOATING
C1769 S.n1582 VSUBS 0.12fF $ **FLOATING
C1770 S.t176 VSUBS 0.02fF
C1771 S.n1583 VSUBS 0.14fF $ **FLOATING
C1772 S.n1585 VSUBS 1.16fF $ **FLOATING
C1773 S.n1586 VSUBS 0.22fF $ **FLOATING
C1774 S.n1587 VSUBS 0.25fF $ **FLOATING
C1775 S.n1588 VSUBS 0.09fF $ **FLOATING
C1776 S.n1589 VSUBS 1.88fF $ **FLOATING
C1777 S.t1278 VSUBS 0.02fF
C1778 S.n1590 VSUBS 0.24fF $ **FLOATING
C1779 S.n1591 VSUBS 0.91fF $ **FLOATING
C1780 S.n1592 VSUBS 0.05fF $ **FLOATING
C1781 S.t1050 VSUBS 0.02fF
C1782 S.n1593 VSUBS 0.12fF $ **FLOATING
C1783 S.n1594 VSUBS 0.14fF $ **FLOATING
C1784 S.n1596 VSUBS 0.78fF $ **FLOATING
C1785 S.n1597 VSUBS 1.94fF $ **FLOATING
C1786 S.n1598 VSUBS 1.88fF $ **FLOATING
C1787 S.n1599 VSUBS 0.12fF $ **FLOATING
C1788 S.t1098 VSUBS 0.02fF
C1789 S.n1600 VSUBS 0.14fF $ **FLOATING
C1790 S.t1775 VSUBS 0.02fF
C1791 S.n1602 VSUBS 0.24fF $ **FLOATING
C1792 S.n1603 VSUBS 0.36fF $ **FLOATING
C1793 S.n1604 VSUBS 0.61fF $ **FLOATING
C1794 S.n1605 VSUBS 1.84fF $ **FLOATING
C1795 S.n1606 VSUBS 2.99fF $ **FLOATING
C1796 S.t2065 VSUBS 0.02fF
C1797 S.n1607 VSUBS 0.24fF $ **FLOATING
C1798 S.n1608 VSUBS 0.91fF $ **FLOATING
C1799 S.n1609 VSUBS 0.05fF $ **FLOATING
C1800 S.t1832 VSUBS 0.02fF
C1801 S.n1610 VSUBS 0.12fF $ **FLOATING
C1802 S.n1611 VSUBS 0.14fF $ **FLOATING
C1803 S.n1613 VSUBS 1.89fF $ **FLOATING
C1804 S.n1614 VSUBS 1.88fF $ **FLOATING
C1805 S.t1508 VSUBS 0.02fF
C1806 S.n1615 VSUBS 0.24fF $ **FLOATING
C1807 S.n1616 VSUBS 0.36fF $ **FLOATING
C1808 S.n1617 VSUBS 0.61fF $ **FLOATING
C1809 S.n1618 VSUBS 0.12fF $ **FLOATING
C1810 S.t692 VSUBS 0.02fF
C1811 S.n1619 VSUBS 0.14fF $ **FLOATING
C1812 S.n1621 VSUBS 1.16fF $ **FLOATING
C1813 S.n1622 VSUBS 0.22fF $ **FLOATING
C1814 S.n1623 VSUBS 0.25fF $ **FLOATING
C1815 S.n1624 VSUBS 0.09fF $ **FLOATING
C1816 S.n1625 VSUBS 1.88fF $ **FLOATING
C1817 S.t1797 VSUBS 0.02fF
C1818 S.n1626 VSUBS 0.24fF $ **FLOATING
C1819 S.n1627 VSUBS 0.91fF $ **FLOATING
C1820 S.n1628 VSUBS 0.05fF $ **FLOATING
C1821 S.t223 VSUBS 0.02fF
C1822 S.n1629 VSUBS 0.12fF $ **FLOATING
C1823 S.n1630 VSUBS 0.14fF $ **FLOATING
C1824 S.n1632 VSUBS 0.78fF $ **FLOATING
C1825 S.n1633 VSUBS 1.94fF $ **FLOATING
C1826 S.n1634 VSUBS 1.88fF $ **FLOATING
C1827 S.n1635 VSUBS 0.12fF $ **FLOATING
C1828 S.t1481 VSUBS 0.02fF
C1829 S.n1636 VSUBS 0.14fF $ **FLOATING
C1830 S.t2294 VSUBS 0.02fF
C1831 S.n1638 VSUBS 0.24fF $ **FLOATING
C1832 S.n1639 VSUBS 0.36fF $ **FLOATING
C1833 S.n1640 VSUBS 0.61fF $ **FLOATING
C1834 S.n1641 VSUBS 1.84fF $ **FLOATING
C1835 S.n1642 VSUBS 2.99fF $ **FLOATING
C1836 S.t2581 VSUBS 0.02fF
C1837 S.n1643 VSUBS 0.24fF $ **FLOATING
C1838 S.n1644 VSUBS 0.91fF $ **FLOATING
C1839 S.n1645 VSUBS 0.05fF $ **FLOATING
C1840 S.t2348 VSUBS 0.02fF
C1841 S.n1646 VSUBS 0.12fF $ **FLOATING
C1842 S.n1647 VSUBS 0.14fF $ **FLOATING
C1843 S.n1649 VSUBS 1.89fF $ **FLOATING
C1844 S.n1650 VSUBS 1.88fF $ **FLOATING
C1845 S.t563 VSUBS 0.02fF
C1846 S.n1651 VSUBS 0.24fF $ **FLOATING
C1847 S.n1652 VSUBS 0.36fF $ **FLOATING
C1848 S.n1653 VSUBS 0.61fF $ **FLOATING
C1849 S.n1654 VSUBS 0.12fF $ **FLOATING
C1850 S.t2264 VSUBS 0.02fF
C1851 S.n1655 VSUBS 0.14fF $ **FLOATING
C1852 S.n1657 VSUBS 1.16fF $ **FLOATING
C1853 S.n1658 VSUBS 0.22fF $ **FLOATING
C1854 S.n1659 VSUBS 0.25fF $ **FLOATING
C1855 S.n1660 VSUBS 0.09fF $ **FLOATING
C1856 S.n1661 VSUBS 1.88fF $ **FLOATING
C1857 S.t843 VSUBS 0.02fF
C1858 S.n1662 VSUBS 0.24fF $ **FLOATING
C1859 S.n1663 VSUBS 0.91fF $ **FLOATING
C1860 S.n1664 VSUBS 0.05fF $ **FLOATING
C1861 S.t612 VSUBS 0.02fF
C1862 S.n1665 VSUBS 0.12fF $ **FLOATING
C1863 S.n1666 VSUBS 0.14fF $ **FLOATING
C1864 S.n1668 VSUBS 0.78fF $ **FLOATING
C1865 S.n1669 VSUBS 1.94fF $ **FLOATING
C1866 S.n1670 VSUBS 1.88fF $ **FLOATING
C1867 S.n1671 VSUBS 0.12fF $ **FLOATING
C1868 S.t537 VSUBS 0.02fF
C1869 S.n1672 VSUBS 0.14fF $ **FLOATING
C1870 S.t1351 VSUBS 0.02fF
C1871 S.n1674 VSUBS 0.24fF $ **FLOATING
C1872 S.n1675 VSUBS 0.36fF $ **FLOATING
C1873 S.n1676 VSUBS 0.61fF $ **FLOATING
C1874 S.n1677 VSUBS 0.06fF $ **FLOATING
C1875 S.n1678 VSUBS 0.90fF $ **FLOATING
C1876 S.n1679 VSUBS 1.11fF $ **FLOATING
C1877 S.n1680 VSUBS 2.98fF $ **FLOATING
C1878 S.t1626 VSUBS 0.02fF
C1879 S.n1681 VSUBS 0.24fF $ **FLOATING
C1880 S.n1682 VSUBS 0.91fF $ **FLOATING
C1881 S.n1683 VSUBS 0.05fF $ **FLOATING
C1882 S.t1402 VSUBS 0.02fF
C1883 S.n1684 VSUBS 0.12fF $ **FLOATING
C1884 S.n1685 VSUBS 0.14fF $ **FLOATING
C1885 S.n1687 VSUBS 0.25fF $ **FLOATING
C1886 S.n1688 VSUBS 0.09fF $ **FLOATING
C1887 S.n1689 VSUBS 1.16fF $ **FLOATING
C1888 S.n1690 VSUBS 0.22fF $ **FLOATING
C1889 S.n1691 VSUBS 1.89fF $ **FLOATING
C1890 S.n1692 VSUBS 0.12fF $ **FLOATING
C1891 S.t1440 VSUBS 0.02fF
C1892 S.n1693 VSUBS 0.14fF $ **FLOATING
C1893 S.t2138 VSUBS 0.02fF
C1894 S.n1695 VSUBS 0.24fF $ **FLOATING
C1895 S.n1696 VSUBS 0.36fF $ **FLOATING
C1896 S.n1697 VSUBS 0.61fF $ **FLOATING
C1897 S.n1698 VSUBS 1.10fF $ **FLOATING
C1898 S.n1699 VSUBS 0.68fF $ **FLOATING
C1899 S.n1700 VSUBS 0.55fF $ **FLOATING
C1900 S.n1701 VSUBS 0.32fF $ **FLOATING
C1901 S.n1702 VSUBS 1.83fF $ **FLOATING
C1902 S.t2413 VSUBS 0.02fF
C1903 S.n1703 VSUBS 0.24fF $ **FLOATING
C1904 S.n1704 VSUBS 0.91fF $ **FLOATING
C1905 S.n1705 VSUBS 0.05fF $ **FLOATING
C1906 S.t2191 VSUBS 0.02fF
C1907 S.n1706 VSUBS 0.12fF $ **FLOATING
C1908 S.n1707 VSUBS 0.14fF $ **FLOATING
C1909 S.n1709 VSUBS 1.88fF $ **FLOATING
C1910 S.n1710 VSUBS 0.48fF $ **FLOATING
C1911 S.n1711 VSUBS 0.09fF $ **FLOATING
C1912 S.n1712 VSUBS 0.33fF $ **FLOATING
C1913 S.n1713 VSUBS 0.30fF $ **FLOATING
C1914 S.n1714 VSUBS 0.77fF $ **FLOATING
C1915 S.n1715 VSUBS 0.59fF $ **FLOATING
C1916 S.t335 VSUBS 0.02fF
C1917 S.n1716 VSUBS 0.24fF $ **FLOATING
C1918 S.n1717 VSUBS 0.36fF $ **FLOATING
C1919 S.n1718 VSUBS 0.61fF $ **FLOATING
C1920 S.n1719 VSUBS 0.12fF $ **FLOATING
C1921 S.t526 VSUBS 0.02fF
C1922 S.n1720 VSUBS 0.14fF $ **FLOATING
C1923 S.n1722 VSUBS 2.61fF $ **FLOATING
C1924 S.n1723 VSUBS 2.15fF $ **FLOATING
C1925 S.t1177 VSUBS 0.02fF
C1926 S.n1724 VSUBS 0.24fF $ **FLOATING
C1927 S.n1725 VSUBS 0.91fF $ **FLOATING
C1928 S.n1726 VSUBS 0.05fF $ **FLOATING
C1929 S.t1393 VSUBS 0.02fF
C1930 S.n1727 VSUBS 0.12fF $ **FLOATING
C1931 S.n1728 VSUBS 0.14fF $ **FLOATING
C1932 S.n1730 VSUBS 1.88fF $ **FLOATING
C1933 S.n1731 VSUBS 0.48fF $ **FLOATING
C1934 S.n1732 VSUBS 0.35fF $ **FLOATING
C1935 S.n1733 VSUBS 0.30fF $ **FLOATING
C1936 S.n1734 VSUBS 1.27fF $ **FLOATING
C1937 S.t1121 VSUBS 0.02fF
C1938 S.n1735 VSUBS 0.24fF $ **FLOATING
C1939 S.n1736 VSUBS 0.36fF $ **FLOATING
C1940 S.n1737 VSUBS 0.61fF $ **FLOATING
C1941 S.n1738 VSUBS 0.12fF $ **FLOATING
C1942 S.t1314 VSUBS 0.02fF
C1943 S.n1739 VSUBS 0.14fF $ **FLOATING
C1944 S.n1741 VSUBS 0.78fF $ **FLOATING
C1945 S.n1742 VSUBS 2.30fF $ **FLOATING
C1946 S.n1743 VSUBS 2.02fF $ **FLOATING
C1947 S.t1960 VSUBS 0.02fF
C1948 S.n1744 VSUBS 0.24fF $ **FLOATING
C1949 S.n1745 VSUBS 0.91fF $ **FLOATING
C1950 S.n1746 VSUBS 0.05fF $ **FLOATING
C1951 S.t2183 VSUBS 0.02fF
C1952 S.n1747 VSUBS 0.12fF $ **FLOATING
C1953 S.n1748 VSUBS 0.14fF $ **FLOATING
C1954 S.n1750 VSUBS 1.89fF $ **FLOATING
C1955 S.n1751 VSUBS 2.68fF $ **FLOATING
C1956 S.t1904 VSUBS 0.02fF
C1957 S.n1752 VSUBS 0.24fF $ **FLOATING
C1958 S.n1753 VSUBS 0.36fF $ **FLOATING
C1959 S.n1754 VSUBS 0.61fF $ **FLOATING
C1960 S.n1755 VSUBS 0.12fF $ **FLOATING
C1961 S.t2100 VSUBS 0.02fF
C1962 S.n1756 VSUBS 0.14fF $ **FLOATING
C1963 S.n1758 VSUBS 1.16fF $ **FLOATING
C1964 S.n1759 VSUBS 0.22fF $ **FLOATING
C1965 S.n1760 VSUBS 0.25fF $ **FLOATING
C1966 S.n1761 VSUBS 0.09fF $ **FLOATING
C1967 S.n1762 VSUBS 1.88fF $ **FLOATING
C1968 S.t220 VSUBS 0.02fF
C1969 S.n1763 VSUBS 0.24fF $ **FLOATING
C1970 S.n1764 VSUBS 0.91fF $ **FLOATING
C1971 S.n1765 VSUBS 0.05fF $ **FLOATING
C1972 S.t447 VSUBS 0.02fF
C1973 S.n1766 VSUBS 0.12fF $ **FLOATING
C1974 S.n1767 VSUBS 0.14fF $ **FLOATING
C1975 S.n1769 VSUBS 20.78fF $ **FLOATING
C1976 S.n1770 VSUBS 2.72fF $ **FLOATING
C1977 S.n1771 VSUBS 1.59fF $ **FLOATING
C1978 S.n1772 VSUBS 0.12fF $ **FLOATING
C1979 S.t1180 VSUBS 0.02fF
C1980 S.n1773 VSUBS 0.14fF $ **FLOATING
C1981 S.t697 VSUBS 0.02fF
C1982 S.n1775 VSUBS 0.24fF $ **FLOATING
C1983 S.n1776 VSUBS 0.36fF $ **FLOATING
C1984 S.n1777 VSUBS 0.61fF $ **FLOATING
C1985 S.n1778 VSUBS 2.36fF $ **FLOATING
C1986 S.n1779 VSUBS 2.30fF $ **FLOATING
C1987 S.t2016 VSUBS 0.02fF
C1988 S.n1780 VSUBS 0.12fF $ **FLOATING
C1989 S.n1781 VSUBS 0.14fF $ **FLOATING
C1990 S.t2112 VSUBS 0.02fF
C1991 S.n1783 VSUBS 0.24fF $ **FLOATING
C1992 S.n1784 VSUBS 0.91fF $ **FLOATING
C1993 S.n1785 VSUBS 0.05fF $ **FLOATING
C1994 S.t175 VSUBS 48.27fF
C1995 S.t1236 VSUBS 0.02fF
C1996 S.n1786 VSUBS 0.12fF $ **FLOATING
C1997 S.n1787 VSUBS 0.14fF $ **FLOATING
C1998 S.t1008 VSUBS 0.02fF
C1999 S.n1789 VSUBS 0.24fF $ **FLOATING
C2000 S.n1790 VSUBS 0.91fF $ **FLOATING
C2001 S.n1791 VSUBS 0.05fF $ **FLOATING
C2002 S.t154 VSUBS 0.02fF
C2003 S.n1792 VSUBS 0.24fF $ **FLOATING
C2004 S.n1793 VSUBS 0.36fF $ **FLOATING
C2005 S.n1794 VSUBS 0.61fF $ **FLOATING
C2006 S.n1795 VSUBS 0.32fF $ **FLOATING
C2007 S.n1796 VSUBS 1.55fF $ **FLOATING
C2008 S.n1797 VSUBS 0.15fF $ **FLOATING
C2009 S.n1798 VSUBS 4.97fF $ **FLOATING
C2010 S.n1799 VSUBS 1.88fF $ **FLOATING
C2011 S.n1800 VSUBS 0.12fF $ **FLOATING
C2012 S.t349 VSUBS 0.02fF
C2013 S.n1801 VSUBS 0.14fF $ **FLOATING
C2014 S.t122 VSUBS 0.02fF
C2015 S.n1803 VSUBS 0.24fF $ **FLOATING
C2016 S.n1804 VSUBS 0.36fF $ **FLOATING
C2017 S.n1805 VSUBS 0.61fF $ **FLOATING
C2018 S.n1806 VSUBS 0.70fF $ **FLOATING
C2019 S.n1807 VSUBS 1.27fF $ **FLOATING
C2020 S.n1808 VSUBS 5.97fF $ **FLOATING
C2021 S.t1217 VSUBS 0.02fF
C2022 S.n1809 VSUBS 0.12fF $ **FLOATING
C2023 S.n1810 VSUBS 0.14fF $ **FLOATING
C2024 S.t980 VSUBS 0.02fF
C2025 S.n1812 VSUBS 0.24fF $ **FLOATING
C2026 S.n1813 VSUBS 0.91fF $ **FLOATING
C2027 S.n1814 VSUBS 0.05fF $ **FLOATING
C2028 S.t72 VSUBS 47.89fF
C2029 S.t2529 VSUBS 0.02fF
C2030 S.n1815 VSUBS 0.01fF $ **FLOATING
C2031 S.n1816 VSUBS 0.26fF $ **FLOATING
C2032 S.t429 VSUBS 0.02fF
C2033 S.n1818 VSUBS 1.19fF $ **FLOATING
C2034 S.n1819 VSUBS 0.05fF $ **FLOATING
C2035 S.t126 VSUBS 0.02fF
C2036 S.n1820 VSUBS 0.64fF $ **FLOATING
C2037 S.n1821 VSUBS 0.61fF $ **FLOATING
C2038 S.n1822 VSUBS 1.50fF $ **FLOATING
C2039 S.n1823 VSUBS 0.35fF $ **FLOATING
C2040 S.n1824 VSUBS 1.30fF $ **FLOATING
C2041 S.n1825 VSUBS 0.16fF $ **FLOATING
C2042 S.n1826 VSUBS 1.66fF $ **FLOATING
C2043 S.n1827 VSUBS 2.64fF $ **FLOATING
C2044 S.n1828 VSUBS 0.24fF $ **FLOATING
C2045 S.n1829 VSUBS 1.50fF $ **FLOATING
C2046 S.n1830 VSUBS 1.31fF $ **FLOATING
C2047 S.n1831 VSUBS 0.28fF $ **FLOATING
C2048 S.n1832 VSUBS 1.89fF $ **FLOATING
C2049 S.n1833 VSUBS 0.06fF $ **FLOATING
C2050 S.n1834 VSUBS 0.03fF $ **FLOATING
C2051 S.n1835 VSUBS 0.04fF $ **FLOATING
C2052 S.n1836 VSUBS 0.99fF $ **FLOATING
C2053 S.n1837 VSUBS 0.02fF $ **FLOATING
C2054 S.n1838 VSUBS 0.01fF $ **FLOATING
C2055 S.n1839 VSUBS 0.02fF $ **FLOATING
C2056 S.n1840 VSUBS 0.08fF $ **FLOATING
C2057 S.n1841 VSUBS 0.36fF $ **FLOATING
C2058 S.n1842 VSUBS 1.85fF $ **FLOATING
C2059 S.t1707 VSUBS 0.02fF
C2060 S.n1843 VSUBS 0.24fF $ **FLOATING
C2061 S.n1844 VSUBS 0.36fF $ **FLOATING
C2062 S.n1845 VSUBS 0.61fF $ **FLOATING
C2063 S.n1846 VSUBS 0.12fF $ **FLOATING
C2064 S.t1194 VSUBS 0.02fF
C2065 S.n1847 VSUBS 0.14fF $ **FLOATING
C2066 S.n1849 VSUBS 0.70fF $ **FLOATING
C2067 S.n1850 VSUBS 0.23fF $ **FLOATING
C2068 S.n1851 VSUBS 0.23fF $ **FLOATING
C2069 S.n1852 VSUBS 0.70fF $ **FLOATING
C2070 S.n1853 VSUBS 1.16fF $ **FLOATING
C2071 S.n1854 VSUBS 0.22fF $ **FLOATING
C2072 S.n1855 VSUBS 0.25fF $ **FLOATING
C2073 S.n1856 VSUBS 0.09fF $ **FLOATING
C2074 S.n1857 VSUBS 1.88fF $ **FLOATING
C2075 S.t2276 VSUBS 0.02fF
C2076 S.n1858 VSUBS 0.24fF $ **FLOATING
C2077 S.n1859 VSUBS 0.91fF $ **FLOATING
C2078 S.n1860 VSUBS 0.05fF $ **FLOATING
C2079 S.t2059 VSUBS 0.02fF
C2080 S.n1861 VSUBS 0.12fF $ **FLOATING
C2081 S.n1862 VSUBS 0.14fF $ **FLOATING
C2082 S.n1864 VSUBS 0.25fF $ **FLOATING
C2083 S.n1865 VSUBS 0.09fF $ **FLOATING
C2084 S.n1866 VSUBS 0.21fF $ **FLOATING
C2085 S.n1867 VSUBS 0.92fF $ **FLOATING
C2086 S.n1868 VSUBS 0.44fF $ **FLOATING
C2087 S.n1869 VSUBS 1.88fF $ **FLOATING
C2088 S.n1870 VSUBS 0.12fF $ **FLOATING
C2089 S.t2097 VSUBS 0.02fF
C2090 S.n1871 VSUBS 0.14fF $ **FLOATING
C2091 S.t74 VSUBS 0.02fF
C2092 S.n1873 VSUBS 0.24fF $ **FLOATING
C2093 S.n1874 VSUBS 0.36fF $ **FLOATING
C2094 S.n1875 VSUBS 0.61fF $ **FLOATING
C2095 S.n1876 VSUBS 0.02fF $ **FLOATING
C2096 S.n1877 VSUBS 0.01fF $ **FLOATING
C2097 S.n1878 VSUBS 0.02fF $ **FLOATING
C2098 S.n1879 VSUBS 0.08fF $ **FLOATING
C2099 S.n1880 VSUBS 0.06fF $ **FLOATING
C2100 S.n1881 VSUBS 0.03fF $ **FLOATING
C2101 S.n1882 VSUBS 0.04fF $ **FLOATING
C2102 S.n1883 VSUBS 1.00fF $ **FLOATING
C2103 S.n1884 VSUBS 0.36fF $ **FLOATING
C2104 S.n1885 VSUBS 1.87fF $ **FLOATING
C2105 S.n1886 VSUBS 1.99fF $ **FLOATING
C2106 S.t666 VSUBS 0.02fF
C2107 S.n1887 VSUBS 0.24fF $ **FLOATING
C2108 S.n1888 VSUBS 0.91fF $ **FLOATING
C2109 S.n1889 VSUBS 0.05fF $ **FLOATING
C2110 S.t444 VSUBS 0.02fF
C2111 S.n1890 VSUBS 0.12fF $ **FLOATING
C2112 S.n1891 VSUBS 0.14fF $ **FLOATING
C2113 S.n1893 VSUBS 1.89fF $ **FLOATING
C2114 S.n1894 VSUBS 0.06fF $ **FLOATING
C2115 S.n1895 VSUBS 0.03fF $ **FLOATING
C2116 S.n1896 VSUBS 0.04fF $ **FLOATING
C2117 S.n1897 VSUBS 0.99fF $ **FLOATING
C2118 S.n1898 VSUBS 0.02fF $ **FLOATING
C2119 S.n1899 VSUBS 0.01fF $ **FLOATING
C2120 S.n1900 VSUBS 0.02fF $ **FLOATING
C2121 S.n1901 VSUBS 0.08fF $ **FLOATING
C2122 S.n1902 VSUBS 0.36fF $ **FLOATING
C2123 S.n1903 VSUBS 1.85fF $ **FLOATING
C2124 S.t2237 VSUBS 0.02fF
C2125 S.n1904 VSUBS 0.24fF $ **FLOATING
C2126 S.n1905 VSUBS 0.36fF $ **FLOATING
C2127 S.n1906 VSUBS 0.61fF $ **FLOATING
C2128 S.n1907 VSUBS 0.12fF $ **FLOATING
C2129 S.t1701 VSUBS 0.02fF
C2130 S.n1908 VSUBS 0.14fF $ **FLOATING
C2131 S.n1910 VSUBS 0.70fF $ **FLOATING
C2132 S.n1911 VSUBS 0.23fF $ **FLOATING
C2133 S.n1912 VSUBS 0.23fF $ **FLOATING
C2134 S.n1913 VSUBS 0.70fF $ **FLOATING
C2135 S.n1914 VSUBS 1.16fF $ **FLOATING
C2136 S.n1915 VSUBS 0.22fF $ **FLOATING
C2137 S.n1916 VSUBS 0.25fF $ **FLOATING
C2138 S.n1917 VSUBS 0.09fF $ **FLOATING
C2139 S.n1918 VSUBS 1.88fF $ **FLOATING
C2140 S.t296 VSUBS 0.02fF
C2141 S.n1919 VSUBS 0.24fF $ **FLOATING
C2142 S.n1920 VSUBS 0.91fF $ **FLOATING
C2143 S.n1921 VSUBS 0.05fF $ **FLOATING
C2144 S.t1235 VSUBS 0.02fF
C2145 S.n1922 VSUBS 0.12fF $ **FLOATING
C2146 S.n1923 VSUBS 0.14fF $ **FLOATING
C2147 S.n1925 VSUBS 0.25fF $ **FLOATING
C2148 S.n1926 VSUBS 0.09fF $ **FLOATING
C2149 S.n1927 VSUBS 0.21fF $ **FLOATING
C2150 S.n1928 VSUBS 0.92fF $ **FLOATING
C2151 S.n1929 VSUBS 0.44fF $ **FLOATING
C2152 S.n1930 VSUBS 1.88fF $ **FLOATING
C2153 S.n1931 VSUBS 0.12fF $ **FLOATING
C2154 S.t2490 VSUBS 0.02fF
C2155 S.n1932 VSUBS 0.14fF $ **FLOATING
C2156 S.t1077 VSUBS 0.02fF
C2157 S.n1934 VSUBS 0.24fF $ **FLOATING
C2158 S.n1935 VSUBS 0.91fF $ **FLOATING
C2159 S.n1936 VSUBS 0.05fF $ **FLOATING
C2160 S.t505 VSUBS 0.02fF
C2161 S.n1937 VSUBS 0.24fF $ **FLOATING
C2162 S.n1938 VSUBS 0.36fF $ **FLOATING
C2163 S.n1939 VSUBS 0.61fF $ **FLOATING
C2164 S.n1940 VSUBS 0.02fF $ **FLOATING
C2165 S.n1941 VSUBS 0.01fF $ **FLOATING
C2166 S.n1942 VSUBS 0.02fF $ **FLOATING
C2167 S.n1943 VSUBS 0.08fF $ **FLOATING
C2168 S.n1944 VSUBS 0.06fF $ **FLOATING
C2169 S.n1945 VSUBS 0.03fF $ **FLOATING
C2170 S.n1946 VSUBS 0.04fF $ **FLOATING
C2171 S.n1947 VSUBS 1.00fF $ **FLOATING
C2172 S.n1948 VSUBS 0.36fF $ **FLOATING
C2173 S.n1949 VSUBS 1.87fF $ **FLOATING
C2174 S.n1950 VSUBS 1.99fF $ **FLOATING
C2175 S.t836 VSUBS 0.02fF
C2176 S.n1951 VSUBS 0.12fF $ **FLOATING
C2177 S.n1952 VSUBS 0.14fF $ **FLOATING
C2178 S.n1954 VSUBS 1.89fF $ **FLOATING
C2179 S.n1955 VSUBS 0.06fF $ **FLOATING
C2180 S.n1956 VSUBS 0.03fF $ **FLOATING
C2181 S.n1957 VSUBS 0.04fF $ **FLOATING
C2182 S.n1958 VSUBS 0.99fF $ **FLOATING
C2183 S.n1959 VSUBS 0.02fF $ **FLOATING
C2184 S.n1960 VSUBS 0.01fF $ **FLOATING
C2185 S.n1961 VSUBS 0.02fF $ **FLOATING
C2186 S.n1962 VSUBS 0.08fF $ **FLOATING
C2187 S.n1963 VSUBS 0.36fF $ **FLOATING
C2188 S.n1964 VSUBS 1.85fF $ **FLOATING
C2189 S.t1289 VSUBS 0.02fF
C2190 S.n1965 VSUBS 0.24fF $ **FLOATING
C2191 S.n1966 VSUBS 0.36fF $ **FLOATING
C2192 S.n1967 VSUBS 0.61fF $ **FLOATING
C2193 S.n1968 VSUBS 0.12fF $ **FLOATING
C2194 S.t744 VSUBS 0.02fF
C2195 S.n1969 VSUBS 0.14fF $ **FLOATING
C2196 S.n1971 VSUBS 0.70fF $ **FLOATING
C2197 S.n1972 VSUBS 0.23fF $ **FLOATING
C2198 S.n1973 VSUBS 0.23fF $ **FLOATING
C2199 S.n1974 VSUBS 0.70fF $ **FLOATING
C2200 S.n1975 VSUBS 1.16fF $ **FLOATING
C2201 S.n1976 VSUBS 0.22fF $ **FLOATING
C2202 S.n1977 VSUBS 0.25fF $ **FLOATING
C2203 S.n1978 VSUBS 0.09fF $ **FLOATING
C2204 S.n1979 VSUBS 1.88fF $ **FLOATING
C2205 S.t1858 VSUBS 0.02fF
C2206 S.n1980 VSUBS 0.24fF $ **FLOATING
C2207 S.n1981 VSUBS 0.91fF $ **FLOATING
C2208 S.n1982 VSUBS 0.05fF $ **FLOATING
C2209 S.t1617 VSUBS 0.02fF
C2210 S.n1983 VSUBS 0.12fF $ **FLOATING
C2211 S.n1984 VSUBS 0.14fF $ **FLOATING
C2212 S.n1986 VSUBS 0.25fF $ **FLOATING
C2213 S.n1987 VSUBS 0.09fF $ **FLOATING
C2214 S.n1988 VSUBS 0.21fF $ **FLOATING
C2215 S.n1989 VSUBS 0.92fF $ **FLOATING
C2216 S.n1990 VSUBS 0.44fF $ **FLOATING
C2217 S.n1991 VSUBS 1.88fF $ **FLOATING
C2218 S.n1992 VSUBS 0.12fF $ **FLOATING
C2219 S.t1536 VSUBS 0.02fF
C2220 S.n1993 VSUBS 0.14fF $ **FLOATING
C2221 S.t2079 VSUBS 0.02fF
C2222 S.n1995 VSUBS 0.24fF $ **FLOATING
C2223 S.n1996 VSUBS 0.36fF $ **FLOATING
C2224 S.n1997 VSUBS 0.61fF $ **FLOATING
C2225 S.n1998 VSUBS 0.02fF $ **FLOATING
C2226 S.n1999 VSUBS 0.01fF $ **FLOATING
C2227 S.n2000 VSUBS 0.02fF $ **FLOATING
C2228 S.n2001 VSUBS 0.08fF $ **FLOATING
C2229 S.n2002 VSUBS 0.06fF $ **FLOATING
C2230 S.n2003 VSUBS 0.03fF $ **FLOATING
C2231 S.n2004 VSUBS 0.04fF $ **FLOATING
C2232 S.n2005 VSUBS 1.00fF $ **FLOATING
C2233 S.n2006 VSUBS 0.36fF $ **FLOATING
C2234 S.n2007 VSUBS 1.87fF $ **FLOATING
C2235 S.n2008 VSUBS 1.99fF $ **FLOATING
C2236 S.t98 VSUBS 0.02fF
C2237 S.n2009 VSUBS 0.24fF $ **FLOATING
C2238 S.n2010 VSUBS 0.91fF $ **FLOATING
C2239 S.n2011 VSUBS 0.05fF $ **FLOATING
C2240 S.t2405 VSUBS 0.02fF
C2241 S.n2012 VSUBS 0.12fF $ **FLOATING
C2242 S.n2013 VSUBS 0.14fF $ **FLOATING
C2243 S.n2015 VSUBS 1.89fF $ **FLOATING
C2244 S.n2016 VSUBS 0.06fF $ **FLOATING
C2245 S.n2017 VSUBS 0.03fF $ **FLOATING
C2246 S.n2018 VSUBS 0.04fF $ **FLOATING
C2247 S.n2019 VSUBS 0.99fF $ **FLOATING
C2248 S.n2020 VSUBS 0.02fF $ **FLOATING
C2249 S.n2021 VSUBS 0.01fF $ **FLOATING
C2250 S.n2022 VSUBS 0.02fF $ **FLOATING
C2251 S.n2023 VSUBS 0.08fF $ **FLOATING
C2252 S.n2024 VSUBS 0.36fF $ **FLOATING
C2253 S.n2025 VSUBS 1.85fF $ **FLOATING
C2254 S.t468 VSUBS 0.02fF
C2255 S.n2026 VSUBS 0.24fF $ **FLOATING
C2256 S.n2027 VSUBS 0.36fF $ **FLOATING
C2257 S.n2028 VSUBS 0.61fF $ **FLOATING
C2258 S.n2029 VSUBS 0.12fF $ **FLOATING
C2259 S.t2444 VSUBS 0.02fF
C2260 S.n2030 VSUBS 0.14fF $ **FLOATING
C2261 S.n2032 VSUBS 0.70fF $ **FLOATING
C2262 S.n2033 VSUBS 0.23fF $ **FLOATING
C2263 S.n2034 VSUBS 0.23fF $ **FLOATING
C2264 S.n2035 VSUBS 0.70fF $ **FLOATING
C2265 S.n2036 VSUBS 1.16fF $ **FLOATING
C2266 S.n2037 VSUBS 0.22fF $ **FLOATING
C2267 S.n2038 VSUBS 0.25fF $ **FLOATING
C2268 S.n2039 VSUBS 0.09fF $ **FLOATING
C2269 S.n2040 VSUBS 1.88fF $ **FLOATING
C2270 S.t1042 VSUBS 0.02fF
C2271 S.n2041 VSUBS 0.24fF $ **FLOATING
C2272 S.n2042 VSUBS 0.91fF $ **FLOATING
C2273 S.n2043 VSUBS 0.05fF $ **FLOATING
C2274 S.t788 VSUBS 0.02fF
C2275 S.n2044 VSUBS 0.12fF $ **FLOATING
C2276 S.n2045 VSUBS 0.14fF $ **FLOATING
C2277 S.n2047 VSUBS 0.25fF $ **FLOATING
C2278 S.n2048 VSUBS 0.09fF $ **FLOATING
C2279 S.n2049 VSUBS 0.21fF $ **FLOATING
C2280 S.n2050 VSUBS 0.92fF $ **FLOATING
C2281 S.n2051 VSUBS 0.44fF $ **FLOATING
C2282 S.n2052 VSUBS 1.88fF $ **FLOATING
C2283 S.n2053 VSUBS 0.12fF $ **FLOATING
C2284 S.t2072 VSUBS 0.02fF
C2285 S.n2054 VSUBS 0.14fF $ **FLOATING
C2286 S.t22 VSUBS 0.02fF
C2287 S.n2056 VSUBS 0.24fF $ **FLOATING
C2288 S.n2057 VSUBS 0.36fF $ **FLOATING
C2289 S.n2058 VSUBS 0.61fF $ **FLOATING
C2290 S.n2059 VSUBS 0.02fF $ **FLOATING
C2291 S.n2060 VSUBS 0.01fF $ **FLOATING
C2292 S.n2061 VSUBS 0.02fF $ **FLOATING
C2293 S.n2062 VSUBS 0.08fF $ **FLOATING
C2294 S.n2063 VSUBS 0.06fF $ **FLOATING
C2295 S.n2064 VSUBS 0.03fF $ **FLOATING
C2296 S.n2065 VSUBS 0.04fF $ **FLOATING
C2297 S.n2066 VSUBS 1.00fF $ **FLOATING
C2298 S.n2067 VSUBS 0.36fF $ **FLOATING
C2299 S.n2068 VSUBS 1.87fF $ **FLOATING
C2300 S.n2069 VSUBS 1.99fF $ **FLOATING
C2301 S.t641 VSUBS 0.02fF
C2302 S.n2070 VSUBS 0.24fF $ **FLOATING
C2303 S.n2071 VSUBS 0.91fF $ **FLOATING
C2304 S.n2072 VSUBS 0.05fF $ **FLOATING
C2305 S.t419 VSUBS 0.02fF
C2306 S.n2073 VSUBS 0.12fF $ **FLOATING
C2307 S.n2074 VSUBS 0.14fF $ **FLOATING
C2308 S.n2076 VSUBS 1.89fF $ **FLOATING
C2309 S.n2077 VSUBS 0.06fF $ **FLOATING
C2310 S.n2078 VSUBS 0.03fF $ **FLOATING
C2311 S.n2079 VSUBS 0.04fF $ **FLOATING
C2312 S.n2080 VSUBS 0.99fF $ **FLOATING
C2313 S.n2081 VSUBS 0.02fF $ **FLOATING
C2314 S.n2082 VSUBS 0.01fF $ **FLOATING
C2315 S.n2083 VSUBS 0.02fF $ **FLOATING
C2316 S.n2084 VSUBS 0.08fF $ **FLOATING
C2317 S.n2085 VSUBS 0.36fF $ **FLOATING
C2318 S.n2086 VSUBS 1.85fF $ **FLOATING
C2319 S.t857 VSUBS 0.02fF
C2320 S.n2087 VSUBS 0.24fF $ **FLOATING
C2321 S.n2088 VSUBS 0.36fF $ **FLOATING
C2322 S.n2089 VSUBS 0.61fF $ **FLOATING
C2323 S.n2090 VSUBS 0.12fF $ **FLOATING
C2324 S.t342 VSUBS 0.02fF
C2325 S.n2091 VSUBS 0.14fF $ **FLOATING
C2326 S.n2093 VSUBS 0.70fF $ **FLOATING
C2327 S.n2094 VSUBS 0.23fF $ **FLOATING
C2328 S.n2095 VSUBS 0.23fF $ **FLOATING
C2329 S.n2096 VSUBS 0.70fF $ **FLOATING
C2330 S.n2097 VSUBS 1.16fF $ **FLOATING
C2331 S.n2098 VSUBS 0.22fF $ **FLOATING
C2332 S.n2099 VSUBS 0.25fF $ **FLOATING
C2333 S.n2100 VSUBS 0.09fF $ **FLOATING
C2334 S.n2101 VSUBS 1.88fF $ **FLOATING
C2335 S.t1428 VSUBS 0.02fF
C2336 S.n2102 VSUBS 0.24fF $ **FLOATING
C2337 S.n2103 VSUBS 0.91fF $ **FLOATING
C2338 S.n2104 VSUBS 0.05fF $ **FLOATING
C2339 S.t1211 VSUBS 0.02fF
C2340 S.n2105 VSUBS 0.12fF $ **FLOATING
C2341 S.n2106 VSUBS 0.14fF $ **FLOATING
C2342 S.n2108 VSUBS 0.25fF $ **FLOATING
C2343 S.n2109 VSUBS 0.09fF $ **FLOATING
C2344 S.n2110 VSUBS 0.21fF $ **FLOATING
C2345 S.n2111 VSUBS 0.92fF $ **FLOATING
C2346 S.n2112 VSUBS 0.44fF $ **FLOATING
C2347 S.n2113 VSUBS 1.88fF $ **FLOATING
C2348 S.n2114 VSUBS 0.12fF $ **FLOATING
C2349 S.t1129 VSUBS 0.02fF
C2350 S.n2115 VSUBS 0.14fF $ **FLOATING
C2351 S.t1641 VSUBS 0.02fF
C2352 S.n2117 VSUBS 0.24fF $ **FLOATING
C2353 S.n2118 VSUBS 0.36fF $ **FLOATING
C2354 S.n2119 VSUBS 0.61fF $ **FLOATING
C2355 S.n2120 VSUBS 0.02fF $ **FLOATING
C2356 S.n2121 VSUBS 0.01fF $ **FLOATING
C2357 S.n2122 VSUBS 0.02fF $ **FLOATING
C2358 S.n2123 VSUBS 0.08fF $ **FLOATING
C2359 S.n2124 VSUBS 0.06fF $ **FLOATING
C2360 S.n2125 VSUBS 0.03fF $ **FLOATING
C2361 S.n2126 VSUBS 0.04fF $ **FLOATING
C2362 S.n2127 VSUBS 1.00fF $ **FLOATING
C2363 S.n2128 VSUBS 0.36fF $ **FLOATING
C2364 S.n2129 VSUBS 1.83fF $ **FLOATING
C2365 S.n2130 VSUBS 1.99fF $ **FLOATING
C2366 S.t2218 VSUBS 0.02fF
C2367 S.n2131 VSUBS 0.24fF $ **FLOATING
C2368 S.n2132 VSUBS 0.91fF $ **FLOATING
C2369 S.n2133 VSUBS 0.05fF $ **FLOATING
C2370 S.t1990 VSUBS 0.02fF
C2371 S.n2134 VSUBS 0.12fF $ **FLOATING
C2372 S.n2135 VSUBS 0.14fF $ **FLOATING
C2373 S.n2137 VSUBS 1.89fF $ **FLOATING
C2374 S.n2138 VSUBS 0.63fF $ **FLOATING
C2375 S.n2139 VSUBS 0.07fF $ **FLOATING
C2376 S.n2140 VSUBS 0.04fF $ **FLOATING
C2377 S.n2141 VSUBS 0.05fF $ **FLOATING
C2378 S.n2142 VSUBS 0.87fF $ **FLOATING
C2379 S.n2143 VSUBS 0.01fF $ **FLOATING
C2380 S.n2144 VSUBS 0.01fF $ **FLOATING
C2381 S.n2145 VSUBS 0.01fF $ **FLOATING
C2382 S.n2146 VSUBS 0.07fF $ **FLOATING
C2383 S.n2147 VSUBS 0.68fF $ **FLOATING
C2384 S.n2148 VSUBS 0.13fF $ **FLOATING
C2385 S.t2425 VSUBS 0.02fF
C2386 S.n2149 VSUBS 0.24fF $ **FLOATING
C2387 S.n2150 VSUBS 0.36fF $ **FLOATING
C2388 S.n2151 VSUBS 0.61fF $ **FLOATING
C2389 S.n2152 VSUBS 0.12fF $ **FLOATING
C2390 S.t1911 VSUBS 0.02fF
C2391 S.n2153 VSUBS 0.14fF $ **FLOATING
C2392 S.n2155 VSUBS 0.70fF $ **FLOATING
C2393 S.n2156 VSUBS 0.23fF $ **FLOATING
C2394 S.n2157 VSUBS 0.23fF $ **FLOATING
C2395 S.n2158 VSUBS 0.70fF $ **FLOATING
C2396 S.n2159 VSUBS 1.16fF $ **FLOATING
C2397 S.n2160 VSUBS 0.22fF $ **FLOATING
C2398 S.n2161 VSUBS 0.25fF $ **FLOATING
C2399 S.n2162 VSUBS 0.09fF $ **FLOATING
C2400 S.n2163 VSUBS 2.31fF $ **FLOATING
C2401 S.t484 VSUBS 0.02fF
C2402 S.n2164 VSUBS 0.24fF $ **FLOATING
C2403 S.n2165 VSUBS 0.91fF $ **FLOATING
C2404 S.n2166 VSUBS 0.05fF $ **FLOATING
C2405 S.t260 VSUBS 0.02fF
C2406 S.n2167 VSUBS 0.12fF $ **FLOATING
C2407 S.n2168 VSUBS 0.14fF $ **FLOATING
C2408 S.n2170 VSUBS 1.88fF $ **FLOATING
C2409 S.n2171 VSUBS 0.46fF $ **FLOATING
C2410 S.n2172 VSUBS 0.22fF $ **FLOATING
C2411 S.n2173 VSUBS 0.38fF $ **FLOATING
C2412 S.n2174 VSUBS 0.16fF $ **FLOATING
C2413 S.n2175 VSUBS 0.28fF $ **FLOATING
C2414 S.n2176 VSUBS 0.21fF $ **FLOATING
C2415 S.n2177 VSUBS 0.30fF $ **FLOATING
C2416 S.n2178 VSUBS 0.42fF $ **FLOATING
C2417 S.n2179 VSUBS 0.21fF $ **FLOATING
C2418 S.t1220 VSUBS 0.02fF
C2419 S.n2180 VSUBS 0.24fF $ **FLOATING
C2420 S.n2181 VSUBS 0.36fF $ **FLOATING
C2421 S.n2182 VSUBS 0.61fF $ **FLOATING
C2422 S.n2183 VSUBS 0.12fF $ **FLOATING
C2423 S.t552 VSUBS 0.02fF
C2424 S.n2184 VSUBS 0.14fF $ **FLOATING
C2425 S.n2186 VSUBS 0.04fF $ **FLOATING
C2426 S.n2187 VSUBS 0.03fF $ **FLOATING
C2427 S.n2188 VSUBS 0.03fF $ **FLOATING
C2428 S.n2189 VSUBS 0.10fF $ **FLOATING
C2429 S.n2190 VSUBS 0.36fF $ **FLOATING
C2430 S.n2191 VSUBS 0.38fF $ **FLOATING
C2431 S.n2192 VSUBS 0.11fF $ **FLOATING
C2432 S.n2193 VSUBS 0.12fF $ **FLOATING
C2433 S.n2194 VSUBS 0.07fF $ **FLOATING
C2434 S.n2195 VSUBS 0.12fF $ **FLOATING
C2435 S.n2196 VSUBS 0.18fF $ **FLOATING
C2436 S.n2197 VSUBS 3.99fF $ **FLOATING
C2437 S.t1207 VSUBS 0.02fF
C2438 S.n2198 VSUBS 0.24fF $ **FLOATING
C2439 S.n2199 VSUBS 0.91fF $ **FLOATING
C2440 S.n2200 VSUBS 0.05fF $ **FLOATING
C2441 S.t1168 VSUBS 0.02fF
C2442 S.n2201 VSUBS 0.12fF $ **FLOATING
C2443 S.n2202 VSUBS 0.14fF $ **FLOATING
C2444 S.n2204 VSUBS 0.25fF $ **FLOATING
C2445 S.n2205 VSUBS 0.09fF $ **FLOATING
C2446 S.n2206 VSUBS 0.21fF $ **FLOATING
C2447 S.n2207 VSUBS 1.28fF $ **FLOATING
C2448 S.n2208 VSUBS 0.53fF $ **FLOATING
C2449 S.n2209 VSUBS 1.88fF $ **FLOATING
C2450 S.n2210 VSUBS 0.12fF $ **FLOATING
C2451 S.t1341 VSUBS 0.02fF
C2452 S.n2211 VSUBS 0.14fF $ **FLOATING
C2453 S.t1997 VSUBS 0.02fF
C2454 S.n2213 VSUBS 0.24fF $ **FLOATING
C2455 S.n2214 VSUBS 0.36fF $ **FLOATING
C2456 S.n2215 VSUBS 0.61fF $ **FLOATING
C2457 S.n2216 VSUBS 0.71fF $ **FLOATING
C2458 S.n2217 VSUBS 1.58fF $ **FLOATING
C2459 S.n2218 VSUBS 2.45fF $ **FLOATING
C2460 S.t1985 VSUBS 0.02fF
C2461 S.n2219 VSUBS 0.24fF $ **FLOATING
C2462 S.n2220 VSUBS 0.91fF $ **FLOATING
C2463 S.n2221 VSUBS 0.05fF $ **FLOATING
C2464 S.t2206 VSUBS 0.02fF
C2465 S.n2222 VSUBS 0.12fF $ **FLOATING
C2466 S.n2223 VSUBS 0.14fF $ **FLOATING
C2467 S.n2225 VSUBS 1.89fF $ **FLOATING
C2468 S.n2226 VSUBS 0.06fF $ **FLOATING
C2469 S.n2227 VSUBS 0.03fF $ **FLOATING
C2470 S.n2228 VSUBS 0.04fF $ **FLOATING
C2471 S.n2229 VSUBS 0.99fF $ **FLOATING
C2472 S.n2230 VSUBS 0.02fF $ **FLOATING
C2473 S.n2231 VSUBS 0.01fF $ **FLOATING
C2474 S.n2232 VSUBS 0.02fF $ **FLOATING
C2475 S.n2233 VSUBS 0.08fF $ **FLOATING
C2476 S.n2234 VSUBS 0.36fF $ **FLOATING
C2477 S.n2235 VSUBS 1.85fF $ **FLOATING
C2478 S.t268 VSUBS 0.02fF
C2479 S.n2236 VSUBS 0.24fF $ **FLOATING
C2480 S.n2237 VSUBS 0.36fF $ **FLOATING
C2481 S.n2238 VSUBS 0.61fF $ **FLOATING
C2482 S.n2239 VSUBS 0.12fF $ **FLOATING
C2483 S.t2127 VSUBS 0.02fF
C2484 S.n2240 VSUBS 0.14fF $ **FLOATING
C2485 S.n2242 VSUBS 0.70fF $ **FLOATING
C2486 S.n2243 VSUBS 0.23fF $ **FLOATING
C2487 S.n2244 VSUBS 0.23fF $ **FLOATING
C2488 S.n2245 VSUBS 0.70fF $ **FLOATING
C2489 S.n2246 VSUBS 1.16fF $ **FLOATING
C2490 S.n2247 VSUBS 0.22fF $ **FLOATING
C2491 S.n2248 VSUBS 0.25fF $ **FLOATING
C2492 S.n2249 VSUBS 0.09fF $ **FLOATING
C2493 S.n2250 VSUBS 1.88fF $ **FLOATING
C2494 S.t251 VSUBS 0.02fF
C2495 S.n2251 VSUBS 0.24fF $ **FLOATING
C2496 S.n2252 VSUBS 0.91fF $ **FLOATING
C2497 S.n2253 VSUBS 0.05fF $ **FLOATING
C2498 S.t472 VSUBS 0.02fF
C2499 S.n2254 VSUBS 0.12fF $ **FLOATING
C2500 S.n2255 VSUBS 0.14fF $ **FLOATING
C2501 S.n2257 VSUBS 20.78fF $ **FLOATING
C2502 S.n2258 VSUBS 0.06fF $ **FLOATING
C2503 S.n2259 VSUBS 0.20fF $ **FLOATING
C2504 S.n2260 VSUBS 0.09fF $ **FLOATING
C2505 S.n2261 VSUBS 0.21fF $ **FLOATING
C2506 S.n2262 VSUBS 0.10fF $ **FLOATING
C2507 S.n2263 VSUBS 0.30fF $ **FLOATING
C2508 S.n2264 VSUBS 0.69fF $ **FLOATING
C2509 S.n2265 VSUBS 0.45fF $ **FLOATING
C2510 S.n2266 VSUBS 2.33fF $ **FLOATING
C2511 S.n2267 VSUBS 0.12fF $ **FLOATING
C2512 S.t404 VSUBS 0.02fF
C2513 S.n2268 VSUBS 0.14fF $ **FLOATING
C2514 S.t930 VSUBS 0.02fF
C2515 S.n2270 VSUBS 0.24fF $ **FLOATING
C2516 S.n2271 VSUBS 0.36fF $ **FLOATING
C2517 S.n2272 VSUBS 0.61fF $ **FLOATING
C2518 S.n2273 VSUBS 1.90fF $ **FLOATING
C2519 S.n2274 VSUBS 0.17fF $ **FLOATING
C2520 S.n2275 VSUBS 0.76fF $ **FLOATING
C2521 S.n2276 VSUBS 0.32fF $ **FLOATING
C2522 S.n2277 VSUBS 0.25fF $ **FLOATING
C2523 S.n2278 VSUBS 0.30fF $ **FLOATING
C2524 S.n2279 VSUBS 0.47fF $ **FLOATING
C2525 S.n2280 VSUBS 0.16fF $ **FLOATING
C2526 S.n2281 VSUBS 1.93fF $ **FLOATING
C2527 S.t1269 VSUBS 0.02fF
C2528 S.n2282 VSUBS 0.12fF $ **FLOATING
C2529 S.n2283 VSUBS 0.14fF $ **FLOATING
C2530 S.t1493 VSUBS 0.02fF
C2531 S.n2285 VSUBS 0.24fF $ **FLOATING
C2532 S.n2286 VSUBS 0.91fF $ **FLOATING
C2533 S.n2287 VSUBS 0.05fF $ **FLOATING
C2534 S.n2288 VSUBS 1.88fF $ **FLOATING
C2535 S.n2289 VSUBS 0.12fF $ **FLOATING
C2536 S.t1273 VSUBS 0.02fF
C2537 S.n2290 VSUBS 0.14fF $ **FLOATING
C2538 S.t2139 VSUBS 0.02fF
C2539 S.n2292 VSUBS 0.12fF $ **FLOATING
C2540 S.n2293 VSUBS 0.14fF $ **FLOATING
C2541 S.t1919 VSUBS 0.02fF
C2542 S.n2295 VSUBS 0.24fF $ **FLOATING
C2543 S.n2296 VSUBS 0.91fF $ **FLOATING
C2544 S.n2297 VSUBS 0.05fF $ **FLOATING
C2545 S.t1076 VSUBS 0.02fF
C2546 S.n2298 VSUBS 0.24fF $ **FLOATING
C2547 S.n2299 VSUBS 0.36fF $ **FLOATING
C2548 S.n2300 VSUBS 0.61fF $ **FLOATING
C2549 S.n2301 VSUBS 0.32fF $ **FLOATING
C2550 S.n2302 VSUBS 1.09fF $ **FLOATING
C2551 S.n2303 VSUBS 0.15fF $ **FLOATING
C2552 S.n2304 VSUBS 2.10fF $ **FLOATING
C2553 S.n2305 VSUBS 2.94fF $ **FLOATING
C2554 S.n2306 VSUBS 1.88fF $ **FLOATING
C2555 S.n2307 VSUBS 0.12fF $ **FLOATING
C2556 S.t393 VSUBS 0.02fF
C2557 S.n2308 VSUBS 0.14fF $ **FLOATING
C2558 S.t1048 VSUBS 0.02fF
C2559 S.n2310 VSUBS 0.24fF $ **FLOATING
C2560 S.n2311 VSUBS 0.36fF $ **FLOATING
C2561 S.n2312 VSUBS 0.61fF $ **FLOATING
C2562 S.n2313 VSUBS 0.92fF $ **FLOATING
C2563 S.n2314 VSUBS 0.32fF $ **FLOATING
C2564 S.n2315 VSUBS 0.92fF $ **FLOATING
C2565 S.n2316 VSUBS 1.09fF $ **FLOATING
C2566 S.n2317 VSUBS 0.15fF $ **FLOATING
C2567 S.n2318 VSUBS 4.68fF $ **FLOATING
C2568 S.t1259 VSUBS 0.02fF
C2569 S.n2319 VSUBS 0.12fF $ **FLOATING
C2570 S.n2320 VSUBS 0.14fF $ **FLOATING
C2571 S.t1036 VSUBS 0.02fF
C2572 S.n2322 VSUBS 0.24fF $ **FLOATING
C2573 S.n2323 VSUBS 0.91fF $ **FLOATING
C2574 S.n2324 VSUBS 0.05fF $ **FLOATING
C2575 S.n2325 VSUBS 1.88fF $ **FLOATING
C2576 S.n2326 VSUBS 2.67fF $ **FLOATING
C2577 S.t1831 VSUBS 0.02fF
C2578 S.n2327 VSUBS 0.24fF $ **FLOATING
C2579 S.n2328 VSUBS 0.36fF $ **FLOATING
C2580 S.n2329 VSUBS 0.61fF $ **FLOATING
C2581 S.n2330 VSUBS 0.12fF $ **FLOATING
C2582 S.t1186 VSUBS 0.02fF
C2583 S.n2331 VSUBS 0.14fF $ **FLOATING
C2584 S.n2333 VSUBS 1.88fF $ **FLOATING
C2585 S.n2334 VSUBS 2.68fF $ **FLOATING
C2586 S.t1857 VSUBS 0.02fF
C2587 S.n2335 VSUBS 0.24fF $ **FLOATING
C2588 S.n2336 VSUBS 0.36fF $ **FLOATING
C2589 S.n2337 VSUBS 0.61fF $ **FLOATING
C2590 S.t1502 VSUBS 0.02fF
C2591 S.n2338 VSUBS 1.22fF $ **FLOATING
C2592 S.n2339 VSUBS 0.36fF $ **FLOATING
C2593 S.n2340 VSUBS 1.22fF $ **FLOATING
C2594 S.n2341 VSUBS 0.61fF $ **FLOATING
C2595 S.n2342 VSUBS 0.35fF $ **FLOATING
C2596 S.n2343 VSUBS 0.63fF $ **FLOATING
C2597 S.n2344 VSUBS 1.15fF $ **FLOATING
C2598 S.n2345 VSUBS 3.00fF $ **FLOATING
C2599 S.n2346 VSUBS 0.59fF $ **FLOATING
C2600 S.n2347 VSUBS 0.01fF $ **FLOATING
C2601 S.n2348 VSUBS 0.97fF $ **FLOATING
C2602 S.t117 VSUBS 21.42fF
C2603 S.n2349 VSUBS 20.29fF $ **FLOATING
C2604 S.n2351 VSUBS 0.38fF $ **FLOATING
C2605 S.n2352 VSUBS 0.23fF $ **FLOATING
C2606 S.n2353 VSUBS 2.79fF $ **FLOATING
C2607 S.n2354 VSUBS 2.46fF $ **FLOATING
C2608 S.n2355 VSUBS 4.00fF $ **FLOATING
C2609 S.n2356 VSUBS 0.25fF $ **FLOATING
C2610 S.n2357 VSUBS 0.01fF $ **FLOATING
C2611 S.t687 VSUBS 0.02fF
C2612 S.n2358 VSUBS 0.26fF $ **FLOATING
C2613 S.t1794 VSUBS 0.02fF
C2614 S.n2359 VSUBS 0.95fF $ **FLOATING
C2615 S.n2360 VSUBS 0.71fF $ **FLOATING
C2616 S.n2361 VSUBS 1.89fF $ **FLOATING
C2617 S.n2362 VSUBS 1.88fF $ **FLOATING
C2618 S.t2291 VSUBS 0.02fF
C2619 S.n2363 VSUBS 0.24fF $ **FLOATING
C2620 S.n2364 VSUBS 0.36fF $ **FLOATING
C2621 S.n2365 VSUBS 0.61fF $ **FLOATING
C2622 S.n2366 VSUBS 0.12fF $ **FLOATING
C2623 S.t1477 VSUBS 0.02fF
C2624 S.n2367 VSUBS 0.14fF $ **FLOATING
C2625 S.n2369 VSUBS 1.16fF $ **FLOATING
C2626 S.n2370 VSUBS 0.22fF $ **FLOATING
C2627 S.n2371 VSUBS 0.25fF $ **FLOATING
C2628 S.n2372 VSUBS 0.09fF $ **FLOATING
C2629 S.n2373 VSUBS 1.88fF $ **FLOATING
C2630 S.t2576 VSUBS 0.02fF
C2631 S.n2374 VSUBS 0.24fF $ **FLOATING
C2632 S.n2375 VSUBS 0.91fF $ **FLOATING
C2633 S.n2376 VSUBS 0.05fF $ **FLOATING
C2634 S.t2345 VSUBS 0.02fF
C2635 S.n2377 VSUBS 0.12fF $ **FLOATING
C2636 S.n2378 VSUBS 0.14fF $ **FLOATING
C2637 S.n2380 VSUBS 0.78fF $ **FLOATING
C2638 S.n2381 VSUBS 1.94fF $ **FLOATING
C2639 S.n2382 VSUBS 1.88fF $ **FLOATING
C2640 S.n2383 VSUBS 0.12fF $ **FLOATING
C2641 S.t2385 VSUBS 0.02fF
C2642 S.n2384 VSUBS 0.14fF $ **FLOATING
C2643 S.t559 VSUBS 0.02fF
C2644 S.n2386 VSUBS 0.24fF $ **FLOATING
C2645 S.n2387 VSUBS 0.36fF $ **FLOATING
C2646 S.n2388 VSUBS 0.61fF $ **FLOATING
C2647 S.n2389 VSUBS 1.84fF $ **FLOATING
C2648 S.n2390 VSUBS 2.99fF $ **FLOATING
C2649 S.t839 VSUBS 0.02fF
C2650 S.n2391 VSUBS 0.24fF $ **FLOATING
C2651 S.n2392 VSUBS 0.91fF $ **FLOATING
C2652 S.n2393 VSUBS 0.05fF $ **FLOATING
C2653 S.t608 VSUBS 0.02fF
C2654 S.n2394 VSUBS 0.12fF $ **FLOATING
C2655 S.n2395 VSUBS 0.14fF $ **FLOATING
C2656 S.n2397 VSUBS 1.89fF $ **FLOATING
C2657 S.n2398 VSUBS 1.88fF $ **FLOATING
C2658 S.t1465 VSUBS 0.02fF
C2659 S.n2399 VSUBS 0.24fF $ **FLOATING
C2660 S.n2400 VSUBS 0.36fF $ **FLOATING
C2661 S.n2401 VSUBS 0.61fF $ **FLOATING
C2662 S.n2402 VSUBS 0.12fF $ **FLOATING
C2663 S.t647 VSUBS 0.02fF
C2664 S.n2403 VSUBS 0.14fF $ **FLOATING
C2665 S.n2405 VSUBS 1.16fF $ **FLOATING
C2666 S.n2406 VSUBS 0.22fF $ **FLOATING
C2667 S.n2407 VSUBS 0.25fF $ **FLOATING
C2668 S.n2408 VSUBS 0.09fF $ **FLOATING
C2669 S.n2409 VSUBS 1.88fF $ **FLOATING
C2670 S.t1756 VSUBS 0.02fF
C2671 S.n2410 VSUBS 0.24fF $ **FLOATING
C2672 S.n2411 VSUBS 0.91fF $ **FLOATING
C2673 S.n2412 VSUBS 0.05fF $ **FLOATING
C2674 S.t1516 VSUBS 0.02fF
C2675 S.n2413 VSUBS 0.12fF $ **FLOATING
C2676 S.n2414 VSUBS 0.14fF $ **FLOATING
C2677 S.n2416 VSUBS 0.78fF $ **FLOATING
C2678 S.n2417 VSUBS 1.94fF $ **FLOATING
C2679 S.n2418 VSUBS 1.88fF $ **FLOATING
C2680 S.n2419 VSUBS 0.12fF $ **FLOATING
C2681 S.t281 VSUBS 0.02fF
C2682 S.n2420 VSUBS 0.14fF $ **FLOATING
C2683 S.t1091 VSUBS 0.02fF
C2684 S.n2422 VSUBS 0.24fF $ **FLOATING
C2685 S.n2423 VSUBS 0.36fF $ **FLOATING
C2686 S.n2424 VSUBS 0.61fF $ **FLOATING
C2687 S.n2425 VSUBS 1.84fF $ **FLOATING
C2688 S.n2426 VSUBS 2.99fF $ **FLOATING
C2689 S.t1371 VSUBS 0.02fF
C2690 S.n2427 VSUBS 0.24fF $ **FLOATING
C2691 S.n2428 VSUBS 0.91fF $ **FLOATING
C2692 S.n2429 VSUBS 0.05fF $ **FLOATING
C2693 S.t1148 VSUBS 0.02fF
C2694 S.n2430 VSUBS 0.12fF $ **FLOATING
C2695 S.n2431 VSUBS 0.14fF $ **FLOATING
C2696 S.n2433 VSUBS 1.89fF $ **FLOATING
C2697 S.n2434 VSUBS 1.88fF $ **FLOATING
C2698 S.t1872 VSUBS 0.02fF
C2699 S.n2435 VSUBS 0.24fF $ **FLOATING
C2700 S.n2436 VSUBS 0.36fF $ **FLOATING
C2701 S.n2437 VSUBS 0.61fF $ **FLOATING
C2702 S.n2438 VSUBS 0.12fF $ **FLOATING
C2703 S.t1062 VSUBS 0.02fF
C2704 S.n2439 VSUBS 0.14fF $ **FLOATING
C2705 S.n2441 VSUBS 1.16fF $ **FLOATING
C2706 S.n2442 VSUBS 0.22fF $ **FLOATING
C2707 S.n2443 VSUBS 0.25fF $ **FLOATING
C2708 S.n2444 VSUBS 0.09fF $ **FLOATING
C2709 S.n2445 VSUBS 1.88fF $ **FLOATING
C2710 S.t2157 VSUBS 0.02fF
C2711 S.n2446 VSUBS 0.24fF $ **FLOATING
C2712 S.n2447 VSUBS 0.91fF $ **FLOATING
C2713 S.n2448 VSUBS 0.05fF $ **FLOATING
C2714 S.t1930 VSUBS 0.02fF
C2715 S.n2449 VSUBS 0.12fF $ **FLOATING
C2716 S.n2450 VSUBS 0.14fF $ **FLOATING
C2717 S.n2452 VSUBS 0.78fF $ **FLOATING
C2718 S.n2453 VSUBS 1.94fF $ **FLOATING
C2719 S.n2454 VSUBS 1.88fF $ **FLOATING
C2720 S.n2455 VSUBS 0.12fF $ **FLOATING
C2721 S.t1846 VSUBS 0.02fF
C2722 S.n2456 VSUBS 0.14fF $ **FLOATING
C2723 S.t118 VSUBS 0.02fF
C2724 S.n2458 VSUBS 0.24fF $ **FLOATING
C2725 S.n2459 VSUBS 0.36fF $ **FLOATING
C2726 S.n2460 VSUBS 0.61fF $ **FLOATING
C2727 S.n2461 VSUBS 1.84fF $ **FLOATING
C2728 S.n2462 VSUBS 2.99fF $ **FLOATING
C2729 S.t425 VSUBS 0.02fF
C2730 S.n2463 VSUBS 0.24fF $ **FLOATING
C2731 S.n2464 VSUBS 0.91fF $ **FLOATING
C2732 S.n2465 VSUBS 0.05fF $ **FLOATING
C2733 S.t188 VSUBS 0.02fF
C2734 S.n2466 VSUBS 0.12fF $ **FLOATING
C2735 S.n2467 VSUBS 0.14fF $ **FLOATING
C2736 S.n2469 VSUBS 1.89fF $ **FLOATING
C2737 S.n2470 VSUBS 1.88fF $ **FLOATING
C2738 S.t919 VSUBS 0.02fF
C2739 S.n2471 VSUBS 0.24fF $ **FLOATING
C2740 S.n2472 VSUBS 0.36fF $ **FLOATING
C2741 S.n2473 VSUBS 0.61fF $ **FLOATING
C2742 S.n2474 VSUBS 0.12fF $ **FLOATING
C2743 S.t237 VSUBS 0.02fF
C2744 S.n2475 VSUBS 0.14fF $ **FLOATING
C2745 S.n2477 VSUBS 1.16fF $ **FLOATING
C2746 S.n2478 VSUBS 0.22fF $ **FLOATING
C2747 S.n2479 VSUBS 0.25fF $ **FLOATING
C2748 S.n2480 VSUBS 0.09fF $ **FLOATING
C2749 S.n2481 VSUBS 1.88fF $ **FLOATING
C2750 S.t1219 VSUBS 0.02fF
C2751 S.n2482 VSUBS 0.24fF $ **FLOATING
C2752 S.n2483 VSUBS 0.91fF $ **FLOATING
C2753 S.n2484 VSUBS 0.05fF $ **FLOATING
C2754 S.t975 VSUBS 0.02fF
C2755 S.n2485 VSUBS 0.12fF $ **FLOATING
C2756 S.n2486 VSUBS 0.14fF $ **FLOATING
C2757 S.n2488 VSUBS 0.78fF $ **FLOATING
C2758 S.n2489 VSUBS 1.94fF $ **FLOATING
C2759 S.n2490 VSUBS 1.88fF $ **FLOATING
C2760 S.n2491 VSUBS 0.12fF $ **FLOATING
C2761 S.t2355 VSUBS 0.02fF
C2762 S.n2492 VSUBS 0.14fF $ **FLOATING
C2763 S.t648 VSUBS 0.02fF
C2764 S.n2494 VSUBS 0.24fF $ **FLOATING
C2765 S.n2495 VSUBS 0.36fF $ **FLOATING
C2766 S.n2496 VSUBS 0.61fF $ **FLOATING
C2767 S.n2497 VSUBS 1.84fF $ **FLOATING
C2768 S.n2498 VSUBS 2.99fF $ **FLOATING
C2769 S.t941 VSUBS 0.02fF
C2770 S.n2499 VSUBS 0.24fF $ **FLOATING
C2771 S.n2500 VSUBS 0.91fF $ **FLOATING
C2772 S.n2501 VSUBS 0.05fF $ **FLOATING
C2773 S.t1889 VSUBS 0.02fF
C2774 S.n2502 VSUBS 0.12fF $ **FLOATING
C2775 S.n2503 VSUBS 0.14fF $ **FLOATING
C2776 S.n2505 VSUBS 1.89fF $ **FLOATING
C2777 S.n2506 VSUBS 1.88fF $ **FLOATING
C2778 S.t1436 VSUBS 0.02fF
C2779 S.n2507 VSUBS 0.24fF $ **FLOATING
C2780 S.n2508 VSUBS 0.36fF $ **FLOATING
C2781 S.n2509 VSUBS 0.61fF $ **FLOATING
C2782 S.n2510 VSUBS 0.12fF $ **FLOATING
C2783 S.t622 VSUBS 0.02fF
C2784 S.n2511 VSUBS 0.14fF $ **FLOATING
C2785 S.n2513 VSUBS 1.16fF $ **FLOATING
C2786 S.n2514 VSUBS 0.22fF $ **FLOATING
C2787 S.n2515 VSUBS 0.25fF $ **FLOATING
C2788 S.n2516 VSUBS 0.09fF $ **FLOATING
C2789 S.n2517 VSUBS 1.88fF $ **FLOATING
C2790 S.t1723 VSUBS 0.02fF
C2791 S.n2518 VSUBS 0.24fF $ **FLOATING
C2792 S.n2519 VSUBS 0.91fF $ **FLOATING
C2793 S.n2520 VSUBS 0.05fF $ **FLOATING
C2794 S.t1491 VSUBS 0.02fF
C2795 S.n2521 VSUBS 0.12fF $ **FLOATING
C2796 S.n2522 VSUBS 0.14fF $ **FLOATING
C2797 S.n2524 VSUBS 0.78fF $ **FLOATING
C2798 S.n2525 VSUBS 1.94fF $ **FLOATING
C2799 S.n2526 VSUBS 1.88fF $ **FLOATING
C2800 S.n2527 VSUBS 0.12fF $ **FLOATING
C2801 S.t1412 VSUBS 0.02fF
C2802 S.n2528 VSUBS 0.14fF $ **FLOATING
C2803 S.t2226 VSUBS 0.02fF
C2804 S.n2530 VSUBS 0.24fF $ **FLOATING
C2805 S.n2531 VSUBS 0.36fF $ **FLOATING
C2806 S.n2532 VSUBS 0.61fF $ **FLOATING
C2807 S.n2533 VSUBS 1.84fF $ **FLOATING
C2808 S.n2534 VSUBS 2.99fF $ **FLOATING
C2809 S.t2511 VSUBS 0.02fF
C2810 S.n2535 VSUBS 0.24fF $ **FLOATING
C2811 S.n2536 VSUBS 0.91fF $ **FLOATING
C2812 S.n2537 VSUBS 0.05fF $ **FLOATING
C2813 S.t2275 VSUBS 0.02fF
C2814 S.n2538 VSUBS 0.12fF $ **FLOATING
C2815 S.n2539 VSUBS 0.14fF $ **FLOATING
C2816 S.n2541 VSUBS 1.89fF $ **FLOATING
C2817 S.n2542 VSUBS 1.75fF $ **FLOATING
C2818 S.t496 VSUBS 0.02fF
C2819 S.n2543 VSUBS 0.24fF $ **FLOATING
C2820 S.n2544 VSUBS 0.36fF $ **FLOATING
C2821 S.n2545 VSUBS 0.61fF $ **FLOATING
C2822 S.n2546 VSUBS 0.12fF $ **FLOATING
C2823 S.t2202 VSUBS 0.02fF
C2824 S.n2547 VSUBS 0.14fF $ **FLOATING
C2825 S.n2549 VSUBS 1.16fF $ **FLOATING
C2826 S.n2550 VSUBS 0.22fF $ **FLOATING
C2827 S.n2551 VSUBS 0.25fF $ **FLOATING
C2828 S.n2552 VSUBS 0.09fF $ **FLOATING
C2829 S.n2553 VSUBS 2.44fF $ **FLOATING
C2830 S.t771 VSUBS 0.02fF
C2831 S.n2554 VSUBS 0.24fF $ **FLOATING
C2832 S.n2555 VSUBS 0.91fF $ **FLOATING
C2833 S.n2556 VSUBS 0.05fF $ **FLOATING
C2834 S.t547 VSUBS 0.02fF
C2835 S.n2557 VSUBS 0.12fF $ **FLOATING
C2836 S.n2558 VSUBS 0.14fF $ **FLOATING
C2837 S.n2560 VSUBS 1.88fF $ **FLOATING
C2838 S.n2561 VSUBS 0.48fF $ **FLOATING
C2839 S.n2562 VSUBS 0.09fF $ **FLOATING
C2840 S.n2563 VSUBS 0.33fF $ **FLOATING
C2841 S.n2564 VSUBS 0.30fF $ **FLOATING
C2842 S.n2565 VSUBS 0.77fF $ **FLOATING
C2843 S.n2566 VSUBS 0.59fF $ **FLOATING
C2844 S.t1284 VSUBS 0.02fF
C2845 S.n2567 VSUBS 0.24fF $ **FLOATING
C2846 S.n2568 VSUBS 0.36fF $ **FLOATING
C2847 S.n2569 VSUBS 0.61fF $ **FLOATING
C2848 S.n2570 VSUBS 0.12fF $ **FLOATING
C2849 S.t585 VSUBS 0.02fF
C2850 S.n2571 VSUBS 0.14fF $ **FLOATING
C2851 S.n2573 VSUBS 2.61fF $ **FLOATING
C2852 S.n2574 VSUBS 2.15fF $ **FLOATING
C2853 S.t1558 VSUBS 0.02fF
C2854 S.n2575 VSUBS 0.24fF $ **FLOATING
C2855 S.n2576 VSUBS 0.91fF $ **FLOATING
C2856 S.n2577 VSUBS 0.05fF $ **FLOATING
C2857 S.t1335 VSUBS 0.02fF
C2858 S.n2578 VSUBS 0.12fF $ **FLOATING
C2859 S.n2579 VSUBS 0.14fF $ **FLOATING
C2860 S.n2581 VSUBS 0.78fF $ **FLOATING
C2861 S.n2582 VSUBS 2.30fF $ **FLOATING
C2862 S.n2583 VSUBS 1.88fF $ **FLOATING
C2863 S.n2584 VSUBS 0.12fF $ **FLOATING
C2864 S.t2219 VSUBS 0.02fF
C2865 S.n2585 VSUBS 0.14fF $ **FLOATING
C2866 S.t2019 VSUBS 0.02fF
C2867 S.n2587 VSUBS 0.24fF $ **FLOATING
C2868 S.n2588 VSUBS 0.36fF $ **FLOATING
C2869 S.n2589 VSUBS 0.61fF $ **FLOATING
C2870 S.n2590 VSUBS 1.39fF $ **FLOATING
C2871 S.n2591 VSUBS 0.71fF $ **FLOATING
C2872 S.n2592 VSUBS 1.14fF $ **FLOATING
C2873 S.n2593 VSUBS 0.35fF $ **FLOATING
C2874 S.n2594 VSUBS 2.02fF $ **FLOATING
C2875 S.t350 VSUBS 0.02fF
C2876 S.n2595 VSUBS 0.24fF $ **FLOATING
C2877 S.n2596 VSUBS 0.91fF $ **FLOATING
C2878 S.n2597 VSUBS 0.05fF $ **FLOATING
C2879 S.t564 VSUBS 0.02fF
C2880 S.n2598 VSUBS 0.12fF $ **FLOATING
C2881 S.n2599 VSUBS 0.14fF $ **FLOATING
C2882 S.n2601 VSUBS 1.89fF $ **FLOATING
C2883 S.n2602 VSUBS 1.88fF $ **FLOATING
C2884 S.t293 VSUBS 0.02fF
C2885 S.n2603 VSUBS 0.24fF $ **FLOATING
C2886 S.n2604 VSUBS 0.36fF $ **FLOATING
C2887 S.n2605 VSUBS 0.61fF $ **FLOATING
C2888 S.n2606 VSUBS 0.12fF $ **FLOATING
C2889 S.t485 VSUBS 0.02fF
C2890 S.n2607 VSUBS 0.14fF $ **FLOATING
C2891 S.n2609 VSUBS 1.16fF $ **FLOATING
C2892 S.n2610 VSUBS 0.22fF $ **FLOATING
C2893 S.n2611 VSUBS 0.25fF $ **FLOATING
C2894 S.n2612 VSUBS 0.09fF $ **FLOATING
C2895 S.n2613 VSUBS 1.88fF $ **FLOATING
C2896 S.t1138 VSUBS 0.02fF
C2897 S.n2614 VSUBS 0.24fF $ **FLOATING
C2898 S.n2615 VSUBS 0.91fF $ **FLOATING
C2899 S.n2616 VSUBS 0.05fF $ **FLOATING
C2900 S.t1352 VSUBS 0.02fF
C2901 S.n2617 VSUBS 0.12fF $ **FLOATING
C2902 S.n2618 VSUBS 0.14fF $ **FLOATING
C2903 S.n2620 VSUBS 20.78fF $ **FLOATING
C2904 S.n2621 VSUBS 2.73fF $ **FLOATING
C2905 S.n2622 VSUBS 1.59fF $ **FLOATING
C2906 S.n2623 VSUBS 0.12fF $ **FLOATING
C2907 S.t331 VSUBS 0.02fF
C2908 S.n2624 VSUBS 0.14fF $ **FLOATING
C2909 S.t1090 VSUBS 0.02fF
C2910 S.n2626 VSUBS 0.24fF $ **FLOATING
C2911 S.n2627 VSUBS 0.36fF $ **FLOATING
C2912 S.n2628 VSUBS 0.61fF $ **FLOATING
C2913 S.n2629 VSUBS 0.07fF $ **FLOATING
C2914 S.n2630 VSUBS 0.01fF $ **FLOATING
C2915 S.n2631 VSUBS 0.24fF $ **FLOATING
C2916 S.n2632 VSUBS 1.16fF $ **FLOATING
C2917 S.n2633 VSUBS 1.35fF $ **FLOATING
C2918 S.n2634 VSUBS 2.30fF $ **FLOATING
C2919 S.t1198 VSUBS 0.02fF
C2920 S.n2635 VSUBS 0.12fF $ **FLOATING
C2921 S.n2636 VSUBS 0.14fF $ **FLOATING
C2922 S.t2479 VSUBS 0.02fF
C2923 S.n2638 VSUBS 0.24fF $ **FLOATING
C2924 S.n2639 VSUBS 0.91fF $ **FLOATING
C2925 S.n2640 VSUBS 0.05fF $ **FLOATING
C2926 S.t187 VSUBS 48.27fF
C2927 S.t173 VSUBS 0.02fF
C2928 S.n2641 VSUBS 0.24fF $ **FLOATING
C2929 S.n2642 VSUBS 0.91fF $ **FLOATING
C2930 S.n2643 VSUBS 0.05fF $ **FLOATING
C2931 S.t407 VSUBS 0.02fF
C2932 S.n2644 VSUBS 0.12fF $ **FLOATING
C2933 S.n2645 VSUBS 0.14fF $ **FLOATING
C2934 S.n2647 VSUBS 0.12fF $ **FLOATING
C2935 S.t2060 VSUBS 0.02fF
C2936 S.n2648 VSUBS 0.14fF $ **FLOATING
C2937 S.n2650 VSUBS 5.17fF $ **FLOATING
C2938 S.n2651 VSUBS 5.45fF $ **FLOATING
C2939 S.t2050 VSUBS 0.02fF
C2940 S.n2652 VSUBS 0.12fF $ **FLOATING
C2941 S.n2653 VSUBS 0.14fF $ **FLOATING
C2942 S.t1814 VSUBS 0.02fF
C2943 S.n2655 VSUBS 0.24fF $ **FLOATING
C2944 S.n2656 VSUBS 0.91fF $ **FLOATING
C2945 S.n2657 VSUBS 0.05fF $ **FLOATING
C2946 S.t259 VSUBS 47.89fF
C2947 S.t2318 VSUBS 0.02fF
C2948 S.n2658 VSUBS 0.01fF $ **FLOATING
C2949 S.n2659 VSUBS 0.26fF $ **FLOATING
C2950 S.t2367 VSUBS 0.02fF
C2951 S.n2661 VSUBS 1.19fF $ **FLOATING
C2952 S.n2662 VSUBS 0.05fF $ **FLOATING
C2953 S.t1805 VSUBS 0.02fF
C2954 S.n2663 VSUBS 0.64fF $ **FLOATING
C2955 S.n2664 VSUBS 0.61fF $ **FLOATING
C2956 S.n2665 VSUBS 8.97fF $ **FLOATING
C2957 S.n2666 VSUBS 8.97fF $ **FLOATING
C2958 S.n2667 VSUBS 0.60fF $ **FLOATING
C2959 S.n2668 VSUBS 0.22fF $ **FLOATING
C2960 S.n2669 VSUBS 0.59fF $ **FLOATING
C2961 S.n2670 VSUBS 3.39fF $ **FLOATING
C2962 S.n2671 VSUBS 0.29fF $ **FLOATING
C2963 S.t21 VSUBS 21.42fF
C2964 S.n2672 VSUBS 21.71fF $ **FLOATING
C2965 S.n2673 VSUBS 0.77fF $ **FLOATING
C2966 S.n2674 VSUBS 0.28fF $ **FLOATING
C2967 S.n2675 VSUBS 4.00fF $ **FLOATING
C2968 S.n2676 VSUBS 1.35fF $ **FLOATING
C2969 S.n2677 VSUBS 0.01fF $ **FLOATING
C2970 S.n2678 VSUBS 0.02fF $ **FLOATING
C2971 S.n2679 VSUBS 0.03fF $ **FLOATING
C2972 S.n2680 VSUBS 0.04fF $ **FLOATING
C2973 S.n2681 VSUBS 0.17fF $ **FLOATING
C2974 S.n2682 VSUBS 0.01fF $ **FLOATING
C2975 S.n2683 VSUBS 0.02fF $ **FLOATING
C2976 S.n2684 VSUBS 0.01fF $ **FLOATING
C2977 S.n2685 VSUBS 0.01fF $ **FLOATING
C2978 S.n2686 VSUBS 0.01fF $ **FLOATING
C2979 S.n2687 VSUBS 0.01fF $ **FLOATING
C2980 S.n2688 VSUBS 0.02fF $ **FLOATING
C2981 S.n2689 VSUBS 0.01fF $ **FLOATING
C2982 S.n2690 VSUBS 0.02fF $ **FLOATING
C2983 S.n2691 VSUBS 0.05fF $ **FLOATING
C2984 S.n2692 VSUBS 0.04fF $ **FLOATING
C2985 S.n2693 VSUBS 0.11fF $ **FLOATING
C2986 S.n2694 VSUBS 0.38fF $ **FLOATING
C2987 S.n2695 VSUBS 0.20fF $ **FLOATING
C2988 S.n2696 VSUBS 4.39fF $ **FLOATING
C2989 S.n2697 VSUBS 0.24fF $ **FLOATING
C2990 S.n2698 VSUBS 1.50fF $ **FLOATING
C2991 S.n2699 VSUBS 1.30fF $ **FLOATING
C2992 S.n2700 VSUBS 0.28fF $ **FLOATING
C2993 S.n2701 VSUBS 0.25fF $ **FLOATING
C2994 S.n2702 VSUBS 0.09fF $ **FLOATING
C2995 S.n2703 VSUBS 0.21fF $ **FLOATING
C2996 S.n2704 VSUBS 0.92fF $ **FLOATING
C2997 S.n2705 VSUBS 0.44fF $ **FLOATING
C2998 S.n2706 VSUBS 1.88fF $ **FLOATING
C2999 S.n2707 VSUBS 0.12fF $ **FLOATING
C3000 S.t1405 VSUBS 0.02fF
C3001 S.n2708 VSUBS 0.14fF $ **FLOATING
C3002 S.t2221 VSUBS 0.02fF
C3003 S.n2710 VSUBS 0.24fF $ **FLOATING
C3004 S.n2711 VSUBS 0.36fF $ **FLOATING
C3005 S.n2712 VSUBS 0.61fF $ **FLOATING
C3006 S.n2713 VSUBS 0.02fF $ **FLOATING
C3007 S.n2714 VSUBS 0.01fF $ **FLOATING
C3008 S.n2715 VSUBS 0.02fF $ **FLOATING
C3009 S.n2716 VSUBS 0.08fF $ **FLOATING
C3010 S.n2717 VSUBS 0.06fF $ **FLOATING
C3011 S.n2718 VSUBS 0.03fF $ **FLOATING
C3012 S.n2719 VSUBS 0.04fF $ **FLOATING
C3013 S.n2720 VSUBS 1.00fF $ **FLOATING
C3014 S.n2721 VSUBS 0.36fF $ **FLOATING
C3015 S.n2722 VSUBS 1.87fF $ **FLOATING
C3016 S.n2723 VSUBS 1.99fF $ **FLOATING
C3017 S.t1425 VSUBS 0.02fF
C3018 S.n2724 VSUBS 0.24fF $ **FLOATING
C3019 S.n2725 VSUBS 0.91fF $ **FLOATING
C3020 S.n2726 VSUBS 0.05fF $ **FLOATING
C3021 S.t2267 VSUBS 0.02fF
C3022 S.n2727 VSUBS 0.12fF $ **FLOATING
C3023 S.n2728 VSUBS 0.14fF $ **FLOATING
C3024 S.n2730 VSUBS 1.89fF $ **FLOATING
C3025 S.n2731 VSUBS 0.06fF $ **FLOATING
C3026 S.n2732 VSUBS 0.03fF $ **FLOATING
C3027 S.n2733 VSUBS 0.04fF $ **FLOATING
C3028 S.n2734 VSUBS 0.99fF $ **FLOATING
C3029 S.n2735 VSUBS 0.02fF $ **FLOATING
C3030 S.n2736 VSUBS 0.01fF $ **FLOATING
C3031 S.n2737 VSUBS 0.02fF $ **FLOATING
C3032 S.n2738 VSUBS 0.08fF $ **FLOATING
C3033 S.n2739 VSUBS 0.36fF $ **FLOATING
C3034 S.n2740 VSUBS 1.85fF $ **FLOATING
C3035 S.t604 VSUBS 0.02fF
C3036 S.n2741 VSUBS 0.24fF $ **FLOATING
C3037 S.n2742 VSUBS 0.36fF $ **FLOATING
C3038 S.n2743 VSUBS 0.61fF $ **FLOATING
C3039 S.n2744 VSUBS 0.12fF $ **FLOATING
C3040 S.t2313 VSUBS 0.02fF
C3041 S.n2745 VSUBS 0.14fF $ **FLOATING
C3042 S.n2747 VSUBS 0.70fF $ **FLOATING
C3043 S.n2748 VSUBS 0.23fF $ **FLOATING
C3044 S.n2749 VSUBS 0.23fF $ **FLOATING
C3045 S.n2750 VSUBS 0.70fF $ **FLOATING
C3046 S.n2751 VSUBS 1.16fF $ **FLOATING
C3047 S.n2752 VSUBS 0.22fF $ **FLOATING
C3048 S.n2753 VSUBS 0.25fF $ **FLOATING
C3049 S.n2754 VSUBS 0.09fF $ **FLOATING
C3050 S.n2755 VSUBS 1.88fF $ **FLOATING
C3051 S.t2333 VSUBS 0.02fF
C3052 S.n2756 VSUBS 0.24fF $ **FLOATING
C3053 S.n2757 VSUBS 0.91fF $ **FLOATING
C3054 S.n2758 VSUBS 0.05fF $ **FLOATING
C3055 S.t655 VSUBS 0.02fF
C3056 S.n2759 VSUBS 0.12fF $ **FLOATING
C3057 S.n2760 VSUBS 0.14fF $ **FLOATING
C3058 S.n2762 VSUBS 0.25fF $ **FLOATING
C3059 S.n2763 VSUBS 0.09fF $ **FLOATING
C3060 S.n2764 VSUBS 0.21fF $ **FLOATING
C3061 S.n2765 VSUBS 0.92fF $ **FLOATING
C3062 S.n2766 VSUBS 0.44fF $ **FLOATING
C3063 S.n2767 VSUBS 1.88fF $ **FLOATING
C3064 S.n2768 VSUBS 0.12fF $ **FLOATING
C3065 S.t1937 VSUBS 0.02fF
C3066 S.n2769 VSUBS 0.14fF $ **FLOATING
C3067 S.t228 VSUBS 0.02fF
C3068 S.n2771 VSUBS 0.24fF $ **FLOATING
C3069 S.n2772 VSUBS 0.36fF $ **FLOATING
C3070 S.n2773 VSUBS 0.61fF $ **FLOATING
C3071 S.n2774 VSUBS 0.02fF $ **FLOATING
C3072 S.n2775 VSUBS 0.01fF $ **FLOATING
C3073 S.n2776 VSUBS 0.02fF $ **FLOATING
C3074 S.n2777 VSUBS 0.08fF $ **FLOATING
C3075 S.n2778 VSUBS 0.06fF $ **FLOATING
C3076 S.n2779 VSUBS 0.03fF $ **FLOATING
C3077 S.n2780 VSUBS 0.04fF $ **FLOATING
C3078 S.n2781 VSUBS 1.00fF $ **FLOATING
C3079 S.n2782 VSUBS 0.36fF $ **FLOATING
C3080 S.n2783 VSUBS 1.87fF $ **FLOATING
C3081 S.n2784 VSUBS 1.99fF $ **FLOATING
C3082 S.t1959 VSUBS 0.02fF
C3083 S.n2785 VSUBS 0.24fF $ **FLOATING
C3084 S.n2786 VSUBS 0.91fF $ **FLOATING
C3085 S.n2787 VSUBS 0.05fF $ **FLOATING
C3086 S.t1447 VSUBS 0.02fF
C3087 S.n2788 VSUBS 0.12fF $ **FLOATING
C3088 S.n2789 VSUBS 0.14fF $ **FLOATING
C3089 S.n2791 VSUBS 1.89fF $ **FLOATING
C3090 S.n2792 VSUBS 0.06fF $ **FLOATING
C3091 S.n2793 VSUBS 0.03fF $ **FLOATING
C3092 S.n2794 VSUBS 0.04fF $ **FLOATING
C3093 S.n2795 VSUBS 0.99fF $ **FLOATING
C3094 S.n2796 VSUBS 0.02fF $ **FLOATING
C3095 S.n2797 VSUBS 0.01fF $ **FLOATING
C3096 S.n2798 VSUBS 0.02fF $ **FLOATING
C3097 S.n2799 VSUBS 0.08fF $ **FLOATING
C3098 S.n2800 VSUBS 0.36fF $ **FLOATING
C3099 S.n2801 VSUBS 1.85fF $ **FLOATING
C3100 S.t1013 VSUBS 0.02fF
C3101 S.n2802 VSUBS 0.24fF $ **FLOATING
C3102 S.n2803 VSUBS 0.36fF $ **FLOATING
C3103 S.n2804 VSUBS 0.61fF $ **FLOATING
C3104 S.n2805 VSUBS 0.12fF $ **FLOATING
C3105 S.t196 VSUBS 0.02fF
C3106 S.n2806 VSUBS 0.14fF $ **FLOATING
C3107 S.n2808 VSUBS 0.70fF $ **FLOATING
C3108 S.n2809 VSUBS 0.23fF $ **FLOATING
C3109 S.n2810 VSUBS 0.23fF $ **FLOATING
C3110 S.n2811 VSUBS 0.70fF $ **FLOATING
C3111 S.n2812 VSUBS 1.16fF $ **FLOATING
C3112 S.n2813 VSUBS 0.22fF $ **FLOATING
C3113 S.n2814 VSUBS 0.25fF $ **FLOATING
C3114 S.n2815 VSUBS 0.09fF $ **FLOATING
C3115 S.n2816 VSUBS 1.88fF $ **FLOATING
C3116 S.t217 VSUBS 0.02fF
C3117 S.n2817 VSUBS 0.24fF $ **FLOATING
C3118 S.n2818 VSUBS 0.91fF $ **FLOATING
C3119 S.n2819 VSUBS 0.05fF $ **FLOATING
C3120 S.t1068 VSUBS 0.02fF
C3121 S.n2820 VSUBS 0.12fF $ **FLOATING
C3122 S.n2821 VSUBS 0.14fF $ **FLOATING
C3123 S.n2823 VSUBS 0.25fF $ **FLOATING
C3124 S.n2824 VSUBS 0.09fF $ **FLOATING
C3125 S.n2825 VSUBS 0.21fF $ **FLOATING
C3126 S.n2826 VSUBS 0.92fF $ **FLOATING
C3127 S.n2827 VSUBS 0.44fF $ **FLOATING
C3128 S.n2828 VSUBS 1.88fF $ **FLOATING
C3129 S.n2829 VSUBS 0.12fF $ **FLOATING
C3130 S.t983 VSUBS 0.02fF
C3131 S.n2830 VSUBS 0.14fF $ **FLOATING
C3132 S.t1791 VSUBS 0.02fF
C3133 S.n2832 VSUBS 0.24fF $ **FLOATING
C3134 S.n2833 VSUBS 0.36fF $ **FLOATING
C3135 S.n2834 VSUBS 0.61fF $ **FLOATING
C3136 S.n2835 VSUBS 0.02fF $ **FLOATING
C3137 S.n2836 VSUBS 0.01fF $ **FLOATING
C3138 S.n2837 VSUBS 0.02fF $ **FLOATING
C3139 S.n2838 VSUBS 0.08fF $ **FLOATING
C3140 S.n2839 VSUBS 0.06fF $ **FLOATING
C3141 S.n2840 VSUBS 0.03fF $ **FLOATING
C3142 S.n2841 VSUBS 0.04fF $ **FLOATING
C3143 S.n2842 VSUBS 1.00fF $ **FLOATING
C3144 S.n2843 VSUBS 0.36fF $ **FLOATING
C3145 S.n2844 VSUBS 1.87fF $ **FLOATING
C3146 S.n2845 VSUBS 1.99fF $ **FLOATING
C3147 S.t1006 VSUBS 0.02fF
C3148 S.n2846 VSUBS 0.24fF $ **FLOATING
C3149 S.n2847 VSUBS 0.91fF $ **FLOATING
C3150 S.n2848 VSUBS 0.05fF $ **FLOATING
C3151 S.t1854 VSUBS 0.02fF
C3152 S.n2849 VSUBS 0.12fF $ **FLOATING
C3153 S.n2850 VSUBS 0.14fF $ **FLOATING
C3154 S.n2852 VSUBS 1.89fF $ **FLOATING
C3155 S.n2853 VSUBS 0.06fF $ **FLOATING
C3156 S.n2854 VSUBS 0.03fF $ **FLOATING
C3157 S.n2855 VSUBS 0.04fF $ **FLOATING
C3158 S.n2856 VSUBS 0.99fF $ **FLOATING
C3159 S.n2857 VSUBS 0.02fF $ **FLOATING
C3160 S.n2858 VSUBS 0.01fF $ **FLOATING
C3161 S.n2859 VSUBS 0.02fF $ **FLOATING
C3162 S.n2860 VSUBS 0.08fF $ **FLOATING
C3163 S.n2861 VSUBS 0.36fF $ **FLOATING
C3164 S.n2862 VSUBS 1.85fF $ **FLOATING
C3165 S.t2574 VSUBS 0.02fF
C3166 S.n2863 VSUBS 0.24fF $ **FLOATING
C3167 S.n2864 VSUBS 0.36fF $ **FLOATING
C3168 S.n2865 VSUBS 0.61fF $ **FLOATING
C3169 S.n2866 VSUBS 0.12fF $ **FLOATING
C3170 S.t1764 VSUBS 0.02fF
C3171 S.n2867 VSUBS 0.14fF $ **FLOATING
C3172 S.n2869 VSUBS 0.70fF $ **FLOATING
C3173 S.n2870 VSUBS 0.23fF $ **FLOATING
C3174 S.n2871 VSUBS 0.23fF $ **FLOATING
C3175 S.n2872 VSUBS 0.70fF $ **FLOATING
C3176 S.n2873 VSUBS 1.16fF $ **FLOATING
C3177 S.n2874 VSUBS 0.22fF $ **FLOATING
C3178 S.n2875 VSUBS 0.25fF $ **FLOATING
C3179 S.n2876 VSUBS 0.09fF $ **FLOATING
C3180 S.n2877 VSUBS 1.88fF $ **FLOATING
C3181 S.t1787 VSUBS 0.02fF
C3182 S.n2878 VSUBS 0.24fF $ **FLOATING
C3183 S.n2879 VSUBS 0.91fF $ **FLOATING
C3184 S.n2880 VSUBS 0.05fF $ **FLOATING
C3185 S.t85 VSUBS 0.02fF
C3186 S.n2881 VSUBS 0.12fF $ **FLOATING
C3187 S.n2882 VSUBS 0.14fF $ **FLOATING
C3188 S.n2884 VSUBS 0.25fF $ **FLOATING
C3189 S.n2885 VSUBS 0.09fF $ **FLOATING
C3190 S.n2886 VSUBS 0.21fF $ **FLOATING
C3191 S.n2887 VSUBS 0.92fF $ **FLOATING
C3192 S.n2888 VSUBS 0.44fF $ **FLOATING
C3193 S.n2889 VSUBS 1.88fF $ **FLOATING
C3194 S.n2890 VSUBS 0.12fF $ **FLOATING
C3195 S.t147 VSUBS 0.02fF
C3196 S.n2891 VSUBS 0.14fF $ **FLOATING
C3197 S.t972 VSUBS 0.02fF
C3198 S.n2893 VSUBS 0.24fF $ **FLOATING
C3199 S.n2894 VSUBS 0.36fF $ **FLOATING
C3200 S.n2895 VSUBS 0.61fF $ **FLOATING
C3201 S.n2896 VSUBS 0.02fF $ **FLOATING
C3202 S.n2897 VSUBS 0.01fF $ **FLOATING
C3203 S.n2898 VSUBS 0.02fF $ **FLOATING
C3204 S.n2899 VSUBS 0.08fF $ **FLOATING
C3205 S.n2900 VSUBS 0.06fF $ **FLOATING
C3206 S.n2901 VSUBS 0.03fF $ **FLOATING
C3207 S.n2902 VSUBS 0.04fF $ **FLOATING
C3208 S.n2903 VSUBS 1.00fF $ **FLOATING
C3209 S.n2904 VSUBS 0.36fF $ **FLOATING
C3210 S.n2905 VSUBS 1.87fF $ **FLOATING
C3211 S.n2906 VSUBS 1.99fF $ **FLOATING
C3212 S.t178 VSUBS 0.02fF
C3213 S.n2907 VSUBS 0.24fF $ **FLOATING
C3214 S.n2908 VSUBS 0.91fF $ **FLOATING
C3215 S.n2909 VSUBS 0.05fF $ **FLOATING
C3216 S.t1028 VSUBS 0.02fF
C3217 S.n2910 VSUBS 0.12fF $ **FLOATING
C3218 S.n2911 VSUBS 0.14fF $ **FLOATING
C3219 S.n2913 VSUBS 1.89fF $ **FLOATING
C3220 S.n2914 VSUBS 0.06fF $ **FLOATING
C3221 S.n2915 VSUBS 0.03fF $ **FLOATING
C3222 S.n2916 VSUBS 0.04fF $ **FLOATING
C3223 S.n2917 VSUBS 0.99fF $ **FLOATING
C3224 S.n2918 VSUBS 0.02fF $ **FLOATING
C3225 S.n2919 VSUBS 0.01fF $ **FLOATING
C3226 S.n2920 VSUBS 0.02fF $ **FLOATING
C3227 S.n2921 VSUBS 0.08fF $ **FLOATING
C3228 S.n2922 VSUBS 0.36fF $ **FLOATING
C3229 S.n2923 VSUBS 1.85fF $ **FLOATING
C3230 S.t580 VSUBS 0.02fF
C3231 S.n2924 VSUBS 0.24fF $ **FLOATING
C3232 S.n2925 VSUBS 0.36fF $ **FLOATING
C3233 S.n2926 VSUBS 0.61fF $ **FLOATING
C3234 S.n2927 VSUBS 0.12fF $ **FLOATING
C3235 S.t2283 VSUBS 0.02fF
C3236 S.n2928 VSUBS 0.14fF $ **FLOATING
C3237 S.n2930 VSUBS 0.70fF $ **FLOATING
C3238 S.n2931 VSUBS 0.23fF $ **FLOATING
C3239 S.n2932 VSUBS 0.23fF $ **FLOATING
C3240 S.n2933 VSUBS 0.70fF $ **FLOATING
C3241 S.n2934 VSUBS 1.16fF $ **FLOATING
C3242 S.n2935 VSUBS 0.22fF $ **FLOATING
C3243 S.n2936 VSUBS 0.25fF $ **FLOATING
C3244 S.n2937 VSUBS 0.09fF $ **FLOATING
C3245 S.n2938 VSUBS 1.88fF $ **FLOATING
C3246 S.t2304 VSUBS 0.02fF
C3247 S.n2939 VSUBS 0.24fF $ **FLOATING
C3248 S.n2940 VSUBS 0.91fF $ **FLOATING
C3249 S.n2941 VSUBS 0.05fF $ **FLOATING
C3250 S.t629 VSUBS 0.02fF
C3251 S.n2942 VSUBS 0.12fF $ **FLOATING
C3252 S.n2943 VSUBS 0.14fF $ **FLOATING
C3253 S.n2945 VSUBS 0.25fF $ **FLOATING
C3254 S.n2946 VSUBS 0.09fF $ **FLOATING
C3255 S.n2947 VSUBS 0.21fF $ **FLOATING
C3256 S.n2948 VSUBS 0.92fF $ **FLOATING
C3257 S.n2949 VSUBS 0.44fF $ **FLOATING
C3258 S.n2950 VSUBS 1.88fF $ **FLOATING
C3259 S.n2951 VSUBS 0.12fF $ **FLOATING
C3260 S.t555 VSUBS 0.02fF
C3261 S.n2952 VSUBS 0.14fF $ **FLOATING
C3262 S.t1370 VSUBS 0.02fF
C3263 S.n2954 VSUBS 0.24fF $ **FLOATING
C3264 S.n2955 VSUBS 0.36fF $ **FLOATING
C3265 S.n2956 VSUBS 0.61fF $ **FLOATING
C3266 S.n2957 VSUBS 0.02fF $ **FLOATING
C3267 S.n2958 VSUBS 0.01fF $ **FLOATING
C3268 S.n2959 VSUBS 0.02fF $ **FLOATING
C3269 S.n2960 VSUBS 0.08fF $ **FLOATING
C3270 S.n2961 VSUBS 0.06fF $ **FLOATING
C3271 S.n2962 VSUBS 0.03fF $ **FLOATING
C3272 S.n2963 VSUBS 0.04fF $ **FLOATING
C3273 S.n2964 VSUBS 1.00fF $ **FLOATING
C3274 S.n2965 VSUBS 0.36fF $ **FLOATING
C3275 S.n2966 VSUBS 1.87fF $ **FLOATING
C3276 S.n2967 VSUBS 1.99fF $ **FLOATING
C3277 S.t574 VSUBS 0.02fF
C3278 S.n2968 VSUBS 0.24fF $ **FLOATING
C3279 S.n2969 VSUBS 0.91fF $ **FLOATING
C3280 S.n2970 VSUBS 0.05fF $ **FLOATING
C3281 S.t1419 VSUBS 0.02fF
C3282 S.n2971 VSUBS 0.12fF $ **FLOATING
C3283 S.n2972 VSUBS 0.14fF $ **FLOATING
C3284 S.n2974 VSUBS 1.89fF $ **FLOATING
C3285 S.n2975 VSUBS 0.04fF $ **FLOATING
C3286 S.n2976 VSUBS 0.07fF $ **FLOATING
C3287 S.n2977 VSUBS 0.05fF $ **FLOATING
C3288 S.n2978 VSUBS 0.87fF $ **FLOATING
C3289 S.n2979 VSUBS 0.01fF $ **FLOATING
C3290 S.n2980 VSUBS 0.01fF $ **FLOATING
C3291 S.n2981 VSUBS 0.01fF $ **FLOATING
C3292 S.n2982 VSUBS 0.07fF $ **FLOATING
C3293 S.n2983 VSUBS 0.68fF $ **FLOATING
C3294 S.n2984 VSUBS 0.72fF $ **FLOATING
C3295 S.t2155 VSUBS 0.02fF
C3296 S.n2985 VSUBS 0.24fF $ **FLOATING
C3297 S.n2986 VSUBS 0.36fF $ **FLOATING
C3298 S.n2987 VSUBS 0.61fF $ **FLOATING
C3299 S.n2988 VSUBS 0.12fF $ **FLOATING
C3300 S.t1343 VSUBS 0.02fF
C3301 S.n2989 VSUBS 0.14fF $ **FLOATING
C3302 S.n2991 VSUBS 0.70fF $ **FLOATING
C3303 S.n2992 VSUBS 0.23fF $ **FLOATING
C3304 S.n2993 VSUBS 0.23fF $ **FLOATING
C3305 S.n2994 VSUBS 0.70fF $ **FLOATING
C3306 S.n2995 VSUBS 1.16fF $ **FLOATING
C3307 S.n2996 VSUBS 0.22fF $ **FLOATING
C3308 S.n2997 VSUBS 0.25fF $ **FLOATING
C3309 S.n2998 VSUBS 0.09fF $ **FLOATING
C3310 S.n2999 VSUBS 2.31fF $ **FLOATING
C3311 S.t1363 VSUBS 0.02fF
C3312 S.n3000 VSUBS 0.24fF $ **FLOATING
C3313 S.n3001 VSUBS 0.91fF $ **FLOATING
C3314 S.n3002 VSUBS 0.05fF $ **FLOATING
C3315 S.t2208 VSUBS 0.02fF
C3316 S.n3003 VSUBS 0.12fF $ **FLOATING
C3317 S.n3004 VSUBS 0.14fF $ **FLOATING
C3318 S.n3006 VSUBS 1.88fF $ **FLOATING
C3319 S.n3007 VSUBS 0.46fF $ **FLOATING
C3320 S.n3008 VSUBS 0.22fF $ **FLOATING
C3321 S.n3009 VSUBS 0.38fF $ **FLOATING
C3322 S.n3010 VSUBS 0.16fF $ **FLOATING
C3323 S.n3011 VSUBS 0.28fF $ **FLOATING
C3324 S.n3012 VSUBS 0.21fF $ **FLOATING
C3325 S.n3013 VSUBS 0.30fF $ **FLOATING
C3326 S.n3014 VSUBS 0.42fF $ **FLOATING
C3327 S.n3015 VSUBS 0.21fF $ **FLOATING
C3328 S.t424 VSUBS 0.02fF
C3329 S.n3016 VSUBS 0.24fF $ **FLOATING
C3330 S.n3017 VSUBS 0.36fF $ **FLOATING
C3331 S.n3018 VSUBS 0.61fF $ **FLOATING
C3332 S.n3019 VSUBS 0.12fF $ **FLOATING
C3333 S.t2130 VSUBS 0.02fF
C3334 S.n3020 VSUBS 0.14fF $ **FLOATING
C3335 S.n3022 VSUBS 0.04fF $ **FLOATING
C3336 S.n3023 VSUBS 0.03fF $ **FLOATING
C3337 S.n3024 VSUBS 0.03fF $ **FLOATING
C3338 S.n3025 VSUBS 0.10fF $ **FLOATING
C3339 S.n3026 VSUBS 0.36fF $ **FLOATING
C3340 S.n3027 VSUBS 0.38fF $ **FLOATING
C3341 S.n3028 VSUBS 0.11fF $ **FLOATING
C3342 S.n3029 VSUBS 0.12fF $ **FLOATING
C3343 S.n3030 VSUBS 0.07fF $ **FLOATING
C3344 S.n3031 VSUBS 0.12fF $ **FLOATING
C3345 S.n3032 VSUBS 0.18fF $ **FLOATING
C3346 S.n3033 VSUBS 3.99fF $ **FLOATING
C3347 S.t2150 VSUBS 0.02fF
C3348 S.n3034 VSUBS 0.24fF $ **FLOATING
C3349 S.n3035 VSUBS 0.91fF $ **FLOATING
C3350 S.n3036 VSUBS 0.05fF $ **FLOATING
C3351 S.t475 VSUBS 0.02fF
C3352 S.n3037 VSUBS 0.12fF $ **FLOATING
C3353 S.n3038 VSUBS 0.14fF $ **FLOATING
C3354 S.n3040 VSUBS 0.25fF $ **FLOATING
C3355 S.n3041 VSUBS 0.09fF $ **FLOATING
C3356 S.n3042 VSUBS 0.21fF $ **FLOATING
C3357 S.n3043 VSUBS 1.28fF $ **FLOATING
C3358 S.n3044 VSUBS 0.53fF $ **FLOATING
C3359 S.n3045 VSUBS 1.88fF $ **FLOATING
C3360 S.n3046 VSUBS 0.12fF $ **FLOATING
C3361 S.t1968 VSUBS 0.02fF
C3362 S.n3047 VSUBS 0.14fF $ **FLOATING
C3363 S.t1757 VSUBS 0.02fF
C3364 S.n3049 VSUBS 0.24fF $ **FLOATING
C3365 S.n3050 VSUBS 0.36fF $ **FLOATING
C3366 S.n3051 VSUBS 0.61fF $ **FLOATING
C3367 S.n3052 VSUBS 1.58fF $ **FLOATING
C3368 S.n3053 VSUBS 2.45fF $ **FLOATING
C3369 S.t371 VSUBS 0.02fF
C3370 S.n3054 VSUBS 0.24fF $ **FLOATING
C3371 S.n3055 VSUBS 0.91fF $ **FLOATING
C3372 S.n3056 VSUBS 0.05fF $ **FLOATING
C3373 S.t1382 VSUBS 0.02fF
C3374 S.n3057 VSUBS 0.12fF $ **FLOATING
C3375 S.n3058 VSUBS 0.14fF $ **FLOATING
C3376 S.n3060 VSUBS 1.89fF $ **FLOATING
C3377 S.n3061 VSUBS 0.06fF $ **FLOATING
C3378 S.n3062 VSUBS 0.03fF $ **FLOATING
C3379 S.n3063 VSUBS 0.04fF $ **FLOATING
C3380 S.n3064 VSUBS 0.99fF $ **FLOATING
C3381 S.n3065 VSUBS 0.02fF $ **FLOATING
C3382 S.n3066 VSUBS 0.01fF $ **FLOATING
C3383 S.n3067 VSUBS 0.02fF $ **FLOATING
C3384 S.n3068 VSUBS 0.08fF $ **FLOATING
C3385 S.n3069 VSUBS 0.36fF $ **FLOATING
C3386 S.n3070 VSUBS 1.85fF $ **FLOATING
C3387 S.t2538 VSUBS 0.02fF
C3388 S.n3071 VSUBS 0.24fF $ **FLOATING
C3389 S.n3072 VSUBS 0.36fF $ **FLOATING
C3390 S.n3073 VSUBS 0.61fF $ **FLOATING
C3391 S.n3074 VSUBS 0.12fF $ **FLOATING
C3392 S.t229 VSUBS 0.02fF
C3393 S.n3075 VSUBS 0.14fF $ **FLOATING
C3394 S.n3077 VSUBS 0.70fF $ **FLOATING
C3395 S.n3078 VSUBS 0.23fF $ **FLOATING
C3396 S.n3079 VSUBS 0.23fF $ **FLOATING
C3397 S.n3080 VSUBS 0.70fF $ **FLOATING
C3398 S.n3081 VSUBS 1.16fF $ **FLOATING
C3399 S.n3082 VSUBS 0.22fF $ **FLOATING
C3400 S.n3083 VSUBS 0.25fF $ **FLOATING
C3401 S.n3084 VSUBS 0.09fF $ **FLOATING
C3402 S.n3085 VSUBS 1.88fF $ **FLOATING
C3403 S.t1159 VSUBS 0.02fF
C3404 S.n3086 VSUBS 0.24fF $ **FLOATING
C3405 S.n3087 VSUBS 0.91fF $ **FLOATING
C3406 S.n3088 VSUBS 0.05fF $ **FLOATING
C3407 S.t1104 VSUBS 0.02fF
C3408 S.n3089 VSUBS 0.12fF $ **FLOATING
C3409 S.n3090 VSUBS 0.14fF $ **FLOATING
C3410 S.n3092 VSUBS 20.78fF $ **FLOATING
C3411 S.n3093 VSUBS 1.72fF $ **FLOATING
C3412 S.n3094 VSUBS 3.05fF $ **FLOATING
C3413 S.t1429 VSUBS 0.02fF
C3414 S.n3095 VSUBS 0.24fF $ **FLOATING
C3415 S.n3096 VSUBS 0.36fF $ **FLOATING
C3416 S.n3097 VSUBS 0.61fF $ **FLOATING
C3417 S.n3098 VSUBS 0.12fF $ **FLOATING
C3418 S.t614 VSUBS 0.02fF
C3419 S.n3099 VSUBS 0.14fF $ **FLOATING
C3420 S.n3101 VSUBS 0.31fF $ **FLOATING
C3421 S.n3102 VSUBS 0.23fF $ **FLOATING
C3422 S.n3103 VSUBS 0.66fF $ **FLOATING
C3423 S.n3104 VSUBS 0.95fF $ **FLOATING
C3424 S.n3105 VSUBS 0.23fF $ **FLOATING
C3425 S.n3106 VSUBS 0.21fF $ **FLOATING
C3426 S.n3107 VSUBS 0.20fF $ **FLOATING
C3427 S.n3108 VSUBS 0.06fF $ **FLOATING
C3428 S.n3109 VSUBS 0.09fF $ **FLOATING
C3429 S.n3110 VSUBS 0.10fF $ **FLOATING
C3430 S.n3111 VSUBS 1.99fF $ **FLOATING
C3431 S.t1483 VSUBS 0.02fF
C3432 S.n3112 VSUBS 0.12fF $ **FLOATING
C3433 S.n3113 VSUBS 0.14fF $ **FLOATING
C3434 S.t638 VSUBS 0.02fF
C3435 S.n3115 VSUBS 0.24fF $ **FLOATING
C3436 S.n3116 VSUBS 0.91fF $ **FLOATING
C3437 S.n3117 VSUBS 0.05fF $ **FLOATING
C3438 S.n3118 VSUBS 1.88fF $ **FLOATING
C3439 S.n3119 VSUBS 0.12fF $ **FLOATING
C3440 S.t1043 VSUBS 0.02fF
C3441 S.n3120 VSUBS 0.14fF $ **FLOATING
C3442 S.t2018 VSUBS 0.02fF
C3443 S.n3122 VSUBS 1.22fF $ **FLOATING
C3444 S.n3123 VSUBS 0.61fF $ **FLOATING
C3445 S.n3124 VSUBS 0.35fF $ **FLOATING
C3446 S.n3125 VSUBS 0.63fF $ **FLOATING
C3447 S.n3126 VSUBS 1.15fF $ **FLOATING
C3448 S.n3127 VSUBS 3.00fF $ **FLOATING
C3449 S.n3128 VSUBS 0.59fF $ **FLOATING
C3450 S.n3129 VSUBS 0.01fF $ **FLOATING
C3451 S.n3130 VSUBS 0.97fF $ **FLOATING
C3452 S.t111 VSUBS 21.42fF
C3453 S.n3131 VSUBS 20.29fF $ **FLOATING
C3454 S.n3133 VSUBS 0.38fF $ **FLOATING
C3455 S.n3134 VSUBS 0.23fF $ **FLOATING
C3456 S.n3135 VSUBS 2.90fF $ **FLOATING
C3457 S.n3136 VSUBS 2.46fF $ **FLOATING
C3458 S.n3137 VSUBS 1.96fF $ **FLOATING
C3459 S.n3138 VSUBS 3.94fF $ **FLOATING
C3460 S.n3139 VSUBS 0.25fF $ **FLOATING
C3461 S.n3140 VSUBS 0.01fF $ **FLOATING
C3462 S.t1214 VSUBS 0.02fF
C3463 S.n3141 VSUBS 0.26fF $ **FLOATING
C3464 S.t2296 VSUBS 0.02fF
C3465 S.n3142 VSUBS 0.95fF $ **FLOATING
C3466 S.n3143 VSUBS 0.71fF $ **FLOATING
C3467 S.n3144 VSUBS 0.78fF $ **FLOATING
C3468 S.n3145 VSUBS 1.93fF $ **FLOATING
C3469 S.n3146 VSUBS 1.88fF $ **FLOATING
C3470 S.n3147 VSUBS 0.12fF $ **FLOATING
C3471 S.t1992 VSUBS 0.02fF
C3472 S.n3148 VSUBS 0.14fF $ **FLOATING
C3473 S.t290 VSUBS 0.02fF
C3474 S.n3150 VSUBS 0.24fF $ **FLOATING
C3475 S.n3151 VSUBS 0.36fF $ **FLOATING
C3476 S.n3152 VSUBS 0.61fF $ **FLOATING
C3477 S.n3153 VSUBS 1.52fF $ **FLOATING
C3478 S.n3154 VSUBS 2.99fF $ **FLOATING
C3479 S.t565 VSUBS 0.02fF
C3480 S.n3155 VSUBS 0.24fF $ **FLOATING
C3481 S.n3156 VSUBS 0.91fF $ **FLOATING
C3482 S.n3157 VSUBS 0.05fF $ **FLOATING
C3483 S.t344 VSUBS 0.02fF
C3484 S.n3158 VSUBS 0.12fF $ **FLOATING
C3485 S.n3159 VSUBS 0.14fF $ **FLOATING
C3486 S.n3161 VSUBS 1.89fF $ **FLOATING
C3487 S.n3162 VSUBS 1.88fF $ **FLOATING
C3488 S.t1075 VSUBS 0.02fF
C3489 S.n3163 VSUBS 0.24fF $ **FLOATING
C3490 S.n3164 VSUBS 0.36fF $ **FLOATING
C3491 S.n3165 VSUBS 0.61fF $ **FLOATING
C3492 S.n3166 VSUBS 0.12fF $ **FLOATING
C3493 S.t384 VSUBS 0.02fF
C3494 S.n3167 VSUBS 0.14fF $ **FLOATING
C3495 S.n3169 VSUBS 1.16fF $ **FLOATING
C3496 S.n3170 VSUBS 0.22fF $ **FLOATING
C3497 S.n3171 VSUBS 0.25fF $ **FLOATING
C3498 S.n3172 VSUBS 0.09fF $ **FLOATING
C3499 S.n3173 VSUBS 1.88fF $ **FLOATING
C3500 S.t1355 VSUBS 0.02fF
C3501 S.n3174 VSUBS 0.24fF $ **FLOATING
C3502 S.n3175 VSUBS 0.91fF $ **FLOATING
C3503 S.n3176 VSUBS 0.05fF $ **FLOATING
C3504 S.t1133 VSUBS 0.02fF
C3505 S.n3177 VSUBS 0.12fF $ **FLOATING
C3506 S.n3178 VSUBS 0.14fF $ **FLOATING
C3507 S.n3180 VSUBS 0.78fF $ **FLOATING
C3508 S.n3181 VSUBS 1.94fF $ **FLOATING
C3509 S.n3182 VSUBS 1.88fF $ **FLOATING
C3510 S.n3183 VSUBS 0.12fF $ **FLOATING
C3511 S.t1175 VSUBS 0.02fF
C3512 S.n3184 VSUBS 0.14fF $ **FLOATING
C3513 S.t1984 VSUBS 0.02fF
C3514 S.n3186 VSUBS 0.24fF $ **FLOATING
C3515 S.n3187 VSUBS 0.36fF $ **FLOATING
C3516 S.n3188 VSUBS 0.61fF $ **FLOATING
C3517 S.n3189 VSUBS 1.84fF $ **FLOATING
C3518 S.n3190 VSUBS 2.99fF $ **FLOATING
C3519 S.t2261 VSUBS 0.02fF
C3520 S.n3191 VSUBS 0.24fF $ **FLOATING
C3521 S.n3192 VSUBS 0.91fF $ **FLOATING
C3522 S.n3193 VSUBS 0.05fF $ **FLOATING
C3523 S.t2034 VSUBS 0.02fF
C3524 S.n3194 VSUBS 0.12fF $ **FLOATING
C3525 S.n3195 VSUBS 0.14fF $ **FLOATING
C3526 S.n3197 VSUBS 1.89fF $ **FLOATING
C3527 S.n3198 VSUBS 1.88fF $ **FLOATING
C3528 S.t1577 VSUBS 0.02fF
C3529 S.n3199 VSUBS 0.24fF $ **FLOATING
C3530 S.n3200 VSUBS 0.36fF $ **FLOATING
C3531 S.n3201 VSUBS 0.61fF $ **FLOATING
C3532 S.n3202 VSUBS 0.12fF $ **FLOATING
C3533 S.t765 VSUBS 0.02fF
C3534 S.n3203 VSUBS 0.14fF $ **FLOATING
C3535 S.n3205 VSUBS 1.16fF $ **FLOATING
C3536 S.n3206 VSUBS 0.22fF $ **FLOATING
C3537 S.n3207 VSUBS 0.25fF $ **FLOATING
C3538 S.n3208 VSUBS 0.09fF $ **FLOATING
C3539 S.n3209 VSUBS 1.88fF $ **FLOATING
C3540 S.t1881 VSUBS 0.02fF
C3541 S.n3210 VSUBS 0.24fF $ **FLOATING
C3542 S.n3211 VSUBS 0.91fF $ **FLOATING
C3543 S.n3212 VSUBS 0.05fF $ **FLOATING
C3544 S.t1636 VSUBS 0.02fF
C3545 S.n3213 VSUBS 0.12fF $ **FLOATING
C3546 S.n3214 VSUBS 0.14fF $ **FLOATING
C3547 S.n3216 VSUBS 0.78fF $ **FLOATING
C3548 S.n3217 VSUBS 1.94fF $ **FLOATING
C3549 S.n3218 VSUBS 1.88fF $ **FLOATING
C3550 S.n3219 VSUBS 0.12fF $ **FLOATING
C3551 S.t1554 VSUBS 0.02fF
C3552 S.n3220 VSUBS 0.14fF $ **FLOATING
C3553 S.t2366 VSUBS 0.02fF
C3554 S.n3222 VSUBS 0.24fF $ **FLOATING
C3555 S.n3223 VSUBS 0.36fF $ **FLOATING
C3556 S.n3224 VSUBS 0.61fF $ **FLOATING
C3557 S.n3225 VSUBS 1.84fF $ **FLOATING
C3558 S.n3226 VSUBS 2.99fF $ **FLOATING
C3559 S.t129 VSUBS 0.02fF
C3560 S.n3227 VSUBS 0.24fF $ **FLOATING
C3561 S.n3228 VSUBS 0.91fF $ **FLOATING
C3562 S.n3229 VSUBS 0.05fF $ **FLOATING
C3563 S.t2420 VSUBS 0.02fF
C3564 S.n3230 VSUBS 0.12fF $ **FLOATING
C3565 S.n3231 VSUBS 0.14fF $ **FLOATING
C3566 S.n3233 VSUBS 1.89fF $ **FLOATING
C3567 S.n3234 VSUBS 1.88fF $ **FLOATING
C3568 S.t635 VSUBS 0.02fF
C3569 S.n3235 VSUBS 0.24fF $ **FLOATING
C3570 S.n3236 VSUBS 0.36fF $ **FLOATING
C3571 S.n3237 VSUBS 0.61fF $ **FLOATING
C3572 S.n3238 VSUBS 0.12fF $ **FLOATING
C3573 S.t2342 VSUBS 0.02fF
C3574 S.n3239 VSUBS 0.14fF $ **FLOATING
C3575 S.n3241 VSUBS 1.16fF $ **FLOATING
C3576 S.n3242 VSUBS 0.22fF $ **FLOATING
C3577 S.n3243 VSUBS 0.25fF $ **FLOATING
C3578 S.n3244 VSUBS 0.09fF $ **FLOATING
C3579 S.n3245 VSUBS 1.88fF $ **FLOATING
C3580 S.t927 VSUBS 0.02fF
C3581 S.n3246 VSUBS 0.24fF $ **FLOATING
C3582 S.n3247 VSUBS 0.91fF $ **FLOATING
C3583 S.n3248 VSUBS 0.05fF $ **FLOATING
C3584 S.t685 VSUBS 0.02fF
C3585 S.n3249 VSUBS 0.12fF $ **FLOATING
C3586 S.n3250 VSUBS 0.14fF $ **FLOATING
C3587 S.n3252 VSUBS 0.78fF $ **FLOATING
C3588 S.n3253 VSUBS 1.94fF $ **FLOATING
C3589 S.n3254 VSUBS 1.88fF $ **FLOATING
C3590 S.n3255 VSUBS 0.12fF $ **FLOATING
C3591 S.t723 VSUBS 0.02fF
C3592 S.n3256 VSUBS 0.14fF $ **FLOATING
C3593 S.t1422 VSUBS 0.02fF
C3594 S.n3258 VSUBS 0.24fF $ **FLOATING
C3595 S.n3259 VSUBS 0.36fF $ **FLOATING
C3596 S.n3260 VSUBS 0.61fF $ **FLOATING
C3597 S.n3261 VSUBS 1.84fF $ **FLOATING
C3598 S.n3262 VSUBS 2.99fF $ **FLOATING
C3599 S.t1704 VSUBS 0.02fF
C3600 S.n3263 VSUBS 0.24fF $ **FLOATING
C3601 S.n3264 VSUBS 0.91fF $ **FLOATING
C3602 S.n3265 VSUBS 0.05fF $ **FLOATING
C3603 S.t1473 VSUBS 0.02fF
C3604 S.n3266 VSUBS 0.12fF $ **FLOATING
C3605 S.n3267 VSUBS 0.14fF $ **FLOATING
C3606 S.n3269 VSUBS 1.89fF $ **FLOATING
C3607 S.n3270 VSUBS 1.88fF $ **FLOATING
C3608 S.t1172 VSUBS 0.02fF
C3609 S.n3271 VSUBS 0.24fF $ **FLOATING
C3610 S.n3272 VSUBS 0.36fF $ **FLOATING
C3611 S.n3273 VSUBS 0.61fF $ **FLOATING
C3612 S.n3274 VSUBS 0.12fF $ **FLOATING
C3613 S.t360 VSUBS 0.02fF
C3614 S.n3275 VSUBS 0.14fF $ **FLOATING
C3615 S.n3277 VSUBS 1.16fF $ **FLOATING
C3616 S.n3278 VSUBS 0.22fF $ **FLOATING
C3617 S.n3279 VSUBS 0.25fF $ **FLOATING
C3618 S.n3280 VSUBS 0.09fF $ **FLOATING
C3619 S.n3281 VSUBS 1.88fF $ **FLOATING
C3620 S.t1446 VSUBS 0.02fF
C3621 S.n3282 VSUBS 0.24fF $ **FLOATING
C3622 S.n3283 VSUBS 0.91fF $ **FLOATING
C3623 S.n3284 VSUBS 0.05fF $ **FLOATING
C3624 S.t2384 VSUBS 0.02fF
C3625 S.n3285 VSUBS 0.12fF $ **FLOATING
C3626 S.n3286 VSUBS 0.14fF $ **FLOATING
C3627 S.n3288 VSUBS 0.78fF $ **FLOATING
C3628 S.n3289 VSUBS 1.94fF $ **FLOATING
C3629 S.n3290 VSUBS 1.88fF $ **FLOATING
C3630 S.n3291 VSUBS 0.12fF $ **FLOATING
C3631 S.t1146 VSUBS 0.02fF
C3632 S.n3292 VSUBS 0.14fF $ **FLOATING
C3633 S.t1957 VSUBS 0.02fF
C3634 S.n3294 VSUBS 0.24fF $ **FLOATING
C3635 S.n3295 VSUBS 0.36fF $ **FLOATING
C3636 S.n3296 VSUBS 0.61fF $ **FLOATING
C3637 S.n3297 VSUBS 1.84fF $ **FLOATING
C3638 S.n3298 VSUBS 2.99fF $ **FLOATING
C3639 S.t2236 VSUBS 0.02fF
C3640 S.n3299 VSUBS 0.24fF $ **FLOATING
C3641 S.n3300 VSUBS 0.91fF $ **FLOATING
C3642 S.n3301 VSUBS 0.05fF $ **FLOATING
C3643 S.t2006 VSUBS 0.02fF
C3644 S.n3302 VSUBS 0.12fF $ **FLOATING
C3645 S.n3303 VSUBS 0.14fF $ **FLOATING
C3646 S.n3305 VSUBS 1.89fF $ **FLOATING
C3647 S.n3306 VSUBS 1.75fF $ **FLOATING
C3648 S.t214 VSUBS 0.02fF
C3649 S.n3307 VSUBS 0.24fF $ **FLOATING
C3650 S.n3308 VSUBS 0.36fF $ **FLOATING
C3651 S.n3309 VSUBS 0.61fF $ **FLOATING
C3652 S.n3310 VSUBS 0.12fF $ **FLOATING
C3653 S.t1928 VSUBS 0.02fF
C3654 S.n3311 VSUBS 0.14fF $ **FLOATING
C3655 S.n3313 VSUBS 1.16fF $ **FLOATING
C3656 S.n3314 VSUBS 0.22fF $ **FLOATING
C3657 S.n3315 VSUBS 0.25fF $ **FLOATING
C3658 S.n3316 VSUBS 0.09fF $ **FLOATING
C3659 S.n3317 VSUBS 2.44fF $ **FLOATING
C3660 S.t503 VSUBS 0.02fF
C3661 S.n3318 VSUBS 0.24fF $ **FLOATING
C3662 S.n3319 VSUBS 0.91fF $ **FLOATING
C3663 S.n3320 VSUBS 0.05fF $ **FLOATING
C3664 S.t279 VSUBS 0.02fF
C3665 S.n3321 VSUBS 0.12fF $ **FLOATING
C3666 S.n3322 VSUBS 0.14fF $ **FLOATING
C3667 S.n3324 VSUBS 1.88fF $ **FLOATING
C3668 S.n3325 VSUBS 0.48fF $ **FLOATING
C3669 S.n3326 VSUBS 0.09fF $ **FLOATING
C3670 S.n3327 VSUBS 0.33fF $ **FLOATING
C3671 S.n3328 VSUBS 0.30fF $ **FLOATING
C3672 S.n3329 VSUBS 0.77fF $ **FLOATING
C3673 S.n3330 VSUBS 0.59fF $ **FLOATING
C3674 S.t1002 VSUBS 0.02fF
C3675 S.n3331 VSUBS 0.24fF $ **FLOATING
C3676 S.n3332 VSUBS 0.36fF $ **FLOATING
C3677 S.n3333 VSUBS 0.61fF $ **FLOATING
C3678 S.n3334 VSUBS 0.12fF $ **FLOATING
C3679 S.t184 VSUBS 0.02fF
C3680 S.n3335 VSUBS 0.14fF $ **FLOATING
C3681 S.n3337 VSUBS 2.61fF $ **FLOATING
C3682 S.n3338 VSUBS 2.15fF $ **FLOATING
C3683 S.t1286 VSUBS 0.02fF
C3684 S.n3339 VSUBS 0.24fF $ **FLOATING
C3685 S.n3340 VSUBS 0.91fF $ **FLOATING
C3686 S.n3341 VSUBS 0.05fF $ **FLOATING
C3687 S.t1059 VSUBS 0.02fF
C3688 S.n3342 VSUBS 0.12fF $ **FLOATING
C3689 S.n3343 VSUBS 0.14fF $ **FLOATING
C3690 S.n3345 VSUBS 0.78fF $ **FLOATING
C3691 S.n3346 VSUBS 2.30fF $ **FLOATING
C3692 S.n3347 VSUBS 1.88fF $ **FLOATING
C3693 S.n3348 VSUBS 0.12fF $ **FLOATING
C3694 S.t1108 VSUBS 0.02fF
C3695 S.n3349 VSUBS 0.14fF $ **FLOATING
C3696 S.t1786 VSUBS 0.02fF
C3697 S.n3351 VSUBS 0.24fF $ **FLOATING
C3698 S.n3352 VSUBS 0.36fF $ **FLOATING
C3699 S.n3353 VSUBS 0.61fF $ **FLOATING
C3700 S.n3354 VSUBS 1.39fF $ **FLOATING
C3701 S.n3355 VSUBS 0.71fF $ **FLOATING
C3702 S.n3356 VSUBS 1.14fF $ **FLOATING
C3703 S.n3357 VSUBS 0.35fF $ **FLOATING
C3704 S.n3358 VSUBS 2.02fF $ **FLOATING
C3705 S.t2077 VSUBS 0.02fF
C3706 S.n3359 VSUBS 0.24fF $ **FLOATING
C3707 S.n3360 VSUBS 0.91fF $ **FLOATING
C3708 S.n3361 VSUBS 0.05fF $ **FLOATING
C3709 S.t1844 VSUBS 0.02fF
C3710 S.n3362 VSUBS 0.12fF $ **FLOATING
C3711 S.n3363 VSUBS 0.14fF $ **FLOATING
C3712 S.n3365 VSUBS 1.89fF $ **FLOATING
C3713 S.n3366 VSUBS 1.88fF $ **FLOATING
C3714 S.t2564 VSUBS 0.02fF
C3715 S.n3367 VSUBS 0.24fF $ **FLOATING
C3716 S.n3368 VSUBS 0.36fF $ **FLOATING
C3717 S.n3369 VSUBS 0.61fF $ **FLOATING
C3718 S.n3370 VSUBS 0.12fF $ **FLOATING
C3719 S.t261 VSUBS 0.02fF
C3720 S.n3371 VSUBS 0.14fF $ **FLOATING
C3721 S.n3373 VSUBS 1.16fF $ **FLOATING
C3722 S.n3374 VSUBS 0.22fF $ **FLOATING
C3723 S.n3375 VSUBS 0.25fF $ **FLOATING
C3724 S.n3376 VSUBS 0.09fF $ **FLOATING
C3725 S.n3377 VSUBS 1.88fF $ **FLOATING
C3726 S.t887 VSUBS 0.02fF
C3727 S.n3378 VSUBS 0.24fF $ **FLOATING
C3728 S.n3379 VSUBS 0.91fF $ **FLOATING
C3729 S.n3380 VSUBS 0.05fF $ **FLOATING
C3730 S.t1130 VSUBS 0.02fF
C3731 S.n3381 VSUBS 0.12fF $ **FLOATING
C3732 S.n3382 VSUBS 0.14fF $ **FLOATING
C3733 S.n3384 VSUBS 20.78fF $ **FLOATING
C3734 S.n3385 VSUBS 1.88fF $ **FLOATING
C3735 S.n3386 VSUBS 2.68fF $ **FLOATING
C3736 S.t2400 VSUBS 0.02fF
C3737 S.n3387 VSUBS 0.24fF $ **FLOATING
C3738 S.n3388 VSUBS 0.36fF $ **FLOATING
C3739 S.n3389 VSUBS 0.61fF $ **FLOATING
C3740 S.n3390 VSUBS 0.12fF $ **FLOATING
C3741 S.t39 VSUBS 0.02fF
C3742 S.n3391 VSUBS 0.14fF $ **FLOATING
C3743 S.n3393 VSUBS 5.17fF $ **FLOATING
C3744 S.t952 VSUBS 0.02fF
C3745 S.n3394 VSUBS 0.12fF $ **FLOATING
C3746 S.n3395 VSUBS 0.14fF $ **FLOATING
C3747 S.t715 VSUBS 0.02fF
C3748 S.n3397 VSUBS 0.24fF $ **FLOATING
C3749 S.n3398 VSUBS 0.91fF $ **FLOATING
C3750 S.n3399 VSUBS 0.05fF $ **FLOATING
C3751 S.n3400 VSUBS 2.74fF $ **FLOATING
C3752 S.n3401 VSUBS 1.58fF $ **FLOATING
C3753 S.n3402 VSUBS 0.12fF $ **FLOATING
C3754 S.t967 VSUBS 0.02fF
C3755 S.n3403 VSUBS 0.14fF $ **FLOATING
C3756 S.t170 VSUBS 0.02fF
C3757 S.n3405 VSUBS 0.24fF $ **FLOATING
C3758 S.n3406 VSUBS 0.36fF $ **FLOATING
C3759 S.n3407 VSUBS 0.61fF $ **FLOATING
C3760 S.n3408 VSUBS 0.07fF $ **FLOATING
C3761 S.n3409 VSUBS 0.01fF $ **FLOATING
C3762 S.n3410 VSUBS 0.24fF $ **FLOATING
C3763 S.n3411 VSUBS 1.16fF $ **FLOATING
C3764 S.n3412 VSUBS 1.34fF $ **FLOATING
C3765 S.n3413 VSUBS 2.30fF $ **FLOATING
C3766 S.t1734 VSUBS 0.02fF
C3767 S.n3414 VSUBS 0.12fF $ **FLOATING
C3768 S.n3415 VSUBS 0.14fF $ **FLOATING
C3769 S.t1561 VSUBS 0.02fF
C3770 S.n3417 VSUBS 0.24fF $ **FLOATING
C3771 S.n3418 VSUBS 0.91fF $ **FLOATING
C3772 S.n3419 VSUBS 0.05fF $ **FLOATING
C3773 S.t38 VSUBS 48.27fF
C3774 S.t1912 VSUBS 0.02fF
C3775 S.n3420 VSUBS 0.12fF $ **FLOATING
C3776 S.n3421 VSUBS 0.14fF $ **FLOATING
C3777 S.t1669 VSUBS 0.02fF
C3778 S.n3423 VSUBS 0.24fF $ **FLOATING
C3779 S.n3424 VSUBS 0.91fF $ **FLOATING
C3780 S.n3425 VSUBS 0.05fF $ **FLOATING
C3781 S.t831 VSUBS 0.02fF
C3782 S.n3426 VSUBS 0.24fF $ **FLOATING
C3783 S.n3427 VSUBS 0.36fF $ **FLOATING
C3784 S.n3428 VSUBS 0.61fF $ **FLOATING
C3785 S.n3429 VSUBS 0.32fF $ **FLOATING
C3786 S.n3430 VSUBS 1.09fF $ **FLOATING
C3787 S.n3431 VSUBS 0.15fF $ **FLOATING
C3788 S.n3432 VSUBS 2.10fF $ **FLOATING
C3789 S.n3433 VSUBS 2.94fF $ **FLOATING
C3790 S.n3434 VSUBS 1.88fF $ **FLOATING
C3791 S.n3435 VSUBS 0.12fF $ **FLOATING
C3792 S.t1014 VSUBS 0.02fF
C3793 S.n3436 VSUBS 0.14fF $ **FLOATING
C3794 S.t803 VSUBS 0.02fF
C3795 S.n3438 VSUBS 0.24fF $ **FLOATING
C3796 S.n3439 VSUBS 0.36fF $ **FLOATING
C3797 S.n3440 VSUBS 0.61fF $ **FLOATING
C3798 S.n3441 VSUBS 0.92fF $ **FLOATING
C3799 S.n3442 VSUBS 0.32fF $ **FLOATING
C3800 S.n3443 VSUBS 0.92fF $ **FLOATING
C3801 S.n3444 VSUBS 1.09fF $ **FLOATING
C3802 S.n3445 VSUBS 0.15fF $ **FLOATING
C3803 S.n3446 VSUBS 4.96fF $ **FLOATING
C3804 S.t1882 VSUBS 0.02fF
C3805 S.n3447 VSUBS 0.12fF $ **FLOATING
C3806 S.n3448 VSUBS 0.14fF $ **FLOATING
C3807 S.t1944 VSUBS 0.02fF
C3808 S.n3450 VSUBS 0.24fF $ **FLOATING
C3809 S.n3451 VSUBS 0.91fF $ **FLOATING
C3810 S.n3452 VSUBS 0.05fF $ **FLOATING
C3811 S.n3453 VSUBS 1.88fF $ **FLOATING
C3812 S.n3454 VSUBS 2.67fF $ **FLOATING
C3813 S.t1582 VSUBS 0.02fF
C3814 S.n3455 VSUBS 0.24fF $ **FLOATING
C3815 S.n3456 VSUBS 0.36fF $ **FLOATING
C3816 S.n3457 VSUBS 0.61fF $ **FLOATING
C3817 S.n3458 VSUBS 0.12fF $ **FLOATING
C3818 S.t1793 VSUBS 0.02fF
C3819 S.n3459 VSUBS 0.14fF $ **FLOATING
C3820 S.n3461 VSUBS 1.88fF $ **FLOATING
C3821 S.n3462 VSUBS 2.67fF $ **FLOATING
C3822 S.t1614 VSUBS 0.02fF
C3823 S.n3463 VSUBS 0.24fF $ **FLOATING
C3824 S.n3464 VSUBS 0.36fF $ **FLOATING
C3825 S.n3465 VSUBS 0.61fF $ **FLOATING
C3826 S.t2457 VSUBS 0.02fF
C3827 S.n3466 VSUBS 0.24fF $ **FLOATING
C3828 S.n3467 VSUBS 0.91fF $ **FLOATING
C3829 S.n3468 VSUBS 0.05fF $ **FLOATING
C3830 S.t164 VSUBS 0.02fF
C3831 S.n3469 VSUBS 0.12fF $ **FLOATING
C3832 S.n3470 VSUBS 0.14fF $ **FLOATING
C3833 S.n3472 VSUBS 0.12fF $ **FLOATING
C3834 S.t1824 VSUBS 0.02fF
C3835 S.n3473 VSUBS 0.14fF $ **FLOATING
C3836 S.n3475 VSUBS 2.30fF $ **FLOATING
C3837 S.n3476 VSUBS 2.94fF $ **FLOATING
C3838 S.n3477 VSUBS 4.88fF $ **FLOATING
C3839 S.t132 VSUBS 0.02fF
C3840 S.n3478 VSUBS 0.12fF $ **FLOATING
C3841 S.n3479 VSUBS 0.14fF $ **FLOATING
C3842 S.t201 VSUBS 0.02fF
C3843 S.n3481 VSUBS 0.24fF $ **FLOATING
C3844 S.n3482 VSUBS 0.91fF $ **FLOATING
C3845 S.n3483 VSUBS 0.05fF $ **FLOATING
C3846 S.n3484 VSUBS 1.88fF $ **FLOATING
C3847 S.n3485 VSUBS 2.67fF $ **FLOATING
C3848 S.t2375 VSUBS 0.02fF
C3849 S.n3486 VSUBS 0.24fF $ **FLOATING
C3850 S.n3487 VSUBS 0.36fF $ **FLOATING
C3851 S.n3488 VSUBS 0.61fF $ **FLOATING
C3852 S.n3489 VSUBS 0.12fF $ **FLOATING
C3853 S.t2575 VSUBS 0.02fF
C3854 S.n3490 VSUBS 0.14fF $ **FLOATING
C3855 S.n3492 VSUBS 5.44fF $ **FLOATING
C3856 S.t929 VSUBS 0.02fF
C3857 S.n3493 VSUBS 0.12fF $ **FLOATING
C3858 S.n3494 VSUBS 0.14fF $ **FLOATING
C3859 S.t990 VSUBS 0.02fF
C3860 S.n3496 VSUBS 0.24fF $ **FLOATING
C3861 S.n3497 VSUBS 0.91fF $ **FLOATING
C3862 S.n3498 VSUBS 0.05fF $ **FLOATING
C3863 S.t84 VSUBS 47.89fF
C3864 S.t2327 VSUBS 0.02fF
C3865 S.n3499 VSUBS 0.01fF $ **FLOATING
C3866 S.n3500 VSUBS 0.26fF $ **FLOATING
C3867 S.t1513 VSUBS 0.02fF
C3868 S.n3502 VSUBS 1.19fF $ **FLOATING
C3869 S.n3503 VSUBS 0.05fF $ **FLOATING
C3870 S.t2306 VSUBS 0.02fF
C3871 S.n3504 VSUBS 0.64fF $ **FLOATING
C3872 S.n3505 VSUBS 0.61fF $ **FLOATING
C3873 S.n3506 VSUBS 8.97fF $ **FLOATING
C3874 S.n3507 VSUBS 0.77fF $ **FLOATING
C3875 S.n3508 VSUBS 0.28fF $ **FLOATING
C3876 S.n3509 VSUBS 0.60fF $ **FLOATING
C3877 S.n3510 VSUBS 0.22fF $ **FLOATING
C3878 S.n3511 VSUBS 0.59fF $ **FLOATING
C3879 S.n3512 VSUBS 3.39fF $ **FLOATING
C3880 S.n3513 VSUBS 0.29fF $ **FLOATING
C3881 S.t128 VSUBS 21.42fF
C3882 S.n3514 VSUBS 21.71fF $ **FLOATING
C3883 S.n3515 VSUBS 8.97fF $ **FLOATING
C3884 S.n3516 VSUBS 4.00fF $ **FLOATING
C3885 S.n3517 VSUBS 1.35fF $ **FLOATING
C3886 S.n3518 VSUBS 0.01fF $ **FLOATING
C3887 S.n3519 VSUBS 0.02fF $ **FLOATING
C3888 S.n3520 VSUBS 0.03fF $ **FLOATING
C3889 S.n3521 VSUBS 0.04fF $ **FLOATING
C3890 S.n3522 VSUBS 0.17fF $ **FLOATING
C3891 S.n3523 VSUBS 0.01fF $ **FLOATING
C3892 S.n3524 VSUBS 0.02fF $ **FLOATING
C3893 S.n3525 VSUBS 0.01fF $ **FLOATING
C3894 S.n3526 VSUBS 0.01fF $ **FLOATING
C3895 S.n3527 VSUBS 0.01fF $ **FLOATING
C3896 S.n3528 VSUBS 0.01fF $ **FLOATING
C3897 S.n3529 VSUBS 0.02fF $ **FLOATING
C3898 S.n3530 VSUBS 0.01fF $ **FLOATING
C3899 S.n3531 VSUBS 0.02fF $ **FLOATING
C3900 S.n3532 VSUBS 0.05fF $ **FLOATING
C3901 S.n3533 VSUBS 0.04fF $ **FLOATING
C3902 S.n3534 VSUBS 0.11fF $ **FLOATING
C3903 S.n3535 VSUBS 0.38fF $ **FLOATING
C3904 S.n3536 VSUBS 0.20fF $ **FLOATING
C3905 S.n3537 VSUBS 4.42fF $ **FLOATING
C3906 S.n3538 VSUBS 0.24fF $ **FLOATING
C3907 S.n3539 VSUBS 1.50fF $ **FLOATING
C3908 S.n3540 VSUBS 1.31fF $ **FLOATING
C3909 S.n3541 VSUBS 0.28fF $ **FLOATING
C3910 S.n3542 VSUBS 1.89fF $ **FLOATING
C3911 S.n3543 VSUBS 0.06fF $ **FLOATING
C3912 S.n3544 VSUBS 0.03fF $ **FLOATING
C3913 S.n3545 VSUBS 0.04fF $ **FLOATING
C3914 S.n3546 VSUBS 0.99fF $ **FLOATING
C3915 S.n3547 VSUBS 0.02fF $ **FLOATING
C3916 S.n3548 VSUBS 0.01fF $ **FLOATING
C3917 S.n3549 VSUBS 0.02fF $ **FLOATING
C3918 S.n3550 VSUBS 0.08fF $ **FLOATING
C3919 S.n3551 VSUBS 0.36fF $ **FLOATING
C3920 S.n3552 VSUBS 1.85fF $ **FLOATING
C3921 S.t1644 VSUBS 0.02fF
C3922 S.n3553 VSUBS 0.24fF $ **FLOATING
C3923 S.n3554 VSUBS 0.36fF $ **FLOATING
C3924 S.n3555 VSUBS 0.61fF $ **FLOATING
C3925 S.n3556 VSUBS 0.12fF $ **FLOATING
C3926 S.t828 VSUBS 0.02fF
C3927 S.n3557 VSUBS 0.14fF $ **FLOATING
C3928 S.n3559 VSUBS 0.70fF $ **FLOATING
C3929 S.n3560 VSUBS 0.23fF $ **FLOATING
C3930 S.n3561 VSUBS 0.23fF $ **FLOATING
C3931 S.n3562 VSUBS 0.70fF $ **FLOATING
C3932 S.n3563 VSUBS 1.16fF $ **FLOATING
C3933 S.n3564 VSUBS 0.22fF $ **FLOATING
C3934 S.n3565 VSUBS 0.25fF $ **FLOATING
C3935 S.n3566 VSUBS 0.09fF $ **FLOATING
C3936 S.n3567 VSUBS 1.88fF $ **FLOATING
C3937 S.t1943 VSUBS 0.02fF
C3938 S.n3568 VSUBS 0.24fF $ **FLOATING
C3939 S.n3569 VSUBS 0.91fF $ **FLOATING
C3940 S.n3570 VSUBS 0.05fF $ **FLOATING
C3941 S.t1693 VSUBS 0.02fF
C3942 S.n3571 VSUBS 0.12fF $ **FLOATING
C3943 S.n3572 VSUBS 0.14fF $ **FLOATING
C3944 S.n3574 VSUBS 0.25fF $ **FLOATING
C3945 S.n3575 VSUBS 0.09fF $ **FLOATING
C3946 S.n3576 VSUBS 0.21fF $ **FLOATING
C3947 S.n3577 VSUBS 0.92fF $ **FLOATING
C3948 S.n3578 VSUBS 0.44fF $ **FLOATING
C3949 S.n3579 VSUBS 1.88fF $ **FLOATING
C3950 S.n3580 VSUBS 0.12fF $ **FLOATING
C3951 S.t1741 VSUBS 0.02fF
C3952 S.n3581 VSUBS 0.14fF $ **FLOATING
C3953 S.t2552 VSUBS 0.02fF
C3954 S.n3583 VSUBS 0.24fF $ **FLOATING
C3955 S.n3584 VSUBS 0.36fF $ **FLOATING
C3956 S.n3585 VSUBS 0.61fF $ **FLOATING
C3957 S.n3586 VSUBS 0.02fF $ **FLOATING
C3958 S.n3587 VSUBS 0.01fF $ **FLOATING
C3959 S.n3588 VSUBS 0.02fF $ **FLOATING
C3960 S.n3589 VSUBS 0.08fF $ **FLOATING
C3961 S.n3590 VSUBS 0.06fF $ **FLOATING
C3962 S.n3591 VSUBS 0.03fF $ **FLOATING
C3963 S.n3592 VSUBS 0.04fF $ **FLOATING
C3964 S.n3593 VSUBS 1.00fF $ **FLOATING
C3965 S.n3594 VSUBS 0.36fF $ **FLOATING
C3966 S.n3595 VSUBS 1.87fF $ **FLOATING
C3967 S.n3596 VSUBS 1.99fF $ **FLOATING
C3968 S.t333 VSUBS 0.02fF
C3969 S.n3597 VSUBS 0.24fF $ **FLOATING
C3970 S.n3598 VSUBS 0.91fF $ **FLOATING
C3971 S.n3599 VSUBS 0.05fF $ **FLOATING
C3972 S.t54 VSUBS 0.02fF
C3973 S.n3600 VSUBS 0.12fF $ **FLOATING
C3974 S.n3601 VSUBS 0.14fF $ **FLOATING
C3975 S.n3603 VSUBS 1.89fF $ **FLOATING
C3976 S.n3604 VSUBS 0.06fF $ **FLOATING
C3977 S.n3605 VSUBS 0.03fF $ **FLOATING
C3978 S.n3606 VSUBS 0.04fF $ **FLOATING
C3979 S.n3607 VSUBS 0.99fF $ **FLOATING
C3980 S.n3608 VSUBS 0.02fF $ **FLOATING
C3981 S.n3609 VSUBS 0.01fF $ **FLOATING
C3982 S.n3610 VSUBS 0.02fF $ **FLOATING
C3983 S.n3611 VSUBS 0.08fF $ **FLOATING
C3984 S.n3612 VSUBS 0.36fF $ **FLOATING
C3985 S.n3613 VSUBS 1.85fF $ **FLOATING
C3986 S.t2173 VSUBS 0.02fF
C3987 S.n3614 VSUBS 0.24fF $ **FLOATING
C3988 S.n3615 VSUBS 0.36fF $ **FLOATING
C3989 S.n3616 VSUBS 0.61fF $ **FLOATING
C3990 S.n3617 VSUBS 0.12fF $ **FLOATING
C3991 S.t1359 VSUBS 0.02fF
C3992 S.n3618 VSUBS 0.14fF $ **FLOATING
C3993 S.n3620 VSUBS 0.70fF $ **FLOATING
C3994 S.n3621 VSUBS 0.23fF $ **FLOATING
C3995 S.n3622 VSUBS 0.23fF $ **FLOATING
C3996 S.n3623 VSUBS 0.70fF $ **FLOATING
C3997 S.n3624 VSUBS 1.16fF $ **FLOATING
C3998 S.n3625 VSUBS 0.22fF $ **FLOATING
C3999 S.n3626 VSUBS 0.25fF $ **FLOATING
C4000 S.n3627 VSUBS 0.09fF $ **FLOATING
C4001 S.n3628 VSUBS 1.88fF $ **FLOATING
C4002 S.t2451 VSUBS 0.02fF
C4003 S.n3629 VSUBS 0.24fF $ **FLOATING
C4004 S.n3630 VSUBS 0.91fF $ **FLOATING
C4005 S.n3631 VSUBS 0.05fF $ **FLOATING
C4006 S.t870 VSUBS 0.02fF
C4007 S.n3632 VSUBS 0.12fF $ **FLOATING
C4008 S.n3633 VSUBS 0.14fF $ **FLOATING
C4009 S.n3635 VSUBS 0.25fF $ **FLOATING
C4010 S.n3636 VSUBS 0.09fF $ **FLOATING
C4011 S.n3637 VSUBS 0.21fF $ **FLOATING
C4012 S.n3638 VSUBS 0.92fF $ **FLOATING
C4013 S.n3639 VSUBS 0.44fF $ **FLOATING
C4014 S.n3640 VSUBS 1.88fF $ **FLOATING
C4015 S.n3641 VSUBS 0.12fF $ **FLOATING
C4016 S.t2143 VSUBS 0.02fF
C4017 S.n3642 VSUBS 0.14fF $ **FLOATING
C4018 S.t438 VSUBS 0.02fF
C4019 S.n3644 VSUBS 0.24fF $ **FLOATING
C4020 S.n3645 VSUBS 0.36fF $ **FLOATING
C4021 S.n3646 VSUBS 0.61fF $ **FLOATING
C4022 S.n3647 VSUBS 0.02fF $ **FLOATING
C4023 S.n3648 VSUBS 0.01fF $ **FLOATING
C4024 S.n3649 VSUBS 0.02fF $ **FLOATING
C4025 S.n3650 VSUBS 0.08fF $ **FLOATING
C4026 S.n3651 VSUBS 0.06fF $ **FLOATING
C4027 S.n3652 VSUBS 0.03fF $ **FLOATING
C4028 S.n3653 VSUBS 0.04fF $ **FLOATING
C4029 S.n3654 VSUBS 1.00fF $ **FLOATING
C4030 S.n3655 VSUBS 0.36fF $ **FLOATING
C4031 S.n3656 VSUBS 1.87fF $ **FLOATING
C4032 S.n3657 VSUBS 1.99fF $ **FLOATING
C4033 S.t708 VSUBS 0.02fF
C4034 S.n3658 VSUBS 0.24fF $ **FLOATING
C4035 S.n3659 VSUBS 0.91fF $ **FLOATING
C4036 S.n3660 VSUBS 0.05fF $ **FLOATING
C4037 S.t490 VSUBS 0.02fF
C4038 S.n3661 VSUBS 0.12fF $ **FLOATING
C4039 S.n3662 VSUBS 0.14fF $ **FLOATING
C4040 S.n3664 VSUBS 1.89fF $ **FLOATING
C4041 S.n3665 VSUBS 0.06fF $ **FLOATING
C4042 S.n3666 VSUBS 0.03fF $ **FLOATING
C4043 S.n3667 VSUBS 0.04fF $ **FLOATING
C4044 S.n3668 VSUBS 0.99fF $ **FLOATING
C4045 S.n3669 VSUBS 0.02fF $ **FLOATING
C4046 S.n3670 VSUBS 0.01fF $ **FLOATING
C4047 S.n3671 VSUBS 0.02fF $ **FLOATING
C4048 S.n3672 VSUBS 0.08fF $ **FLOATING
C4049 S.n3673 VSUBS 0.36fF $ **FLOATING
C4050 S.n3674 VSUBS 1.85fF $ **FLOATING
C4051 S.t1231 VSUBS 0.02fF
C4052 S.n3675 VSUBS 0.24fF $ **FLOATING
C4053 S.n3676 VSUBS 0.36fF $ **FLOATING
C4054 S.n3677 VSUBS 0.61fF $ **FLOATING
C4055 S.n3678 VSUBS 0.12fF $ **FLOATING
C4056 S.t413 VSUBS 0.02fF
C4057 S.n3679 VSUBS 0.14fF $ **FLOATING
C4058 S.n3681 VSUBS 0.70fF $ **FLOATING
C4059 S.n3682 VSUBS 0.23fF $ **FLOATING
C4060 S.n3683 VSUBS 0.23fF $ **FLOATING
C4061 S.n3684 VSUBS 0.70fF $ **FLOATING
C4062 S.n3685 VSUBS 1.16fF $ **FLOATING
C4063 S.n3686 VSUBS 0.22fF $ **FLOATING
C4064 S.n3687 VSUBS 0.25fF $ **FLOATING
C4065 S.n3688 VSUBS 0.09fF $ **FLOATING
C4066 S.n3689 VSUBS 1.88fF $ **FLOATING
C4067 S.t1501 VSUBS 0.02fF
C4068 S.n3690 VSUBS 0.24fF $ **FLOATING
C4069 S.n3691 VSUBS 0.91fF $ **FLOATING
C4070 S.n3692 VSUBS 0.05fF $ **FLOATING
C4071 S.t1276 VSUBS 0.02fF
C4072 S.n3693 VSUBS 0.12fF $ **FLOATING
C4073 S.n3694 VSUBS 0.14fF $ **FLOATING
C4074 S.n3696 VSUBS 0.25fF $ **FLOATING
C4075 S.n3697 VSUBS 0.09fF $ **FLOATING
C4076 S.n3698 VSUBS 0.21fF $ **FLOATING
C4077 S.n3699 VSUBS 0.92fF $ **FLOATING
C4078 S.n3700 VSUBS 0.44fF $ **FLOATING
C4079 S.n3701 VSUBS 1.88fF $ **FLOATING
C4080 S.n3702 VSUBS 0.12fF $ **FLOATING
C4081 S.t1205 VSUBS 0.02fF
C4082 S.n3703 VSUBS 0.14fF $ **FLOATING
C4083 S.t2012 VSUBS 0.02fF
C4084 S.n3705 VSUBS 0.24fF $ **FLOATING
C4085 S.n3706 VSUBS 0.36fF $ **FLOATING
C4086 S.n3707 VSUBS 0.61fF $ **FLOATING
C4087 S.n3708 VSUBS 0.02fF $ **FLOATING
C4088 S.n3709 VSUBS 0.01fF $ **FLOATING
C4089 S.n3710 VSUBS 0.02fF $ **FLOATING
C4090 S.n3711 VSUBS 0.08fF $ **FLOATING
C4091 S.n3712 VSUBS 0.06fF $ **FLOATING
C4092 S.n3713 VSUBS 0.03fF $ **FLOATING
C4093 S.n3714 VSUBS 0.04fF $ **FLOATING
C4094 S.n3715 VSUBS 1.00fF $ **FLOATING
C4095 S.n3716 VSUBS 0.36fF $ **FLOATING
C4096 S.n3717 VSUBS 1.87fF $ **FLOATING
C4097 S.n3718 VSUBS 1.99fF $ **FLOATING
C4098 S.t2288 VSUBS 0.02fF
C4099 S.n3719 VSUBS 0.24fF $ **FLOATING
C4100 S.n3720 VSUBS 0.91fF $ **FLOATING
C4101 S.n3721 VSUBS 0.05fF $ **FLOATING
C4102 S.t2066 VSUBS 0.02fF
C4103 S.n3722 VSUBS 0.12fF $ **FLOATING
C4104 S.n3723 VSUBS 0.14fF $ **FLOATING
C4105 S.n3725 VSUBS 1.89fF $ **FLOATING
C4106 S.n3726 VSUBS 0.06fF $ **FLOATING
C4107 S.n3727 VSUBS 0.03fF $ **FLOATING
C4108 S.n3728 VSUBS 0.04fF $ **FLOATING
C4109 S.n3729 VSUBS 0.99fF $ **FLOATING
C4110 S.n3730 VSUBS 0.02fF $ **FLOATING
C4111 S.n3731 VSUBS 0.01fF $ **FLOATING
C4112 S.n3732 VSUBS 0.02fF $ **FLOATING
C4113 S.n3733 VSUBS 0.08fF $ **FLOATING
C4114 S.n3734 VSUBS 0.36fF $ **FLOATING
C4115 S.n3735 VSUBS 1.85fF $ **FLOATING
C4116 S.t406 VSUBS 0.02fF
C4117 S.n3736 VSUBS 0.24fF $ **FLOATING
C4118 S.n3737 VSUBS 0.36fF $ **FLOATING
C4119 S.n3738 VSUBS 0.61fF $ **FLOATING
C4120 S.n3739 VSUBS 0.12fF $ **FLOATING
C4121 S.t2110 VSUBS 0.02fF
C4122 S.n3740 VSUBS 0.14fF $ **FLOATING
C4123 S.n3742 VSUBS 0.70fF $ **FLOATING
C4124 S.n3743 VSUBS 0.23fF $ **FLOATING
C4125 S.n3744 VSUBS 0.23fF $ **FLOATING
C4126 S.n3745 VSUBS 0.70fF $ **FLOATING
C4127 S.n3746 VSUBS 1.16fF $ **FLOATING
C4128 S.n3747 VSUBS 0.22fF $ **FLOATING
C4129 S.n3748 VSUBS 0.25fF $ **FLOATING
C4130 S.n3749 VSUBS 0.09fF $ **FLOATING
C4131 S.n3750 VSUBS 1.88fF $ **FLOATING
C4132 S.t676 VSUBS 0.02fF
C4133 S.n3751 VSUBS 0.24fF $ **FLOATING
C4134 S.n3752 VSUBS 0.91fF $ **FLOATING
C4135 S.n3753 VSUBS 0.05fF $ **FLOATING
C4136 S.t454 VSUBS 0.02fF
C4137 S.n3754 VSUBS 0.12fF $ **FLOATING
C4138 S.n3755 VSUBS 0.14fF $ **FLOATING
C4139 S.n3757 VSUBS 0.25fF $ **FLOATING
C4140 S.n3758 VSUBS 0.09fF $ **FLOATING
C4141 S.n3759 VSUBS 0.21fF $ **FLOATING
C4142 S.n3760 VSUBS 0.92fF $ **FLOATING
C4143 S.n3761 VSUBS 0.44fF $ **FLOATING
C4144 S.n3762 VSUBS 1.88fF $ **FLOATING
C4145 S.n3763 VSUBS 0.12fF $ **FLOATING
C4146 S.t1710 VSUBS 0.02fF
C4147 S.n3764 VSUBS 0.14fF $ **FLOATING
C4148 S.t2523 VSUBS 0.02fF
C4149 S.n3766 VSUBS 0.24fF $ **FLOATING
C4150 S.n3767 VSUBS 0.36fF $ **FLOATING
C4151 S.n3768 VSUBS 0.61fF $ **FLOATING
C4152 S.n3769 VSUBS 0.02fF $ **FLOATING
C4153 S.n3770 VSUBS 0.01fF $ **FLOATING
C4154 S.n3771 VSUBS 0.02fF $ **FLOATING
C4155 S.n3772 VSUBS 0.08fF $ **FLOATING
C4156 S.n3773 VSUBS 0.06fF $ **FLOATING
C4157 S.n3774 VSUBS 0.03fF $ **FLOATING
C4158 S.n3775 VSUBS 0.04fF $ **FLOATING
C4159 S.n3776 VSUBS 1.00fF $ **FLOATING
C4160 S.n3777 VSUBS 0.36fF $ **FLOATING
C4161 S.n3778 VSUBS 1.87fF $ **FLOATING
C4162 S.n3779 VSUBS 1.99fF $ **FLOATING
C4163 S.t304 VSUBS 0.02fF
C4164 S.n3780 VSUBS 0.24fF $ **FLOATING
C4165 S.n3781 VSUBS 0.91fF $ **FLOATING
C4166 S.n3782 VSUBS 0.05fF $ **FLOATING
C4167 S.t2580 VSUBS 0.02fF
C4168 S.n3783 VSUBS 0.12fF $ **FLOATING
C4169 S.n3784 VSUBS 0.14fF $ **FLOATING
C4170 S.n3786 VSUBS 1.89fF $ **FLOATING
C4171 S.n3787 VSUBS 0.07fF $ **FLOATING
C4172 S.n3788 VSUBS 0.04fF $ **FLOATING
C4173 S.n3789 VSUBS 0.05fF $ **FLOATING
C4174 S.n3790 VSUBS 0.87fF $ **FLOATING
C4175 S.n3791 VSUBS 0.01fF $ **FLOATING
C4176 S.n3792 VSUBS 0.01fF $ **FLOATING
C4177 S.n3793 VSUBS 0.01fF $ **FLOATING
C4178 S.n3794 VSUBS 0.07fF $ **FLOATING
C4179 S.n3795 VSUBS 0.68fF $ **FLOATING
C4180 S.n3796 VSUBS 0.72fF $ **FLOATING
C4181 S.t783 VSUBS 0.02fF
C4182 S.n3797 VSUBS 0.24fF $ **FLOATING
C4183 S.n3798 VSUBS 0.36fF $ **FLOATING
C4184 S.n3799 VSUBS 0.61fF $ **FLOATING
C4185 S.n3800 VSUBS 0.12fF $ **FLOATING
C4186 S.t2497 VSUBS 0.02fF
C4187 S.n3801 VSUBS 0.14fF $ **FLOATING
C4188 S.n3803 VSUBS 0.70fF $ **FLOATING
C4189 S.n3804 VSUBS 0.23fF $ **FLOATING
C4190 S.n3805 VSUBS 0.23fF $ **FLOATING
C4191 S.n3806 VSUBS 0.70fF $ **FLOATING
C4192 S.n3807 VSUBS 1.16fF $ **FLOATING
C4193 S.n3808 VSUBS 0.22fF $ **FLOATING
C4194 S.n3809 VSUBS 0.25fF $ **FLOATING
C4195 S.n3810 VSUBS 0.09fF $ **FLOATING
C4196 S.n3811 VSUBS 2.31fF $ **FLOATING
C4197 S.t1088 VSUBS 0.02fF
C4198 S.n3812 VSUBS 0.24fF $ **FLOATING
C4199 S.n3813 VSUBS 0.91fF $ **FLOATING
C4200 S.n3814 VSUBS 0.05fF $ **FLOATING
C4201 S.t842 VSUBS 0.02fF
C4202 S.n3815 VSUBS 0.12fF $ **FLOATING
C4203 S.n3816 VSUBS 0.14fF $ **FLOATING
C4204 S.n3818 VSUBS 1.88fF $ **FLOATING
C4205 S.n3819 VSUBS 0.46fF $ **FLOATING
C4206 S.n3820 VSUBS 0.22fF $ **FLOATING
C4207 S.n3821 VSUBS 0.38fF $ **FLOATING
C4208 S.n3822 VSUBS 0.16fF $ **FLOATING
C4209 S.n3823 VSUBS 0.28fF $ **FLOATING
C4210 S.n3824 VSUBS 0.21fF $ **FLOATING
C4211 S.n3825 VSUBS 0.30fF $ **FLOATING
C4212 S.n3826 VSUBS 0.42fF $ **FLOATING
C4213 S.n3827 VSUBS 0.21fF $ **FLOATING
C4214 S.t1568 VSUBS 0.02fF
C4215 S.n3828 VSUBS 0.24fF $ **FLOATING
C4216 S.n3829 VSUBS 0.36fF $ **FLOATING
C4217 S.n3830 VSUBS 0.61fF $ **FLOATING
C4218 S.n3831 VSUBS 0.12fF $ **FLOATING
C4219 S.t753 VSUBS 0.02fF
C4220 S.n3832 VSUBS 0.14fF $ **FLOATING
C4221 S.n3834 VSUBS 0.04fF $ **FLOATING
C4222 S.n3835 VSUBS 0.03fF $ **FLOATING
C4223 S.n3836 VSUBS 0.03fF $ **FLOATING
C4224 S.n3837 VSUBS 0.10fF $ **FLOATING
C4225 S.n3838 VSUBS 0.36fF $ **FLOATING
C4226 S.n3839 VSUBS 0.38fF $ **FLOATING
C4227 S.n3840 VSUBS 0.11fF $ **FLOATING
C4228 S.n3841 VSUBS 0.12fF $ **FLOATING
C4229 S.n3842 VSUBS 0.07fF $ **FLOATING
C4230 S.n3843 VSUBS 0.12fF $ **FLOATING
C4231 S.n3844 VSUBS 0.18fF $ **FLOATING
C4232 S.n3845 VSUBS 3.99fF $ **FLOATING
C4233 S.t1868 VSUBS 0.02fF
C4234 S.n3846 VSUBS 0.24fF $ **FLOATING
C4235 S.n3847 VSUBS 0.91fF $ **FLOATING
C4236 S.n3848 VSUBS 0.05fF $ **FLOATING
C4237 S.t1625 VSUBS 0.02fF
C4238 S.n3849 VSUBS 0.12fF $ **FLOATING
C4239 S.n3850 VSUBS 0.14fF $ **FLOATING
C4240 S.n3852 VSUBS 0.25fF $ **FLOATING
C4241 S.n3853 VSUBS 0.09fF $ **FLOATING
C4242 S.n3854 VSUBS 0.21fF $ **FLOATING
C4243 S.n3855 VSUBS 1.28fF $ **FLOATING
C4244 S.n3856 VSUBS 0.53fF $ **FLOATING
C4245 S.n3857 VSUBS 1.88fF $ **FLOATING
C4246 S.n3858 VSUBS 0.12fF $ **FLOATING
C4247 S.t1546 VSUBS 0.02fF
C4248 S.n3859 VSUBS 0.14fF $ **FLOATING
C4249 S.t2358 VSUBS 0.02fF
C4250 S.n3861 VSUBS 0.24fF $ **FLOATING
C4251 S.n3862 VSUBS 0.36fF $ **FLOATING
C4252 S.n3863 VSUBS 0.61fF $ **FLOATING
C4253 S.n3864 VSUBS 1.58fF $ **FLOATING
C4254 S.n3865 VSUBS 2.45fF $ **FLOATING
C4255 S.t112 VSUBS 0.02fF
C4256 S.n3866 VSUBS 0.24fF $ **FLOATING
C4257 S.n3867 VSUBS 0.91fF $ **FLOATING
C4258 S.n3868 VSUBS 0.05fF $ **FLOATING
C4259 S.t2412 VSUBS 0.02fF
C4260 S.n3869 VSUBS 0.12fF $ **FLOATING
C4261 S.n3870 VSUBS 0.14fF $ **FLOATING
C4262 S.n3872 VSUBS 1.89fF $ **FLOATING
C4263 S.n3873 VSUBS 0.06fF $ **FLOATING
C4264 S.n3874 VSUBS 0.03fF $ **FLOATING
C4265 S.n3875 VSUBS 0.04fF $ **FLOATING
C4266 S.n3876 VSUBS 0.99fF $ **FLOATING
C4267 S.n3877 VSUBS 0.02fF $ **FLOATING
C4268 S.n3878 VSUBS 0.01fF $ **FLOATING
C4269 S.n3879 VSUBS 0.02fF $ **FLOATING
C4270 S.n3880 VSUBS 0.08fF $ **FLOATING
C4271 S.n3881 VSUBS 0.36fF $ **FLOATING
C4272 S.n3882 VSUBS 1.85fF $ **FLOATING
C4273 S.t20 VSUBS 0.02fF
C4274 S.n3883 VSUBS 0.24fF $ **FLOATING
C4275 S.n3884 VSUBS 0.36fF $ **FLOATING
C4276 S.n3885 VSUBS 0.61fF $ **FLOATING
C4277 S.n3886 VSUBS 0.12fF $ **FLOATING
C4278 S.t286 VSUBS 0.02fF
C4279 S.n3887 VSUBS 0.14fF $ **FLOATING
C4280 S.n3889 VSUBS 0.70fF $ **FLOATING
C4281 S.n3890 VSUBS 0.23fF $ **FLOATING
C4282 S.n3891 VSUBS 0.23fF $ **FLOATING
C4283 S.n3892 VSUBS 0.70fF $ **FLOATING
C4284 S.n3893 VSUBS 1.16fF $ **FLOATING
C4285 S.n3894 VSUBS 0.22fF $ **FLOATING
C4286 S.n3895 VSUBS 0.25fF $ **FLOATING
C4287 S.n3896 VSUBS 0.09fF $ **FLOATING
C4288 S.n3897 VSUBS 1.88fF $ **FLOATING
C4289 S.t916 VSUBS 0.02fF
C4290 S.n3898 VSUBS 0.24fF $ **FLOATING
C4291 S.n3899 VSUBS 0.91fF $ **FLOATING
C4292 S.n3900 VSUBS 0.05fF $ **FLOATING
C4293 S.t809 VSUBS 0.02fF
C4294 S.n3901 VSUBS 0.12fF $ **FLOATING
C4295 S.n3902 VSUBS 0.14fF $ **FLOATING
C4296 S.n3904 VSUBS 20.78fF $ **FLOATING
C4297 S.n3905 VSUBS 0.06fF $ **FLOATING
C4298 S.n3906 VSUBS 0.20fF $ **FLOATING
C4299 S.n3907 VSUBS 0.09fF $ **FLOATING
C4300 S.n3908 VSUBS 0.21fF $ **FLOATING
C4301 S.n3909 VSUBS 0.10fF $ **FLOATING
C4302 S.n3910 VSUBS 0.30fF $ **FLOATING
C4303 S.n3911 VSUBS 0.69fF $ **FLOATING
C4304 S.n3912 VSUBS 0.45fF $ **FLOATING
C4305 S.n3913 VSUBS 2.33fF $ **FLOATING
C4306 S.n3914 VSUBS 0.12fF $ **FLOATING
C4307 S.t2562 VSUBS 0.02fF
C4308 S.n3915 VSUBS 0.14fF $ **FLOATING
C4309 S.t860 VSUBS 0.02fF
C4310 S.n3917 VSUBS 0.24fF $ **FLOATING
C4311 S.n3918 VSUBS 0.36fF $ **FLOATING
C4312 S.n3919 VSUBS 0.61fF $ **FLOATING
C4313 S.n3920 VSUBS 1.90fF $ **FLOATING
C4314 S.n3921 VSUBS 0.17fF $ **FLOATING
C4315 S.n3922 VSUBS 0.76fF $ **FLOATING
C4316 S.n3923 VSUBS 0.25fF $ **FLOATING
C4317 S.n3924 VSUBS 0.30fF $ **FLOATING
C4318 S.n3925 VSUBS 0.32fF $ **FLOATING
C4319 S.n3926 VSUBS 0.47fF $ **FLOATING
C4320 S.n3927 VSUBS 0.16fF $ **FLOATING
C4321 S.n3928 VSUBS 1.93fF $ **FLOATING
C4322 S.t914 VSUBS 0.02fF
C4323 S.n3929 VSUBS 0.12fF $ **FLOATING
C4324 S.n3930 VSUBS 0.14fF $ **FLOATING
C4325 S.t1158 VSUBS 0.02fF
C4326 S.n3932 VSUBS 0.24fF $ **FLOATING
C4327 S.n3933 VSUBS 0.91fF $ **FLOATING
C4328 S.n3934 VSUBS 0.05fF $ **FLOATING
C4329 S.n3935 VSUBS 1.88fF $ **FLOATING
C4330 S.n3936 VSUBS 0.12fF $ **FLOATING
C4331 S.t1094 VSUBS 0.02fF
C4332 S.n3937 VSUBS 0.14fF $ **FLOATING
C4333 S.t1962 VSUBS 0.02fF
C4334 S.n3939 VSUBS 0.12fF $ **FLOATING
C4335 S.n3940 VSUBS 0.14fF $ **FLOATING
C4336 S.t1722 VSUBS 0.02fF
C4337 S.n3942 VSUBS 0.24fF $ **FLOATING
C4338 S.n3943 VSUBS 0.91fF $ **FLOATING
C4339 S.n3944 VSUBS 0.05fF $ **FLOATING
C4340 S.t882 VSUBS 0.02fF
C4341 S.n3945 VSUBS 0.24fF $ **FLOATING
C4342 S.n3946 VSUBS 0.36fF $ **FLOATING
C4343 S.n3947 VSUBS 0.61fF $ **FLOATING
C4344 S.n3948 VSUBS 0.32fF $ **FLOATING
C4345 S.n3949 VSUBS 1.09fF $ **FLOATING
C4346 S.n3950 VSUBS 0.15fF $ **FLOATING
C4347 S.n3951 VSUBS 2.10fF $ **FLOATING
C4348 S.n3952 VSUBS 2.94fF $ **FLOATING
C4349 S.n3953 VSUBS 1.88fF $ **FLOATING
C4350 S.n3954 VSUBS 0.12fF $ **FLOATING
C4351 S.t1067 VSUBS 0.02fF
C4352 S.n3955 VSUBS 0.14fF $ **FLOATING
C4353 S.t858 VSUBS 0.02fF
C4354 S.n3957 VSUBS 0.24fF $ **FLOATING
C4355 S.n3958 VSUBS 0.36fF $ **FLOATING
C4356 S.n3959 VSUBS 0.61fF $ **FLOATING
C4357 S.n3960 VSUBS 0.92fF $ **FLOATING
C4358 S.n3961 VSUBS 0.32fF $ **FLOATING
C4359 S.n3962 VSUBS 0.92fF $ **FLOATING
C4360 S.n3963 VSUBS 1.09fF $ **FLOATING
C4361 S.n3964 VSUBS 0.15fF $ **FLOATING
C4362 S.n3965 VSUBS 4.96fF $ **FLOATING
C4363 S.t1936 VSUBS 0.02fF
C4364 S.n3966 VSUBS 0.12fF $ **FLOATING
C4365 S.n3967 VSUBS 0.14fF $ **FLOATING
C4366 S.t1695 VSUBS 0.02fF
C4367 S.n3969 VSUBS 0.24fF $ **FLOATING
C4368 S.n3970 VSUBS 0.91fF $ **FLOATING
C4369 S.n3971 VSUBS 0.05fF $ **FLOATING
C4370 S.n3972 VSUBS 1.88fF $ **FLOATING
C4371 S.n3973 VSUBS 2.67fF $ **FLOATING
C4372 S.t1640 VSUBS 0.02fF
C4373 S.n3974 VSUBS 0.24fF $ **FLOATING
C4374 S.n3975 VSUBS 0.36fF $ **FLOATING
C4375 S.n3976 VSUBS 0.61fF $ **FLOATING
C4376 S.n3977 VSUBS 0.12fF $ **FLOATING
C4377 S.t1851 VSUBS 0.02fF
C4378 S.n3978 VSUBS 0.14fF $ **FLOATING
C4379 S.n3980 VSUBS 1.88fF $ **FLOATING
C4380 S.n3981 VSUBS 2.67fF $ **FLOATING
C4381 S.t1664 VSUBS 0.02fF
C4382 S.n3982 VSUBS 0.24fF $ **FLOATING
C4383 S.n3983 VSUBS 0.36fF $ **FLOATING
C4384 S.n3984 VSUBS 0.61fF $ **FLOATING
C4385 S.t2510 VSUBS 0.02fF
C4386 S.n3985 VSUBS 0.24fF $ **FLOATING
C4387 S.n3986 VSUBS 0.91fF $ **FLOATING
C4388 S.n3987 VSUBS 0.05fF $ **FLOATING
C4389 S.t219 VSUBS 0.02fF
C4390 S.n3988 VSUBS 0.12fF $ **FLOATING
C4391 S.n3989 VSUBS 0.14fF $ **FLOATING
C4392 S.n3991 VSUBS 0.12fF $ **FLOATING
C4393 S.t1875 VSUBS 0.02fF
C4394 S.n3992 VSUBS 0.14fF $ **FLOATING
C4395 S.n3994 VSUBS 2.30fF $ **FLOATING
C4396 S.n3995 VSUBS 2.94fF $ **FLOATING
C4397 S.n3996 VSUBS 5.16fF $ **FLOATING
C4398 S.t193 VSUBS 0.02fF
C4399 S.n3997 VSUBS 0.12fF $ **FLOATING
C4400 S.n3998 VSUBS 0.14fF $ **FLOATING
C4401 S.t2486 VSUBS 0.02fF
C4402 S.n4000 VSUBS 0.24fF $ **FLOATING
C4403 S.n4001 VSUBS 0.91fF $ **FLOATING
C4404 S.n4002 VSUBS 0.05fF $ **FLOATING
C4405 S.n4003 VSUBS 1.88fF $ **FLOATING
C4406 S.n4004 VSUBS 2.67fF $ **FLOATING
C4407 S.t2424 VSUBS 0.02fF
C4408 S.n4005 VSUBS 0.24fF $ **FLOATING
C4409 S.n4006 VSUBS 0.36fF $ **FLOATING
C4410 S.n4007 VSUBS 0.61fF $ **FLOATING
C4411 S.n4008 VSUBS 0.12fF $ **FLOATING
C4412 S.t83 VSUBS 0.02fF
C4413 S.n4009 VSUBS 0.14fF $ **FLOATING
C4414 S.n4011 VSUBS 4.89fF $ **FLOATING
C4415 S.t981 VSUBS 0.02fF
C4416 S.n4012 VSUBS 0.12fF $ **FLOATING
C4417 S.n4013 VSUBS 0.14fF $ **FLOATING
C4418 S.t740 VSUBS 0.02fF
C4419 S.n4015 VSUBS 0.24fF $ **FLOATING
C4420 S.n4016 VSUBS 0.91fF $ **FLOATING
C4421 S.n4017 VSUBS 0.05fF $ **FLOATING
C4422 S.n4018 VSUBS 1.88fF $ **FLOATING
C4423 S.n4019 VSUBS 0.12fF $ **FLOATING
C4424 S.t925 VSUBS 0.02fF
C4425 S.n4020 VSUBS 0.14fF $ **FLOATING
C4426 S.t1438 VSUBS 0.02fF
C4427 S.n4022 VSUBS 1.22fF $ **FLOATING
C4428 S.n4023 VSUBS 0.36fF $ **FLOATING
C4429 S.n4024 VSUBS 1.22fF $ **FLOATING
C4430 S.n4025 VSUBS 0.61fF $ **FLOATING
C4431 S.n4026 VSUBS 0.35fF $ **FLOATING
C4432 S.n4027 VSUBS 0.63fF $ **FLOATING
C4433 S.n4028 VSUBS 1.15fF $ **FLOATING
C4434 S.n4029 VSUBS 3.00fF $ **FLOATING
C4435 S.n4030 VSUBS 0.59fF $ **FLOATING
C4436 S.n4031 VSUBS 0.01fF $ **FLOATING
C4437 S.n4032 VSUBS 0.97fF $ **FLOATING
C4438 S.t2 VSUBS 21.42fF
C4439 S.n4033 VSUBS 20.29fF $ **FLOATING
C4440 S.n4035 VSUBS 0.38fF $ **FLOATING
C4441 S.n4036 VSUBS 0.23fF $ **FLOATING
C4442 S.n4037 VSUBS 2.79fF $ **FLOATING
C4443 S.n4038 VSUBS 2.46fF $ **FLOATING
C4444 S.n4039 VSUBS 4.00fF $ **FLOATING
C4445 S.n4040 VSUBS 0.25fF $ **FLOATING
C4446 S.n4041 VSUBS 0.01fF $ **FLOATING
C4447 S.t624 VSUBS 0.02fF
C4448 S.n4042 VSUBS 0.26fF $ **FLOATING
C4449 S.t1726 VSUBS 0.02fF
C4450 S.n4043 VSUBS 0.95fF $ **FLOATING
C4451 S.n4044 VSUBS 0.71fF $ **FLOATING
C4452 S.n4045 VSUBS 1.89fF $ **FLOATING
C4453 S.n4046 VSUBS 1.88fF $ **FLOATING
C4454 S.t2230 VSUBS 0.02fF
C4455 S.n4047 VSUBS 0.24fF $ **FLOATING
C4456 S.n4048 VSUBS 0.36fF $ **FLOATING
C4457 S.n4049 VSUBS 0.61fF $ **FLOATING
C4458 S.n4050 VSUBS 0.12fF $ **FLOATING
C4459 S.t1413 VSUBS 0.02fF
C4460 S.n4051 VSUBS 0.14fF $ **FLOATING
C4461 S.n4053 VSUBS 1.16fF $ **FLOATING
C4462 S.n4054 VSUBS 0.22fF $ **FLOATING
C4463 S.n4055 VSUBS 0.25fF $ **FLOATING
C4464 S.n4056 VSUBS 0.09fF $ **FLOATING
C4465 S.n4057 VSUBS 1.88fF $ **FLOATING
C4466 S.t2513 VSUBS 0.02fF
C4467 S.n4058 VSUBS 0.24fF $ **FLOATING
C4468 S.n4059 VSUBS 0.91fF $ **FLOATING
C4469 S.n4060 VSUBS 0.05fF $ **FLOATING
C4470 S.t2277 VSUBS 0.02fF
C4471 S.n4061 VSUBS 0.12fF $ **FLOATING
C4472 S.n4062 VSUBS 0.14fF $ **FLOATING
C4473 S.n4064 VSUBS 0.78fF $ **FLOATING
C4474 S.n4065 VSUBS 1.94fF $ **FLOATING
C4475 S.n4066 VSUBS 1.88fF $ **FLOATING
C4476 S.n4067 VSUBS 0.12fF $ **FLOATING
C4477 S.t2323 VSUBS 0.02fF
C4478 S.n4068 VSUBS 0.14fF $ **FLOATING
C4479 S.t497 VSUBS 0.02fF
C4480 S.n4070 VSUBS 0.24fF $ **FLOATING
C4481 S.n4071 VSUBS 0.36fF $ **FLOATING
C4482 S.n4072 VSUBS 0.61fF $ **FLOATING
C4483 S.n4073 VSUBS 1.84fF $ **FLOATING
C4484 S.n4074 VSUBS 2.99fF $ **FLOATING
C4485 S.t774 VSUBS 0.02fF
C4486 S.n4075 VSUBS 0.24fF $ **FLOATING
C4487 S.n4076 VSUBS 0.91fF $ **FLOATING
C4488 S.n4077 VSUBS 0.05fF $ **FLOATING
C4489 S.t548 VSUBS 0.02fF
C4490 S.n4078 VSUBS 0.12fF $ **FLOATING
C4491 S.n4079 VSUBS 0.14fF $ **FLOATING
C4492 S.n4081 VSUBS 1.89fF $ **FLOATING
C4493 S.n4082 VSUBS 1.88fF $ **FLOATING
C4494 S.t1407 VSUBS 0.02fF
C4495 S.n4083 VSUBS 0.24fF $ **FLOATING
C4496 S.n4084 VSUBS 0.36fF $ **FLOATING
C4497 S.n4085 VSUBS 0.61fF $ **FLOATING
C4498 S.n4086 VSUBS 0.12fF $ **FLOATING
C4499 S.t586 VSUBS 0.02fF
C4500 S.n4087 VSUBS 0.14fF $ **FLOATING
C4501 S.n4089 VSUBS 1.16fF $ **FLOATING
C4502 S.n4090 VSUBS 0.22fF $ **FLOATING
C4503 S.n4091 VSUBS 0.25fF $ **FLOATING
C4504 S.n4092 VSUBS 0.09fF $ **FLOATING
C4505 S.n4093 VSUBS 1.88fF $ **FLOATING
C4506 S.t1684 VSUBS 0.02fF
C4507 S.n4094 VSUBS 0.24fF $ **FLOATING
C4508 S.n4095 VSUBS 0.91fF $ **FLOATING
C4509 S.n4096 VSUBS 0.05fF $ **FLOATING
C4510 S.t1454 VSUBS 0.02fF
C4511 S.n4097 VSUBS 0.12fF $ **FLOATING
C4512 S.n4098 VSUBS 0.14fF $ **FLOATING
C4513 S.n4100 VSUBS 0.78fF $ **FLOATING
C4514 S.n4101 VSUBS 1.94fF $ **FLOATING
C4515 S.n4102 VSUBS 1.88fF $ **FLOATING
C4516 S.n4103 VSUBS 0.12fF $ **FLOATING
C4517 S.t203 VSUBS 0.02fF
C4518 S.n4104 VSUBS 0.14fF $ **FLOATING
C4519 S.t1022 VSUBS 0.02fF
C4520 S.n4106 VSUBS 0.24fF $ **FLOATING
C4521 S.n4107 VSUBS 0.36fF $ **FLOATING
C4522 S.n4108 VSUBS 0.61fF $ **FLOATING
C4523 S.n4109 VSUBS 1.84fF $ **FLOATING
C4524 S.n4110 VSUBS 2.99fF $ **FLOATING
C4525 S.t1305 VSUBS 0.02fF
C4526 S.n4111 VSUBS 0.24fF $ **FLOATING
C4527 S.n4112 VSUBS 0.91fF $ **FLOATING
C4528 S.n4113 VSUBS 0.05fF $ **FLOATING
C4529 S.t1078 VSUBS 0.02fF
C4530 S.n4114 VSUBS 0.12fF $ **FLOATING
C4531 S.n4115 VSUBS 0.14fF $ **FLOATING
C4532 S.n4117 VSUBS 1.89fF $ **FLOATING
C4533 S.n4118 VSUBS 1.88fF $ **FLOATING
C4534 S.t1801 VSUBS 0.02fF
C4535 S.n4119 VSUBS 0.24fF $ **FLOATING
C4536 S.n4120 VSUBS 0.36fF $ **FLOATING
C4537 S.n4121 VSUBS 0.61fF $ **FLOATING
C4538 S.n4122 VSUBS 0.12fF $ **FLOATING
C4539 S.t992 VSUBS 0.02fF
C4540 S.n4123 VSUBS 0.14fF $ **FLOATING
C4541 S.n4125 VSUBS 1.16fF $ **FLOATING
C4542 S.n4126 VSUBS 0.22fF $ **FLOATING
C4543 S.n4127 VSUBS 0.25fF $ **FLOATING
C4544 S.n4128 VSUBS 0.09fF $ **FLOATING
C4545 S.n4129 VSUBS 1.88fF $ **FLOATING
C4546 S.t2092 VSUBS 0.02fF
C4547 S.n4130 VSUBS 0.24fF $ **FLOATING
C4548 S.n4131 VSUBS 0.91fF $ **FLOATING
C4549 S.n4132 VSUBS 0.05fF $ **FLOATING
C4550 S.t1859 VSUBS 0.02fF
C4551 S.n4133 VSUBS 0.12fF $ **FLOATING
C4552 S.n4134 VSUBS 0.14fF $ **FLOATING
C4553 S.n4136 VSUBS 0.78fF $ **FLOATING
C4554 S.n4137 VSUBS 1.94fF $ **FLOATING
C4555 S.n4138 VSUBS 1.88fF $ **FLOATING
C4556 S.n4139 VSUBS 0.12fF $ **FLOATING
C4557 S.t1774 VSUBS 0.02fF
C4558 S.n4140 VSUBS 0.14fF $ **FLOATING
C4559 S.t3 VSUBS 0.02fF
C4560 S.n4142 VSUBS 0.24fF $ **FLOATING
C4561 S.n4143 VSUBS 0.36fF $ **FLOATING
C4562 S.n4144 VSUBS 0.61fF $ **FLOATING
C4563 S.n4145 VSUBS 1.84fF $ **FLOATING
C4564 S.n4146 VSUBS 2.99fF $ **FLOATING
C4565 S.t364 VSUBS 0.02fF
C4566 S.n4147 VSUBS 0.24fF $ **FLOATING
C4567 S.n4148 VSUBS 0.91fF $ **FLOATING
C4568 S.n4149 VSUBS 0.05fF $ **FLOATING
C4569 S.t95 VSUBS 0.02fF
C4570 S.n4150 VSUBS 0.12fF $ **FLOATING
C4571 S.n4151 VSUBS 0.14fF $ **FLOATING
C4572 S.n4153 VSUBS 1.89fF $ **FLOATING
C4573 S.n4154 VSUBS 1.88fF $ **FLOATING
C4574 S.t849 VSUBS 0.02fF
C4575 S.n4155 VSUBS 0.24fF $ **FLOATING
C4576 S.n4156 VSUBS 0.36fF $ **FLOATING
C4577 S.n4157 VSUBS 0.61fF $ **FLOATING
C4578 S.n4158 VSUBS 0.12fF $ **FLOATING
C4579 S.t161 VSUBS 0.02fF
C4580 S.n4159 VSUBS 0.14fF $ **FLOATING
C4581 S.n4161 VSUBS 1.16fF $ **FLOATING
C4582 S.n4162 VSUBS 0.22fF $ **FLOATING
C4583 S.n4163 VSUBS 0.25fF $ **FLOATING
C4584 S.n4164 VSUBS 0.09fF $ **FLOATING
C4585 S.n4165 VSUBS 1.88fF $ **FLOATING
C4586 S.t1151 VSUBS 0.02fF
C4587 S.n4166 VSUBS 0.24fF $ **FLOATING
C4588 S.n4167 VSUBS 0.91fF $ **FLOATING
C4589 S.n4168 VSUBS 0.05fF $ **FLOATING
C4590 S.t908 VSUBS 0.02fF
C4591 S.n4169 VSUBS 0.12fF $ **FLOATING
C4592 S.n4170 VSUBS 0.14fF $ **FLOATING
C4593 S.n4172 VSUBS 0.78fF $ **FLOATING
C4594 S.n4173 VSUBS 1.94fF $ **FLOATING
C4595 S.n4174 VSUBS 1.88fF $ **FLOATING
C4596 S.n4175 VSUBS 0.12fF $ **FLOATING
C4597 S.t2293 VSUBS 0.02fF
C4598 S.n4176 VSUBS 0.14fF $ **FLOATING
C4599 S.t587 VSUBS 0.02fF
C4600 S.n4178 VSUBS 0.24fF $ **FLOATING
C4601 S.n4179 VSUBS 0.36fF $ **FLOATING
C4602 S.n4180 VSUBS 0.61fF $ **FLOATING
C4603 S.n4181 VSUBS 1.84fF $ **FLOATING
C4604 S.n4182 VSUBS 2.99fF $ **FLOATING
C4605 S.t872 VSUBS 0.02fF
C4606 S.n4183 VSUBS 0.24fF $ **FLOATING
C4607 S.n4184 VSUBS 0.91fF $ **FLOATING
C4608 S.n4185 VSUBS 0.05fF $ **FLOATING
C4609 S.t1821 VSUBS 0.02fF
C4610 S.n4186 VSUBS 0.12fF $ **FLOATING
C4611 S.n4187 VSUBS 0.14fF $ **FLOATING
C4612 S.n4189 VSUBS 1.89fF $ **FLOATING
C4613 S.n4190 VSUBS 1.75fF $ **FLOATING
C4614 S.t1379 VSUBS 0.02fF
C4615 S.n4191 VSUBS 0.24fF $ **FLOATING
C4616 S.n4192 VSUBS 0.36fF $ **FLOATING
C4617 S.n4193 VSUBS 0.61fF $ **FLOATING
C4618 S.n4194 VSUBS 0.12fF $ **FLOATING
C4619 S.t562 VSUBS 0.02fF
C4620 S.n4195 VSUBS 0.14fF $ **FLOATING
C4621 S.n4197 VSUBS 1.16fF $ **FLOATING
C4622 S.n4198 VSUBS 0.22fF $ **FLOATING
C4623 S.n4199 VSUBS 0.25fF $ **FLOATING
C4624 S.n4200 VSUBS 0.09fF $ **FLOATING
C4625 S.n4201 VSUBS 2.44fF $ **FLOATING
C4626 S.t1653 VSUBS 0.02fF
C4627 S.n4202 VSUBS 0.24fF $ **FLOATING
C4628 S.n4203 VSUBS 0.91fF $ **FLOATING
C4629 S.n4204 VSUBS 0.05fF $ **FLOATING
C4630 S.t1427 VSUBS 0.02fF
C4631 S.n4205 VSUBS 0.12fF $ **FLOATING
C4632 S.n4206 VSUBS 0.14fF $ **FLOATING
C4633 S.n4208 VSUBS 1.88fF $ **FLOATING
C4634 S.n4209 VSUBS 0.48fF $ **FLOATING
C4635 S.n4210 VSUBS 0.09fF $ **FLOATING
C4636 S.n4211 VSUBS 0.33fF $ **FLOATING
C4637 S.n4212 VSUBS 0.30fF $ **FLOATING
C4638 S.n4213 VSUBS 0.77fF $ **FLOATING
C4639 S.n4214 VSUBS 0.59fF $ **FLOATING
C4640 S.t2164 VSUBS 0.02fF
C4641 S.n4215 VSUBS 0.24fF $ **FLOATING
C4642 S.n4216 VSUBS 0.36fF $ **FLOATING
C4643 S.n4217 VSUBS 0.61fF $ **FLOATING
C4644 S.n4218 VSUBS 0.12fF $ **FLOATING
C4645 S.t1350 VSUBS 0.02fF
C4646 S.n4219 VSUBS 0.14fF $ **FLOATING
C4647 S.n4221 VSUBS 2.61fF $ **FLOATING
C4648 S.n4222 VSUBS 2.15fF $ **FLOATING
C4649 S.t2440 VSUBS 0.02fF
C4650 S.n4223 VSUBS 0.24fF $ **FLOATING
C4651 S.n4224 VSUBS 0.91fF $ **FLOATING
C4652 S.n4225 VSUBS 0.05fF $ **FLOATING
C4653 S.t2217 VSUBS 0.02fF
C4654 S.n4226 VSUBS 0.12fF $ **FLOATING
C4655 S.n4227 VSUBS 0.14fF $ **FLOATING
C4656 S.n4229 VSUBS 0.78fF $ **FLOATING
C4657 S.n4230 VSUBS 2.30fF $ **FLOATING
C4658 S.n4231 VSUBS 1.88fF $ **FLOATING
C4659 S.n4232 VSUBS 0.12fF $ **FLOATING
C4660 S.t2137 VSUBS 0.02fF
C4661 S.n4233 VSUBS 0.14fF $ **FLOATING
C4662 S.t433 VSUBS 0.02fF
C4663 S.n4235 VSUBS 0.24fF $ **FLOATING
C4664 S.n4236 VSUBS 0.36fF $ **FLOATING
C4665 S.n4237 VSUBS 0.61fF $ **FLOATING
C4666 S.n4238 VSUBS 1.39fF $ **FLOATING
C4667 S.n4239 VSUBS 0.71fF $ **FLOATING
C4668 S.n4240 VSUBS 1.14fF $ **FLOATING
C4669 S.n4241 VSUBS 0.35fF $ **FLOATING
C4670 S.n4242 VSUBS 2.02fF $ **FLOATING
C4671 S.t700 VSUBS 0.02fF
C4672 S.n4243 VSUBS 0.24fF $ **FLOATING
C4673 S.n4244 VSUBS 0.91fF $ **FLOATING
C4674 S.n4245 VSUBS 0.05fF $ **FLOATING
C4675 S.t483 VSUBS 0.02fF
C4676 S.n4246 VSUBS 0.12fF $ **FLOATING
C4677 S.n4247 VSUBS 0.14fF $ **FLOATING
C4678 S.n4249 VSUBS 1.89fF $ **FLOATING
C4679 S.n4250 VSUBS 1.88fF $ **FLOATING
C4680 S.t1228 VSUBS 0.02fF
C4681 S.n4251 VSUBS 0.24fF $ **FLOATING
C4682 S.n4252 VSUBS 0.36fF $ **FLOATING
C4683 S.n4253 VSUBS 0.61fF $ **FLOATING
C4684 S.n4254 VSUBS 0.12fF $ **FLOATING
C4685 S.t528 VSUBS 0.02fF
C4686 S.n4255 VSUBS 0.14fF $ **FLOATING
C4687 S.n4257 VSUBS 1.16fF $ **FLOATING
C4688 S.n4258 VSUBS 0.22fF $ **FLOATING
C4689 S.n4259 VSUBS 0.25fF $ **FLOATING
C4690 S.n4260 VSUBS 0.09fF $ **FLOATING
C4691 S.n4261 VSUBS 1.88fF $ **FLOATING
C4692 S.t1495 VSUBS 0.02fF
C4693 S.n4262 VSUBS 0.24fF $ **FLOATING
C4694 S.n4263 VSUBS 0.91fF $ **FLOATING
C4695 S.n4264 VSUBS 0.05fF $ **FLOATING
C4696 S.t1271 VSUBS 0.02fF
C4697 S.n4265 VSUBS 0.12fF $ **FLOATING
C4698 S.n4266 VSUBS 0.14fF $ **FLOATING
C4699 S.n4268 VSUBS 20.78fF $ **FLOATING
C4700 S.n4269 VSUBS 1.88fF $ **FLOATING
C4701 S.n4270 VSUBS 2.67fF $ **FLOATING
C4702 S.t2449 VSUBS 0.02fF
C4703 S.n4271 VSUBS 0.24fF $ **FLOATING
C4704 S.n4272 VSUBS 0.36fF $ **FLOATING
C4705 S.n4273 VSUBS 0.61fF $ **FLOATING
C4706 S.n4274 VSUBS 0.12fF $ **FLOATING
C4707 S.t123 VSUBS 0.02fF
C4708 S.n4275 VSUBS 0.14fF $ **FLOATING
C4709 S.n4277 VSUBS 2.80fF $ **FLOATING
C4710 S.n4278 VSUBS 2.30fF $ **FLOATING
C4711 S.t1010 VSUBS 0.02fF
C4712 S.n4279 VSUBS 0.12fF $ **FLOATING
C4713 S.n4280 VSUBS 0.14fF $ **FLOATING
C4714 S.t769 VSUBS 0.02fF
C4715 S.n4282 VSUBS 0.24fF $ **FLOATING
C4716 S.n4283 VSUBS 0.91fF $ **FLOATING
C4717 S.n4284 VSUBS 0.05fF $ **FLOATING
C4718 S.n4285 VSUBS 2.73fF $ **FLOATING
C4719 S.n4286 VSUBS 1.59fF $ **FLOATING
C4720 S.n4287 VSUBS 0.12fF $ **FLOATING
C4721 S.t741 VSUBS 0.02fF
C4722 S.n4288 VSUBS 0.14fF $ **FLOATING
C4723 S.t2408 VSUBS 0.02fF
C4724 S.n4290 VSUBS 0.24fF $ **FLOATING
C4725 S.n4291 VSUBS 0.36fF $ **FLOATING
C4726 S.n4292 VSUBS 0.61fF $ **FLOATING
C4727 S.n4293 VSUBS 0.07fF $ **FLOATING
C4728 S.n4294 VSUBS 0.01fF $ **FLOATING
C4729 S.n4295 VSUBS 0.24fF $ **FLOATING
C4730 S.n4296 VSUBS 1.16fF $ **FLOATING
C4731 S.n4297 VSUBS 1.35fF $ **FLOATING
C4732 S.n4298 VSUBS 2.30fF $ **FLOATING
C4733 S.t2572 VSUBS 0.02fF
C4734 S.n4299 VSUBS 0.12fF $ **FLOATING
C4735 S.n4300 VSUBS 0.14fF $ **FLOATING
C4736 S.t1296 VSUBS 0.02fF
C4737 S.n4302 VSUBS 0.24fF $ **FLOATING
C4738 S.n4303 VSUBS 0.91fF $ **FLOATING
C4739 S.n4304 VSUBS 0.05fF $ **FLOATING
C4740 S.t94 VSUBS 48.27fF
C4741 S.t1790 VSUBS 0.02fF
C4742 S.n4305 VSUBS 0.12fF $ **FLOATING
C4743 S.n4306 VSUBS 0.14fF $ **FLOATING
C4744 S.t1557 VSUBS 0.02fF
C4745 S.n4308 VSUBS 0.24fF $ **FLOATING
C4746 S.n4309 VSUBS 0.91fF $ **FLOATING
C4747 S.n4310 VSUBS 0.05fF $ **FLOATING
C4748 S.t710 VSUBS 0.02fF
C4749 S.n4311 VSUBS 0.24fF $ **FLOATING
C4750 S.n4312 VSUBS 0.36fF $ **FLOATING
C4751 S.n4313 VSUBS 0.61fF $ **FLOATING
C4752 S.n4314 VSUBS 2.67fF $ **FLOATING
C4753 S.n4315 VSUBS 5.17fF $ **FLOATING
C4754 S.n4316 VSUBS 1.88fF $ **FLOATING
C4755 S.n4317 VSUBS 0.12fF $ **FLOATING
C4756 S.t896 VSUBS 0.02fF
C4757 S.n4318 VSUBS 0.14fF $ **FLOATING
C4758 S.t690 VSUBS 0.02fF
C4759 S.n4320 VSUBS 0.24fF $ **FLOATING
C4760 S.n4321 VSUBS 0.36fF $ **FLOATING
C4761 S.n4322 VSUBS 0.61fF $ **FLOATING
C4762 S.n4323 VSUBS 2.67fF $ **FLOATING
C4763 S.n4324 VSUBS 5.44fF $ **FLOATING
C4764 S.t1765 VSUBS 0.02fF
C4765 S.n4325 VSUBS 0.12fF $ **FLOATING
C4766 S.n4326 VSUBS 0.14fF $ **FLOATING
C4767 S.t1532 VSUBS 0.02fF
C4768 S.n4328 VSUBS 0.24fF $ **FLOATING
C4769 S.n4329 VSUBS 0.91fF $ **FLOATING
C4770 S.n4330 VSUBS 0.05fF $ **FLOATING
C4771 S.t53 VSUBS 47.89fF
C4772 S.t2124 VSUBS 0.02fF
C4773 S.n4331 VSUBS 0.01fF $ **FLOATING
C4774 S.n4332 VSUBS 0.26fF $ **FLOATING
C4775 S.t2029 VSUBS 0.02fF
C4776 S.n4334 VSUBS 1.19fF $ **FLOATING
C4777 S.n4335 VSUBS 0.05fF $ **FLOATING
C4778 S.t1735 VSUBS 0.02fF
C4779 S.n4336 VSUBS 0.64fF $ **FLOATING
C4780 S.n4337 VSUBS 0.61fF $ **FLOATING
C4781 S.n4338 VSUBS 8.97fF $ **FLOATING
C4782 S.n4339 VSUBS 8.97fF $ **FLOATING
C4783 S.n4340 VSUBS 0.60fF $ **FLOATING
C4784 S.n4341 VSUBS 0.22fF $ **FLOATING
C4785 S.n4342 VSUBS 0.59fF $ **FLOATING
C4786 S.n4343 VSUBS 3.39fF $ **FLOATING
C4787 S.n4344 VSUBS 0.29fF $ **FLOATING
C4788 S.t19 VSUBS 21.42fF
C4789 S.n4345 VSUBS 21.71fF $ **FLOATING
C4790 S.n4346 VSUBS 0.77fF $ **FLOATING
C4791 S.n4347 VSUBS 0.28fF $ **FLOATING
C4792 S.n4348 VSUBS 4.00fF $ **FLOATING
C4793 S.n4349 VSUBS 1.35fF $ **FLOATING
C4794 S.n4350 VSUBS 0.01fF $ **FLOATING
C4795 S.n4351 VSUBS 0.02fF $ **FLOATING
C4796 S.n4352 VSUBS 0.03fF $ **FLOATING
C4797 S.n4353 VSUBS 0.04fF $ **FLOATING
C4798 S.n4354 VSUBS 0.17fF $ **FLOATING
C4799 S.n4355 VSUBS 0.01fF $ **FLOATING
C4800 S.n4356 VSUBS 0.02fF $ **FLOATING
C4801 S.n4357 VSUBS 0.01fF $ **FLOATING
C4802 S.n4358 VSUBS 0.01fF $ **FLOATING
C4803 S.n4359 VSUBS 0.01fF $ **FLOATING
C4804 S.n4360 VSUBS 0.01fF $ **FLOATING
C4805 S.n4361 VSUBS 0.02fF $ **FLOATING
C4806 S.n4362 VSUBS 0.01fF $ **FLOATING
C4807 S.n4363 VSUBS 0.02fF $ **FLOATING
C4808 S.n4364 VSUBS 0.05fF $ **FLOATING
C4809 S.n4365 VSUBS 0.04fF $ **FLOATING
C4810 S.n4366 VSUBS 0.11fF $ **FLOATING
C4811 S.n4367 VSUBS 0.38fF $ **FLOATING
C4812 S.n4368 VSUBS 0.20fF $ **FLOATING
C4813 S.n4369 VSUBS 4.39fF $ **FLOATING
C4814 S.n4370 VSUBS 0.24fF $ **FLOATING
C4815 S.n4371 VSUBS 1.50fF $ **FLOATING
C4816 S.n4372 VSUBS 1.31fF $ **FLOATING
C4817 S.n4373 VSUBS 0.28fF $ **FLOATING
C4818 S.n4374 VSUBS 0.25fF $ **FLOATING
C4819 S.n4375 VSUBS 0.09fF $ **FLOATING
C4820 S.n4376 VSUBS 0.21fF $ **FLOATING
C4821 S.n4377 VSUBS 0.92fF $ **FLOATING
C4822 S.n4378 VSUBS 0.44fF $ **FLOATING
C4823 S.n4379 VSUBS 1.88fF $ **FLOATING
C4824 S.n4380 VSUBS 0.12fF $ **FLOATING
C4825 S.t272 VSUBS 0.02fF
C4826 S.n4381 VSUBS 0.14fF $ **FLOATING
C4827 S.t1083 VSUBS 0.02fF
C4828 S.n4383 VSUBS 0.24fF $ **FLOATING
C4829 S.n4384 VSUBS 0.36fF $ **FLOATING
C4830 S.n4385 VSUBS 0.61fF $ **FLOATING
C4831 S.n4386 VSUBS 0.02fF $ **FLOATING
C4832 S.n4387 VSUBS 0.01fF $ **FLOATING
C4833 S.n4388 VSUBS 0.02fF $ **FLOATING
C4834 S.n4389 VSUBS 0.08fF $ **FLOATING
C4835 S.n4390 VSUBS 0.06fF $ **FLOATING
C4836 S.n4391 VSUBS 0.03fF $ **FLOATING
C4837 S.n4392 VSUBS 0.04fF $ **FLOATING
C4838 S.n4393 VSUBS 1.00fF $ **FLOATING
C4839 S.n4394 VSUBS 0.36fF $ **FLOATING
C4840 S.n4395 VSUBS 1.87fF $ **FLOATING
C4841 S.n4396 VSUBS 1.99fF $ **FLOATING
C4842 S.t1364 VSUBS 0.02fF
C4843 S.n4397 VSUBS 0.24fF $ **FLOATING
C4844 S.n4398 VSUBS 0.91fF $ **FLOATING
C4845 S.n4399 VSUBS 0.05fF $ **FLOATING
C4846 S.t1141 VSUBS 0.02fF
C4847 S.n4400 VSUBS 0.12fF $ **FLOATING
C4848 S.n4401 VSUBS 0.14fF $ **FLOATING
C4849 S.n4403 VSUBS 1.89fF $ **FLOATING
C4850 S.n4404 VSUBS 0.06fF $ **FLOATING
C4851 S.n4405 VSUBS 0.03fF $ **FLOATING
C4852 S.n4406 VSUBS 0.04fF $ **FLOATING
C4853 S.n4407 VSUBS 0.99fF $ **FLOATING
C4854 S.n4408 VSUBS 0.02fF $ **FLOATING
C4855 S.n4409 VSUBS 0.01fF $ **FLOATING
C4856 S.n4410 VSUBS 0.02fF $ **FLOATING
C4857 S.n4411 VSUBS 0.08fF $ **FLOATING
C4858 S.n4412 VSUBS 0.36fF $ **FLOATING
C4859 S.n4413 VSUBS 1.85fF $ **FLOATING
C4860 S.t1995 VSUBS 0.02fF
C4861 S.n4414 VSUBS 0.24fF $ **FLOATING
C4862 S.n4415 VSUBS 0.36fF $ **FLOATING
C4863 S.n4416 VSUBS 0.61fF $ **FLOATING
C4864 S.n4417 VSUBS 0.12fF $ **FLOATING
C4865 S.t1187 VSUBS 0.02fF
C4866 S.n4418 VSUBS 0.14fF $ **FLOATING
C4867 S.n4420 VSUBS 0.70fF $ **FLOATING
C4868 S.n4421 VSUBS 0.23fF $ **FLOATING
C4869 S.n4422 VSUBS 0.23fF $ **FLOATING
C4870 S.n4423 VSUBS 0.70fF $ **FLOATING
C4871 S.n4424 VSUBS 1.16fF $ **FLOATING
C4872 S.n4425 VSUBS 0.22fF $ **FLOATING
C4873 S.n4426 VSUBS 0.25fF $ **FLOATING
C4874 S.n4427 VSUBS 0.09fF $ **FLOATING
C4875 S.n4428 VSUBS 1.88fF $ **FLOATING
C4876 S.t2270 VSUBS 0.02fF
C4877 S.n4429 VSUBS 0.24fF $ **FLOATING
C4878 S.n4430 VSUBS 0.91fF $ **FLOATING
C4879 S.n4431 VSUBS 0.05fF $ **FLOATING
C4880 S.t2051 VSUBS 0.02fF
C4881 S.n4432 VSUBS 0.12fF $ **FLOATING
C4882 S.n4433 VSUBS 0.14fF $ **FLOATING
C4883 S.n4435 VSUBS 0.25fF $ **FLOATING
C4884 S.n4436 VSUBS 0.09fF $ **FLOATING
C4885 S.n4437 VSUBS 0.21fF $ **FLOATING
C4886 S.n4438 VSUBS 0.92fF $ **FLOATING
C4887 S.n4439 VSUBS 0.44fF $ **FLOATING
C4888 S.n4440 VSUBS 1.88fF $ **FLOATING
C4889 S.n4441 VSUBS 0.12fF $ **FLOATING
C4890 S.t776 VSUBS 0.02fF
C4891 S.n4442 VSUBS 0.14fF $ **FLOATING
C4892 S.t1588 VSUBS 0.02fF
C4893 S.n4444 VSUBS 0.24fF $ **FLOATING
C4894 S.n4445 VSUBS 0.36fF $ **FLOATING
C4895 S.n4446 VSUBS 0.61fF $ **FLOATING
C4896 S.n4447 VSUBS 0.02fF $ **FLOATING
C4897 S.n4448 VSUBS 0.01fF $ **FLOATING
C4898 S.n4449 VSUBS 0.02fF $ **FLOATING
C4899 S.n4450 VSUBS 0.08fF $ **FLOATING
C4900 S.n4451 VSUBS 0.06fF $ **FLOATING
C4901 S.n4452 VSUBS 0.03fF $ **FLOATING
C4902 S.n4453 VSUBS 0.04fF $ **FLOATING
C4903 S.n4454 VSUBS 1.00fF $ **FLOATING
C4904 S.n4455 VSUBS 0.36fF $ **FLOATING
C4905 S.n4456 VSUBS 1.87fF $ **FLOATING
C4906 S.n4457 VSUBS 1.99fF $ **FLOATING
C4907 S.t1890 VSUBS 0.02fF
C4908 S.n4458 VSUBS 0.24fF $ **FLOATING
C4909 S.n4459 VSUBS 0.91fF $ **FLOATING
C4910 S.n4460 VSUBS 0.05fF $ **FLOATING
C4911 S.t315 VSUBS 0.02fF
C4912 S.n4461 VSUBS 0.12fF $ **FLOATING
C4913 S.n4462 VSUBS 0.14fF $ **FLOATING
C4914 S.n4464 VSUBS 1.89fF $ **FLOATING
C4915 S.n4465 VSUBS 0.06fF $ **FLOATING
C4916 S.n4466 VSUBS 0.03fF $ **FLOATING
C4917 S.n4467 VSUBS 0.04fF $ **FLOATING
C4918 S.n4468 VSUBS 0.99fF $ **FLOATING
C4919 S.n4469 VSUBS 0.02fF $ **FLOATING
C4920 S.n4470 VSUBS 0.01fF $ **FLOATING
C4921 S.n4471 VSUBS 0.02fF $ **FLOATING
C4922 S.n4472 VSUBS 0.08fF $ **FLOATING
C4923 S.n4473 VSUBS 0.36fF $ **FLOATING
C4924 S.n4474 VSUBS 1.85fF $ **FLOATING
C4925 S.t2379 VSUBS 0.02fF
C4926 S.n4475 VSUBS 0.24fF $ **FLOATING
C4927 S.n4476 VSUBS 0.36fF $ **FLOATING
C4928 S.n4477 VSUBS 0.61fF $ **FLOATING
C4929 S.n4478 VSUBS 0.12fF $ **FLOATING
C4930 S.t1560 VSUBS 0.02fF
C4931 S.n4479 VSUBS 0.14fF $ **FLOATING
C4932 S.n4481 VSUBS 0.70fF $ **FLOATING
C4933 S.n4482 VSUBS 0.23fF $ **FLOATING
C4934 S.n4483 VSUBS 0.23fF $ **FLOATING
C4935 S.n4484 VSUBS 0.70fF $ **FLOATING
C4936 S.n4485 VSUBS 1.16fF $ **FLOATING
C4937 S.n4486 VSUBS 0.22fF $ **FLOATING
C4938 S.n4487 VSUBS 0.25fF $ **FLOATING
C4939 S.n4488 VSUBS 0.09fF $ **FLOATING
C4940 S.n4489 VSUBS 1.88fF $ **FLOATING
C4941 S.t139 VSUBS 0.02fF
C4942 S.n4490 VSUBS 0.24fF $ **FLOATING
C4943 S.n4491 VSUBS 0.91fF $ **FLOATING
C4944 S.n4492 VSUBS 0.05fF $ **FLOATING
C4945 S.t2430 VSUBS 0.02fF
C4946 S.n4493 VSUBS 0.12fF $ **FLOATING
C4947 S.n4494 VSUBS 0.14fF $ **FLOATING
C4948 S.n4496 VSUBS 0.25fF $ **FLOATING
C4949 S.n4497 VSUBS 0.09fF $ **FLOATING
C4950 S.n4498 VSUBS 0.21fF $ **FLOATING
C4951 S.n4499 VSUBS 0.92fF $ **FLOATING
C4952 S.n4500 VSUBS 0.44fF $ **FLOATING
C4953 S.n4501 VSUBS 1.88fF $ **FLOATING
C4954 S.n4502 VSUBS 0.12fF $ **FLOATING
C4955 S.t2351 VSUBS 0.02fF
C4956 S.n4503 VSUBS 0.14fF $ **FLOATING
C4957 S.t644 VSUBS 0.02fF
C4958 S.n4505 VSUBS 0.24fF $ **FLOATING
C4959 S.n4506 VSUBS 0.36fF $ **FLOATING
C4960 S.n4507 VSUBS 0.61fF $ **FLOATING
C4961 S.n4508 VSUBS 0.02fF $ **FLOATING
C4962 S.n4509 VSUBS 0.01fF $ **FLOATING
C4963 S.n4510 VSUBS 0.02fF $ **FLOATING
C4964 S.n4511 VSUBS 0.08fF $ **FLOATING
C4965 S.n4512 VSUBS 0.06fF $ **FLOATING
C4966 S.n4513 VSUBS 0.03fF $ **FLOATING
C4967 S.n4514 VSUBS 0.04fF $ **FLOATING
C4968 S.n4515 VSUBS 1.00fF $ **FLOATING
C4969 S.n4516 VSUBS 0.36fF $ **FLOATING
C4970 S.n4517 VSUBS 1.87fF $ **FLOATING
C4971 S.n4518 VSUBS 1.99fF $ **FLOATING
C4972 S.t935 VSUBS 0.02fF
C4973 S.n4519 VSUBS 0.24fF $ **FLOATING
C4974 S.n4520 VSUBS 0.91fF $ **FLOATING
C4975 S.n4521 VSUBS 0.05fF $ **FLOATING
C4976 S.t694 VSUBS 0.02fF
C4977 S.n4522 VSUBS 0.12fF $ **FLOATING
C4978 S.n4523 VSUBS 0.14fF $ **FLOATING
C4979 S.n4525 VSUBS 1.89fF $ **FLOATING
C4980 S.n4526 VSUBS 0.06fF $ **FLOATING
C4981 S.n4527 VSUBS 0.03fF $ **FLOATING
C4982 S.n4528 VSUBS 0.04fF $ **FLOATING
C4983 S.n4529 VSUBS 0.99fF $ **FLOATING
C4984 S.n4530 VSUBS 0.02fF $ **FLOATING
C4985 S.n4531 VSUBS 0.01fF $ **FLOATING
C4986 S.n4532 VSUBS 0.02fF $ **FLOATING
C4987 S.n4533 VSUBS 0.08fF $ **FLOATING
C4988 S.n4534 VSUBS 0.36fF $ **FLOATING
C4989 S.n4535 VSUBS 1.85fF $ **FLOATING
C4990 S.t1430 VSUBS 0.02fF
C4991 S.n4536 VSUBS 0.24fF $ **FLOATING
C4992 S.n4537 VSUBS 0.36fF $ **FLOATING
C4993 S.n4538 VSUBS 0.61fF $ **FLOATING
C4994 S.n4539 VSUBS 0.12fF $ **FLOATING
C4995 S.t618 VSUBS 0.02fF
C4996 S.n4540 VSUBS 0.14fF $ **FLOATING
C4997 S.n4542 VSUBS 0.70fF $ **FLOATING
C4998 S.n4543 VSUBS 0.23fF $ **FLOATING
C4999 S.n4544 VSUBS 0.23fF $ **FLOATING
C5000 S.n4545 VSUBS 0.70fF $ **FLOATING
C5001 S.n4546 VSUBS 1.16fF $ **FLOATING
C5002 S.n4547 VSUBS 0.22fF $ **FLOATING
C5003 S.n4548 VSUBS 0.25fF $ **FLOATING
C5004 S.n4549 VSUBS 0.09fF $ **FLOATING
C5005 S.n4550 VSUBS 1.88fF $ **FLOATING
C5006 S.t1717 VSUBS 0.02fF
C5007 S.n4551 VSUBS 0.24fF $ **FLOATING
C5008 S.n4552 VSUBS 0.91fF $ **FLOATING
C5009 S.n4553 VSUBS 0.05fF $ **FLOATING
C5010 S.t1486 VSUBS 0.02fF
C5011 S.n4554 VSUBS 0.12fF $ **FLOATING
C5012 S.n4555 VSUBS 0.14fF $ **FLOATING
C5013 S.n4557 VSUBS 0.25fF $ **FLOATING
C5014 S.n4558 VSUBS 0.09fF $ **FLOATING
C5015 S.n4559 VSUBS 0.21fF $ **FLOATING
C5016 S.n4560 VSUBS 0.92fF $ **FLOATING
C5017 S.n4561 VSUBS 0.44fF $ **FLOATING
C5018 S.n4562 VSUBS 1.88fF $ **FLOATING
C5019 S.n4563 VSUBS 0.12fF $ **FLOATING
C5020 S.t1527 VSUBS 0.02fF
C5021 S.n4564 VSUBS 0.14fF $ **FLOATING
C5022 S.t2344 VSUBS 0.02fF
C5023 S.n4566 VSUBS 0.24fF $ **FLOATING
C5024 S.n4567 VSUBS 0.36fF $ **FLOATING
C5025 S.n4568 VSUBS 0.61fF $ **FLOATING
C5026 S.n4569 VSUBS 0.02fF $ **FLOATING
C5027 S.n4570 VSUBS 0.01fF $ **FLOATING
C5028 S.n4571 VSUBS 0.02fF $ **FLOATING
C5029 S.n4572 VSUBS 0.08fF $ **FLOATING
C5030 S.n4573 VSUBS 0.06fF $ **FLOATING
C5031 S.n4574 VSUBS 0.03fF $ **FLOATING
C5032 S.n4575 VSUBS 0.04fF $ **FLOATING
C5033 S.n4576 VSUBS 1.00fF $ **FLOATING
C5034 S.n4577 VSUBS 0.36fF $ **FLOATING
C5035 S.n4578 VSUBS 1.87fF $ **FLOATING
C5036 S.n4579 VSUBS 1.99fF $ **FLOATING
C5037 S.t89 VSUBS 0.02fF
C5038 S.n4580 VSUBS 0.24fF $ **FLOATING
C5039 S.n4581 VSUBS 0.91fF $ **FLOATING
C5040 S.n4582 VSUBS 0.05fF $ **FLOATING
C5041 S.t2394 VSUBS 0.02fF
C5042 S.n4583 VSUBS 0.12fF $ **FLOATING
C5043 S.n4584 VSUBS 0.14fF $ **FLOATING
C5044 S.n4586 VSUBS 1.89fF $ **FLOATING
C5045 S.n4587 VSUBS 0.04fF $ **FLOATING
C5046 S.n4588 VSUBS 0.07fF $ **FLOATING
C5047 S.n4589 VSUBS 0.05fF $ **FLOATING
C5048 S.n4590 VSUBS 0.87fF $ **FLOATING
C5049 S.n4591 VSUBS 0.01fF $ **FLOATING
C5050 S.n4592 VSUBS 0.01fF $ **FLOATING
C5051 S.n4593 VSUBS 0.01fF $ **FLOATING
C5052 S.n4594 VSUBS 0.07fF $ **FLOATING
C5053 S.n4595 VSUBS 0.68fF $ **FLOATING
C5054 S.n4596 VSUBS 0.72fF $ **FLOATING
C5055 S.t1969 VSUBS 0.02fF
C5056 S.n4597 VSUBS 0.24fF $ **FLOATING
C5057 S.n4598 VSUBS 0.36fF $ **FLOATING
C5058 S.n4599 VSUBS 0.61fF $ **FLOATING
C5059 S.n4600 VSUBS 0.12fF $ **FLOATING
C5060 S.t1156 VSUBS 0.02fF
C5061 S.n4601 VSUBS 0.14fF $ **FLOATING
C5062 S.n4603 VSUBS 0.70fF $ **FLOATING
C5063 S.n4604 VSUBS 0.23fF $ **FLOATING
C5064 S.n4605 VSUBS 0.23fF $ **FLOATING
C5065 S.n4606 VSUBS 0.70fF $ **FLOATING
C5066 S.n4607 VSUBS 1.16fF $ **FLOATING
C5067 S.n4608 VSUBS 0.22fF $ **FLOATING
C5068 S.n4609 VSUBS 0.25fF $ **FLOATING
C5069 S.n4610 VSUBS 0.09fF $ **FLOATING
C5070 S.n4611 VSUBS 2.31fF $ **FLOATING
C5071 S.t2242 VSUBS 0.02fF
C5072 S.n4612 VSUBS 0.24fF $ **FLOATING
C5073 S.n4613 VSUBS 0.91fF $ **FLOATING
C5074 S.n4614 VSUBS 0.05fF $ **FLOATING
C5075 S.t2015 VSUBS 0.02fF
C5076 S.n4615 VSUBS 0.12fF $ **FLOATING
C5077 S.n4616 VSUBS 0.14fF $ **FLOATING
C5078 S.n4618 VSUBS 1.88fF $ **FLOATING
C5079 S.n4619 VSUBS 0.46fF $ **FLOATING
C5080 S.n4620 VSUBS 0.22fF $ **FLOATING
C5081 S.n4621 VSUBS 0.38fF $ **FLOATING
C5082 S.n4622 VSUBS 0.16fF $ **FLOATING
C5083 S.n4623 VSUBS 0.28fF $ **FLOATING
C5084 S.n4624 VSUBS 0.21fF $ **FLOATING
C5085 S.n4625 VSUBS 0.30fF $ **FLOATING
C5086 S.n4626 VSUBS 0.42fF $ **FLOATING
C5087 S.n4627 VSUBS 0.21fF $ **FLOATING
C5088 S.t231 VSUBS 0.02fF
C5089 S.n4628 VSUBS 0.24fF $ **FLOATING
C5090 S.n4629 VSUBS 0.36fF $ **FLOATING
C5091 S.n4630 VSUBS 0.61fF $ **FLOATING
C5092 S.n4631 VSUBS 0.12fF $ **FLOATING
C5093 S.t1940 VSUBS 0.02fF
C5094 S.n4632 VSUBS 0.14fF $ **FLOATING
C5095 S.n4634 VSUBS 0.04fF $ **FLOATING
C5096 S.n4635 VSUBS 0.03fF $ **FLOATING
C5097 S.n4636 VSUBS 0.03fF $ **FLOATING
C5098 S.n4637 VSUBS 0.10fF $ **FLOATING
C5099 S.n4638 VSUBS 0.36fF $ **FLOATING
C5100 S.n4639 VSUBS 0.38fF $ **FLOATING
C5101 S.n4640 VSUBS 0.11fF $ **FLOATING
C5102 S.n4641 VSUBS 0.12fF $ **FLOATING
C5103 S.n4642 VSUBS 0.07fF $ **FLOATING
C5104 S.n4643 VSUBS 0.12fF $ **FLOATING
C5105 S.n4644 VSUBS 0.18fF $ **FLOATING
C5106 S.n4645 VSUBS 3.99fF $ **FLOATING
C5107 S.t512 VSUBS 0.02fF
C5108 S.n4646 VSUBS 0.24fF $ **FLOATING
C5109 S.n4647 VSUBS 0.91fF $ **FLOATING
C5110 S.n4648 VSUBS 0.05fF $ **FLOATING
C5111 S.t288 VSUBS 0.02fF
C5112 S.n4649 VSUBS 0.12fF $ **FLOATING
C5113 S.n4650 VSUBS 0.14fF $ **FLOATING
C5114 S.n4652 VSUBS 0.25fF $ **FLOATING
C5115 S.n4653 VSUBS 0.09fF $ **FLOATING
C5116 S.n4654 VSUBS 0.21fF $ **FLOATING
C5117 S.n4655 VSUBS 1.28fF $ **FLOATING
C5118 S.n4656 VSUBS 0.53fF $ **FLOATING
C5119 S.n4657 VSUBS 1.88fF $ **FLOATING
C5120 S.n4658 VSUBS 0.12fF $ **FLOATING
C5121 S.t198 VSUBS 0.02fF
C5122 S.n4659 VSUBS 0.14fF $ **FLOATING
C5123 S.t1017 VSUBS 0.02fF
C5124 S.n4661 VSUBS 0.24fF $ **FLOATING
C5125 S.n4662 VSUBS 0.36fF $ **FLOATING
C5126 S.n4663 VSUBS 0.61fF $ **FLOATING
C5127 S.n4664 VSUBS 1.58fF $ **FLOATING
C5128 S.n4665 VSUBS 2.45fF $ **FLOATING
C5129 S.t1298 VSUBS 0.02fF
C5130 S.n4666 VSUBS 0.24fF $ **FLOATING
C5131 S.n4667 VSUBS 0.91fF $ **FLOATING
C5132 S.n4668 VSUBS 0.05fF $ **FLOATING
C5133 S.t1071 VSUBS 0.02fF
C5134 S.n4669 VSUBS 0.12fF $ **FLOATING
C5135 S.n4670 VSUBS 0.14fF $ **FLOATING
C5136 S.n4672 VSUBS 1.89fF $ **FLOATING
C5137 S.n4673 VSUBS 0.06fF $ **FLOATING
C5138 S.n4674 VSUBS 0.03fF $ **FLOATING
C5139 S.n4675 VSUBS 0.04fF $ **FLOATING
C5140 S.n4676 VSUBS 0.99fF $ **FLOATING
C5141 S.n4677 VSUBS 0.02fF $ **FLOATING
C5142 S.n4678 VSUBS 0.01fF $ **FLOATING
C5143 S.n4679 VSUBS 0.02fF $ **FLOATING
C5144 S.n4680 VSUBS 0.08fF $ **FLOATING
C5145 S.n4681 VSUBS 0.36fF $ **FLOATING
C5146 S.n4682 VSUBS 1.85fF $ **FLOATING
C5147 S.t1795 VSUBS 0.02fF
C5148 S.n4683 VSUBS 0.24fF $ **FLOATING
C5149 S.n4684 VSUBS 0.36fF $ **FLOATING
C5150 S.n4685 VSUBS 0.61fF $ **FLOATING
C5151 S.n4686 VSUBS 0.12fF $ **FLOATING
C5152 S.t985 VSUBS 0.02fF
C5153 S.n4687 VSUBS 0.14fF $ **FLOATING
C5154 S.n4689 VSUBS 0.70fF $ **FLOATING
C5155 S.n4690 VSUBS 0.23fF $ **FLOATING
C5156 S.n4691 VSUBS 0.23fF $ **FLOATING
C5157 S.n4692 VSUBS 0.70fF $ **FLOATING
C5158 S.n4693 VSUBS 1.16fF $ **FLOATING
C5159 S.n4694 VSUBS 0.22fF $ **FLOATING
C5160 S.n4695 VSUBS 0.25fF $ **FLOATING
C5161 S.n4696 VSUBS 0.09fF $ **FLOATING
C5162 S.n4697 VSUBS 1.88fF $ **FLOATING
C5163 S.t2086 VSUBS 0.02fF
C5164 S.n4698 VSUBS 0.24fF $ **FLOATING
C5165 S.n4699 VSUBS 0.91fF $ **FLOATING
C5166 S.n4700 VSUBS 0.05fF $ **FLOATING
C5167 S.t1856 VSUBS 0.02fF
C5168 S.n4701 VSUBS 0.12fF $ **FLOATING
C5169 S.n4702 VSUBS 0.14fF $ **FLOATING
C5170 S.n4704 VSUBS 20.78fF $ **FLOATING
C5171 S.n4705 VSUBS 1.72fF $ **FLOATING
C5172 S.n4706 VSUBS 3.05fF $ **FLOATING
C5173 S.t298 VSUBS 0.02fF
C5174 S.n4707 VSUBS 0.24fF $ **FLOATING
C5175 S.n4708 VSUBS 0.36fF $ **FLOATING
C5176 S.n4709 VSUBS 0.61fF $ **FLOATING
C5177 S.n4710 VSUBS 0.12fF $ **FLOATING
C5178 S.t2002 VSUBS 0.02fF
C5179 S.n4711 VSUBS 0.14fF $ **FLOATING
C5180 S.n4713 VSUBS 0.31fF $ **FLOATING
C5181 S.n4714 VSUBS 0.23fF $ **FLOATING
C5182 S.n4715 VSUBS 0.66fF $ **FLOATING
C5183 S.n4716 VSUBS 0.95fF $ **FLOATING
C5184 S.n4717 VSUBS 0.23fF $ **FLOATING
C5185 S.n4718 VSUBS 0.21fF $ **FLOATING
C5186 S.n4719 VSUBS 0.20fF $ **FLOATING
C5187 S.n4720 VSUBS 0.06fF $ **FLOATING
C5188 S.n4721 VSUBS 0.09fF $ **FLOATING
C5189 S.n4722 VSUBS 0.10fF $ **FLOATING
C5190 S.n4723 VSUBS 1.99fF $ **FLOATING
C5191 S.t355 VSUBS 0.02fF
C5192 S.n4724 VSUBS 0.12fF $ **FLOATING
C5193 S.n4725 VSUBS 0.14fF $ **FLOATING
C5194 S.t575 VSUBS 0.02fF
C5195 S.n4727 VSUBS 0.24fF $ **FLOATING
C5196 S.n4728 VSUBS 0.91fF $ **FLOATING
C5197 S.n4729 VSUBS 0.05fF $ **FLOATING
C5198 S.n4730 VSUBS 1.88fF $ **FLOATING
C5199 S.n4731 VSUBS 0.12fF $ **FLOATING
C5200 S.t2467 VSUBS 0.02fF
C5201 S.n4732 VSUBS 0.14fF $ **FLOATING
C5202 S.t688 VSUBS 0.02fF
C5203 S.n4734 VSUBS 0.12fF $ **FLOATING
C5204 S.n4735 VSUBS 0.14fF $ **FLOATING
C5205 S.t931 VSUBS 0.02fF
C5206 S.n4737 VSUBS 0.24fF $ **FLOATING
C5207 S.n4738 VSUBS 0.91fF $ **FLOATING
C5208 S.n4739 VSUBS 0.05fF $ **FLOATING
C5209 S.t639 VSUBS 0.02fF
C5210 S.n4740 VSUBS 0.24fF $ **FLOATING
C5211 S.n4741 VSUBS 0.36fF $ **FLOATING
C5212 S.n4742 VSUBS 0.61fF $ **FLOATING
C5213 S.n4743 VSUBS 0.32fF $ **FLOATING
C5214 S.n4744 VSUBS 1.09fF $ **FLOATING
C5215 S.n4745 VSUBS 0.15fF $ **FLOATING
C5216 S.n4746 VSUBS 2.10fF $ **FLOATING
C5217 S.n4747 VSUBS 2.94fF $ **FLOATING
C5218 S.n4748 VSUBS 1.88fF $ **FLOATING
C5219 S.n4749 VSUBS 0.12fF $ **FLOATING
C5220 S.t1122 VSUBS 0.02fF
C5221 S.n4750 VSUBS 0.14fF $ **FLOATING
C5222 S.t911 VSUBS 0.02fF
C5223 S.n4752 VSUBS 0.24fF $ **FLOATING
C5224 S.n4753 VSUBS 0.36fF $ **FLOATING
C5225 S.n4754 VSUBS 0.61fF $ **FLOATING
C5226 S.n4755 VSUBS 0.92fF $ **FLOATING
C5227 S.n4756 VSUBS 0.32fF $ **FLOATING
C5228 S.n4757 VSUBS 0.92fF $ **FLOATING
C5229 S.n4758 VSUBS 1.09fF $ **FLOATING
C5230 S.n4759 VSUBS 0.15fF $ **FLOATING
C5231 S.n4760 VSUBS 4.96fF $ **FLOATING
C5232 S.t246 VSUBS 0.02fF
C5233 S.n4761 VSUBS 0.12fF $ **FLOATING
C5234 S.n4762 VSUBS 0.14fF $ **FLOATING
C5235 S.t1749 VSUBS 0.02fF
C5236 S.n4764 VSUBS 0.24fF $ **FLOATING
C5237 S.n4765 VSUBS 0.91fF $ **FLOATING
C5238 S.n4766 VSUBS 0.05fF $ **FLOATING
C5239 S.n4767 VSUBS 1.88fF $ **FLOATING
C5240 S.n4768 VSUBS 2.67fF $ **FLOATING
C5241 S.t1691 VSUBS 0.02fF
C5242 S.n4769 VSUBS 0.24fF $ **FLOATING
C5243 S.n4770 VSUBS 0.36fF $ **FLOATING
C5244 S.n4771 VSUBS 0.61fF $ **FLOATING
C5245 S.n4772 VSUBS 0.12fF $ **FLOATING
C5246 S.t1903 VSUBS 0.02fF
C5247 S.n4773 VSUBS 0.14fF $ **FLOATING
C5248 S.n4775 VSUBS 1.88fF $ **FLOATING
C5249 S.n4776 VSUBS 2.67fF $ **FLOATING
C5250 S.t1719 VSUBS 0.02fF
C5251 S.n4777 VSUBS 0.24fF $ **FLOATING
C5252 S.n4778 VSUBS 0.36fF $ **FLOATING
C5253 S.n4779 VSUBS 0.61fF $ **FLOATING
C5254 S.t2560 VSUBS 0.02fF
C5255 S.n4780 VSUBS 0.24fF $ **FLOATING
C5256 S.n4781 VSUBS 0.91fF $ **FLOATING
C5257 S.n4782 VSUBS 0.05fF $ **FLOATING
C5258 S.t282 VSUBS 0.02fF
C5259 S.n4783 VSUBS 0.12fF $ **FLOATING
C5260 S.n4784 VSUBS 0.14fF $ **FLOATING
C5261 S.n4786 VSUBS 0.12fF $ **FLOATING
C5262 S.t1931 VSUBS 0.02fF
C5263 S.n4787 VSUBS 0.14fF $ **FLOATING
C5264 S.n4789 VSUBS 2.30fF $ **FLOATING
C5265 S.n4790 VSUBS 2.94fF $ **FLOATING
C5266 S.n4791 VSUBS 5.16fF $ **FLOATING
C5267 S.t252 VSUBS 0.02fF
C5268 S.n4792 VSUBS 0.12fF $ **FLOATING
C5269 S.n4793 VSUBS 0.14fF $ **FLOATING
C5270 S.t2532 VSUBS 0.02fF
C5271 S.n4795 VSUBS 0.24fF $ **FLOATING
C5272 S.n4796 VSUBS 0.91fF $ **FLOATING
C5273 S.n4797 VSUBS 0.05fF $ **FLOATING
C5274 S.n4798 VSUBS 1.88fF $ **FLOATING
C5275 S.n4799 VSUBS 2.67fF $ **FLOATING
C5276 S.t2478 VSUBS 0.02fF
C5277 S.n4800 VSUBS 0.24fF $ **FLOATING
C5278 S.n4801 VSUBS 0.36fF $ **FLOATING
C5279 S.n4802 VSUBS 0.61fF $ **FLOATING
C5280 S.n4803 VSUBS 0.12fF $ **FLOATING
C5281 S.t155 VSUBS 0.02fF
C5282 S.n4804 VSUBS 0.14fF $ **FLOATING
C5283 S.n4806 VSUBS 5.17fF $ **FLOATING
C5284 S.t1035 VSUBS 0.02fF
C5285 S.n4807 VSUBS 0.12fF $ **FLOATING
C5286 S.n4808 VSUBS 0.14fF $ **FLOATING
C5287 S.t795 VSUBS 0.02fF
C5288 S.n4810 VSUBS 0.24fF $ **FLOATING
C5289 S.n4811 VSUBS 0.91fF $ **FLOATING
C5290 S.n4812 VSUBS 0.05fF $ **FLOATING
C5291 S.n4813 VSUBS 1.88fF $ **FLOATING
C5292 S.n4814 VSUBS 0.12fF $ **FLOATING
C5293 S.t948 VSUBS 0.02fF
C5294 S.n4815 VSUBS 0.14fF $ **FLOATING
C5295 S.t737 VSUBS 0.02fF
C5296 S.n4817 VSUBS 0.24fF $ **FLOATING
C5297 S.n4818 VSUBS 0.36fF $ **FLOATING
C5298 S.n4819 VSUBS 0.61fF $ **FLOATING
C5299 S.n4820 VSUBS 2.67fF $ **FLOATING
C5300 S.n4821 VSUBS 4.90fF $ **FLOATING
C5301 S.t1817 VSUBS 0.02fF
C5302 S.n4822 VSUBS 0.12fF $ **FLOATING
C5303 S.n4823 VSUBS 0.14fF $ **FLOATING
C5304 S.t1575 VSUBS 0.02fF
C5305 S.n4825 VSUBS 0.24fF $ **FLOATING
C5306 S.n4826 VSUBS 0.91fF $ **FLOATING
C5307 S.n4827 VSUBS 0.05fF $ **FLOATING
C5308 S.n4828 VSUBS 1.88fF $ **FLOATING
C5309 S.n4829 VSUBS 2.67fF $ **FLOATING
C5310 S.t1529 VSUBS 0.02fF
C5311 S.n4830 VSUBS 0.24fF $ **FLOATING
C5312 S.n4831 VSUBS 0.36fF $ **FLOATING
C5313 S.n4832 VSUBS 0.61fF $ **FLOATING
C5314 S.n4833 VSUBS 0.12fF $ **FLOATING
C5315 S.t1731 VSUBS 0.02fF
C5316 S.n4834 VSUBS 0.14fF $ **FLOATING
C5317 S.n4836 VSUBS 1.88fF $ **FLOATING
C5318 S.n4837 VSUBS 2.68fF $ **FLOATING
C5319 S.t1552 VSUBS 0.02fF
C5320 S.n4838 VSUBS 0.24fF $ **FLOATING
C5321 S.n4839 VSUBS 0.36fF $ **FLOATING
C5322 S.n4840 VSUBS 0.61fF $ **FLOATING
C5323 S.t865 VSUBS 0.02fF
C5324 S.n4841 VSUBS 1.22fF $ **FLOATING
C5325 S.n4842 VSUBS 0.61fF $ **FLOATING
C5326 S.n4843 VSUBS 0.35fF $ **FLOATING
C5327 S.n4844 VSUBS 0.63fF $ **FLOATING
C5328 S.n4845 VSUBS 1.15fF $ **FLOATING
C5329 S.n4846 VSUBS 3.00fF $ **FLOATING
C5330 S.n4847 VSUBS 0.59fF $ **FLOATING
C5331 S.n4848 VSUBS 0.01fF $ **FLOATING
C5332 S.n4849 VSUBS 0.97fF $ **FLOATING
C5333 S.t9 VSUBS 21.42fF
C5334 S.n4850 VSUBS 20.29fF $ **FLOATING
C5335 S.n4852 VSUBS 0.38fF $ **FLOATING
C5336 S.n4853 VSUBS 0.23fF $ **FLOATING
C5337 S.n4854 VSUBS 2.90fF $ **FLOATING
C5338 S.n4855 VSUBS 2.46fF $ **FLOATING
C5339 S.n4856 VSUBS 1.96fF $ **FLOATING
C5340 S.n4857 VSUBS 3.94fF $ **FLOATING
C5341 S.n4858 VSUBS 0.25fF $ **FLOATING
C5342 S.n4859 VSUBS 0.01fF $ **FLOATING
C5343 S.t2573 VSUBS 0.02fF
C5344 S.n4860 VSUBS 0.26fF $ **FLOATING
C5345 S.t1164 VSUBS 0.02fF
C5346 S.n4861 VSUBS 0.95fF $ **FLOATING
C5347 S.n4862 VSUBS 0.71fF $ **FLOATING
C5348 S.n4863 VSUBS 0.78fF $ **FLOATING
C5349 S.n4864 VSUBS 1.93fF $ **FLOATING
C5350 S.n4865 VSUBS 1.88fF $ **FLOATING
C5351 S.n4866 VSUBS 0.12fF $ **FLOATING
C5352 S.t838 VSUBS 0.02fF
C5353 S.n4867 VSUBS 0.14fF $ **FLOATING
C5354 S.t1648 VSUBS 0.02fF
C5355 S.n4869 VSUBS 0.24fF $ **FLOATING
C5356 S.n4870 VSUBS 0.36fF $ **FLOATING
C5357 S.n4871 VSUBS 0.61fF $ **FLOATING
C5358 S.n4872 VSUBS 1.52fF $ **FLOATING
C5359 S.n4873 VSUBS 2.99fF $ **FLOATING
C5360 S.t1951 VSUBS 0.02fF
C5361 S.n4874 VSUBS 0.24fF $ **FLOATING
C5362 S.n4875 VSUBS 0.91fF $ **FLOATING
C5363 S.n4876 VSUBS 0.05fF $ **FLOATING
C5364 S.t1703 VSUBS 0.02fF
C5365 S.n4877 VSUBS 0.12fF $ **FLOATING
C5366 S.n4878 VSUBS 0.14fF $ **FLOATING
C5367 S.n4880 VSUBS 1.89fF $ **FLOATING
C5368 S.n4881 VSUBS 1.88fF $ **FLOATING
C5369 S.t2435 VSUBS 0.02fF
C5370 S.n4882 VSUBS 0.24fF $ **FLOATING
C5371 S.n4883 VSUBS 0.36fF $ **FLOATING
C5372 S.n4884 VSUBS 0.61fF $ **FLOATING
C5373 S.n4885 VSUBS 0.12fF $ **FLOATING
C5374 S.t1754 VSUBS 0.02fF
C5375 S.n4886 VSUBS 0.14fF $ **FLOATING
C5376 S.n4888 VSUBS 1.16fF $ **FLOATING
C5377 S.n4889 VSUBS 0.22fF $ **FLOATING
C5378 S.n4890 VSUBS 0.25fF $ **FLOATING
C5379 S.n4891 VSUBS 0.09fF $ **FLOATING
C5380 S.n4892 VSUBS 1.88fF $ **FLOATING
C5381 S.t209 VSUBS 0.02fF
C5382 S.n4893 VSUBS 0.24fF $ **FLOATING
C5383 S.n4894 VSUBS 0.91fF $ **FLOATING
C5384 S.n4895 VSUBS 0.05fF $ **FLOATING
C5385 S.t2493 VSUBS 0.02fF
C5386 S.n4896 VSUBS 0.12fF $ **FLOATING
C5387 S.n4897 VSUBS 0.14fF $ **FLOATING
C5388 S.n4899 VSUBS 0.78fF $ **FLOATING
C5389 S.n4900 VSUBS 1.94fF $ **FLOATING
C5390 S.n4901 VSUBS 1.88fF $ **FLOATING
C5391 S.n4902 VSUBS 0.12fF $ **FLOATING
C5392 S.t2536 VSUBS 0.02fF
C5393 S.n4903 VSUBS 0.14fF $ **FLOATING
C5394 S.t832 VSUBS 0.02fF
C5395 S.n4905 VSUBS 0.24fF $ **FLOATING
C5396 S.n4906 VSUBS 0.36fF $ **FLOATING
C5397 S.n4907 VSUBS 0.61fF $ **FLOATING
C5398 S.n4908 VSUBS 1.84fF $ **FLOATING
C5399 S.n4909 VSUBS 2.99fF $ **FLOATING
C5400 S.t1135 VSUBS 0.02fF
C5401 S.n4910 VSUBS 0.24fF $ **FLOATING
C5402 S.n4911 VSUBS 0.91fF $ **FLOATING
C5403 S.n4912 VSUBS 0.05fF $ **FLOATING
C5404 S.t886 VSUBS 0.02fF
C5405 S.n4913 VSUBS 0.12fF $ **FLOATING
C5406 S.n4914 VSUBS 0.14fF $ **FLOATING
C5407 S.n4916 VSUBS 1.89fF $ **FLOATING
C5408 S.n4917 VSUBS 1.88fF $ **FLOATING
C5409 S.t448 VSUBS 0.02fF
C5410 S.n4918 VSUBS 0.24fF $ **FLOATING
C5411 S.n4919 VSUBS 0.36fF $ **FLOATING
C5412 S.n4920 VSUBS 0.61fF $ **FLOATING
C5413 S.n4921 VSUBS 0.12fF $ **FLOATING
C5414 S.t2154 VSUBS 0.02fF
C5415 S.n4922 VSUBS 0.14fF $ **FLOATING
C5416 S.n4924 VSUBS 1.16fF $ **FLOATING
C5417 S.n4925 VSUBS 0.22fF $ **FLOATING
C5418 S.n4926 VSUBS 0.25fF $ **FLOATING
C5419 S.n4927 VSUBS 0.09fF $ **FLOATING
C5420 S.n4928 VSUBS 1.88fF $ **FLOATING
C5421 S.t719 VSUBS 0.02fF
C5422 S.n4929 VSUBS 0.24fF $ **FLOATING
C5423 S.n4930 VSUBS 0.91fF $ **FLOATING
C5424 S.n4931 VSUBS 0.05fF $ **FLOATING
C5425 S.t502 VSUBS 0.02fF
C5426 S.n4932 VSUBS 0.12fF $ **FLOATING
C5427 S.n4933 VSUBS 0.14fF $ **FLOATING
C5428 S.n4935 VSUBS 0.78fF $ **FLOATING
C5429 S.n4936 VSUBS 1.94fF $ **FLOATING
C5430 S.n4937 VSUBS 1.88fF $ **FLOATING
C5431 S.n4938 VSUBS 0.12fF $ **FLOATING
C5432 S.t423 VSUBS 0.02fF
C5433 S.n4939 VSUBS 0.14fF $ **FLOATING
C5434 S.t1238 VSUBS 0.02fF
C5435 S.n4941 VSUBS 0.24fF $ **FLOATING
C5436 S.n4942 VSUBS 0.36fF $ **FLOATING
C5437 S.n4943 VSUBS 0.61fF $ **FLOATING
C5438 S.n4944 VSUBS 1.84fF $ **FLOATING
C5439 S.n4945 VSUBS 2.99fF $ **FLOATING
C5440 S.t1511 VSUBS 0.02fF
C5441 S.n4946 VSUBS 0.24fF $ **FLOATING
C5442 S.n4947 VSUBS 0.91fF $ **FLOATING
C5443 S.n4948 VSUBS 0.05fF $ **FLOATING
C5444 S.t1288 VSUBS 0.02fF
C5445 S.n4949 VSUBS 0.12fF $ **FLOATING
C5446 S.n4950 VSUBS 0.14fF $ **FLOATING
C5447 S.n4952 VSUBS 1.89fF $ **FLOATING
C5448 S.n4953 VSUBS 1.88fF $ **FLOATING
C5449 S.t2022 VSUBS 0.02fF
C5450 S.n4954 VSUBS 0.24fF $ **FLOATING
C5451 S.n4955 VSUBS 0.36fF $ **FLOATING
C5452 S.n4956 VSUBS 0.61fF $ **FLOATING
C5453 S.n4957 VSUBS 0.12fF $ **FLOATING
C5454 S.t1218 VSUBS 0.02fF
C5455 S.n4958 VSUBS 0.14fF $ **FLOATING
C5456 S.n4960 VSUBS 1.16fF $ **FLOATING
C5457 S.n4961 VSUBS 0.22fF $ **FLOATING
C5458 S.n4962 VSUBS 0.25fF $ **FLOATING
C5459 S.n4963 VSUBS 0.09fF $ **FLOATING
C5460 S.n4964 VSUBS 1.88fF $ **FLOATING
C5461 S.t2297 VSUBS 0.02fF
C5462 S.n4965 VSUBS 0.24fF $ **FLOATING
C5463 S.n4966 VSUBS 0.91fF $ **FLOATING
C5464 S.n4967 VSUBS 0.05fF $ **FLOATING
C5465 S.t2076 VSUBS 0.02fF
C5466 S.n4968 VSUBS 0.12fF $ **FLOATING
C5467 S.n4969 VSUBS 0.14fF $ **FLOATING
C5468 S.n4971 VSUBS 0.78fF $ **FLOATING
C5469 S.n4972 VSUBS 1.94fF $ **FLOATING
C5470 S.n4973 VSUBS 1.88fF $ **FLOATING
C5471 S.n4974 VSUBS 0.12fF $ **FLOATING
C5472 S.t2119 VSUBS 0.02fF
C5473 S.n4975 VSUBS 0.14fF $ **FLOATING
C5474 S.t291 VSUBS 0.02fF
C5475 S.n4977 VSUBS 0.24fF $ **FLOATING
C5476 S.n4978 VSUBS 0.36fF $ **FLOATING
C5477 S.n4979 VSUBS 0.61fF $ **FLOATING
C5478 S.n4980 VSUBS 1.84fF $ **FLOATING
C5479 S.n4981 VSUBS 2.99fF $ **FLOATING
C5480 S.t568 VSUBS 0.02fF
C5481 S.n4982 VSUBS 0.24fF $ **FLOATING
C5482 S.n4983 VSUBS 0.91fF $ **FLOATING
C5483 S.n4984 VSUBS 0.05fF $ **FLOATING
C5484 S.t347 VSUBS 0.02fF
C5485 S.n4985 VSUBS 0.12fF $ **FLOATING
C5486 S.n4986 VSUBS 0.14fF $ **FLOATING
C5487 S.n4988 VSUBS 1.89fF $ **FLOATING
C5488 S.n4989 VSUBS 1.75fF $ **FLOATING
C5489 S.t2535 VSUBS 0.02fF
C5490 S.n4990 VSUBS 0.24fF $ **FLOATING
C5491 S.n4991 VSUBS 0.36fF $ **FLOATING
C5492 S.n4992 VSUBS 0.61fF $ **FLOATING
C5493 S.n4993 VSUBS 0.12fF $ **FLOATING
C5494 S.t1721 VSUBS 0.02fF
C5495 S.n4994 VSUBS 0.14fF $ **FLOATING
C5496 S.n4996 VSUBS 1.16fF $ **FLOATING
C5497 S.n4997 VSUBS 0.22fF $ **FLOATING
C5498 S.n4998 VSUBS 0.25fF $ **FLOATING
C5499 S.n4999 VSUBS 0.09fF $ **FLOATING
C5500 S.n5000 VSUBS 2.44fF $ **FLOATING
C5501 S.t316 VSUBS 0.02fF
C5502 S.n5001 VSUBS 0.24fF $ **FLOATING
C5503 S.n5002 VSUBS 0.91fF $ **FLOATING
C5504 S.n5003 VSUBS 0.05fF $ **FLOATING
C5505 S.t1252 VSUBS 0.02fF
C5506 S.n5004 VSUBS 0.12fF $ **FLOATING
C5507 S.n5005 VSUBS 0.14fF $ **FLOATING
C5508 S.n5007 VSUBS 1.88fF $ **FLOATING
C5509 S.n5008 VSUBS 0.48fF $ **FLOATING
C5510 S.n5009 VSUBS 0.09fF $ **FLOATING
C5511 S.n5010 VSUBS 0.33fF $ **FLOATING
C5512 S.n5011 VSUBS 0.30fF $ **FLOATING
C5513 S.n5012 VSUBS 0.77fF $ **FLOATING
C5514 S.n5013 VSUBS 0.59fF $ **FLOATING
C5515 S.t799 VSUBS 0.02fF
C5516 S.n5014 VSUBS 0.24fF $ **FLOATING
C5517 S.n5015 VSUBS 0.36fF $ **FLOATING
C5518 S.n5016 VSUBS 0.61fF $ **FLOATING
C5519 S.n5017 VSUBS 0.12fF $ **FLOATING
C5520 S.t2508 VSUBS 0.02fF
C5521 S.n5018 VSUBS 0.14fF $ **FLOATING
C5522 S.n5020 VSUBS 2.61fF $ **FLOATING
C5523 S.n5021 VSUBS 2.15fF $ **FLOATING
C5524 S.t1105 VSUBS 0.02fF
C5525 S.n5022 VSUBS 0.24fF $ **FLOATING
C5526 S.n5023 VSUBS 0.91fF $ **FLOATING
C5527 S.n5024 VSUBS 0.05fF $ **FLOATING
C5528 S.t856 VSUBS 0.02fF
C5529 S.n5025 VSUBS 0.12fF $ **FLOATING
C5530 S.n5026 VSUBS 0.14fF $ **FLOATING
C5531 S.n5028 VSUBS 0.78fF $ **FLOATING
C5532 S.n5029 VSUBS 2.30fF $ **FLOATING
C5533 S.n5030 VSUBS 1.88fF $ **FLOATING
C5534 S.n5031 VSUBS 0.12fF $ **FLOATING
C5535 S.t768 VSUBS 0.02fF
C5536 S.n5032 VSUBS 0.14fF $ **FLOATING
C5537 S.t1580 VSUBS 0.02fF
C5538 S.n5034 VSUBS 0.24fF $ **FLOATING
C5539 S.n5035 VSUBS 0.36fF $ **FLOATING
C5540 S.n5036 VSUBS 0.61fF $ **FLOATING
C5541 S.n5037 VSUBS 1.39fF $ **FLOATING
C5542 S.n5038 VSUBS 0.71fF $ **FLOATING
C5543 S.n5039 VSUBS 1.14fF $ **FLOATING
C5544 S.n5040 VSUBS 0.35fF $ **FLOATING
C5545 S.n5041 VSUBS 2.02fF $ **FLOATING
C5546 S.t1885 VSUBS 0.02fF
C5547 S.n5042 VSUBS 0.24fF $ **FLOATING
C5548 S.n5043 VSUBS 0.91fF $ **FLOATING
C5549 S.n5044 VSUBS 0.05fF $ **FLOATING
C5550 S.t1639 VSUBS 0.02fF
C5551 S.n5045 VSUBS 0.12fF $ **FLOATING
C5552 S.n5046 VSUBS 0.14fF $ **FLOATING
C5553 S.n5048 VSUBS 1.89fF $ **FLOATING
C5554 S.n5049 VSUBS 1.88fF $ **FLOATING
C5555 S.t2371 VSUBS 0.02fF
C5556 S.n5050 VSUBS 0.24fF $ **FLOATING
C5557 S.n5051 VSUBS 0.36fF $ **FLOATING
C5558 S.n5052 VSUBS 0.61fF $ **FLOATING
C5559 S.n5053 VSUBS 0.12fF $ **FLOATING
C5560 S.t1556 VSUBS 0.02fF
C5561 S.n5054 VSUBS 0.14fF $ **FLOATING
C5562 S.n5056 VSUBS 1.16fF $ **FLOATING
C5563 S.n5057 VSUBS 0.22fF $ **FLOATING
C5564 S.n5058 VSUBS 0.25fF $ **FLOATING
C5565 S.n5059 VSUBS 0.09fF $ **FLOATING
C5566 S.n5060 VSUBS 1.88fF $ **FLOATING
C5567 S.t134 VSUBS 0.02fF
C5568 S.n5061 VSUBS 0.24fF $ **FLOATING
C5569 S.n5062 VSUBS 0.91fF $ **FLOATING
C5570 S.n5063 VSUBS 0.05fF $ **FLOATING
C5571 S.t2423 VSUBS 0.02fF
C5572 S.n5064 VSUBS 0.12fF $ **FLOATING
C5573 S.n5065 VSUBS 0.14fF $ **FLOATING
C5574 S.n5067 VSUBS 20.78fF $ **FLOATING
C5575 S.n5068 VSUBS 1.88fF $ **FLOATING
C5576 S.n5069 VSUBS 2.67fF $ **FLOATING
C5577 S.t2504 VSUBS 0.02fF
C5578 S.n5070 VSUBS 0.24fF $ **FLOATING
C5579 S.n5071 VSUBS 0.36fF $ **FLOATING
C5580 S.n5072 VSUBS 0.61fF $ **FLOATING
C5581 S.n5073 VSUBS 0.12fF $ **FLOATING
C5582 S.t189 VSUBS 0.02fF
C5583 S.n5074 VSUBS 0.14fF $ **FLOATING
C5584 S.n5076 VSUBS 2.80fF $ **FLOATING
C5585 S.n5077 VSUBS 2.30fF $ **FLOATING
C5586 S.t1063 VSUBS 0.02fF
C5587 S.n5078 VSUBS 0.12fF $ **FLOATING
C5588 S.n5079 VSUBS 0.14fF $ **FLOATING
C5589 S.t826 VSUBS 0.02fF
C5590 S.n5081 VSUBS 0.24fF $ **FLOATING
C5591 S.n5082 VSUBS 0.91fF $ **FLOATING
C5592 S.n5083 VSUBS 0.05fF $ **FLOATING
C5593 S.n5084 VSUBS 2.80fF $ **FLOATING
C5594 S.n5085 VSUBS 1.88fF $ **FLOATING
C5595 S.n5086 VSUBS 0.12fF $ **FLOATING
C5596 S.t977 VSUBS 0.02fF
C5597 S.n5087 VSUBS 0.14fF $ **FLOATING
C5598 S.t762 VSUBS 0.02fF
C5599 S.n5089 VSUBS 0.24fF $ **FLOATING
C5600 S.n5090 VSUBS 0.36fF $ **FLOATING
C5601 S.n5091 VSUBS 0.61fF $ **FLOATING
C5602 S.n5092 VSUBS 2.67fF $ **FLOATING
C5603 S.n5093 VSUBS 2.30fF $ **FLOATING
C5604 S.t1848 VSUBS 0.02fF
C5605 S.n5094 VSUBS 0.12fF $ **FLOATING
C5606 S.n5095 VSUBS 0.14fF $ **FLOATING
C5607 S.t1608 VSUBS 0.02fF
C5608 S.n5097 VSUBS 0.24fF $ **FLOATING
C5609 S.n5098 VSUBS 0.91fF $ **FLOATING
C5610 S.n5099 VSUBS 0.05fF $ **FLOATING
C5611 S.n5100 VSUBS 2.73fF $ **FLOATING
C5612 S.n5101 VSUBS 1.59fF $ **FLOATING
C5613 S.n5102 VSUBS 0.12fF $ **FLOATING
C5614 S.t542 VSUBS 0.02fF
C5615 S.n5103 VSUBS 0.14fF $ **FLOATING
C5616 S.t2140 VSUBS 0.02fF
C5617 S.n5105 VSUBS 0.24fF $ **FLOATING
C5618 S.n5106 VSUBS 0.36fF $ **FLOATING
C5619 S.n5107 VSUBS 0.61fF $ **FLOATING
C5620 S.n5108 VSUBS 0.07fF $ **FLOATING
C5621 S.n5109 VSUBS 0.01fF $ **FLOATING
C5622 S.n5110 VSUBS 0.24fF $ **FLOATING
C5623 S.n5111 VSUBS 1.16fF $ **FLOATING
C5624 S.n5112 VSUBS 1.35fF $ **FLOATING
C5625 S.n5113 VSUBS 2.30fF $ **FLOATING
C5626 S.t889 VSUBS 0.02fF
C5627 S.n5114 VSUBS 0.12fF $ **FLOATING
C5628 S.n5115 VSUBS 0.14fF $ **FLOATING
C5629 S.t1021 VSUBS 0.02fF
C5630 S.n5117 VSUBS 0.24fF $ **FLOATING
C5631 S.n5118 VSUBS 0.91fF $ **FLOATING
C5632 S.n5119 VSUBS 0.05fF $ **FLOATING
C5633 S.t77 VSUBS 48.27fF
C5634 S.t2398 VSUBS 0.02fF
C5635 S.n5120 VSUBS 0.24fF $ **FLOATING
C5636 S.n5121 VSUBS 0.91fF $ **FLOATING
C5637 S.n5122 VSUBS 0.05fF $ **FLOATING
C5638 S.t78 VSUBS 0.02fF
C5639 S.n5123 VSUBS 0.12fF $ **FLOATING
C5640 S.n5124 VSUBS 0.14fF $ **FLOATING
C5641 S.n5126 VSUBS 0.12fF $ **FLOATING
C5642 S.t1759 VSUBS 0.02fF
C5643 S.n5127 VSUBS 0.14fF $ **FLOATING
C5644 S.n5129 VSUBS 5.17fF $ **FLOATING
C5645 S.n5130 VSUBS 5.44fF $ **FLOATING
C5646 S.t34 VSUBS 0.02fF
C5647 S.n5131 VSUBS 0.12fF $ **FLOATING
C5648 S.n5132 VSUBS 0.14fF $ **FLOATING
C5649 S.t2368 VSUBS 0.02fF
C5650 S.n5134 VSUBS 0.24fF $ **FLOATING
C5651 S.n5135 VSUBS 0.91fF $ **FLOATING
C5652 S.n5136 VSUBS 0.05fF $ **FLOATING
C5653 S.t33 VSUBS 47.89fF
C5654 S.t1917 VSUBS 0.02fF
C5655 S.n5137 VSUBS 0.01fF $ **FLOATING
C5656 S.n5138 VSUBS 0.26fF $ **FLOATING
C5657 S.t1450 VSUBS 0.02fF
C5658 S.n5140 VSUBS 1.19fF $ **FLOATING
C5659 S.n5141 VSUBS 0.05fF $ **FLOATING
C5660 S.t1179 VSUBS 0.02fF
C5661 S.n5142 VSUBS 0.64fF $ **FLOATING
C5662 S.n5143 VSUBS 0.61fF $ **FLOATING
C5663 S.n5144 VSUBS 8.97fF $ **FLOATING
C5664 S.n5145 VSUBS 8.97fF $ **FLOATING
C5665 S.n5146 VSUBS 0.60fF $ **FLOATING
C5666 S.n5147 VSUBS 0.22fF $ **FLOATING
C5667 S.n5148 VSUBS 0.59fF $ **FLOATING
C5668 S.n5149 VSUBS 3.39fF $ **FLOATING
C5669 S.n5150 VSUBS 0.29fF $ **FLOATING
C5670 S.t133 VSUBS 21.42fF
C5671 S.n5151 VSUBS 21.71fF $ **FLOATING
C5672 S.n5152 VSUBS 0.77fF $ **FLOATING
C5673 S.n5153 VSUBS 0.28fF $ **FLOATING
C5674 S.n5154 VSUBS 4.00fF $ **FLOATING
C5675 S.n5155 VSUBS 1.35fF $ **FLOATING
C5676 S.n5156 VSUBS 0.01fF $ **FLOATING
C5677 S.n5157 VSUBS 0.02fF $ **FLOATING
C5678 S.n5158 VSUBS 0.03fF $ **FLOATING
C5679 S.n5159 VSUBS 0.04fF $ **FLOATING
C5680 S.n5160 VSUBS 0.17fF $ **FLOATING
C5681 S.n5161 VSUBS 0.01fF $ **FLOATING
C5682 S.n5162 VSUBS 0.02fF $ **FLOATING
C5683 S.n5163 VSUBS 0.01fF $ **FLOATING
C5684 S.n5164 VSUBS 0.01fF $ **FLOATING
C5685 S.n5165 VSUBS 0.01fF $ **FLOATING
C5686 S.n5166 VSUBS 0.01fF $ **FLOATING
C5687 S.n5167 VSUBS 0.02fF $ **FLOATING
C5688 S.n5168 VSUBS 0.01fF $ **FLOATING
C5689 S.n5169 VSUBS 0.02fF $ **FLOATING
C5690 S.n5170 VSUBS 0.05fF $ **FLOATING
C5691 S.n5171 VSUBS 0.04fF $ **FLOATING
C5692 S.n5172 VSUBS 0.11fF $ **FLOATING
C5693 S.n5173 VSUBS 0.38fF $ **FLOATING
C5694 S.n5174 VSUBS 0.20fF $ **FLOATING
C5695 S.n5175 VSUBS 4.39fF $ **FLOATING
C5696 S.n5176 VSUBS 0.24fF $ **FLOATING
C5697 S.n5177 VSUBS 1.50fF $ **FLOATING
C5698 S.n5178 VSUBS 1.31fF $ **FLOATING
C5699 S.n5179 VSUBS 0.28fF $ **FLOATING
C5700 S.n5180 VSUBS 1.89fF $ **FLOATING
C5701 S.n5181 VSUBS 0.06fF $ **FLOATING
C5702 S.n5182 VSUBS 0.03fF $ **FLOATING
C5703 S.n5183 VSUBS 0.04fF $ **FLOATING
C5704 S.n5184 VSUBS 0.99fF $ **FLOATING
C5705 S.n5185 VSUBS 0.02fF $ **FLOATING
C5706 S.n5186 VSUBS 0.01fF $ **FLOATING
C5707 S.n5187 VSUBS 0.02fF $ **FLOATING
C5708 S.n5188 VSUBS 0.08fF $ **FLOATING
C5709 S.n5189 VSUBS 0.36fF $ **FLOATING
C5710 S.n5190 VSUBS 1.85fF $ **FLOATING
C5711 S.t507 VSUBS 0.02fF
C5712 S.n5191 VSUBS 0.24fF $ **FLOATING
C5713 S.n5192 VSUBS 0.36fF $ **FLOATING
C5714 S.n5193 VSUBS 0.61fF $ **FLOATING
C5715 S.n5194 VSUBS 0.12fF $ **FLOATING
C5716 S.t2213 VSUBS 0.02fF
C5717 S.n5195 VSUBS 0.14fF $ **FLOATING
C5718 S.n5197 VSUBS 0.70fF $ **FLOATING
C5719 S.n5198 VSUBS 0.23fF $ **FLOATING
C5720 S.n5199 VSUBS 0.23fF $ **FLOATING
C5721 S.n5200 VSUBS 0.70fF $ **FLOATING
C5722 S.n5201 VSUBS 1.16fF $ **FLOATING
C5723 S.n5202 VSUBS 0.22fF $ **FLOATING
C5724 S.n5203 VSUBS 0.25fF $ **FLOATING
C5725 S.n5204 VSUBS 0.09fF $ **FLOATING
C5726 S.n5205 VSUBS 1.88fF $ **FLOATING
C5727 S.t781 VSUBS 0.02fF
C5728 S.n5206 VSUBS 0.24fF $ **FLOATING
C5729 S.n5207 VSUBS 0.91fF $ **FLOATING
C5730 S.n5208 VSUBS 0.05fF $ **FLOATING
C5731 S.t558 VSUBS 0.02fF
C5732 S.n5209 VSUBS 0.12fF $ **FLOATING
C5733 S.n5210 VSUBS 0.14fF $ **FLOATING
C5734 S.n5212 VSUBS 0.25fF $ **FLOATING
C5735 S.n5213 VSUBS 0.09fF $ **FLOATING
C5736 S.n5214 VSUBS 0.21fF $ **FLOATING
C5737 S.n5215 VSUBS 0.92fF $ **FLOATING
C5738 S.n5216 VSUBS 0.44fF $ **FLOATING
C5739 S.n5217 VSUBS 1.88fF $ **FLOATING
C5740 S.n5218 VSUBS 0.12fF $ **FLOATING
C5741 S.t596 VSUBS 0.02fF
C5742 S.n5219 VSUBS 0.14fF $ **FLOATING
C5743 S.t1415 VSUBS 0.02fF
C5744 S.n5221 VSUBS 0.24fF $ **FLOATING
C5745 S.n5222 VSUBS 0.36fF $ **FLOATING
C5746 S.n5223 VSUBS 0.61fF $ **FLOATING
C5747 S.n5224 VSUBS 0.02fF $ **FLOATING
C5748 S.n5225 VSUBS 0.01fF $ **FLOATING
C5749 S.n5226 VSUBS 0.02fF $ **FLOATING
C5750 S.n5227 VSUBS 0.08fF $ **FLOATING
C5751 S.n5228 VSUBS 0.06fF $ **FLOATING
C5752 S.n5229 VSUBS 0.03fF $ **FLOATING
C5753 S.n5230 VSUBS 0.04fF $ **FLOATING
C5754 S.n5231 VSUBS 1.00fF $ **FLOATING
C5755 S.n5232 VSUBS 0.36fF $ **FLOATING
C5756 S.n5233 VSUBS 1.87fF $ **FLOATING
C5757 S.n5234 VSUBS 1.99fF $ **FLOATING
C5758 S.t1696 VSUBS 0.02fF
C5759 S.n5235 VSUBS 0.24fF $ **FLOATING
C5760 S.n5236 VSUBS 0.91fF $ **FLOATING
C5761 S.n5237 VSUBS 0.05fF $ **FLOATING
C5762 S.t1463 VSUBS 0.02fF
C5763 S.n5238 VSUBS 0.12fF $ **FLOATING
C5764 S.n5239 VSUBS 0.14fF $ **FLOATING
C5765 S.n5241 VSUBS 1.89fF $ **FLOATING
C5766 S.n5242 VSUBS 0.06fF $ **FLOATING
C5767 S.n5243 VSUBS 0.03fF $ **FLOATING
C5768 S.n5244 VSUBS 0.04fF $ **FLOATING
C5769 S.n5245 VSUBS 0.99fF $ **FLOATING
C5770 S.n5246 VSUBS 0.02fF $ **FLOATING
C5771 S.n5247 VSUBS 0.01fF $ **FLOATING
C5772 S.n5248 VSUBS 0.02fF $ **FLOATING
C5773 S.n5249 VSUBS 0.08fF $ **FLOATING
C5774 S.n5250 VSUBS 0.36fF $ **FLOATING
C5775 S.n5251 VSUBS 1.85fF $ **FLOATING
C5776 S.t1033 VSUBS 0.02fF
C5777 S.n5252 VSUBS 0.24fF $ **FLOATING
C5778 S.n5253 VSUBS 0.36fF $ **FLOATING
C5779 S.n5254 VSUBS 0.61fF $ **FLOATING
C5780 S.n5255 VSUBS 0.12fF $ **FLOATING
C5781 S.t213 VSUBS 0.02fF
C5782 S.n5256 VSUBS 0.14fF $ **FLOATING
C5783 S.n5258 VSUBS 0.70fF $ **FLOATING
C5784 S.n5259 VSUBS 0.23fF $ **FLOATING
C5785 S.n5260 VSUBS 0.23fF $ **FLOATING
C5786 S.n5261 VSUBS 0.70fF $ **FLOATING
C5787 S.n5262 VSUBS 1.16fF $ **FLOATING
C5788 S.n5263 VSUBS 0.22fF $ **FLOATING
C5789 S.n5264 VSUBS 0.25fF $ **FLOATING
C5790 S.n5265 VSUBS 0.09fF $ **FLOATING
C5791 S.n5266 VSUBS 1.88fF $ **FLOATING
C5792 S.t1315 VSUBS 0.02fF
C5793 S.n5267 VSUBS 0.24fF $ **FLOATING
C5794 S.n5268 VSUBS 0.91fF $ **FLOATING
C5795 S.n5269 VSUBS 0.05fF $ **FLOATING
C5796 S.t2251 VSUBS 0.02fF
C5797 S.n5270 VSUBS 0.12fF $ **FLOATING
C5798 S.n5271 VSUBS 0.14fF $ **FLOATING
C5799 S.n5273 VSUBS 0.25fF $ **FLOATING
C5800 S.n5274 VSUBS 0.09fF $ **FLOATING
C5801 S.n5275 VSUBS 0.21fF $ **FLOATING
C5802 S.n5276 VSUBS 0.92fF $ **FLOATING
C5803 S.n5277 VSUBS 0.44fF $ **FLOATING
C5804 S.n5278 VSUBS 1.88fF $ **FLOATING
C5805 S.n5279 VSUBS 0.12fF $ **FLOATING
C5806 S.t1001 VSUBS 0.02fF
C5807 S.n5280 VSUBS 0.14fF $ **FLOATING
C5808 S.t1812 VSUBS 0.02fF
C5809 S.n5282 VSUBS 0.24fF $ **FLOATING
C5810 S.n5283 VSUBS 0.36fF $ **FLOATING
C5811 S.n5284 VSUBS 0.61fF $ **FLOATING
C5812 S.n5285 VSUBS 0.02fF $ **FLOATING
C5813 S.n5286 VSUBS 0.01fF $ **FLOATING
C5814 S.n5287 VSUBS 0.02fF $ **FLOATING
C5815 S.n5288 VSUBS 0.08fF $ **FLOATING
C5816 S.n5289 VSUBS 0.06fF $ **FLOATING
C5817 S.n5290 VSUBS 0.03fF $ **FLOATING
C5818 S.n5291 VSUBS 0.04fF $ **FLOATING
C5819 S.n5292 VSUBS 1.00fF $ **FLOATING
C5820 S.n5293 VSUBS 0.36fF $ **FLOATING
C5821 S.n5294 VSUBS 1.87fF $ **FLOATING
C5822 S.n5295 VSUBS 1.99fF $ **FLOATING
C5823 S.t2101 VSUBS 0.02fF
C5824 S.n5296 VSUBS 0.24fF $ **FLOATING
C5825 S.n5297 VSUBS 0.91fF $ **FLOATING
C5826 S.n5298 VSUBS 0.05fF $ **FLOATING
C5827 S.t1867 VSUBS 0.02fF
C5828 S.n5299 VSUBS 0.12fF $ **FLOATING
C5829 S.n5300 VSUBS 0.14fF $ **FLOATING
C5830 S.n5302 VSUBS 1.89fF $ **FLOATING
C5831 S.n5303 VSUBS 0.06fF $ **FLOATING
C5832 S.n5304 VSUBS 0.03fF $ **FLOATING
C5833 S.n5305 VSUBS 0.04fF $ **FLOATING
C5834 S.n5306 VSUBS 0.99fF $ **FLOATING
C5835 S.n5307 VSUBS 0.02fF $ **FLOATING
C5836 S.n5308 VSUBS 0.01fF $ **FLOATING
C5837 S.n5309 VSUBS 0.02fF $ **FLOATING
C5838 S.n5310 VSUBS 0.08fF $ **FLOATING
C5839 S.n5311 VSUBS 0.36fF $ **FLOATING
C5840 S.n5312 VSUBS 1.85fF $ **FLOATING
C5841 S.t30 VSUBS 0.02fF
C5842 S.n5313 VSUBS 0.24fF $ **FLOATING
C5843 S.n5314 VSUBS 0.36fF $ **FLOATING
C5844 S.n5315 VSUBS 0.61fF $ **FLOATING
C5845 S.n5316 VSUBS 0.12fF $ **FLOATING
C5846 S.t1785 VSUBS 0.02fF
C5847 S.n5317 VSUBS 0.14fF $ **FLOATING
C5848 S.n5319 VSUBS 0.70fF $ **FLOATING
C5849 S.n5320 VSUBS 0.23fF $ **FLOATING
C5850 S.n5321 VSUBS 0.23fF $ **FLOATING
C5851 S.n5322 VSUBS 0.70fF $ **FLOATING
C5852 S.n5323 VSUBS 1.16fF $ **FLOATING
C5853 S.n5324 VSUBS 0.22fF $ **FLOATING
C5854 S.n5325 VSUBS 0.25fF $ **FLOATING
C5855 S.n5326 VSUBS 0.09fF $ **FLOATING
C5856 S.n5327 VSUBS 1.88fF $ **FLOATING
C5857 S.t373 VSUBS 0.02fF
C5858 S.n5328 VSUBS 0.24fF $ **FLOATING
C5859 S.n5329 VSUBS 0.91fF $ **FLOATING
C5860 S.n5330 VSUBS 0.05fF $ **FLOATING
C5861 S.t110 VSUBS 0.02fF
C5862 S.n5331 VSUBS 0.12fF $ **FLOATING
C5863 S.n5332 VSUBS 0.14fF $ **FLOATING
C5864 S.n5334 VSUBS 0.25fF $ **FLOATING
C5865 S.n5335 VSUBS 0.09fF $ **FLOATING
C5866 S.n5336 VSUBS 0.21fF $ **FLOATING
C5867 S.n5337 VSUBS 0.92fF $ **FLOATING
C5868 S.n5338 VSUBS 0.44fF $ **FLOATING
C5869 S.n5339 VSUBS 1.88fF $ **FLOATING
C5870 S.n5340 VSUBS 0.12fF $ **FLOATING
C5871 S.t2567 VSUBS 0.02fF
C5872 S.n5341 VSUBS 0.14fF $ **FLOATING
C5873 S.t862 VSUBS 0.02fF
C5874 S.n5343 VSUBS 0.24fF $ **FLOATING
C5875 S.n5344 VSUBS 0.36fF $ **FLOATING
C5876 S.n5345 VSUBS 0.61fF $ **FLOATING
C5877 S.n5346 VSUBS 0.02fF $ **FLOATING
C5878 S.n5347 VSUBS 0.01fF $ **FLOATING
C5879 S.n5348 VSUBS 0.02fF $ **FLOATING
C5880 S.n5349 VSUBS 0.08fF $ **FLOATING
C5881 S.n5350 VSUBS 0.06fF $ **FLOATING
C5882 S.n5351 VSUBS 0.03fF $ **FLOATING
C5883 S.n5352 VSUBS 0.04fF $ **FLOATING
C5884 S.n5353 VSUBS 1.00fF $ **FLOATING
C5885 S.n5354 VSUBS 0.36fF $ **FLOATING
C5886 S.n5355 VSUBS 1.87fF $ **FLOATING
C5887 S.n5356 VSUBS 1.99fF $ **FLOATING
C5888 S.t1160 VSUBS 0.02fF
C5889 S.n5357 VSUBS 0.24fF $ **FLOATING
C5890 S.n5358 VSUBS 0.91fF $ **FLOATING
C5891 S.n5359 VSUBS 0.05fF $ **FLOATING
C5892 S.t918 VSUBS 0.02fF
C5893 S.n5360 VSUBS 0.12fF $ **FLOATING
C5894 S.n5361 VSUBS 0.14fF $ **FLOATING
C5895 S.n5363 VSUBS 1.89fF $ **FLOATING
C5896 S.n5364 VSUBS 0.07fF $ **FLOATING
C5897 S.n5365 VSUBS 0.04fF $ **FLOATING
C5898 S.n5366 VSUBS 0.05fF $ **FLOATING
C5899 S.n5367 VSUBS 0.87fF $ **FLOATING
C5900 S.n5368 VSUBS 0.01fF $ **FLOATING
C5901 S.n5369 VSUBS 0.01fF $ **FLOATING
C5902 S.n5370 VSUBS 0.01fF $ **FLOATING
C5903 S.n5371 VSUBS 0.07fF $ **FLOATING
C5904 S.n5372 VSUBS 0.68fF $ **FLOATING
C5905 S.n5373 VSUBS 0.72fF $ **FLOATING
C5906 S.t1777 VSUBS 0.02fF
C5907 S.n5374 VSUBS 0.24fF $ **FLOATING
C5908 S.n5375 VSUBS 0.36fF $ **FLOATING
C5909 S.n5376 VSUBS 0.61fF $ **FLOATING
C5910 S.n5377 VSUBS 0.12fF $ **FLOATING
C5911 S.t962 VSUBS 0.02fF
C5912 S.n5378 VSUBS 0.14fF $ **FLOATING
C5913 S.n5380 VSUBS 0.70fF $ **FLOATING
C5914 S.n5381 VSUBS 0.23fF $ **FLOATING
C5915 S.n5382 VSUBS 0.23fF $ **FLOATING
C5916 S.n5383 VSUBS 0.70fF $ **FLOATING
C5917 S.n5384 VSUBS 1.16fF $ **FLOATING
C5918 S.n5385 VSUBS 0.22fF $ **FLOATING
C5919 S.n5386 VSUBS 0.25fF $ **FLOATING
C5920 S.n5387 VSUBS 0.09fF $ **FLOATING
C5921 S.n5388 VSUBS 2.31fF $ **FLOATING
C5922 S.t2069 VSUBS 0.02fF
C5923 S.n5389 VSUBS 0.24fF $ **FLOATING
C5924 S.n5390 VSUBS 0.91fF $ **FLOATING
C5925 S.n5391 VSUBS 0.05fF $ **FLOATING
C5926 S.t1835 VSUBS 0.02fF
C5927 S.n5392 VSUBS 0.12fF $ **FLOATING
C5928 S.n5393 VSUBS 0.14fF $ **FLOATING
C5929 S.n5395 VSUBS 1.88fF $ **FLOATING
C5930 S.n5396 VSUBS 0.46fF $ **FLOATING
C5931 S.n5397 VSUBS 0.22fF $ **FLOATING
C5932 S.n5398 VSUBS 0.38fF $ **FLOATING
C5933 S.n5399 VSUBS 0.16fF $ **FLOATING
C5934 S.n5400 VSUBS 0.28fF $ **FLOATING
C5935 S.n5401 VSUBS 0.21fF $ **FLOATING
C5936 S.n5402 VSUBS 0.30fF $ **FLOATING
C5937 S.n5403 VSUBS 0.42fF $ **FLOATING
C5938 S.n5404 VSUBS 0.21fF $ **FLOATING
C5939 S.t1388 VSUBS 0.02fF
C5940 S.n5405 VSUBS 0.24fF $ **FLOATING
C5941 S.n5406 VSUBS 0.36fF $ **FLOATING
C5942 S.n5407 VSUBS 0.61fF $ **FLOATING
C5943 S.n5408 VSUBS 0.12fF $ **FLOATING
C5944 S.t572 VSUBS 0.02fF
C5945 S.n5409 VSUBS 0.14fF $ **FLOATING
C5946 S.n5411 VSUBS 0.04fF $ **FLOATING
C5947 S.n5412 VSUBS 0.03fF $ **FLOATING
C5948 S.n5413 VSUBS 0.03fF $ **FLOATING
C5949 S.n5414 VSUBS 0.10fF $ **FLOATING
C5950 S.n5415 VSUBS 0.36fF $ **FLOATING
C5951 S.n5416 VSUBS 0.38fF $ **FLOATING
C5952 S.n5417 VSUBS 0.11fF $ **FLOATING
C5953 S.n5418 VSUBS 0.12fF $ **FLOATING
C5954 S.n5419 VSUBS 0.07fF $ **FLOATING
C5955 S.n5420 VSUBS 0.12fF $ **FLOATING
C5956 S.n5421 VSUBS 0.18fF $ **FLOATING
C5957 S.n5422 VSUBS 3.99fF $ **FLOATING
C5958 S.t1665 VSUBS 0.02fF
C5959 S.n5423 VSUBS 0.24fF $ **FLOATING
C5960 S.n5424 VSUBS 0.91fF $ **FLOATING
C5961 S.n5425 VSUBS 0.05fF $ **FLOATING
C5962 S.t1434 VSUBS 0.02fF
C5963 S.n5426 VSUBS 0.12fF $ **FLOATING
C5964 S.n5427 VSUBS 0.14fF $ **FLOATING
C5965 S.n5429 VSUBS 0.25fF $ **FLOATING
C5966 S.n5430 VSUBS 0.09fF $ **FLOATING
C5967 S.n5431 VSUBS 0.21fF $ **FLOATING
C5968 S.n5432 VSUBS 1.28fF $ **FLOATING
C5969 S.n5433 VSUBS 0.53fF $ **FLOATING
C5970 S.n5434 VSUBS 1.88fF $ **FLOATING
C5971 S.n5435 VSUBS 0.12fF $ **FLOATING
C5972 S.t1361 VSUBS 0.02fF
C5973 S.n5436 VSUBS 0.14fF $ **FLOATING
C5974 S.t2175 VSUBS 0.02fF
C5975 S.n5438 VSUBS 0.24fF $ **FLOATING
C5976 S.n5439 VSUBS 0.36fF $ **FLOATING
C5977 S.n5440 VSUBS 0.61fF $ **FLOATING
C5978 S.n5441 VSUBS 1.58fF $ **FLOATING
C5979 S.n5442 VSUBS 2.45fF $ **FLOATING
C5980 S.t2455 VSUBS 0.02fF
C5981 S.n5443 VSUBS 0.24fF $ **FLOATING
C5982 S.n5444 VSUBS 0.91fF $ **FLOATING
C5983 S.n5445 VSUBS 0.05fF $ **FLOATING
C5984 S.t2225 VSUBS 0.02fF
C5985 S.n5446 VSUBS 0.12fF $ **FLOATING
C5986 S.n5447 VSUBS 0.14fF $ **FLOATING
C5987 S.n5449 VSUBS 1.89fF $ **FLOATING
C5988 S.n5450 VSUBS 0.06fF $ **FLOATING
C5989 S.n5451 VSUBS 0.03fF $ **FLOATING
C5990 S.n5452 VSUBS 0.04fF $ **FLOATING
C5991 S.n5453 VSUBS 0.99fF $ **FLOATING
C5992 S.n5454 VSUBS 0.02fF $ **FLOATING
C5993 S.n5455 VSUBS 0.01fF $ **FLOATING
C5994 S.n5456 VSUBS 0.02fF $ **FLOATING
C5995 S.n5457 VSUBS 0.08fF $ **FLOATING
C5996 S.n5458 VSUBS 0.36fF $ **FLOATING
C5997 S.n5459 VSUBS 1.85fF $ **FLOATING
C5998 S.t440 VSUBS 0.02fF
C5999 S.n5460 VSUBS 0.24fF $ **FLOATING
C6000 S.n5461 VSUBS 0.36fF $ **FLOATING
C6001 S.n5462 VSUBS 0.61fF $ **FLOATING
C6002 S.n5463 VSUBS 0.12fF $ **FLOATING
C6003 S.t2147 VSUBS 0.02fF
C6004 S.n5464 VSUBS 0.14fF $ **FLOATING
C6005 S.n5466 VSUBS 0.70fF $ **FLOATING
C6006 S.n5467 VSUBS 0.23fF $ **FLOATING
C6007 S.n5468 VSUBS 0.23fF $ **FLOATING
C6008 S.n5469 VSUBS 0.70fF $ **FLOATING
C6009 S.n5470 VSUBS 1.16fF $ **FLOATING
C6010 S.n5471 VSUBS 0.22fF $ **FLOATING
C6011 S.n5472 VSUBS 0.25fF $ **FLOATING
C6012 S.n5473 VSUBS 0.09fF $ **FLOATING
C6013 S.n5474 VSUBS 1.88fF $ **FLOATING
C6014 S.t712 VSUBS 0.02fF
C6015 S.n5475 VSUBS 0.24fF $ **FLOATING
C6016 S.n5476 VSUBS 0.91fF $ **FLOATING
C6017 S.n5477 VSUBS 0.05fF $ **FLOATING
C6018 S.t493 VSUBS 0.02fF
C6019 S.n5478 VSUBS 0.12fF $ **FLOATING
C6020 S.n5479 VSUBS 0.14fF $ **FLOATING
C6021 S.n5481 VSUBS 20.78fF $ **FLOATING
C6022 S.n5482 VSUBS 0.06fF $ **FLOATING
C6023 S.n5483 VSUBS 0.20fF $ **FLOATING
C6024 S.n5484 VSUBS 0.09fF $ **FLOATING
C6025 S.n5485 VSUBS 0.21fF $ **FLOATING
C6026 S.n5486 VSUBS 0.10fF $ **FLOATING
C6027 S.n5487 VSUBS 0.30fF $ **FLOATING
C6028 S.n5488 VSUBS 0.69fF $ **FLOATING
C6029 S.n5489 VSUBS 0.45fF $ **FLOATING
C6030 S.n5490 VSUBS 2.33fF $ **FLOATING
C6031 S.n5491 VSUBS 0.12fF $ **FLOATING
C6032 S.t1421 VSUBS 0.02fF
C6033 S.n5492 VSUBS 0.14fF $ **FLOATING
C6034 S.t2239 VSUBS 0.02fF
C6035 S.n5494 VSUBS 0.24fF $ **FLOATING
C6036 S.n5495 VSUBS 0.36fF $ **FLOATING
C6037 S.n5496 VSUBS 0.61fF $ **FLOATING
C6038 S.n5497 VSUBS 1.90fF $ **FLOATING
C6039 S.n5498 VSUBS 0.17fF $ **FLOATING
C6040 S.n5499 VSUBS 0.76fF $ **FLOATING
C6041 S.n5500 VSUBS 0.32fF $ **FLOATING
C6042 S.n5501 VSUBS 0.25fF $ **FLOATING
C6043 S.n5502 VSUBS 0.30fF $ **FLOATING
C6044 S.n5503 VSUBS 0.47fF $ **FLOATING
C6045 S.n5504 VSUBS 0.16fF $ **FLOATING
C6046 S.n5505 VSUBS 1.93fF $ **FLOATING
C6047 S.t2286 VSUBS 0.02fF
C6048 S.n5506 VSUBS 0.12fF $ **FLOATING
C6049 S.n5507 VSUBS 0.14fF $ **FLOATING
C6050 S.t2519 VSUBS 0.02fF
C6051 S.n5509 VSUBS 0.24fF $ **FLOATING
C6052 S.n5510 VSUBS 0.91fF $ **FLOATING
C6053 S.n5511 VSUBS 0.05fF $ **FLOATING
C6054 S.n5512 VSUBS 1.88fF $ **FLOATING
C6055 S.n5513 VSUBS 0.12fF $ **FLOATING
C6056 S.t995 VSUBS 0.02fF
C6057 S.n5514 VSUBS 0.14fF $ **FLOATING
C6058 S.t1860 VSUBS 0.02fF
C6059 S.n5516 VSUBS 0.12fF $ **FLOATING
C6060 S.n5517 VSUBS 0.14fF $ **FLOATING
C6061 S.t2094 VSUBS 0.02fF
C6062 S.n5519 VSUBS 0.24fF $ **FLOATING
C6063 S.n5520 VSUBS 0.91fF $ **FLOATING
C6064 S.n5521 VSUBS 0.05fF $ **FLOATING
C6065 S.t1803 VSUBS 0.02fF
C6066 S.n5522 VSUBS 0.24fF $ **FLOATING
C6067 S.n5523 VSUBS 0.36fF $ **FLOATING
C6068 S.n5524 VSUBS 0.61fF $ **FLOATING
C6069 S.n5525 VSUBS 0.32fF $ **FLOATING
C6070 S.n5526 VSUBS 1.09fF $ **FLOATING
C6071 S.n5527 VSUBS 0.15fF $ **FLOATING
C6072 S.n5528 VSUBS 2.10fF $ **FLOATING
C6073 S.n5529 VSUBS 2.94fF $ **FLOATING
C6074 S.n5530 VSUBS 1.88fF $ **FLOATING
C6075 S.n5531 VSUBS 0.12fF $ **FLOATING
C6076 S.t415 VSUBS 0.02fF
C6077 S.n5532 VSUBS 0.14fF $ **FLOATING
C6078 S.t1233 VSUBS 0.02fF
C6079 S.n5534 VSUBS 0.24fF $ **FLOATING
C6080 S.n5535 VSUBS 0.36fF $ **FLOATING
C6081 S.n5536 VSUBS 0.61fF $ **FLOATING
C6082 S.n5537 VSUBS 0.92fF $ **FLOATING
C6083 S.n5538 VSUBS 0.32fF $ **FLOATING
C6084 S.n5539 VSUBS 0.92fF $ **FLOATING
C6085 S.n5540 VSUBS 1.09fF $ **FLOATING
C6086 S.n5541 VSUBS 0.15fF $ **FLOATING
C6087 S.n5542 VSUBS 4.96fF $ **FLOATING
C6088 S.t1280 VSUBS 0.02fF
C6089 S.n5543 VSUBS 0.12fF $ **FLOATING
C6090 S.n5544 VSUBS 0.14fF $ **FLOATING
C6091 S.t1505 VSUBS 0.02fF
C6092 S.n5546 VSUBS 0.24fF $ **FLOATING
C6093 S.n5547 VSUBS 0.91fF $ **FLOATING
C6094 S.n5548 VSUBS 0.05fF $ **FLOATING
C6095 S.n5549 VSUBS 1.88fF $ **FLOATING
C6096 S.n5550 VSUBS 2.67fF $ **FLOATING
C6097 S.t1743 VSUBS 0.02fF
C6098 S.n5551 VSUBS 0.24fF $ **FLOATING
C6099 S.n5552 VSUBS 0.36fF $ **FLOATING
C6100 S.n5553 VSUBS 0.61fF $ **FLOATING
C6101 S.n5554 VSUBS 0.12fF $ **FLOATING
C6102 S.t1956 VSUBS 0.02fF
C6103 S.n5555 VSUBS 0.14fF $ **FLOATING
C6104 S.n5557 VSUBS 1.88fF $ **FLOATING
C6105 S.n5558 VSUBS 2.67fF $ **FLOATING
C6106 S.t14 VSUBS 0.02fF
C6107 S.n5559 VSUBS 0.24fF $ **FLOATING
C6108 S.n5560 VSUBS 0.36fF $ **FLOATING
C6109 S.n5561 VSUBS 0.61fF $ **FLOATING
C6110 S.t367 VSUBS 0.02fF
C6111 S.n5562 VSUBS 0.24fF $ **FLOATING
C6112 S.n5563 VSUBS 0.91fF $ **FLOATING
C6113 S.n5564 VSUBS 0.05fF $ **FLOATING
C6114 S.t99 VSUBS 0.02fF
C6115 S.n5565 VSUBS 0.12fF $ **FLOATING
C6116 S.n5566 VSUBS 0.14fF $ **FLOATING
C6117 S.n5568 VSUBS 0.12fF $ **FLOATING
C6118 S.t1914 VSUBS 0.02fF
C6119 S.n5569 VSUBS 0.14fF $ **FLOATING
C6120 S.n5571 VSUBS 2.30fF $ **FLOATING
C6121 S.n5572 VSUBS 2.94fF $ **FLOATING
C6122 S.n5573 VSUBS 5.16fF $ **FLOATING
C6123 S.t2192 VSUBS 0.02fF
C6124 S.n5574 VSUBS 0.12fF $ **FLOATING
C6125 S.n5575 VSUBS 0.14fF $ **FLOATING
C6126 S.t10 VSUBS 0.02fF
C6127 S.n5577 VSUBS 0.24fF $ **FLOATING
C6128 S.n5578 VSUBS 0.91fF $ **FLOATING
C6129 S.n5579 VSUBS 0.05fF $ **FLOATING
C6130 S.n5580 VSUBS 1.88fF $ **FLOATING
C6131 S.n5581 VSUBS 2.67fF $ **FLOATING
C6132 S.t2526 VSUBS 0.02fF
C6133 S.n5582 VSUBS 0.24fF $ **FLOATING
C6134 S.n5583 VSUBS 0.36fF $ **FLOATING
C6135 S.n5584 VSUBS 0.61fF $ **FLOATING
C6136 S.n5585 VSUBS 0.12fF $ **FLOATING
C6137 S.t212 VSUBS 0.02fF
C6138 S.n5586 VSUBS 0.14fF $ **FLOATING
C6139 S.n5588 VSUBS 5.17fF $ **FLOATING
C6140 S.t1087 VSUBS 0.02fF
C6141 S.n5589 VSUBS 0.12fF $ **FLOATING
C6142 S.n5590 VSUBS 0.14fF $ **FLOATING
C6143 S.t853 VSUBS 0.02fF
C6144 S.n5592 VSUBS 0.24fF $ **FLOATING
C6145 S.n5593 VSUBS 0.91fF $ **FLOATING
C6146 S.n5594 VSUBS 0.05fF $ **FLOATING
C6147 S.n5595 VSUBS 1.88fF $ **FLOATING
C6148 S.n5596 VSUBS 0.12fF $ **FLOATING
C6149 S.t1004 VSUBS 0.02fF
C6150 S.n5597 VSUBS 0.14fF $ **FLOATING
C6151 S.t786 VSUBS 0.02fF
C6152 S.n5599 VSUBS 0.24fF $ **FLOATING
C6153 S.n5600 VSUBS 0.36fF $ **FLOATING
C6154 S.n5601 VSUBS 0.61fF $ **FLOATING
C6155 S.n5602 VSUBS 2.67fF $ **FLOATING
C6156 S.n5603 VSUBS 5.17fF $ **FLOATING
C6157 S.t1870 VSUBS 0.02fF
C6158 S.n5604 VSUBS 0.12fF $ **FLOATING
C6159 S.n5605 VSUBS 0.14fF $ **FLOATING
C6160 S.t1633 VSUBS 0.02fF
C6161 S.n5607 VSUBS 0.24fF $ **FLOATING
C6162 S.n5608 VSUBS 0.91fF $ **FLOATING
C6163 S.n5609 VSUBS 0.05fF $ **FLOATING
C6164 S.n5610 VSUBS 1.88fF $ **FLOATING
C6165 S.n5611 VSUBS 2.67fF $ **FLOATING
C6166 S.t1572 VSUBS 0.02fF
C6167 S.n5612 VSUBS 0.24fF $ **FLOATING
C6168 S.n5613 VSUBS 0.36fF $ **FLOATING
C6169 S.n5614 VSUBS 0.61fF $ **FLOATING
C6170 S.n5615 VSUBS 0.12fF $ **FLOATING
C6171 S.t1784 VSUBS 0.02fF
C6172 S.n5616 VSUBS 0.14fF $ **FLOATING
C6173 S.n5618 VSUBS 4.89fF $ **FLOATING
C6174 S.t114 VSUBS 0.02fF
C6175 S.n5619 VSUBS 0.12fF $ **FLOATING
C6176 S.n5620 VSUBS 0.14fF $ **FLOATING
C6177 S.t2418 VSUBS 0.02fF
C6178 S.n5622 VSUBS 0.24fF $ **FLOATING
C6179 S.n5623 VSUBS 0.91fF $ **FLOATING
C6180 S.n5624 VSUBS 0.05fF $ **FLOATING
C6181 S.n5625 VSUBS 1.88fF $ **FLOATING
C6182 S.n5626 VSUBS 2.67fF $ **FLOATING
C6183 S.t2363 VSUBS 0.02fF
C6184 S.n5627 VSUBS 0.24fF $ **FLOATING
C6185 S.n5628 VSUBS 0.36fF $ **FLOATING
C6186 S.n5629 VSUBS 0.61fF $ **FLOATING
C6187 S.n5630 VSUBS 0.12fF $ **FLOATING
C6188 S.t2566 VSUBS 0.02fF
C6189 S.n5631 VSUBS 0.14fF $ **FLOATING
C6190 S.n5633 VSUBS 1.88fF $ **FLOATING
C6191 S.n5634 VSUBS 2.68fF $ **FLOATING
C6192 S.t2391 VSUBS 0.02fF
C6193 S.n5635 VSUBS 0.24fF $ **FLOATING
C6194 S.n5636 VSUBS 0.36fF $ **FLOATING
C6195 S.n5637 VSUBS 0.61fF $ **FLOATING
C6196 S.t310 VSUBS 0.02fF
C6197 S.n5638 VSUBS 1.22fF $ **FLOATING
C6198 S.n5639 VSUBS 0.36fF $ **FLOATING
C6199 S.n5640 VSUBS 1.22fF $ **FLOATING
C6200 S.n5641 VSUBS 0.61fF $ **FLOATING
C6201 S.n5642 VSUBS 0.35fF $ **FLOATING
C6202 S.n5643 VSUBS 0.63fF $ **FLOATING
C6203 S.n5644 VSUBS 1.15fF $ **FLOATING
C6204 S.n5645 VSUBS 3.00fF $ **FLOATING
C6205 S.n5646 VSUBS 0.59fF $ **FLOATING
C6206 S.n5647 VSUBS 0.01fF $ **FLOATING
C6207 S.n5648 VSUBS 0.97fF $ **FLOATING
C6208 S.t13 VSUBS 21.42fF
C6209 S.n5649 VSUBS 20.29fF $ **FLOATING
C6210 S.n5651 VSUBS 0.38fF $ **FLOATING
C6211 S.n5652 VSUBS 0.23fF $ **FLOATING
C6212 S.n5653 VSUBS 2.79fF $ **FLOATING
C6213 S.n5654 VSUBS 2.46fF $ **FLOATING
C6214 S.n5655 VSUBS 4.00fF $ **FLOATING
C6215 S.n5656 VSUBS 0.25fF $ **FLOATING
C6216 S.n5657 VSUBS 0.01fF $ **FLOATING
C6217 S.t2011 VSUBS 0.02fF
C6218 S.n5658 VSUBS 0.26fF $ **FLOATING
C6219 S.t581 VSUBS 0.02fF
C6220 S.n5659 VSUBS 0.95fF $ **FLOATING
C6221 S.n5660 VSUBS 0.71fF $ **FLOATING
C6222 S.n5661 VSUBS 1.89fF $ **FLOATING
C6223 S.n5662 VSUBS 1.88fF $ **FLOATING
C6224 S.t1096 VSUBS 0.02fF
C6225 S.n5663 VSUBS 0.24fF $ **FLOATING
C6226 S.n5664 VSUBS 0.36fF $ **FLOATING
C6227 S.n5665 VSUBS 0.61fF $ **FLOATING
C6228 S.n5666 VSUBS 0.12fF $ **FLOATING
C6229 S.t284 VSUBS 0.02fF
C6230 S.n5667 VSUBS 0.14fF $ **FLOATING
C6231 S.n5669 VSUBS 1.16fF $ **FLOATING
C6232 S.n5670 VSUBS 0.22fF $ **FLOATING
C6233 S.n5671 VSUBS 0.25fF $ **FLOATING
C6234 S.n5672 VSUBS 0.09fF $ **FLOATING
C6235 S.n5673 VSUBS 1.88fF $ **FLOATING
C6236 S.t1373 VSUBS 0.02fF
C6237 S.n5674 VSUBS 0.24fF $ **FLOATING
C6238 S.n5675 VSUBS 0.91fF $ **FLOATING
C6239 S.n5676 VSUBS 0.05fF $ **FLOATING
C6240 S.t1150 VSUBS 0.02fF
C6241 S.n5677 VSUBS 0.12fF $ **FLOATING
C6242 S.n5678 VSUBS 0.14fF $ **FLOATING
C6243 S.n5680 VSUBS 0.78fF $ **FLOATING
C6244 S.n5681 VSUBS 1.94fF $ **FLOATING
C6245 S.n5682 VSUBS 1.88fF $ **FLOATING
C6246 S.n5683 VSUBS 0.12fF $ **FLOATING
C6247 S.t1196 VSUBS 0.02fF
C6248 S.n5684 VSUBS 0.14fF $ **FLOATING
C6249 S.t1877 VSUBS 0.02fF
C6250 S.n5686 VSUBS 0.24fF $ **FLOATING
C6251 S.n5687 VSUBS 0.36fF $ **FLOATING
C6252 S.n5688 VSUBS 0.61fF $ **FLOATING
C6253 S.n5689 VSUBS 1.84fF $ **FLOATING
C6254 S.n5690 VSUBS 2.99fF $ **FLOATING
C6255 S.t2162 VSUBS 0.02fF
C6256 S.n5691 VSUBS 0.24fF $ **FLOATING
C6257 S.n5692 VSUBS 0.91fF $ **FLOATING
C6258 S.n5693 VSUBS 0.05fF $ **FLOATING
C6259 S.t1933 VSUBS 0.02fF
C6260 S.n5694 VSUBS 0.12fF $ **FLOATING
C6261 S.n5695 VSUBS 0.14fF $ **FLOATING
C6262 S.n5697 VSUBS 1.89fF $ **FLOATING
C6263 S.n5698 VSUBS 1.88fF $ **FLOATING
C6264 S.t273 VSUBS 0.02fF
C6265 S.n5699 VSUBS 0.24fF $ **FLOATING
C6266 S.n5700 VSUBS 0.36fF $ **FLOATING
C6267 S.n5701 VSUBS 0.61fF $ **FLOATING
C6268 S.n5702 VSUBS 0.12fF $ **FLOATING
C6269 S.t1975 VSUBS 0.02fF
C6270 S.n5703 VSUBS 0.14fF $ **FLOATING
C6271 S.n5705 VSUBS 1.16fF $ **FLOATING
C6272 S.n5706 VSUBS 0.22fF $ **FLOATING
C6273 S.n5707 VSUBS 0.25fF $ **FLOATING
C6274 S.n5708 VSUBS 0.09fF $ **FLOATING
C6275 S.n5709 VSUBS 1.88fF $ **FLOATING
C6276 S.t550 VSUBS 0.02fF
C6277 S.n5710 VSUBS 0.24fF $ **FLOATING
C6278 S.n5711 VSUBS 0.91fF $ **FLOATING
C6279 S.n5712 VSUBS 0.05fF $ **FLOATING
C6280 S.t324 VSUBS 0.02fF
C6281 S.n5713 VSUBS 0.12fF $ **FLOATING
C6282 S.n5714 VSUBS 0.14fF $ **FLOATING
C6283 S.n5716 VSUBS 0.78fF $ **FLOATING
C6284 S.n5717 VSUBS 1.94fF $ **FLOATING
C6285 S.n5718 VSUBS 1.88fF $ **FLOATING
C6286 S.n5719 VSUBS 0.12fF $ **FLOATING
C6287 S.t1567 VSUBS 0.02fF
C6288 S.n5720 VSUBS 0.14fF $ **FLOATING
C6289 S.t2387 VSUBS 0.02fF
C6290 S.n5722 VSUBS 0.24fF $ **FLOATING
C6291 S.n5723 VSUBS 0.36fF $ **FLOATING
C6292 S.n5724 VSUBS 0.61fF $ **FLOATING
C6293 S.n5725 VSUBS 1.84fF $ **FLOATING
C6294 S.n5726 VSUBS 2.99fF $ **FLOATING
C6295 S.t152 VSUBS 0.02fF
C6296 S.n5727 VSUBS 0.24fF $ **FLOATING
C6297 S.n5728 VSUBS 0.91fF $ **FLOATING
C6298 S.n5729 VSUBS 0.05fF $ **FLOATING
C6299 S.t2439 VSUBS 0.02fF
C6300 S.n5730 VSUBS 0.12fF $ **FLOATING
C6301 S.n5731 VSUBS 0.14fF $ **FLOATING
C6302 S.n5733 VSUBS 1.89fF $ **FLOATING
C6303 S.n5734 VSUBS 1.88fF $ **FLOATING
C6304 S.t650 VSUBS 0.02fF
C6305 S.n5735 VSUBS 0.24fF $ **FLOATING
C6306 S.n5736 VSUBS 0.36fF $ **FLOATING
C6307 S.n5737 VSUBS 0.61fF $ **FLOATING
C6308 S.n5738 VSUBS 0.12fF $ **FLOATING
C6309 S.t2357 VSUBS 0.02fF
C6310 S.n5739 VSUBS 0.14fF $ **FLOATING
C6311 S.n5741 VSUBS 1.16fF $ **FLOATING
C6312 S.n5742 VSUBS 0.22fF $ **FLOATING
C6313 S.n5743 VSUBS 0.25fF $ **FLOATING
C6314 S.n5744 VSUBS 0.09fF $ **FLOATING
C6315 S.n5745 VSUBS 1.88fF $ **FLOATING
C6316 S.t944 VSUBS 0.02fF
C6317 S.n5746 VSUBS 0.24fF $ **FLOATING
C6318 S.n5747 VSUBS 0.91fF $ **FLOATING
C6319 S.n5748 VSUBS 0.05fF $ **FLOATING
C6320 S.t699 VSUBS 0.02fF
C6321 S.n5749 VSUBS 0.12fF $ **FLOATING
C6322 S.n5750 VSUBS 0.14fF $ **FLOATING
C6323 S.n5752 VSUBS 0.78fF $ **FLOATING
C6324 S.n5753 VSUBS 1.94fF $ **FLOATING
C6325 S.n5754 VSUBS 1.88fF $ **FLOATING
C6326 S.n5755 VSUBS 0.12fF $ **FLOATING
C6327 S.t627 VSUBS 0.02fF
C6328 S.n5756 VSUBS 0.14fF $ **FLOATING
C6329 S.t1442 VSUBS 0.02fF
C6330 S.n5758 VSUBS 0.24fF $ **FLOATING
C6331 S.n5759 VSUBS 0.36fF $ **FLOATING
C6332 S.n5760 VSUBS 0.61fF $ **FLOATING
C6333 S.n5761 VSUBS 1.84fF $ **FLOATING
C6334 S.n5762 VSUBS 2.99fF $ **FLOATING
C6335 S.t1729 VSUBS 0.02fF
C6336 S.n5763 VSUBS 0.24fF $ **FLOATING
C6337 S.n5764 VSUBS 0.91fF $ **FLOATING
C6338 S.n5765 VSUBS 0.05fF $ **FLOATING
C6339 S.t1494 VSUBS 0.02fF
C6340 S.n5766 VSUBS 0.12fF $ **FLOATING
C6341 S.n5767 VSUBS 0.14fF $ **FLOATING
C6342 S.n5769 VSUBS 1.89fF $ **FLOATING
C6343 S.n5770 VSUBS 1.75fF $ **FLOATING
C6344 S.t2232 VSUBS 0.02fF
C6345 S.n5771 VSUBS 0.24fF $ **FLOATING
C6346 S.n5772 VSUBS 0.36fF $ **FLOATING
C6347 S.n5773 VSUBS 0.61fF $ **FLOATING
C6348 S.n5774 VSUBS 0.12fF $ **FLOATING
C6349 S.t1537 VSUBS 0.02fF
C6350 S.n5775 VSUBS 0.14fF $ **FLOATING
C6351 S.n5777 VSUBS 1.16fF $ **FLOATING
C6352 S.n5778 VSUBS 0.22fF $ **FLOATING
C6353 S.n5779 VSUBS 0.25fF $ **FLOATING
C6354 S.n5780 VSUBS 0.09fF $ **FLOATING
C6355 S.n5781 VSUBS 2.44fF $ **FLOATING
C6356 S.t2514 VSUBS 0.02fF
C6357 S.n5782 VSUBS 0.24fF $ **FLOATING
C6358 S.n5783 VSUBS 0.91fF $ **FLOATING
C6359 S.n5784 VSUBS 0.05fF $ **FLOATING
C6360 S.t2281 VSUBS 0.02fF
C6361 S.n5785 VSUBS 0.12fF $ **FLOATING
C6362 S.n5786 VSUBS 0.14fF $ **FLOATING
C6363 S.n5788 VSUBS 1.88fF $ **FLOATING
C6364 S.n5789 VSUBS 0.48fF $ **FLOATING
C6365 S.n5790 VSUBS 0.09fF $ **FLOATING
C6366 S.n5791 VSUBS 0.33fF $ **FLOATING
C6367 S.n5792 VSUBS 0.30fF $ **FLOATING
C6368 S.n5793 VSUBS 0.77fF $ **FLOATING
C6369 S.n5794 VSUBS 0.59fF $ **FLOATING
C6370 S.t1976 VSUBS 0.02fF
C6371 S.n5795 VSUBS 0.24fF $ **FLOATING
C6372 S.n5796 VSUBS 0.36fF $ **FLOATING
C6373 S.n5797 VSUBS 0.61fF $ **FLOATING
C6374 S.n5798 VSUBS 0.12fF $ **FLOATING
C6375 S.t1163 VSUBS 0.02fF
C6376 S.n5799 VSUBS 0.14fF $ **FLOATING
C6377 S.n5801 VSUBS 2.61fF $ **FLOATING
C6378 S.n5802 VSUBS 2.15fF $ **FLOATING
C6379 S.t2252 VSUBS 0.02fF
C6380 S.n5803 VSUBS 0.24fF $ **FLOATING
C6381 S.n5804 VSUBS 0.91fF $ **FLOATING
C6382 S.n5805 VSUBS 0.05fF $ **FLOATING
C6383 S.t668 VSUBS 0.02fF
C6384 S.n5806 VSUBS 0.12fF $ **FLOATING
C6385 S.n5807 VSUBS 0.14fF $ **FLOATING
C6386 S.n5809 VSUBS 0.78fF $ **FLOATING
C6387 S.n5810 VSUBS 2.30fF $ **FLOATING
C6388 S.n5811 VSUBS 1.88fF $ **FLOATING
C6389 S.n5812 VSUBS 0.12fF $ **FLOATING
C6390 S.t1947 VSUBS 0.02fF
C6391 S.n5813 VSUBS 0.14fF $ **FLOATING
C6392 S.t239 VSUBS 0.02fF
C6393 S.n5815 VSUBS 0.24fF $ **FLOATING
C6394 S.n5816 VSUBS 0.36fF $ **FLOATING
C6395 S.n5817 VSUBS 0.61fF $ **FLOATING
C6396 S.n5818 VSUBS 1.39fF $ **FLOATING
C6397 S.n5819 VSUBS 0.71fF $ **FLOATING
C6398 S.n5820 VSUBS 1.14fF $ **FLOATING
C6399 S.n5821 VSUBS 0.35fF $ **FLOATING
C6400 S.n5822 VSUBS 2.02fF $ **FLOATING
C6401 S.t520 VSUBS 0.02fF
C6402 S.n5823 VSUBS 0.24fF $ **FLOATING
C6403 S.n5824 VSUBS 0.91fF $ **FLOATING
C6404 S.n5825 VSUBS 0.05fF $ **FLOATING
C6405 S.t297 VSUBS 0.02fF
C6406 S.n5826 VSUBS 0.12fF $ **FLOATING
C6407 S.n5827 VSUBS 0.14fF $ **FLOATING
C6408 S.n5829 VSUBS 1.89fF $ **FLOATING
C6409 S.n5830 VSUBS 1.88fF $ **FLOATING
C6410 S.t1024 VSUBS 0.02fF
C6411 S.n5831 VSUBS 0.24fF $ **FLOATING
C6412 S.n5832 VSUBS 0.36fF $ **FLOATING
C6413 S.n5833 VSUBS 0.61fF $ **FLOATING
C6414 S.n5834 VSUBS 0.12fF $ **FLOATING
C6415 S.t204 VSUBS 0.02fF
C6416 S.n5835 VSUBS 0.14fF $ **FLOATING
C6417 S.n5837 VSUBS 1.16fF $ **FLOATING
C6418 S.n5838 VSUBS 0.22fF $ **FLOATING
C6419 S.n5839 VSUBS 0.25fF $ **FLOATING
C6420 S.n5840 VSUBS 0.09fF $ **FLOATING
C6421 S.n5841 VSUBS 1.88fF $ **FLOATING
C6422 S.t1307 VSUBS 0.02fF
C6423 S.n5842 VSUBS 0.24fF $ **FLOATING
C6424 S.n5843 VSUBS 0.91fF $ **FLOATING
C6425 S.n5844 VSUBS 0.05fF $ **FLOATING
C6426 S.t1079 VSUBS 0.02fF
C6427 S.n5845 VSUBS 0.12fF $ **FLOATING
C6428 S.n5846 VSUBS 0.14fF $ **FLOATING
C6429 S.n5848 VSUBS 20.78fF $ **FLOATING
C6430 S.n5849 VSUBS 1.88fF $ **FLOATING
C6431 S.n5850 VSUBS 2.67fF $ **FLOATING
C6432 S.t2555 VSUBS 0.02fF
C6433 S.n5851 VSUBS 0.24fF $ **FLOATING
C6434 S.n5852 VSUBS 0.36fF $ **FLOATING
C6435 S.n5853 VSUBS 0.61fF $ **FLOATING
C6436 S.n5854 VSUBS 0.12fF $ **FLOATING
C6437 S.t247 VSUBS 0.02fF
C6438 S.n5855 VSUBS 0.14fF $ **FLOATING
C6439 S.n5857 VSUBS 2.80fF $ **FLOATING
C6440 S.n5858 VSUBS 2.30fF $ **FLOATING
C6441 S.t1117 VSUBS 0.02fF
C6442 S.n5859 VSUBS 0.12fF $ **FLOATING
C6443 S.n5860 VSUBS 0.14fF $ **FLOATING
C6444 S.t876 VSUBS 0.02fF
C6445 S.n5862 VSUBS 0.24fF $ **FLOATING
C6446 S.n5863 VSUBS 0.91fF $ **FLOATING
C6447 S.n5864 VSUBS 0.05fF $ **FLOATING
C6448 S.n5865 VSUBS 2.80fF $ **FLOATING
C6449 S.n5866 VSUBS 1.88fF $ **FLOATING
C6450 S.n5867 VSUBS 0.12fF $ **FLOATING
C6451 S.t1031 VSUBS 0.02fF
C6452 S.n5868 VSUBS 0.14fF $ **FLOATING
C6453 S.t818 VSUBS 0.02fF
C6454 S.n5870 VSUBS 0.24fF $ **FLOATING
C6455 S.n5871 VSUBS 0.36fF $ **FLOATING
C6456 S.n5872 VSUBS 0.61fF $ **FLOATING
C6457 S.n5873 VSUBS 2.67fF $ **FLOATING
C6458 S.n5874 VSUBS 2.30fF $ **FLOATING
C6459 S.t1898 VSUBS 0.02fF
C6460 S.n5875 VSUBS 0.12fF $ **FLOATING
C6461 S.n5876 VSUBS 0.14fF $ **FLOATING
C6462 S.t1657 VSUBS 0.02fF
C6463 S.n5878 VSUBS 0.24fF $ **FLOATING
C6464 S.n5879 VSUBS 0.91fF $ **FLOATING
C6465 S.n5880 VSUBS 0.05fF $ **FLOATING
C6466 S.n5881 VSUBS 1.88fF $ **FLOATING
C6467 S.n5882 VSUBS 2.67fF $ **FLOATING
C6468 S.t1599 VSUBS 0.02fF
C6469 S.n5883 VSUBS 0.24fF $ **FLOATING
C6470 S.n5884 VSUBS 0.36fF $ **FLOATING
C6471 S.n5885 VSUBS 0.61fF $ **FLOATING
C6472 S.n5886 VSUBS 0.12fF $ **FLOATING
C6473 S.t1810 VSUBS 0.02fF
C6474 S.n5887 VSUBS 0.14fF $ **FLOATING
C6475 S.n5889 VSUBS 2.80fF $ **FLOATING
C6476 S.n5890 VSUBS 2.30fF $ **FLOATING
C6477 S.t150 VSUBS 0.02fF
C6478 S.n5891 VSUBS 0.12fF $ **FLOATING
C6479 S.n5892 VSUBS 0.14fF $ **FLOATING
C6480 S.t2441 VSUBS 0.02fF
C6481 S.n5894 VSUBS 0.24fF $ **FLOATING
C6482 S.n5895 VSUBS 0.91fF $ **FLOATING
C6483 S.n5896 VSUBS 0.05fF $ **FLOATING
C6484 S.n5897 VSUBS 2.73fF $ **FLOATING
C6485 S.n5898 VSUBS 1.59fF $ **FLOATING
C6486 S.n5899 VSUBS 0.12fF $ **FLOATING
C6487 S.t338 VSUBS 0.02fF
C6488 S.n5900 VSUBS 0.14fF $ **FLOATING
C6489 S.t1863 VSUBS 0.02fF
C6490 S.n5902 VSUBS 0.24fF $ **FLOATING
C6491 S.n5903 VSUBS 0.36fF $ **FLOATING
C6492 S.n5904 VSUBS 0.61fF $ **FLOATING
C6493 S.n5905 VSUBS 0.07fF $ **FLOATING
C6494 S.n5906 VSUBS 0.01fF $ **FLOATING
C6495 S.n5907 VSUBS 0.24fF $ **FLOATING
C6496 S.n5908 VSUBS 1.16fF $ **FLOATING
C6497 S.n5909 VSUBS 1.35fF $ **FLOATING
C6498 S.n5910 VSUBS 2.30fF $ **FLOATING
C6499 S.t1725 VSUBS 0.02fF
C6500 S.n5911 VSUBS 0.12fF $ **FLOATING
C6501 S.n5912 VSUBS 0.14fF $ **FLOATING
C6502 S.t727 VSUBS 0.02fF
C6503 S.n5914 VSUBS 0.24fF $ **FLOATING
C6504 S.n5915 VSUBS 0.91fF $ **FLOATING
C6505 S.n5916 VSUBS 0.05fF $ **FLOATING
C6506 S.t25 VSUBS 48.27fF
C6507 S.t704 VSUBS 0.02fF
C6508 S.n5917 VSUBS 0.24fF $ **FLOATING
C6509 S.n5918 VSUBS 0.91fF $ **FLOATING
C6510 S.n5919 VSUBS 0.05fF $ **FLOATING
C6511 S.t943 VSUBS 0.02fF
C6512 S.n5920 VSUBS 0.12fF $ **FLOATING
C6513 S.n5921 VSUBS 0.14fF $ **FLOATING
C6514 S.n5923 VSUBS 0.12fF $ **FLOATING
C6515 S.t26 VSUBS 0.02fF
C6516 S.n5924 VSUBS 0.14fF $ **FLOATING
C6517 S.n5926 VSUBS 5.17fF $ **FLOATING
C6518 S.n5927 VSUBS 5.44fF $ **FLOATING
C6519 S.t917 VSUBS 0.02fF
C6520 S.n5928 VSUBS 0.12fF $ **FLOATING
C6521 S.n5929 VSUBS 0.14fF $ **FLOATING
C6522 S.t682 VSUBS 0.02fF
C6523 S.n5931 VSUBS 0.24fF $ **FLOATING
C6524 S.n5932 VSUBS 0.91fF $ **FLOATING
C6525 S.n5933 VSUBS 0.05fF $ **FLOATING
C6526 S.t109 VSUBS 47.89fF
C6527 S.t1688 VSUBS 0.02fF
C6528 S.n5934 VSUBS 0.01fF $ **FLOATING
C6529 S.n5935 VSUBS 0.26fF $ **FLOATING
C6530 S.t878 VSUBS 0.02fF
C6531 S.n5937 VSUBS 1.19fF $ **FLOATING
C6532 S.n5938 VSUBS 0.05fF $ **FLOATING
C6533 S.t591 VSUBS 0.02fF
C6534 S.n5939 VSUBS 0.64fF $ **FLOATING
C6535 S.n5940 VSUBS 0.61fF $ **FLOATING
C6536 S.n5941 VSUBS 8.97fF $ **FLOATING
C6537 S.n5942 VSUBS 8.97fF $ **FLOATING
C6538 S.n5943 VSUBS 0.60fF $ **FLOATING
C6539 S.n5944 VSUBS 0.22fF $ **FLOATING
C6540 S.n5945 VSUBS 0.59fF $ **FLOATING
C6541 S.n5946 VSUBS 3.39fF $ **FLOATING
C6542 S.n5947 VSUBS 0.29fF $ **FLOATING
C6543 S.t29 VSUBS 21.42fF
C6544 S.n5948 VSUBS 21.71fF $ **FLOATING
C6545 S.n5949 VSUBS 0.77fF $ **FLOATING
C6546 S.n5950 VSUBS 0.28fF $ **FLOATING
C6547 S.n5951 VSUBS 4.00fF $ **FLOATING
C6548 S.n5952 VSUBS 1.35fF $ **FLOATING
C6549 S.n5953 VSUBS 0.01fF $ **FLOATING
C6550 S.n5954 VSUBS 0.02fF $ **FLOATING
C6551 S.n5955 VSUBS 0.03fF $ **FLOATING
C6552 S.n5956 VSUBS 0.04fF $ **FLOATING
C6553 S.n5957 VSUBS 0.17fF $ **FLOATING
C6554 S.n5958 VSUBS 0.01fF $ **FLOATING
C6555 S.n5959 VSUBS 0.02fF $ **FLOATING
C6556 S.n5960 VSUBS 0.01fF $ **FLOATING
C6557 S.n5961 VSUBS 0.01fF $ **FLOATING
C6558 S.n5962 VSUBS 0.01fF $ **FLOATING
C6559 S.n5963 VSUBS 0.01fF $ **FLOATING
C6560 S.n5964 VSUBS 0.02fF $ **FLOATING
C6561 S.n5965 VSUBS 0.01fF $ **FLOATING
C6562 S.n5966 VSUBS 0.02fF $ **FLOATING
C6563 S.n5967 VSUBS 0.05fF $ **FLOATING
C6564 S.n5968 VSUBS 0.04fF $ **FLOATING
C6565 S.n5969 VSUBS 0.11fF $ **FLOATING
C6566 S.n5970 VSUBS 0.38fF $ **FLOATING
C6567 S.n5971 VSUBS 0.20fF $ **FLOATING
C6568 S.n5972 VSUBS 4.39fF $ **FLOATING
C6569 S.n5973 VSUBS 0.24fF $ **FLOATING
C6570 S.n5974 VSUBS 1.50fF $ **FLOATING
C6571 S.n5975 VSUBS 1.31fF $ **FLOATING
C6572 S.n5976 VSUBS 0.28fF $ **FLOATING
C6573 S.n5977 VSUBS 0.25fF $ **FLOATING
C6574 S.n5978 VSUBS 0.09fF $ **FLOATING
C6575 S.n5979 VSUBS 0.21fF $ **FLOATING
C6576 S.n5980 VSUBS 0.92fF $ **FLOATING
C6577 S.n5981 VSUBS 0.44fF $ **FLOATING
C6578 S.n5982 VSUBS 1.88fF $ **FLOATING
C6579 S.n5983 VSUBS 0.12fF $ **FLOATING
C6580 S.t1631 VSUBS 0.02fF
C6581 S.n5984 VSUBS 0.14fF $ **FLOATING
C6582 S.t2170 VSUBS 0.02fF
C6583 S.n5986 VSUBS 0.24fF $ **FLOATING
C6584 S.n5987 VSUBS 0.36fF $ **FLOATING
C6585 S.n5988 VSUBS 0.61fF $ **FLOATING
C6586 S.n5989 VSUBS 0.02fF $ **FLOATING
C6587 S.n5990 VSUBS 0.01fF $ **FLOATING
C6588 S.n5991 VSUBS 0.02fF $ **FLOATING
C6589 S.n5992 VSUBS 0.08fF $ **FLOATING
C6590 S.n5993 VSUBS 0.06fF $ **FLOATING
C6591 S.n5994 VSUBS 0.03fF $ **FLOATING
C6592 S.n5995 VSUBS 0.04fF $ **FLOATING
C6593 S.n5996 VSUBS 1.00fF $ **FLOATING
C6594 S.n5997 VSUBS 0.36fF $ **FLOATING
C6595 S.n5998 VSUBS 1.87fF $ **FLOATING
C6596 S.n5999 VSUBS 1.99fF $ **FLOATING
C6597 S.t221 VSUBS 0.02fF
C6598 S.n6000 VSUBS 0.24fF $ **FLOATING
C6599 S.n6001 VSUBS 0.91fF $ **FLOATING
C6600 S.n6002 VSUBS 0.05fF $ **FLOATING
C6601 S.t2503 VSUBS 0.02fF
C6602 S.n6003 VSUBS 0.12fF $ **FLOATING
C6603 S.n6004 VSUBS 0.14fF $ **FLOATING
C6604 S.n6006 VSUBS 1.89fF $ **FLOATING
C6605 S.n6007 VSUBS 0.06fF $ **FLOATING
C6606 S.n6008 VSUBS 0.03fF $ **FLOATING
C6607 S.n6009 VSUBS 0.04fF $ **FLOATING
C6608 S.n6010 VSUBS 0.99fF $ **FLOATING
C6609 S.n6011 VSUBS 0.02fF $ **FLOATING
C6610 S.n6012 VSUBS 0.01fF $ **FLOATING
C6611 S.n6013 VSUBS 0.02fF $ **FLOATING
C6612 S.n6014 VSUBS 0.08fF $ **FLOATING
C6613 S.n6015 VSUBS 0.36fF $ **FLOATING
C6614 S.n6016 VSUBS 1.85fF $ **FLOATING
C6615 S.t560 VSUBS 0.02fF
C6616 S.n6017 VSUBS 0.24fF $ **FLOATING
C6617 S.n6018 VSUBS 0.36fF $ **FLOATING
C6618 S.n6019 VSUBS 0.61fF $ **FLOATING
C6619 S.n6020 VSUBS 0.12fF $ **FLOATING
C6620 S.t2545 VSUBS 0.02fF
C6621 S.n6021 VSUBS 0.14fF $ **FLOATING
C6622 S.n6023 VSUBS 0.70fF $ **FLOATING
C6623 S.n6024 VSUBS 0.23fF $ **FLOATING
C6624 S.n6025 VSUBS 0.23fF $ **FLOATING
C6625 S.n6026 VSUBS 0.70fF $ **FLOATING
C6626 S.n6027 VSUBS 1.16fF $ **FLOATING
C6627 S.n6028 VSUBS 0.22fF $ **FLOATING
C6628 S.n6029 VSUBS 0.25fF $ **FLOATING
C6629 S.n6030 VSUBS 0.09fF $ **FLOATING
C6630 S.n6031 VSUBS 1.88fF $ **FLOATING
C6631 S.t1142 VSUBS 0.02fF
C6632 S.n6032 VSUBS 0.24fF $ **FLOATING
C6633 S.n6033 VSUBS 0.91fF $ **FLOATING
C6634 S.n6034 VSUBS 0.05fF $ **FLOATING
C6635 S.t898 VSUBS 0.02fF
C6636 S.n6035 VSUBS 0.12fF $ **FLOATING
C6637 S.n6036 VSUBS 0.14fF $ **FLOATING
C6638 S.n6038 VSUBS 0.25fF $ **FLOATING
C6639 S.n6039 VSUBS 0.09fF $ **FLOATING
C6640 S.n6040 VSUBS 0.21fF $ **FLOATING
C6641 S.n6041 VSUBS 0.92fF $ **FLOATING
C6642 S.n6042 VSUBS 0.44fF $ **FLOATING
C6643 S.n6043 VSUBS 1.88fF $ **FLOATING
C6644 S.n6044 VSUBS 0.12fF $ **FLOATING
C6645 S.t2165 VSUBS 0.02fF
C6646 S.n6045 VSUBS 0.14fF $ **FLOATING
C6647 S.t169 VSUBS 0.02fF
C6648 S.n6047 VSUBS 0.24fF $ **FLOATING
C6649 S.n6048 VSUBS 0.36fF $ **FLOATING
C6650 S.n6049 VSUBS 0.61fF $ **FLOATING
C6651 S.n6050 VSUBS 0.02fF $ **FLOATING
C6652 S.n6051 VSUBS 0.01fF $ **FLOATING
C6653 S.n6052 VSUBS 0.02fF $ **FLOATING
C6654 S.n6053 VSUBS 0.08fF $ **FLOATING
C6655 S.n6054 VSUBS 0.06fF $ **FLOATING
C6656 S.n6055 VSUBS 0.03fF $ **FLOATING
C6657 S.n6056 VSUBS 0.04fF $ **FLOATING
C6658 S.n6057 VSUBS 1.00fF $ **FLOATING
C6659 S.n6058 VSUBS 0.36fF $ **FLOATING
C6660 S.n6059 VSUBS 1.87fF $ **FLOATING
C6661 S.n6060 VSUBS 1.99fF $ **FLOATING
C6662 S.t728 VSUBS 0.02fF
C6663 S.n6061 VSUBS 0.24fF $ **FLOATING
C6664 S.n6062 VSUBS 0.91fF $ **FLOATING
C6665 S.n6063 VSUBS 0.05fF $ **FLOATING
C6666 S.t1677 VSUBS 0.02fF
C6667 S.n6064 VSUBS 0.12fF $ **FLOATING
C6668 S.n6065 VSUBS 0.14fF $ **FLOATING
C6669 S.n6067 VSUBS 1.89fF $ **FLOATING
C6670 S.n6068 VSUBS 0.06fF $ **FLOATING
C6671 S.n6069 VSUBS 0.03fF $ **FLOATING
C6672 S.n6070 VSUBS 0.04fF $ **FLOATING
C6673 S.n6071 VSUBS 0.99fF $ **FLOATING
C6674 S.n6072 VSUBS 0.02fF $ **FLOATING
C6675 S.n6073 VSUBS 0.01fF $ **FLOATING
C6676 S.n6074 VSUBS 0.02fF $ **FLOATING
C6677 S.n6075 VSUBS 0.08fF $ **FLOATING
C6678 S.n6076 VSUBS 0.36fF $ **FLOATING
C6679 S.n6077 VSUBS 1.85fF $ **FLOATING
C6680 S.t955 VSUBS 0.02fF
C6681 S.n6078 VSUBS 0.24fF $ **FLOATING
C6682 S.n6079 VSUBS 0.36fF $ **FLOATING
C6683 S.n6080 VSUBS 0.61fF $ **FLOATING
C6684 S.n6081 VSUBS 0.12fF $ **FLOATING
C6685 S.t431 VSUBS 0.02fF
C6686 S.n6082 VSUBS 0.14fF $ **FLOATING
C6687 S.n6084 VSUBS 0.70fF $ **FLOATING
C6688 S.n6085 VSUBS 0.23fF $ **FLOATING
C6689 S.n6086 VSUBS 0.23fF $ **FLOATING
C6690 S.n6087 VSUBS 0.70fF $ **FLOATING
C6691 S.n6088 VSUBS 1.16fF $ **FLOATING
C6692 S.n6089 VSUBS 0.22fF $ **FLOATING
C6693 S.n6090 VSUBS 0.25fF $ **FLOATING
C6694 S.n6091 VSUBS 0.09fF $ **FLOATING
C6695 S.n6092 VSUBS 1.88fF $ **FLOATING
C6696 S.t1519 VSUBS 0.02fF
C6697 S.n6093 VSUBS 0.24fF $ **FLOATING
C6698 S.n6094 VSUBS 0.91fF $ **FLOATING
C6699 S.n6095 VSUBS 0.05fF $ **FLOATING
C6700 S.t1297 VSUBS 0.02fF
C6701 S.n6096 VSUBS 0.12fF $ **FLOATING
C6702 S.n6097 VSUBS 0.14fF $ **FLOATING
C6703 S.n6099 VSUBS 0.25fF $ **FLOATING
C6704 S.n6100 VSUBS 0.09fF $ **FLOATING
C6705 S.n6101 VSUBS 0.21fF $ **FLOATING
C6706 S.n6102 VSUBS 0.92fF $ **FLOATING
C6707 S.n6103 VSUBS 0.44fF $ **FLOATING
C6708 S.n6104 VSUBS 1.88fF $ **FLOATING
C6709 S.n6105 VSUBS 0.12fF $ **FLOATING
C6710 S.t1226 VSUBS 0.02fF
C6711 S.n6106 VSUBS 0.14fF $ **FLOATING
C6712 S.t1738 VSUBS 0.02fF
C6713 S.n6108 VSUBS 0.24fF $ **FLOATING
C6714 S.n6109 VSUBS 0.36fF $ **FLOATING
C6715 S.n6110 VSUBS 0.61fF $ **FLOATING
C6716 S.n6111 VSUBS 0.02fF $ **FLOATING
C6717 S.n6112 VSUBS 0.01fF $ **FLOATING
C6718 S.n6113 VSUBS 0.02fF $ **FLOATING
C6719 S.n6114 VSUBS 0.08fF $ **FLOATING
C6720 S.n6115 VSUBS 0.06fF $ **FLOATING
C6721 S.n6116 VSUBS 0.03fF $ **FLOATING
C6722 S.n6117 VSUBS 0.04fF $ **FLOATING
C6723 S.n6118 VSUBS 1.00fF $ **FLOATING
C6724 S.n6119 VSUBS 0.36fF $ **FLOATING
C6725 S.n6120 VSUBS 1.87fF $ **FLOATING
C6726 S.n6121 VSUBS 1.99fF $ **FLOATING
C6727 S.t2307 VSUBS 0.02fF
C6728 S.n6122 VSUBS 0.24fF $ **FLOATING
C6729 S.n6123 VSUBS 0.91fF $ **FLOATING
C6730 S.n6124 VSUBS 0.05fF $ **FLOATING
C6731 S.t2084 VSUBS 0.02fF
C6732 S.n6125 VSUBS 0.12fF $ **FLOATING
C6733 S.n6126 VSUBS 0.14fF $ **FLOATING
C6734 S.n6128 VSUBS 1.89fF $ **FLOATING
C6735 S.n6129 VSUBS 0.07fF $ **FLOATING
C6736 S.n6130 VSUBS 0.04fF $ **FLOATING
C6737 S.n6131 VSUBS 0.05fF $ **FLOATING
C6738 S.n6132 VSUBS 0.87fF $ **FLOATING
C6739 S.n6133 VSUBS 0.01fF $ **FLOATING
C6740 S.n6134 VSUBS 0.01fF $ **FLOATING
C6741 S.n6135 VSUBS 0.01fF $ **FLOATING
C6742 S.n6136 VSUBS 0.07fF $ **FLOATING
C6743 S.n6137 VSUBS 0.68fF $ **FLOATING
C6744 S.n6138 VSUBS 0.72fF $ **FLOATING
C6745 S.t2522 VSUBS 0.02fF
C6746 S.n6139 VSUBS 0.24fF $ **FLOATING
C6747 S.n6140 VSUBS 0.36fF $ **FLOATING
C6748 S.n6141 VSUBS 0.61fF $ **FLOATING
C6749 S.n6142 VSUBS 0.12fF $ **FLOATING
C6750 S.t2004 VSUBS 0.02fF
C6751 S.n6143 VSUBS 0.14fF $ **FLOATING
C6752 S.n6145 VSUBS 0.70fF $ **FLOATING
C6753 S.n6146 VSUBS 0.23fF $ **FLOATING
C6754 S.n6147 VSUBS 0.23fF $ **FLOATING
C6755 S.n6148 VSUBS 0.70fF $ **FLOATING
C6756 S.n6149 VSUBS 1.16fF $ **FLOATING
C6757 S.n6150 VSUBS 0.22fF $ **FLOATING
C6758 S.n6151 VSUBS 0.25fF $ **FLOATING
C6759 S.n6152 VSUBS 0.09fF $ **FLOATING
C6760 S.n6153 VSUBS 2.31fF $ **FLOATING
C6761 S.t578 VSUBS 0.02fF
C6762 S.n6154 VSUBS 0.24fF $ **FLOATING
C6763 S.n6155 VSUBS 0.91fF $ **FLOATING
C6764 S.n6156 VSUBS 0.05fF $ **FLOATING
C6765 S.t356 VSUBS 0.02fF
C6766 S.n6157 VSUBS 0.12fF $ **FLOATING
C6767 S.n6158 VSUBS 0.14fF $ **FLOATING
C6768 S.n6160 VSUBS 1.88fF $ **FLOATING
C6769 S.n6161 VSUBS 0.46fF $ **FLOATING
C6770 S.n6162 VSUBS 0.22fF $ **FLOATING
C6771 S.n6163 VSUBS 0.38fF $ **FLOATING
C6772 S.n6164 VSUBS 0.16fF $ **FLOATING
C6773 S.n6165 VSUBS 0.28fF $ **FLOATING
C6774 S.n6166 VSUBS 0.21fF $ **FLOATING
C6775 S.n6167 VSUBS 0.30fF $ **FLOATING
C6776 S.n6168 VSUBS 0.42fF $ **FLOATING
C6777 S.n6169 VSUBS 0.21fF $ **FLOATING
C6778 S.t920 VSUBS 0.02fF
C6779 S.n6170 VSUBS 0.24fF $ **FLOATING
C6780 S.n6171 VSUBS 0.36fF $ **FLOATING
C6781 S.n6172 VSUBS 0.61fF $ **FLOATING
C6782 S.n6173 VSUBS 0.12fF $ **FLOATING
C6783 S.t396 VSUBS 0.02fF
C6784 S.n6174 VSUBS 0.14fF $ **FLOATING
C6785 S.n6176 VSUBS 0.04fF $ **FLOATING
C6786 S.n6177 VSUBS 0.03fF $ **FLOATING
C6787 S.n6178 VSUBS 0.03fF $ **FLOATING
C6788 S.n6179 VSUBS 0.10fF $ **FLOATING
C6789 S.n6180 VSUBS 0.36fF $ **FLOATING
C6790 S.n6181 VSUBS 0.38fF $ **FLOATING
C6791 S.n6182 VSUBS 0.11fF $ **FLOATING
C6792 S.n6183 VSUBS 0.12fF $ **FLOATING
C6793 S.n6184 VSUBS 0.07fF $ **FLOATING
C6794 S.n6185 VSUBS 0.12fF $ **FLOATING
C6795 S.n6186 VSUBS 0.18fF $ **FLOATING
C6796 S.n6187 VSUBS 3.99fF $ **FLOATING
C6797 S.t1487 VSUBS 0.02fF
C6798 S.n6188 VSUBS 0.24fF $ **FLOATING
C6799 S.n6189 VSUBS 0.91fF $ **FLOATING
C6800 S.n6190 VSUBS 0.05fF $ **FLOATING
C6801 S.t1262 VSUBS 0.02fF
C6802 S.n6191 VSUBS 0.12fF $ **FLOATING
C6803 S.n6192 VSUBS 0.14fF $ **FLOATING
C6804 S.n6194 VSUBS 0.25fF $ **FLOATING
C6805 S.n6195 VSUBS 0.09fF $ **FLOATING
C6806 S.n6196 VSUBS 0.21fF $ **FLOATING
C6807 S.n6197 VSUBS 1.28fF $ **FLOATING
C6808 S.n6198 VSUBS 0.53fF $ **FLOATING
C6809 S.n6199 VSUBS 1.88fF $ **FLOATING
C6810 S.n6200 VSUBS 0.12fF $ **FLOATING
C6811 S.t2518 VSUBS 0.02fF
C6812 S.n6201 VSUBS 0.14fF $ **FLOATING
C6813 S.t532 VSUBS 0.02fF
C6814 S.n6203 VSUBS 0.24fF $ **FLOATING
C6815 S.n6204 VSUBS 0.36fF $ **FLOATING
C6816 S.n6205 VSUBS 0.61fF $ **FLOATING
C6817 S.n6206 VSUBS 1.58fF $ **FLOATING
C6818 S.n6207 VSUBS 2.45fF $ **FLOATING
C6819 S.t1112 VSUBS 0.02fF
C6820 S.n6208 VSUBS 0.24fF $ **FLOATING
C6821 S.n6209 VSUBS 0.91fF $ **FLOATING
C6822 S.n6210 VSUBS 0.05fF $ **FLOATING
C6823 S.t864 VSUBS 0.02fF
C6824 S.n6211 VSUBS 0.12fF $ **FLOATING
C6825 S.n6212 VSUBS 0.14fF $ **FLOATING
C6826 S.n6214 VSUBS 1.89fF $ **FLOATING
C6827 S.n6215 VSUBS 0.06fF $ **FLOATING
C6828 S.n6216 VSUBS 0.03fF $ **FLOATING
C6829 S.n6217 VSUBS 0.04fF $ **FLOATING
C6830 S.n6218 VSUBS 0.99fF $ **FLOATING
C6831 S.n6219 VSUBS 0.02fF $ **FLOATING
C6832 S.n6220 VSUBS 0.01fF $ **FLOATING
C6833 S.n6221 VSUBS 0.02fF $ **FLOATING
C6834 S.n6222 VSUBS 0.08fF $ **FLOATING
C6835 S.n6223 VSUBS 0.36fF $ **FLOATING
C6836 S.n6224 VSUBS 1.85fF $ **FLOATING
C6837 S.t1318 VSUBS 0.02fF
C6838 S.n6225 VSUBS 0.24fF $ **FLOATING
C6839 S.n6226 VSUBS 0.36fF $ **FLOATING
C6840 S.n6227 VSUBS 0.61fF $ **FLOATING
C6841 S.n6228 VSUBS 0.12fF $ **FLOATING
C6842 S.t777 VSUBS 0.02fF
C6843 S.n6229 VSUBS 0.14fF $ **FLOATING
C6844 S.n6231 VSUBS 0.70fF $ **FLOATING
C6845 S.n6232 VSUBS 0.23fF $ **FLOATING
C6846 S.n6233 VSUBS 0.23fF $ **FLOATING
C6847 S.n6234 VSUBS 0.70fF $ **FLOATING
C6848 S.n6235 VSUBS 1.16fF $ **FLOATING
C6849 S.n6236 VSUBS 0.22fF $ **FLOATING
C6850 S.n6237 VSUBS 0.25fF $ **FLOATING
C6851 S.n6238 VSUBS 0.09fF $ **FLOATING
C6852 S.n6239 VSUBS 1.88fF $ **FLOATING
C6853 S.t1892 VSUBS 0.02fF
C6854 S.n6240 VSUBS 0.24fF $ **FLOATING
C6855 S.n6241 VSUBS 0.91fF $ **FLOATING
C6856 S.n6242 VSUBS 0.05fF $ **FLOATING
C6857 S.t1647 VSUBS 0.02fF
C6858 S.n6243 VSUBS 0.12fF $ **FLOATING
C6859 S.n6244 VSUBS 0.14fF $ **FLOATING
C6860 S.n6246 VSUBS 20.78fF $ **FLOATING
C6861 S.n6247 VSUBS 1.72fF $ **FLOATING
C6862 S.n6248 VSUBS 3.05fF $ **FLOATING
C6863 S.t1385 VSUBS 0.02fF
C6864 S.n6249 VSUBS 0.24fF $ **FLOATING
C6865 S.n6250 VSUBS 0.36fF $ **FLOATING
C6866 S.n6251 VSUBS 0.61fF $ **FLOATING
C6867 S.n6252 VSUBS 0.12fF $ **FLOATING
C6868 S.t848 VSUBS 0.02fF
C6869 S.n6253 VSUBS 0.14fF $ **FLOATING
C6870 S.n6255 VSUBS 0.31fF $ **FLOATING
C6871 S.n6256 VSUBS 0.23fF $ **FLOATING
C6872 S.n6257 VSUBS 0.66fF $ **FLOATING
C6873 S.n6258 VSUBS 0.95fF $ **FLOATING
C6874 S.n6259 VSUBS 0.23fF $ **FLOATING
C6875 S.n6260 VSUBS 0.21fF $ **FLOATING
C6876 S.n6261 VSUBS 0.20fF $ **FLOATING
C6877 S.n6262 VSUBS 0.06fF $ **FLOATING
C6878 S.n6263 VSUBS 0.09fF $ **FLOATING
C6879 S.n6264 VSUBS 0.10fF $ **FLOATING
C6880 S.n6265 VSUBS 1.99fF $ **FLOATING
C6881 S.t1716 VSUBS 0.02fF
C6882 S.n6266 VSUBS 0.12fF $ **FLOATING
C6883 S.n6267 VSUBS 0.14fF $ **FLOATING
C6884 S.t1963 VSUBS 0.02fF
C6885 S.n6269 VSUBS 0.24fF $ **FLOATING
C6886 S.n6270 VSUBS 0.91fF $ **FLOATING
C6887 S.n6271 VSUBS 0.05fF $ **FLOATING
C6888 S.n6272 VSUBS 1.88fF $ **FLOATING
C6889 S.n6273 VSUBS 0.12fF $ **FLOATING
C6890 S.t430 VSUBS 0.02fF
C6891 S.n6274 VSUBS 0.14fF $ **FLOATING
C6892 S.t1295 VSUBS 0.02fF
C6893 S.n6276 VSUBS 0.12fF $ **FLOATING
C6894 S.n6277 VSUBS 0.14fF $ **FLOATING
C6895 S.t451 VSUBS 0.02fF
C6896 S.n6279 VSUBS 0.24fF $ **FLOATING
C6897 S.n6280 VSUBS 0.91fF $ **FLOATING
C6898 S.n6281 VSUBS 0.05fF $ **FLOATING
C6899 S.t1246 VSUBS 0.02fF
C6900 S.n6282 VSUBS 0.24fF $ **FLOATING
C6901 S.n6283 VSUBS 0.36fF $ **FLOATING
C6902 S.n6284 VSUBS 0.61fF $ **FLOATING
C6903 S.n6285 VSUBS 0.32fF $ **FLOATING
C6904 S.n6286 VSUBS 1.09fF $ **FLOATING
C6905 S.n6287 VSUBS 0.15fF $ **FLOATING
C6906 S.n6288 VSUBS 2.10fF $ **FLOATING
C6907 S.n6289 VSUBS 2.94fF $ **FLOATING
C6908 S.n6290 VSUBS 1.88fF $ **FLOATING
C6909 S.n6291 VSUBS 0.12fF $ **FLOATING
C6910 S.t1562 VSUBS 0.02fF
C6911 S.n6292 VSUBS 0.14fF $ **FLOATING
C6912 S.t2107 VSUBS 0.02fF
C6913 S.n6294 VSUBS 0.24fF $ **FLOATING
C6914 S.n6295 VSUBS 0.36fF $ **FLOATING
C6915 S.n6296 VSUBS 0.61fF $ **FLOATING
C6916 S.n6297 VSUBS 0.92fF $ **FLOATING
C6917 S.n6298 VSUBS 0.32fF $ **FLOATING
C6918 S.n6299 VSUBS 0.92fF $ **FLOATING
C6919 S.n6300 VSUBS 1.09fF $ **FLOATING
C6920 S.n6301 VSUBS 0.15fF $ **FLOATING
C6921 S.n6302 VSUBS 4.96fF $ **FLOATING
C6922 S.t2431 VSUBS 0.02fF
C6923 S.n6303 VSUBS 0.12fF $ **FLOATING
C6924 S.n6304 VSUBS 0.14fF $ **FLOATING
C6925 S.t141 VSUBS 0.02fF
C6926 S.n6306 VSUBS 0.24fF $ **FLOATING
C6927 S.n6307 VSUBS 0.91fF $ **FLOATING
C6928 S.n6308 VSUBS 0.05fF $ **FLOATING
C6929 S.n6309 VSUBS 1.88fF $ **FLOATING
C6930 S.n6310 VSUBS 2.67fF $ **FLOATING
C6931 S.t378 VSUBS 0.02fF
C6932 S.n6311 VSUBS 0.24fF $ **FLOATING
C6933 S.n6312 VSUBS 0.36fF $ **FLOATING
C6934 S.n6313 VSUBS 0.61fF $ **FLOATING
C6935 S.n6314 VSUBS 0.12fF $ **FLOATING
C6936 S.t2352 VSUBS 0.02fF
C6937 S.n6315 VSUBS 0.14fF $ **FLOATING
C6938 S.n6317 VSUBS 1.88fF $ **FLOATING
C6939 S.n6318 VSUBS 2.67fF $ **FLOATING
C6940 S.t2031 VSUBS 0.02fF
C6941 S.n6319 VSUBS 0.24fF $ **FLOATING
C6942 S.n6320 VSUBS 0.36fF $ **FLOATING
C6943 S.n6321 VSUBS 0.61fF $ **FLOATING
C6944 S.t1242 VSUBS 0.02fF
C6945 S.n6322 VSUBS 0.24fF $ **FLOATING
C6946 S.n6323 VSUBS 0.91fF $ **FLOATING
C6947 S.n6324 VSUBS 0.05fF $ **FLOATING
C6948 S.t2083 VSUBS 0.02fF
C6949 S.n6325 VSUBS 0.12fF $ **FLOATING
C6950 S.n6326 VSUBS 0.14fF $ **FLOATING
C6951 S.n6328 VSUBS 0.12fF $ **FLOATING
C6952 S.t1227 VSUBS 0.02fF
C6953 S.n6329 VSUBS 0.14fF $ **FLOATING
C6954 S.n6331 VSUBS 2.30fF $ **FLOATING
C6955 S.n6332 VSUBS 2.94fF $ **FLOATING
C6956 S.n6333 VSUBS 5.16fF $ **FLOATING
C6957 S.t695 VSUBS 0.02fF
C6958 S.n6334 VSUBS 0.12fF $ **FLOATING
C6959 S.n6335 VSUBS 0.14fF $ **FLOATING
C6960 S.t938 VSUBS 0.02fF
C6961 S.n6337 VSUBS 0.24fF $ **FLOATING
C6962 S.n6338 VSUBS 0.91fF $ **FLOATING
C6963 S.n6339 VSUBS 0.05fF $ **FLOATING
C6964 S.n6340 VSUBS 1.88fF $ **FLOATING
C6965 S.n6341 VSUBS 2.67fF $ **FLOATING
C6966 S.t921 VSUBS 0.02fF
C6967 S.n6342 VSUBS 0.24fF $ **FLOATING
C6968 S.n6343 VSUBS 0.36fF $ **FLOATING
C6969 S.n6344 VSUBS 0.61fF $ **FLOATING
C6970 S.n6345 VSUBS 0.12fF $ **FLOATING
C6971 S.t275 VSUBS 0.02fF
C6972 S.n6346 VSUBS 0.14fF $ **FLOATING
C6973 S.n6348 VSUBS 5.17fF $ **FLOATING
C6974 S.t1611 VSUBS 0.02fF
C6975 S.n6349 VSUBS 0.12fF $ **FLOATING
C6976 S.n6350 VSUBS 0.14fF $ **FLOATING
C6977 S.t905 VSUBS 0.02fF
C6978 S.n6352 VSUBS 0.24fF $ **FLOATING
C6979 S.n6353 VSUBS 0.91fF $ **FLOATING
C6980 S.n6354 VSUBS 0.05fF $ **FLOATING
C6981 S.n6355 VSUBS 1.88fF $ **FLOATING
C6982 S.n6356 VSUBS 0.12fF $ **FLOATING
C6983 S.t1054 VSUBS 0.02fF
C6984 S.n6357 VSUBS 0.14fF $ **FLOATING
C6985 S.t1699 VSUBS 0.02fF
C6986 S.n6359 VSUBS 0.24fF $ **FLOATING
C6987 S.n6360 VSUBS 0.36fF $ **FLOATING
C6988 S.n6361 VSUBS 0.61fF $ **FLOATING
C6989 S.n6362 VSUBS 2.67fF $ **FLOATING
C6990 S.n6363 VSUBS 5.17fF $ **FLOATING
C6991 S.t1924 VSUBS 0.02fF
C6992 S.n6364 VSUBS 0.12fF $ **FLOATING
C6993 S.n6365 VSUBS 0.14fF $ **FLOATING
C6994 S.t1685 VSUBS 0.02fF
C6995 S.n6367 VSUBS 0.24fF $ **FLOATING
C6996 S.n6368 VSUBS 0.91fF $ **FLOATING
C6997 S.n6369 VSUBS 0.05fF $ **FLOATING
C6998 S.n6370 VSUBS 1.88fF $ **FLOATING
C6999 S.n6371 VSUBS 2.67fF $ **FLOATING
C7000 S.t2488 VSUBS 0.02fF
C7001 S.n6372 VSUBS 0.24fF $ **FLOATING
C7002 S.n6373 VSUBS 0.36fF $ **FLOATING
C7003 S.n6374 VSUBS 0.61fF $ **FLOATING
C7004 S.n6375 VSUBS 0.12fF $ **FLOATING
C7005 S.t1840 VSUBS 0.02fF
C7006 S.n6376 VSUBS 0.14fF $ **FLOATING
C7007 S.n6378 VSUBS 5.17fF $ **FLOATING
C7008 S.t181 VSUBS 0.02fF
C7009 S.n6379 VSUBS 0.12fF $ **FLOATING
C7010 S.n6380 VSUBS 0.14fF $ **FLOATING
C7011 S.t2471 VSUBS 0.02fF
C7012 S.n6382 VSUBS 0.24fF $ **FLOATING
C7013 S.n6383 VSUBS 0.91fF $ **FLOATING
C7014 S.n6384 VSUBS 0.05fF $ **FLOATING
C7015 S.n6385 VSUBS 1.88fF $ **FLOATING
C7016 S.n6386 VSUBS 2.67fF $ **FLOATING
C7017 S.t743 VSUBS 0.02fF
C7018 S.n6387 VSUBS 0.24fF $ **FLOATING
C7019 S.n6388 VSUBS 0.36fF $ **FLOATING
C7020 S.n6389 VSUBS 0.61fF $ **FLOATING
C7021 S.n6390 VSUBS 0.12fF $ **FLOATING
C7022 S.t70 VSUBS 0.02fF
C7023 S.n6391 VSUBS 0.14fF $ **FLOATING
C7024 S.n6393 VSUBS 4.89fF $ **FLOATING
C7025 S.t970 VSUBS 0.02fF
C7026 S.n6394 VSUBS 0.12fF $ **FLOATING
C7027 S.n6395 VSUBS 0.14fF $ **FLOATING
C7028 S.t732 VSUBS 0.02fF
C7029 S.n6397 VSUBS 0.24fF $ **FLOATING
C7030 S.n6398 VSUBS 0.91fF $ **FLOATING
C7031 S.n6399 VSUBS 0.05fF $ **FLOATING
C7032 S.n6400 VSUBS 1.88fF $ **FLOATING
C7033 S.n6401 VSUBS 2.67fF $ **FLOATING
C7034 S.t1535 VSUBS 0.02fF
C7035 S.n6402 VSUBS 0.24fF $ **FLOATING
C7036 S.n6403 VSUBS 0.36fF $ **FLOATING
C7037 S.n6404 VSUBS 0.61fF $ **FLOATING
C7038 S.n6405 VSUBS 0.12fF $ **FLOATING
C7039 S.t885 VSUBS 0.02fF
C7040 S.n6406 VSUBS 0.14fF $ **FLOATING
C7041 S.n6408 VSUBS 1.88fF $ **FLOATING
C7042 S.n6409 VSUBS 2.68fF $ **FLOATING
C7043 S.t1285 VSUBS 0.02fF
C7044 S.n6410 VSUBS 0.24fF $ **FLOATING
C7045 S.n6411 VSUBS 0.36fF $ **FLOATING
C7046 S.n6412 VSUBS 0.61fF $ **FLOATING
C7047 S.t522 VSUBS 0.02fF
C7048 S.n6413 VSUBS 1.22fF $ **FLOATING
C7049 S.n6414 VSUBS 0.61fF $ **FLOATING
C7050 S.n6415 VSUBS 0.35fF $ **FLOATING
C7051 S.n6416 VSUBS 0.63fF $ **FLOATING
C7052 S.n6417 VSUBS 1.15fF $ **FLOATING
C7053 S.n6418 VSUBS 3.00fF $ **FLOATING
C7054 S.n6419 VSUBS 0.59fF $ **FLOATING
C7055 S.n6420 VSUBS 0.01fF $ **FLOATING
C7056 S.n6421 VSUBS 0.97fF $ **FLOATING
C7057 S.t59 VSUBS 21.42fF
C7058 S.n6422 VSUBS 20.29fF $ **FLOATING
C7059 S.n6424 VSUBS 0.38fF $ **FLOATING
C7060 S.n6425 VSUBS 0.23fF $ **FLOATING
C7061 S.n6426 VSUBS 2.90fF $ **FLOATING
C7062 S.n6427 VSUBS 2.46fF $ **FLOATING
C7063 S.n6428 VSUBS 1.96fF $ **FLOATING
C7064 S.n6429 VSUBS 3.94fF $ **FLOATING
C7065 S.n6430 VSUBS 0.25fF $ **FLOATING
C7066 S.n6431 VSUBS 0.01fF $ **FLOATING
C7067 S.t2228 VSUBS 0.02fF
C7068 S.n6432 VSUBS 0.26fF $ **FLOATING
C7069 S.t2247 VSUBS 0.02fF
C7070 S.n6433 VSUBS 0.95fF $ **FLOATING
C7071 S.n6434 VSUBS 0.71fF $ **FLOATING
C7072 S.n6435 VSUBS 0.78fF $ **FLOATING
C7073 S.n6436 VSUBS 1.93fF $ **FLOATING
C7074 S.n6437 VSUBS 1.88fF $ **FLOATING
C7075 S.n6438 VSUBS 0.12fF $ **FLOATING
C7076 S.t498 VSUBS 0.02fF
C7077 S.n6439 VSUBS 0.14fF $ **FLOATING
C7078 S.t1310 VSUBS 0.02fF
C7079 S.n6441 VSUBS 0.24fF $ **FLOATING
C7080 S.n6442 VSUBS 0.36fF $ **FLOATING
C7081 S.n6443 VSUBS 0.61fF $ **FLOATING
C7082 S.n6444 VSUBS 1.52fF $ **FLOATING
C7083 S.n6445 VSUBS 2.99fF $ **FLOATING
C7084 S.t517 VSUBS 0.02fF
C7085 S.n6446 VSUBS 0.24fF $ **FLOATING
C7086 S.n6447 VSUBS 0.91fF $ **FLOATING
C7087 S.n6448 VSUBS 0.05fF $ **FLOATING
C7088 S.t1365 VSUBS 0.02fF
C7089 S.n6449 VSUBS 0.12fF $ **FLOATING
C7090 S.n6450 VSUBS 0.14fF $ **FLOATING
C7091 S.n6452 VSUBS 1.89fF $ **FLOATING
C7092 S.n6453 VSUBS 1.88fF $ **FLOATING
C7093 S.t2098 VSUBS 0.02fF
C7094 S.n6454 VSUBS 0.24fF $ **FLOATING
C7095 S.n6455 VSUBS 0.36fF $ **FLOATING
C7096 S.n6456 VSUBS 0.61fF $ **FLOATING
C7097 S.n6457 VSUBS 0.12fF $ **FLOATING
C7098 S.t1404 VSUBS 0.02fF
C7099 S.n6458 VSUBS 0.14fF $ **FLOATING
C7100 S.n6460 VSUBS 1.16fF $ **FLOATING
C7101 S.n6461 VSUBS 0.22fF $ **FLOATING
C7102 S.n6462 VSUBS 0.25fF $ **FLOATING
C7103 S.n6463 VSUBS 0.09fF $ **FLOATING
C7104 S.n6464 VSUBS 1.88fF $ **FLOATING
C7105 S.t1303 VSUBS 0.02fF
C7106 S.n6465 VSUBS 0.24fF $ **FLOATING
C7107 S.n6466 VSUBS 0.91fF $ **FLOATING
C7108 S.n6467 VSUBS 0.05fF $ **FLOATING
C7109 S.t2151 VSUBS 0.02fF
C7110 S.n6468 VSUBS 0.12fF $ **FLOATING
C7111 S.n6469 VSUBS 0.14fF $ **FLOATING
C7112 S.n6471 VSUBS 0.78fF $ **FLOATING
C7113 S.n6472 VSUBS 1.94fF $ **FLOATING
C7114 S.n6473 VSUBS 1.88fF $ **FLOATING
C7115 S.n6474 VSUBS 0.12fF $ **FLOATING
C7116 S.t2195 VSUBS 0.02fF
C7117 S.n6475 VSUBS 0.14fF $ **FLOATING
C7118 S.t487 VSUBS 0.02fF
C7119 S.n6477 VSUBS 0.24fF $ **FLOATING
C7120 S.n6478 VSUBS 0.36fF $ **FLOATING
C7121 S.n6479 VSUBS 0.61fF $ **FLOATING
C7122 S.n6480 VSUBS 1.84fF $ **FLOATING
C7123 S.n6481 VSUBS 2.99fF $ **FLOATING
C7124 S.t2215 VSUBS 0.02fF
C7125 S.n6482 VSUBS 0.24fF $ **FLOATING
C7126 S.n6483 VSUBS 0.91fF $ **FLOATING
C7127 S.n6484 VSUBS 0.05fF $ **FLOATING
C7128 S.t540 VSUBS 0.02fF
C7129 S.n6485 VSUBS 0.12fF $ **FLOATING
C7130 S.n6486 VSUBS 0.14fF $ **FLOATING
C7131 S.n6488 VSUBS 1.89fF $ **FLOATING
C7132 S.n6489 VSUBS 1.88fF $ **FLOATING
C7133 S.t60 VSUBS 0.02fF
C7134 S.n6490 VSUBS 0.24fF $ **FLOATING
C7135 S.n6491 VSUBS 0.36fF $ **FLOATING
C7136 S.n6492 VSUBS 0.61fF $ **FLOATING
C7137 S.n6493 VSUBS 0.12fF $ **FLOATING
C7138 S.t1800 VSUBS 0.02fF
C7139 S.n6494 VSUBS 0.14fF $ **FLOATING
C7140 S.n6496 VSUBS 1.16fF $ **FLOATING
C7141 S.n6497 VSUBS 0.22fF $ **FLOATING
C7142 S.n6498 VSUBS 0.25fF $ **FLOATING
C7143 S.n6499 VSUBS 0.09fF $ **FLOATING
C7144 S.n6500 VSUBS 1.88fF $ **FLOATING
C7145 S.t1828 VSUBS 0.02fF
C7146 S.n6501 VSUBS 0.24fF $ **FLOATING
C7147 S.n6502 VSUBS 0.91fF $ **FLOATING
C7148 S.n6503 VSUBS 0.05fF $ **FLOATING
C7149 S.t138 VSUBS 0.02fF
C7150 S.n6504 VSUBS 0.12fF $ **FLOATING
C7151 S.n6505 VSUBS 0.14fF $ **FLOATING
C7152 S.n6507 VSUBS 0.78fF $ **FLOATING
C7153 S.n6508 VSUBS 1.94fF $ **FLOATING
C7154 S.n6509 VSUBS 1.88fF $ **FLOATING
C7155 S.n6510 VSUBS 0.12fF $ **FLOATING
C7156 S.t5 VSUBS 0.02fF
C7157 S.n6511 VSUBS 0.14fF $ **FLOATING
C7158 S.t879 VSUBS 0.02fF
C7159 S.n6513 VSUBS 0.24fF $ **FLOATING
C7160 S.n6514 VSUBS 0.36fF $ **FLOATING
C7161 S.n6515 VSUBS 0.61fF $ **FLOATING
C7162 S.n6516 VSUBS 1.84fF $ **FLOATING
C7163 S.n6517 VSUBS 2.99fF $ **FLOATING
C7164 S.t45 VSUBS 0.02fF
C7165 S.n6518 VSUBS 0.24fF $ **FLOATING
C7166 S.n6519 VSUBS 0.91fF $ **FLOATING
C7167 S.n6520 VSUBS 0.05fF $ **FLOATING
C7168 S.t936 VSUBS 0.02fF
C7169 S.n6521 VSUBS 0.12fF $ **FLOATING
C7170 S.n6522 VSUBS 0.14fF $ **FLOATING
C7171 S.n6524 VSUBS 1.89fF $ **FLOATING
C7172 S.n6525 VSUBS 1.75fF $ **FLOATING
C7173 S.t1660 VSUBS 0.02fF
C7174 S.n6526 VSUBS 0.24fF $ **FLOATING
C7175 S.n6527 VSUBS 0.36fF $ **FLOATING
C7176 S.n6528 VSUBS 0.61fF $ **FLOATING
C7177 S.n6529 VSUBS 0.12fF $ **FLOATING
C7178 S.t847 VSUBS 0.02fF
C7179 S.n6530 VSUBS 0.14fF $ **FLOATING
C7180 S.n6532 VSUBS 1.16fF $ **FLOATING
C7181 S.n6533 VSUBS 0.22fF $ **FLOATING
C7182 S.n6534 VSUBS 0.25fF $ **FLOATING
C7183 S.n6535 VSUBS 0.09fF $ **FLOATING
C7184 S.n6536 VSUBS 2.44fF $ **FLOATING
C7185 S.t868 VSUBS 0.02fF
C7186 S.n6537 VSUBS 0.24fF $ **FLOATING
C7187 S.n6538 VSUBS 0.91fF $ **FLOATING
C7188 S.n6539 VSUBS 0.05fF $ **FLOATING
C7189 S.t1714 VSUBS 0.02fF
C7190 S.n6540 VSUBS 0.12fF $ **FLOATING
C7191 S.n6541 VSUBS 0.14fF $ **FLOATING
C7192 S.n6543 VSUBS 1.88fF $ **FLOATING
C7193 S.n6544 VSUBS 0.48fF $ **FLOATING
C7194 S.n6545 VSUBS 0.09fF $ **FLOATING
C7195 S.n6546 VSUBS 0.33fF $ **FLOATING
C7196 S.n6547 VSUBS 0.30fF $ **FLOATING
C7197 S.n6548 VSUBS 0.77fF $ **FLOATING
C7198 S.n6549 VSUBS 0.59fF $ **FLOATING
C7199 S.t2443 VSUBS 0.02fF
C7200 S.n6550 VSUBS 0.24fF $ **FLOATING
C7201 S.n6551 VSUBS 0.36fF $ **FLOATING
C7202 S.n6552 VSUBS 0.61fF $ **FLOATING
C7203 S.n6553 VSUBS 0.12fF $ **FLOATING
C7204 S.t1767 VSUBS 0.02fF
C7205 S.n6554 VSUBS 0.14fF $ **FLOATING
C7206 S.n6556 VSUBS 2.61fF $ **FLOATING
C7207 S.n6557 VSUBS 2.15fF $ **FLOATING
C7208 S.t1652 VSUBS 0.02fF
C7209 S.n6558 VSUBS 0.24fF $ **FLOATING
C7210 S.n6559 VSUBS 0.91fF $ **FLOATING
C7211 S.n6560 VSUBS 0.05fF $ **FLOATING
C7212 S.t2502 VSUBS 0.02fF
C7213 S.n6561 VSUBS 0.12fF $ **FLOATING
C7214 S.n6562 VSUBS 0.14fF $ **FLOATING
C7215 S.n6564 VSUBS 0.78fF $ **FLOATING
C7216 S.n6565 VSUBS 2.30fF $ **FLOATING
C7217 S.n6566 VSUBS 1.88fF $ **FLOATING
C7218 S.n6567 VSUBS 0.12fF $ **FLOATING
C7219 S.t1378 VSUBS 0.02fF
C7220 S.n6568 VSUBS 0.14fF $ **FLOATING
C7221 S.t2194 VSUBS 0.02fF
C7222 S.n6570 VSUBS 0.24fF $ **FLOATING
C7223 S.n6571 VSUBS 0.36fF $ **FLOATING
C7224 S.n6572 VSUBS 0.61fF $ **FLOATING
C7225 S.n6573 VSUBS 1.39fF $ **FLOATING
C7226 S.n6574 VSUBS 0.71fF $ **FLOATING
C7227 S.n6575 VSUBS 1.14fF $ **FLOATING
C7228 S.n6576 VSUBS 0.35fF $ **FLOATING
C7229 S.n6577 VSUBS 2.02fF $ **FLOATING
C7230 S.t1398 VSUBS 0.02fF
C7231 S.n6578 VSUBS 0.24fF $ **FLOATING
C7232 S.n6579 VSUBS 0.91fF $ **FLOATING
C7233 S.n6580 VSUBS 0.05fF $ **FLOATING
C7234 S.t897 VSUBS 0.02fF
C7235 S.n6581 VSUBS 0.12fF $ **FLOATING
C7236 S.n6582 VSUBS 0.14fF $ **FLOATING
C7237 S.n6584 VSUBS 1.89fF $ **FLOATING
C7238 S.n6585 VSUBS 1.88fF $ **FLOATING
C7239 S.t460 VSUBS 0.02fF
C7240 S.n6586 VSUBS 0.24fF $ **FLOATING
C7241 S.n6587 VSUBS 0.36fF $ **FLOATING
C7242 S.n6588 VSUBS 0.61fF $ **FLOATING
C7243 S.n6589 VSUBS 0.12fF $ **FLOATING
C7244 S.t2163 VSUBS 0.02fF
C7245 S.n6590 VSUBS 0.14fF $ **FLOATING
C7246 S.n6592 VSUBS 1.16fF $ **FLOATING
C7247 S.n6593 VSUBS 0.22fF $ **FLOATING
C7248 S.n6594 VSUBS 0.25fF $ **FLOATING
C7249 S.n6595 VSUBS 0.09fF $ **FLOATING
C7250 S.n6596 VSUBS 1.88fF $ **FLOATING
C7251 S.t2186 VSUBS 0.02fF
C7252 S.n6597 VSUBS 0.24fF $ **FLOATING
C7253 S.n6598 VSUBS 0.91fF $ **FLOATING
C7254 S.n6599 VSUBS 0.05fF $ **FLOATING
C7255 S.t511 VSUBS 0.02fF
C7256 S.n6600 VSUBS 0.12fF $ **FLOATING
C7257 S.n6601 VSUBS 0.14fF $ **FLOATING
C7258 S.n6603 VSUBS 20.78fF $ **FLOATING
C7259 S.n6604 VSUBS 1.88fF $ **FLOATING
C7260 S.n6605 VSUBS 2.67fF $ **FLOATING
C7261 S.t302 VSUBS 0.02fF
C7262 S.n6606 VSUBS 0.24fF $ **FLOATING
C7263 S.n6607 VSUBS 0.36fF $ **FLOATING
C7264 S.n6608 VSUBS 0.61fF $ **FLOATING
C7265 S.n6609 VSUBS 0.12fF $ **FLOATING
C7266 S.t2131 VSUBS 0.02fF
C7267 S.n6610 VSUBS 0.14fF $ **FLOATING
C7268 S.n6612 VSUBS 2.80fF $ **FLOATING
C7269 S.n6613 VSUBS 2.30fF $ **FLOATING
C7270 S.t357 VSUBS 0.02fF
C7271 S.n6614 VSUBS 0.12fF $ **FLOATING
C7272 S.n6615 VSUBS 0.14fF $ **FLOATING
C7273 S.t2027 VSUBS 0.02fF
C7274 S.n6617 VSUBS 0.24fF $ **FLOATING
C7275 S.n6618 VSUBS 0.91fF $ **FLOATING
C7276 S.n6619 VSUBS 0.05fF $ **FLOATING
C7277 S.n6620 VSUBS 2.80fF $ **FLOATING
C7278 S.n6621 VSUBS 1.88fF $ **FLOATING
C7279 S.n6622 VSUBS 0.12fF $ **FLOATING
C7280 S.t1642 VSUBS 0.02fF
C7281 S.n6623 VSUBS 0.14fF $ **FLOATING
C7282 S.t1441 VSUBS 0.02fF
C7283 S.n6625 VSUBS 0.24fF $ **FLOATING
C7284 S.n6626 VSUBS 0.36fF $ **FLOATING
C7285 S.n6627 VSUBS 0.61fF $ **FLOATING
C7286 S.n6628 VSUBS 2.67fF $ **FLOATING
C7287 S.n6629 VSUBS 2.30fF $ **FLOATING
C7288 S.t2509 VSUBS 0.02fF
C7289 S.n6630 VSUBS 0.12fF $ **FLOATING
C7290 S.n6631 VSUBS 0.14fF $ **FLOATING
C7291 S.t2569 VSUBS 0.02fF
C7292 S.n6633 VSUBS 0.24fF $ **FLOATING
C7293 S.n6634 VSUBS 0.91fF $ **FLOATING
C7294 S.n6635 VSUBS 0.05fF $ **FLOATING
C7295 S.n6636 VSUBS 1.88fF $ **FLOATING
C7296 S.n6637 VSUBS 2.67fF $ **FLOATING
C7297 S.t2234 VSUBS 0.02fF
C7298 S.n6638 VSUBS 0.24fF $ **FLOATING
C7299 S.n6639 VSUBS 0.36fF $ **FLOATING
C7300 S.n6640 VSUBS 0.61fF $ **FLOATING
C7301 S.n6641 VSUBS 0.12fF $ **FLOATING
C7302 S.t2426 VSUBS 0.02fF
C7303 S.n6642 VSUBS 0.14fF $ **FLOATING
C7304 S.n6644 VSUBS 2.80fF $ **FLOATING
C7305 S.n6645 VSUBS 2.30fF $ **FLOATING
C7306 S.t772 VSUBS 0.02fF
C7307 S.n6646 VSUBS 0.12fF $ **FLOATING
C7308 S.n6647 VSUBS 0.14fF $ **FLOATING
C7309 S.t834 VSUBS 0.02fF
C7310 S.n6649 VSUBS 0.24fF $ **FLOATING
C7311 S.n6650 VSUBS 0.91fF $ **FLOATING
C7312 S.n6651 VSUBS 0.05fF $ **FLOATING
C7313 S.n6652 VSUBS 1.88fF $ **FLOATING
C7314 S.n6653 VSUBS 2.67fF $ **FLOATING
C7315 S.t501 VSUBS 0.02fF
C7316 S.n6654 VSUBS 0.24fF $ **FLOATING
C7317 S.n6655 VSUBS 0.36fF $ **FLOATING
C7318 S.n6656 VSUBS 0.61fF $ **FLOATING
C7319 S.n6657 VSUBS 0.12fF $ **FLOATING
C7320 S.t691 VSUBS 0.02fF
C7321 S.n6658 VSUBS 0.14fF $ **FLOATING
C7322 S.n6660 VSUBS 2.80fF $ **FLOATING
C7323 S.n6661 VSUBS 2.30fF $ **FLOATING
C7324 S.t1559 VSUBS 0.02fF
C7325 S.n6662 VSUBS 0.12fF $ **FLOATING
C7326 S.n6663 VSUBS 0.14fF $ **FLOATING
C7327 S.t1616 VSUBS 0.02fF
C7328 S.n6665 VSUBS 0.24fF $ **FLOATING
C7329 S.n6666 VSUBS 0.91fF $ **FLOATING
C7330 S.n6667 VSUBS 0.05fF $ **FLOATING
C7331 S.n6668 VSUBS 2.73fF $ **FLOATING
C7332 S.n6669 VSUBS 1.59fF $ **FLOATING
C7333 S.n6670 VSUBS 0.12fF $ **FLOATING
C7334 S.t351 VSUBS 0.02fF
C7335 S.n6671 VSUBS 0.14fF $ **FLOATING
C7336 S.t1591 VSUBS 0.02fF
C7337 S.n6673 VSUBS 0.24fF $ **FLOATING
C7338 S.n6674 VSUBS 0.36fF $ **FLOATING
C7339 S.n6675 VSUBS 0.61fF $ **FLOATING
C7340 S.n6676 VSUBS 0.07fF $ **FLOATING
C7341 S.n6677 VSUBS 0.01fF $ **FLOATING
C7342 S.n6678 VSUBS 0.24fF $ **FLOATING
C7343 S.n6679 VSUBS 1.16fF $ **FLOATING
C7344 S.n6680 VSUBS 1.35fF $ **FLOATING
C7345 S.n6681 VSUBS 2.30fF $ **FLOATING
C7346 S.t611 VSUBS 0.02fF
C7347 S.n6682 VSUBS 0.12fF $ **FLOATING
C7348 S.n6683 VSUBS 0.14fF $ **FLOATING
C7349 S.t1128 VSUBS 0.02fF
C7350 S.n6685 VSUBS 0.24fF $ **FLOATING
C7351 S.n6686 VSUBS 0.91fF $ **FLOATING
C7352 S.n6687 VSUBS 0.05fF $ **FLOATING
C7353 S.t4 VSUBS 48.27fF
C7354 S.t2403 VSUBS 0.02fF
C7355 S.n6688 VSUBS 0.24fF $ **FLOATING
C7356 S.n6689 VSUBS 0.91fF $ **FLOATING
C7357 S.n6690 VSUBS 0.05fF $ **FLOATING
C7358 S.t2347 VSUBS 0.02fF
C7359 S.n6691 VSUBS 0.12fF $ **FLOATING
C7360 S.n6692 VSUBS 0.14fF $ **FLOATING
C7361 S.n6694 VSUBS 0.12fF $ **FLOATING
C7362 S.t1480 VSUBS 0.02fF
C7363 S.n6695 VSUBS 0.14fF $ **FLOATING
C7364 S.n6697 VSUBS 5.17fF $ **FLOATING
C7365 S.n6698 VSUBS 5.44fF $ **FLOATING
C7366 S.t1753 VSUBS 0.02fF
C7367 S.n6699 VSUBS 0.12fF $ **FLOATING
C7368 S.n6700 VSUBS 0.14fF $ **FLOATING
C7369 S.t1521 VSUBS 0.02fF
C7370 S.n6702 VSUBS 0.24fF $ **FLOATING
C7371 S.n6703 VSUBS 0.91fF $ **FLOATING
C7372 S.n6704 VSUBS 0.05fF $ **FLOATING
C7373 S.t69 VSUBS 47.89fF
C7374 S.t1479 VSUBS 0.02fF
C7375 S.n6705 VSUBS 0.01fF $ **FLOATING
C7376 S.n6706 VSUBS 0.26fF $ **FLOATING
C7377 S.t319 VSUBS 0.02fF
C7378 S.n6708 VSUBS 1.19fF $ **FLOATING
C7379 S.n6709 VSUBS 0.05fF $ **FLOATING
C7380 S.t2258 VSUBS 0.02fF
C7381 S.n6710 VSUBS 0.64fF $ **FLOATING
C7382 S.n6711 VSUBS 0.61fF $ **FLOATING
C7383 S.n6712 VSUBS 8.97fF $ **FLOATING
C7384 S.n6713 VSUBS 8.97fF $ **FLOATING
C7385 S.n6714 VSUBS 0.60fF $ **FLOATING
C7386 S.n6715 VSUBS 0.22fF $ **FLOATING
C7387 S.n6716 VSUBS 0.59fF $ **FLOATING
C7388 S.n6717 VSUBS 3.39fF $ **FLOATING
C7389 S.n6718 VSUBS 0.29fF $ **FLOATING
C7390 S.t44 VSUBS 21.42fF
C7391 S.n6719 VSUBS 21.71fF $ **FLOATING
C7392 S.n6720 VSUBS 0.77fF $ **FLOATING
C7393 S.n6721 VSUBS 0.28fF $ **FLOATING
C7394 S.n6722 VSUBS 4.00fF $ **FLOATING
C7395 S.n6723 VSUBS 1.35fF $ **FLOATING
C7396 S.n6724 VSUBS 0.01fF $ **FLOATING
C7397 S.n6725 VSUBS 0.02fF $ **FLOATING
C7398 S.n6726 VSUBS 0.03fF $ **FLOATING
C7399 S.n6727 VSUBS 0.04fF $ **FLOATING
C7400 S.n6728 VSUBS 0.17fF $ **FLOATING
C7401 S.n6729 VSUBS 0.01fF $ **FLOATING
C7402 S.n6730 VSUBS 0.02fF $ **FLOATING
C7403 S.n6731 VSUBS 0.01fF $ **FLOATING
C7404 S.n6732 VSUBS 0.01fF $ **FLOATING
C7405 S.n6733 VSUBS 0.01fF $ **FLOATING
C7406 S.n6734 VSUBS 0.01fF $ **FLOATING
C7407 S.n6735 VSUBS 0.02fF $ **FLOATING
C7408 S.n6736 VSUBS 0.01fF $ **FLOATING
C7409 S.n6737 VSUBS 0.02fF $ **FLOATING
C7410 S.n6738 VSUBS 0.05fF $ **FLOATING
C7411 S.n6739 VSUBS 0.04fF $ **FLOATING
C7412 S.n6740 VSUBS 0.11fF $ **FLOATING
C7413 S.n6741 VSUBS 0.38fF $ **FLOATING
C7414 S.n6742 VSUBS 0.20fF $ **FLOATING
C7415 S.n6743 VSUBS 4.39fF $ **FLOATING
C7416 S.n6744 VSUBS 0.24fF $ **FLOATING
C7417 S.n6745 VSUBS 1.50fF $ **FLOATING
C7418 S.n6746 VSUBS 1.31fF $ **FLOATING
C7419 S.n6747 VSUBS 0.28fF $ **FLOATING
C7420 S.n6748 VSUBS 1.89fF $ **FLOATING
C7421 S.n6749 VSUBS 0.06fF $ **FLOATING
C7422 S.n6750 VSUBS 0.03fF $ **FLOATING
C7423 S.n6751 VSUBS 0.04fF $ **FLOATING
C7424 S.n6752 VSUBS 0.99fF $ **FLOATING
C7425 S.n6753 VSUBS 0.02fF $ **FLOATING
C7426 S.n6754 VSUBS 0.01fF $ **FLOATING
C7427 S.n6755 VSUBS 0.02fF $ **FLOATING
C7428 S.n6756 VSUBS 0.08fF $ **FLOATING
C7429 S.n6757 VSUBS 0.36fF $ **FLOATING
C7430 S.n6758 VSUBS 1.85fF $ **FLOATING
C7431 S.t148 VSUBS 0.02fF
C7432 S.n6759 VSUBS 0.24fF $ **FLOATING
C7433 S.n6760 VSUBS 0.36fF $ **FLOATING
C7434 S.n6761 VSUBS 0.61fF $ **FLOATING
C7435 S.n6762 VSUBS 0.12fF $ **FLOATING
C7436 S.t1864 VSUBS 0.02fF
C7437 S.n6763 VSUBS 0.14fF $ **FLOATING
C7438 S.n6765 VSUBS 0.70fF $ **FLOATING
C7439 S.n6766 VSUBS 0.23fF $ **FLOATING
C7440 S.n6767 VSUBS 0.23fF $ **FLOATING
C7441 S.n6768 VSUBS 0.70fF $ **FLOATING
C7442 S.n6769 VSUBS 1.16fF $ **FLOATING
C7443 S.n6770 VSUBS 0.22fF $ **FLOATING
C7444 S.n6771 VSUBS 0.25fF $ **FLOATING
C7445 S.n6772 VSUBS 0.09fF $ **FLOATING
C7446 S.n6773 VSUBS 1.88fF $ **FLOATING
C7447 S.t445 VSUBS 0.02fF
C7448 S.n6774 VSUBS 0.24fF $ **FLOATING
C7449 S.n6775 VSUBS 0.91fF $ **FLOATING
C7450 S.n6776 VSUBS 0.05fF $ **FLOATING
C7451 S.t207 VSUBS 0.02fF
C7452 S.n6777 VSUBS 0.12fF $ **FLOATING
C7453 S.n6778 VSUBS 0.14fF $ **FLOATING
C7454 S.n6780 VSUBS 0.25fF $ **FLOATING
C7455 S.n6781 VSUBS 0.09fF $ **FLOATING
C7456 S.n6782 VSUBS 0.21fF $ **FLOATING
C7457 S.n6783 VSUBS 0.92fF $ **FLOATING
C7458 S.n6784 VSUBS 0.44fF $ **FLOATING
C7459 S.n6785 VSUBS 1.88fF $ **FLOATING
C7460 S.n6786 VSUBS 0.12fF $ **FLOATING
C7461 S.t263 VSUBS 0.02fF
C7462 S.n6787 VSUBS 0.14fF $ **FLOATING
C7463 S.t1074 VSUBS 0.02fF
C7464 S.n6789 VSUBS 0.24fF $ **FLOATING
C7465 S.n6790 VSUBS 0.36fF $ **FLOATING
C7466 S.n6791 VSUBS 0.61fF $ **FLOATING
C7467 S.n6792 VSUBS 0.02fF $ **FLOATING
C7468 S.n6793 VSUBS 0.01fF $ **FLOATING
C7469 S.n6794 VSUBS 0.02fF $ **FLOATING
C7470 S.n6795 VSUBS 0.08fF $ **FLOATING
C7471 S.n6796 VSUBS 0.06fF $ **FLOATING
C7472 S.n6797 VSUBS 0.03fF $ **FLOATING
C7473 S.n6798 VSUBS 0.04fF $ **FLOATING
C7474 S.n6799 VSUBS 1.00fF $ **FLOATING
C7475 S.n6800 VSUBS 0.36fF $ **FLOATING
C7476 S.n6801 VSUBS 1.87fF $ **FLOATING
C7477 S.n6802 VSUBS 1.99fF $ **FLOATING
C7478 S.t1354 VSUBS 0.02fF
C7479 S.n6803 VSUBS 0.24fF $ **FLOATING
C7480 S.n6804 VSUBS 0.91fF $ **FLOATING
C7481 S.n6805 VSUBS 0.05fF $ **FLOATING
C7482 S.t1132 VSUBS 0.02fF
C7483 S.n6806 VSUBS 0.12fF $ **FLOATING
C7484 S.n6807 VSUBS 0.14fF $ **FLOATING
C7485 S.n6809 VSUBS 1.89fF $ **FLOATING
C7486 S.n6810 VSUBS 0.06fF $ **FLOATING
C7487 S.n6811 VSUBS 0.03fF $ **FLOATING
C7488 S.n6812 VSUBS 0.04fF $ **FLOATING
C7489 S.n6813 VSUBS 0.99fF $ **FLOATING
C7490 S.n6814 VSUBS 0.02fF $ **FLOATING
C7491 S.n6815 VSUBS 0.01fF $ **FLOATING
C7492 S.n6816 VSUBS 0.02fF $ **FLOATING
C7493 S.n6817 VSUBS 0.08fF $ **FLOATING
C7494 S.n6818 VSUBS 0.36fF $ **FLOATING
C7495 S.n6819 VSUBS 1.85fF $ **FLOATING
C7496 S.t670 VSUBS 0.02fF
C7497 S.n6820 VSUBS 0.24fF $ **FLOATING
C7498 S.n6821 VSUBS 0.36fF $ **FLOATING
C7499 S.n6822 VSUBS 0.61fF $ **FLOATING
C7500 S.n6823 VSUBS 0.12fF $ **FLOATING
C7501 S.t2378 VSUBS 0.02fF
C7502 S.n6824 VSUBS 0.14fF $ **FLOATING
C7503 S.n6826 VSUBS 0.70fF $ **FLOATING
C7504 S.n6827 VSUBS 0.23fF $ **FLOATING
C7505 S.n6828 VSUBS 0.23fF $ **FLOATING
C7506 S.n6829 VSUBS 0.70fF $ **FLOATING
C7507 S.n6830 VSUBS 1.16fF $ **FLOATING
C7508 S.n6831 VSUBS 0.22fF $ **FLOATING
C7509 S.n6832 VSUBS 0.25fF $ **FLOATING
C7510 S.n6833 VSUBS 0.09fF $ **FLOATING
C7511 S.n6834 VSUBS 1.88fF $ **FLOATING
C7512 S.t965 VSUBS 0.02fF
C7513 S.n6835 VSUBS 0.24fF $ **FLOATING
C7514 S.n6836 VSUBS 0.91fF $ **FLOATING
C7515 S.n6837 VSUBS 0.05fF $ **FLOATING
C7516 S.t1916 VSUBS 0.02fF
C7517 S.n6838 VSUBS 0.12fF $ **FLOATING
C7518 S.n6839 VSUBS 0.14fF $ **FLOATING
C7519 S.n6841 VSUBS 0.25fF $ **FLOATING
C7520 S.n6842 VSUBS 0.09fF $ **FLOATING
C7521 S.n6843 VSUBS 0.21fF $ **FLOATING
C7522 S.n6844 VSUBS 0.92fF $ **FLOATING
C7523 S.n6845 VSUBS 0.44fF $ **FLOATING
C7524 S.n6846 VSUBS 1.88fF $ **FLOATING
C7525 S.n6847 VSUBS 0.12fF $ **FLOATING
C7526 S.t643 VSUBS 0.02fF
C7527 S.n6848 VSUBS 0.14fF $ **FLOATING
C7528 S.t1457 VSUBS 0.02fF
C7529 S.n6850 VSUBS 0.24fF $ **FLOATING
C7530 S.n6851 VSUBS 0.36fF $ **FLOATING
C7531 S.n6852 VSUBS 0.61fF $ **FLOATING
C7532 S.n6853 VSUBS 0.02fF $ **FLOATING
C7533 S.n6854 VSUBS 0.01fF $ **FLOATING
C7534 S.n6855 VSUBS 0.02fF $ **FLOATING
C7535 S.n6856 VSUBS 0.08fF $ **FLOATING
C7536 S.n6857 VSUBS 0.06fF $ **FLOATING
C7537 S.n6858 VSUBS 0.03fF $ **FLOATING
C7538 S.n6859 VSUBS 0.04fF $ **FLOATING
C7539 S.n6860 VSUBS 1.00fF $ **FLOATING
C7540 S.n6861 VSUBS 0.36fF $ **FLOATING
C7541 S.n6862 VSUBS 1.87fF $ **FLOATING
C7542 S.n6863 VSUBS 1.99fF $ **FLOATING
C7543 S.t1746 VSUBS 0.02fF
C7544 S.n6864 VSUBS 0.24fF $ **FLOATING
C7545 S.n6865 VSUBS 0.91fF $ **FLOATING
C7546 S.n6866 VSUBS 0.05fF $ **FLOATING
C7547 S.t1510 VSUBS 0.02fF
C7548 S.n6867 VSUBS 0.12fF $ **FLOATING
C7549 S.n6868 VSUBS 0.14fF $ **FLOATING
C7550 S.n6870 VSUBS 1.89fF $ **FLOATING
C7551 S.n6871 VSUBS 0.04fF $ **FLOATING
C7552 S.n6872 VSUBS 0.07fF $ **FLOATING
C7553 S.n6873 VSUBS 0.05fF $ **FLOATING
C7554 S.n6874 VSUBS 0.87fF $ **FLOATING
C7555 S.n6875 VSUBS 0.01fF $ **FLOATING
C7556 S.n6876 VSUBS 0.01fF $ **FLOATING
C7557 S.n6877 VSUBS 0.01fF $ **FLOATING
C7558 S.n6878 VSUBS 0.07fF $ **FLOATING
C7559 S.n6879 VSUBS 0.68fF $ **FLOATING
C7560 S.n6880 VSUBS 0.72fF $ **FLOATING
C7561 S.t2246 VSUBS 0.02fF
C7562 S.n6881 VSUBS 0.24fF $ **FLOATING
C7563 S.n6882 VSUBS 0.36fF $ **FLOATING
C7564 S.n6883 VSUBS 0.61fF $ **FLOATING
C7565 S.n6884 VSUBS 0.12fF $ **FLOATING
C7566 S.t1431 VSUBS 0.02fF
C7567 S.n6885 VSUBS 0.14fF $ **FLOATING
C7568 S.n6887 VSUBS 0.70fF $ **FLOATING
C7569 S.n6888 VSUBS 0.23fF $ **FLOATING
C7570 S.n6889 VSUBS 0.23fF $ **FLOATING
C7571 S.n6890 VSUBS 0.70fF $ **FLOATING
C7572 S.n6891 VSUBS 1.16fF $ **FLOATING
C7573 S.n6892 VSUBS 0.22fF $ **FLOATING
C7574 S.n6893 VSUBS 0.25fF $ **FLOATING
C7575 S.n6894 VSUBS 0.09fF $ **FLOATING
C7576 S.n6895 VSUBS 2.31fF $ **FLOATING
C7577 S.t2528 VSUBS 0.02fF
C7578 S.n6896 VSUBS 0.24fF $ **FLOATING
C7579 S.n6897 VSUBS 0.91fF $ **FLOATING
C7580 S.n6898 VSUBS 0.05fF $ **FLOATING
C7581 S.t2298 VSUBS 0.02fF
C7582 S.n6899 VSUBS 0.12fF $ **FLOATING
C7583 S.n6900 VSUBS 0.14fF $ **FLOATING
C7584 S.n6902 VSUBS 1.88fF $ **FLOATING
C7585 S.n6903 VSUBS 0.46fF $ **FLOATING
C7586 S.n6904 VSUBS 0.22fF $ **FLOATING
C7587 S.n6905 VSUBS 0.38fF $ **FLOATING
C7588 S.n6906 VSUBS 0.16fF $ **FLOATING
C7589 S.n6907 VSUBS 0.28fF $ **FLOATING
C7590 S.n6908 VSUBS 0.21fF $ **FLOATING
C7591 S.n6909 VSUBS 0.30fF $ **FLOATING
C7592 S.n6910 VSUBS 0.42fF $ **FLOATING
C7593 S.n6911 VSUBS 0.21fF $ **FLOATING
C7594 S.t516 VSUBS 0.02fF
C7595 S.n6912 VSUBS 0.24fF $ **FLOATING
C7596 S.n6913 VSUBS 0.36fF $ **FLOATING
C7597 S.n6914 VSUBS 0.61fF $ **FLOATING
C7598 S.n6915 VSUBS 0.12fF $ **FLOATING
C7599 S.t2222 VSUBS 0.02fF
C7600 S.n6916 VSUBS 0.14fF $ **FLOATING
C7601 S.n6918 VSUBS 0.04fF $ **FLOATING
C7602 S.n6919 VSUBS 0.03fF $ **FLOATING
C7603 S.n6920 VSUBS 0.03fF $ **FLOATING
C7604 S.n6921 VSUBS 0.10fF $ **FLOATING
C7605 S.n6922 VSUBS 0.36fF $ **FLOATING
C7606 S.n6923 VSUBS 0.38fF $ **FLOATING
C7607 S.n6924 VSUBS 0.11fF $ **FLOATING
C7608 S.n6925 VSUBS 0.12fF $ **FLOATING
C7609 S.n6926 VSUBS 0.07fF $ **FLOATING
C7610 S.n6927 VSUBS 0.12fF $ **FLOATING
C7611 S.n6928 VSUBS 0.18fF $ **FLOATING
C7612 S.n6929 VSUBS 3.99fF $ **FLOATING
C7613 S.t792 VSUBS 0.02fF
C7614 S.n6930 VSUBS 0.24fF $ **FLOATING
C7615 S.n6931 VSUBS 0.91fF $ **FLOATING
C7616 S.n6932 VSUBS 0.05fF $ **FLOATING
C7617 S.t567 VSUBS 0.02fF
C7618 S.n6933 VSUBS 0.12fF $ **FLOATING
C7619 S.n6934 VSUBS 0.14fF $ **FLOATING
C7620 S.n6936 VSUBS 0.25fF $ **FLOATING
C7621 S.n6937 VSUBS 0.09fF $ **FLOATING
C7622 S.n6938 VSUBS 0.21fF $ **FLOATING
C7623 S.n6939 VSUBS 1.28fF $ **FLOATING
C7624 S.n6940 VSUBS 0.53fF $ **FLOATING
C7625 S.n6941 VSUBS 1.88fF $ **FLOATING
C7626 S.n6942 VSUBS 0.12fF $ **FLOATING
C7627 S.t607 VSUBS 0.02fF
C7628 S.n6943 VSUBS 0.14fF $ **FLOATING
C7629 S.t1424 VSUBS 0.02fF
C7630 S.n6945 VSUBS 0.24fF $ **FLOATING
C7631 S.n6946 VSUBS 0.36fF $ **FLOATING
C7632 S.n6947 VSUBS 0.61fF $ **FLOATING
C7633 S.n6948 VSUBS 1.58fF $ **FLOATING
C7634 S.n6949 VSUBS 2.45fF $ **FLOATING
C7635 S.t1706 VSUBS 0.02fF
C7636 S.n6950 VSUBS 0.24fF $ **FLOATING
C7637 S.n6951 VSUBS 0.91fF $ **FLOATING
C7638 S.n6952 VSUBS 0.05fF $ **FLOATING
C7639 S.t1476 VSUBS 0.02fF
C7640 S.n6953 VSUBS 0.12fF $ **FLOATING
C7641 S.n6954 VSUBS 0.14fF $ **FLOATING
C7642 S.n6956 VSUBS 1.89fF $ **FLOATING
C7643 S.n6957 VSUBS 0.06fF $ **FLOATING
C7644 S.n6958 VSUBS 0.03fF $ **FLOATING
C7645 S.n6959 VSUBS 0.04fF $ **FLOATING
C7646 S.n6960 VSUBS 0.99fF $ **FLOATING
C7647 S.n6961 VSUBS 0.02fF $ **FLOATING
C7648 S.n6962 VSUBS 0.01fF $ **FLOATING
C7649 S.n6963 VSUBS 0.02fF $ **FLOATING
C7650 S.n6964 VSUBS 0.08fF $ **FLOATING
C7651 S.n6965 VSUBS 0.36fF $ **FLOATING
C7652 S.n6966 VSUBS 1.85fF $ **FLOATING
C7653 S.t1046 VSUBS 0.02fF
C7654 S.n6967 VSUBS 0.24fF $ **FLOATING
C7655 S.n6968 VSUBS 0.36fF $ **FLOATING
C7656 S.n6969 VSUBS 0.61fF $ **FLOATING
C7657 S.n6970 VSUBS 0.12fF $ **FLOATING
C7658 S.t230 VSUBS 0.02fF
C7659 S.n6971 VSUBS 0.14fF $ **FLOATING
C7660 S.n6973 VSUBS 0.70fF $ **FLOATING
C7661 S.n6974 VSUBS 0.23fF $ **FLOATING
C7662 S.n6975 VSUBS 0.23fF $ **FLOATING
C7663 S.n6976 VSUBS 0.70fF $ **FLOATING
C7664 S.n6977 VSUBS 1.16fF $ **FLOATING
C7665 S.n6978 VSUBS 0.22fF $ **FLOATING
C7666 S.n6979 VSUBS 0.25fF $ **FLOATING
C7667 S.n6980 VSUBS 0.09fF $ **FLOATING
C7668 S.n6981 VSUBS 1.88fF $ **FLOATING
C7669 S.t1326 VSUBS 0.02fF
C7670 S.n6982 VSUBS 0.24fF $ **FLOATING
C7671 S.n6983 VSUBS 0.91fF $ **FLOATING
C7672 S.n6984 VSUBS 0.05fF $ **FLOATING
C7673 S.t1103 VSUBS 0.02fF
C7674 S.n6985 VSUBS 0.12fF $ **FLOATING
C7675 S.n6986 VSUBS 0.14fF $ **FLOATING
C7676 S.n6988 VSUBS 20.78fF $ **FLOATING
C7677 S.n6989 VSUBS 0.06fF $ **FLOATING
C7678 S.n6990 VSUBS 0.20fF $ **FLOATING
C7679 S.n6991 VSUBS 0.09fF $ **FLOATING
C7680 S.n6992 VSUBS 0.21fF $ **FLOATING
C7681 S.n6993 VSUBS 0.10fF $ **FLOATING
C7682 S.n6994 VSUBS 0.30fF $ **FLOATING
C7683 S.n6995 VSUBS 0.69fF $ **FLOATING
C7684 S.n6996 VSUBS 0.45fF $ **FLOATING
C7685 S.n6997 VSUBS 2.33fF $ **FLOATING
C7686 S.n6998 VSUBS 0.12fF $ **FLOATING
C7687 S.t1081 VSUBS 0.02fF
C7688 S.n6999 VSUBS 0.14fF $ **FLOATING
C7689 S.t1895 VSUBS 0.02fF
C7690 S.n7001 VSUBS 0.24fF $ **FLOATING
C7691 S.n7002 VSUBS 0.36fF $ **FLOATING
C7692 S.n7003 VSUBS 0.61fF $ **FLOATING
C7693 S.n7004 VSUBS 1.90fF $ **FLOATING
C7694 S.n7005 VSUBS 0.17fF $ **FLOATING
C7695 S.n7006 VSUBS 0.76fF $ **FLOATING
C7696 S.n7007 VSUBS 0.25fF $ **FLOATING
C7697 S.n7008 VSUBS 0.30fF $ **FLOATING
C7698 S.n7009 VSUBS 0.32fF $ **FLOATING
C7699 S.n7010 VSUBS 0.47fF $ **FLOATING
C7700 S.n7011 VSUBS 0.16fF $ **FLOATING
C7701 S.n7012 VSUBS 1.93fF $ **FLOATING
C7702 S.t1949 VSUBS 0.02fF
C7703 S.n7013 VSUBS 0.12fF $ **FLOATING
C7704 S.n7014 VSUBS 0.14fF $ **FLOATING
C7705 S.t2177 VSUBS 0.02fF
C7706 S.n7016 VSUBS 0.24fF $ **FLOATING
C7707 S.n7017 VSUBS 0.91fF $ **FLOATING
C7708 S.n7018 VSUBS 0.05fF $ **FLOATING
C7709 S.n7019 VSUBS 1.88fF $ **FLOATING
C7710 S.n7020 VSUBS 0.12fF $ **FLOATING
C7711 S.t1578 VSUBS 0.02fF
C7712 S.n7021 VSUBS 0.14fF $ **FLOATING
C7713 S.t2452 VSUBS 0.02fF
C7714 S.n7023 VSUBS 0.12fF $ **FLOATING
C7715 S.n7024 VSUBS 0.14fF $ **FLOATING
C7716 S.t168 VSUBS 0.02fF
C7717 S.n7026 VSUBS 0.24fF $ **FLOATING
C7718 S.n7027 VSUBS 0.91fF $ **FLOATING
C7719 S.n7028 VSUBS 0.05fF $ **FLOATING
C7720 S.t2399 VSUBS 0.02fF
C7721 S.n7029 VSUBS 0.24fF $ **FLOATING
C7722 S.n7030 VSUBS 0.36fF $ **FLOATING
C7723 S.n7031 VSUBS 0.61fF $ **FLOATING
C7724 S.n7032 VSUBS 0.32fF $ **FLOATING
C7725 S.n7033 VSUBS 1.09fF $ **FLOATING
C7726 S.n7034 VSUBS 0.15fF $ **FLOATING
C7727 S.n7035 VSUBS 2.10fF $ **FLOATING
C7728 S.n7036 VSUBS 2.94fF $ **FLOATING
C7729 S.n7037 VSUBS 1.88fF $ **FLOATING
C7730 S.n7038 VSUBS 0.12fF $ **FLOATING
C7731 S.t1016 VSUBS 0.02fF
C7732 S.n7039 VSUBS 0.14fF $ **FLOATING
C7733 S.t1826 VSUBS 0.02fF
C7734 S.n7041 VSUBS 0.24fF $ **FLOATING
C7735 S.n7042 VSUBS 0.36fF $ **FLOATING
C7736 S.n7043 VSUBS 0.61fF $ **FLOATING
C7737 S.n7044 VSUBS 0.92fF $ **FLOATING
C7738 S.n7045 VSUBS 0.32fF $ **FLOATING
C7739 S.n7046 VSUBS 0.92fF $ **FLOATING
C7740 S.n7047 VSUBS 1.09fF $ **FLOATING
C7741 S.n7048 VSUBS 0.15fF $ **FLOATING
C7742 S.n7049 VSUBS 4.96fF $ **FLOATING
C7743 S.t1884 VSUBS 0.02fF
C7744 S.n7050 VSUBS 0.12fF $ **FLOATING
C7745 S.n7051 VSUBS 0.14fF $ **FLOATING
C7746 S.t2113 VSUBS 0.02fF
C7747 S.n7053 VSUBS 0.24fF $ **FLOATING
C7748 S.n7054 VSUBS 0.91fF $ **FLOATING
C7749 S.n7055 VSUBS 0.05fF $ **FLOATING
C7750 S.n7056 VSUBS 1.88fF $ **FLOATING
C7751 S.n7057 VSUBS 2.67fF $ **FLOATING
C7752 S.t43 VSUBS 0.02fF
C7753 S.n7058 VSUBS 0.24fF $ **FLOATING
C7754 S.n7059 VSUBS 0.36fF $ **FLOATING
C7755 S.n7060 VSUBS 0.61fF $ **FLOATING
C7756 S.n7061 VSUBS 0.12fF $ **FLOATING
C7757 S.t1792 VSUBS 0.02fF
C7758 S.n7062 VSUBS 0.14fF $ **FLOATING
C7759 S.n7064 VSUBS 1.88fF $ **FLOATING
C7760 S.n7065 VSUBS 2.67fF $ **FLOATING
C7761 S.t662 VSUBS 0.02fF
C7762 S.n7066 VSUBS 0.24fF $ **FLOATING
C7763 S.n7067 VSUBS 0.36fF $ **FLOATING
C7764 S.n7068 VSUBS 0.61fF $ **FLOATING
C7765 S.t954 VSUBS 0.02fF
C7766 S.n7069 VSUBS 0.24fF $ **FLOATING
C7767 S.n7070 VSUBS 0.91fF $ **FLOATING
C7768 S.n7071 VSUBS 0.05fF $ **FLOATING
C7769 S.t711 VSUBS 0.02fF
C7770 S.n7072 VSUBS 0.12fF $ **FLOATING
C7771 S.n7073 VSUBS 0.14fF $ **FLOATING
C7772 S.n7075 VSUBS 0.12fF $ **FLOATING
C7773 S.t2370 VSUBS 0.02fF
C7774 S.n7076 VSUBS 0.14fF $ **FLOATING
C7775 S.n7078 VSUBS 2.30fF $ **FLOATING
C7776 S.n7079 VSUBS 2.94fF $ **FLOATING
C7777 S.n7080 VSUBS 5.16fF $ **FLOATING
C7778 S.t131 VSUBS 0.02fF
C7779 S.n7081 VSUBS 0.12fF $ **FLOATING
C7780 S.n7082 VSUBS 0.14fF $ **FLOATING
C7781 S.t381 VSUBS 0.02fF
C7782 S.n7084 VSUBS 0.24fF $ **FLOATING
C7783 S.n7085 VSUBS 0.91fF $ **FLOATING
C7784 S.n7086 VSUBS 0.05fF $ **FLOATING
C7785 S.n7087 VSUBS 1.88fF $ **FLOATING
C7786 S.n7088 VSUBS 2.67fF $ **FLOATING
C7787 S.t866 VSUBS 0.02fF
C7788 S.n7089 VSUBS 0.24fF $ **FLOATING
C7789 S.n7090 VSUBS 0.36fF $ **FLOATING
C7790 S.n7091 VSUBS 0.61fF $ **FLOATING
C7791 S.n7092 VSUBS 0.12fF $ **FLOATING
C7792 S.t2577 VSUBS 0.02fF
C7793 S.n7093 VSUBS 0.14fF $ **FLOATING
C7794 S.n7095 VSUBS 5.17fF $ **FLOATING
C7795 S.t928 VSUBS 0.02fF
C7796 S.n7096 VSUBS 0.12fF $ **FLOATING
C7797 S.n7097 VSUBS 0.14fF $ **FLOATING
C7798 S.t1167 VSUBS 0.02fF
C7799 S.n7099 VSUBS 0.24fF $ **FLOATING
C7800 S.n7100 VSUBS 0.91fF $ **FLOATING
C7801 S.n7101 VSUBS 0.05fF $ **FLOATING
C7802 S.n7102 VSUBS 1.88fF $ **FLOATING
C7803 S.n7103 VSUBS 0.12fF $ **FLOATING
C7804 S.t1663 VSUBS 0.02fF
C7805 S.n7104 VSUBS 0.14fF $ **FLOATING
C7806 S.t1466 VSUBS 0.02fF
C7807 S.n7106 VSUBS 0.24fF $ **FLOATING
C7808 S.n7107 VSUBS 0.36fF $ **FLOATING
C7809 S.n7108 VSUBS 0.61fF $ **FLOATING
C7810 S.n7109 VSUBS 2.67fF $ **FLOATING
C7811 S.n7110 VSUBS 5.17fF $ **FLOATING
C7812 S.t1845 VSUBS 0.02fF
C7813 S.n7111 VSUBS 0.12fF $ **FLOATING
C7814 S.n7112 VSUBS 0.14fF $ **FLOATING
C7815 S.t2309 VSUBS 0.02fF
C7816 S.n7114 VSUBS 0.24fF $ **FLOATING
C7817 S.n7115 VSUBS 0.91fF $ **FLOATING
C7818 S.n7116 VSUBS 0.05fF $ **FLOATING
C7819 S.n7117 VSUBS 1.88fF $ **FLOATING
C7820 S.n7118 VSUBS 2.67fF $ **FLOATING
C7821 S.t2254 VSUBS 0.02fF
C7822 S.n7119 VSUBS 0.24fF $ **FLOATING
C7823 S.n7120 VSUBS 0.36fF $ **FLOATING
C7824 S.n7121 VSUBS 0.61fF $ **FLOATING
C7825 S.n7122 VSUBS 0.12fF $ **FLOATING
C7826 S.t2453 VSUBS 0.02fF
C7827 S.n7123 VSUBS 0.14fF $ **FLOATING
C7828 S.n7125 VSUBS 5.17fF $ **FLOATING
C7829 S.t797 VSUBS 0.02fF
C7830 S.n7126 VSUBS 0.12fF $ **FLOATING
C7831 S.n7127 VSUBS 0.14fF $ **FLOATING
C7832 S.t577 VSUBS 0.02fF
C7833 S.n7129 VSUBS 0.24fF $ **FLOATING
C7834 S.n7130 VSUBS 0.91fF $ **FLOATING
C7835 S.n7131 VSUBS 0.05fF $ **FLOATING
C7836 S.n7132 VSUBS 1.88fF $ **FLOATING
C7837 S.n7133 VSUBS 2.67fF $ **FLOATING
C7838 S.t524 VSUBS 0.02fF
C7839 S.n7134 VSUBS 0.24fF $ **FLOATING
C7840 S.n7135 VSUBS 0.36fF $ **FLOATING
C7841 S.n7136 VSUBS 0.61fF $ **FLOATING
C7842 S.n7137 VSUBS 0.12fF $ **FLOATING
C7843 S.t709 VSUBS 0.02fF
C7844 S.n7138 VSUBS 0.14fF $ **FLOATING
C7845 S.n7140 VSUBS 5.17fF $ **FLOATING
C7846 S.t1579 VSUBS 0.02fF
C7847 S.n7141 VSUBS 0.12fF $ **FLOATING
C7848 S.n7142 VSUBS 0.14fF $ **FLOATING
C7849 S.t1368 VSUBS 0.02fF
C7850 S.n7144 VSUBS 0.24fF $ **FLOATING
C7851 S.n7145 VSUBS 0.91fF $ **FLOATING
C7852 S.n7146 VSUBS 0.05fF $ **FLOATING
C7853 S.n7147 VSUBS 1.88fF $ **FLOATING
C7854 S.n7148 VSUBS 2.67fF $ **FLOATING
C7855 S.t1309 VSUBS 0.02fF
C7856 S.n7149 VSUBS 0.24fF $ **FLOATING
C7857 S.n7150 VSUBS 0.36fF $ **FLOATING
C7858 S.n7151 VSUBS 0.61fF $ **FLOATING
C7859 S.n7152 VSUBS 0.12fF $ **FLOATING
C7860 S.t1504 VSUBS 0.02fF
C7861 S.n7153 VSUBS 0.14fF $ **FLOATING
C7862 S.n7155 VSUBS 4.89fF $ **FLOATING
C7863 S.t2369 VSUBS 0.02fF
C7864 S.n7156 VSUBS 0.12fF $ **FLOATING
C7865 S.n7157 VSUBS 0.14fF $ **FLOATING
C7866 S.t2153 VSUBS 0.02fF
C7867 S.n7159 VSUBS 0.24fF $ **FLOATING
C7868 S.n7160 VSUBS 0.91fF $ **FLOATING
C7869 S.n7161 VSUBS 0.05fF $ **FLOATING
C7870 S.n7162 VSUBS 1.88fF $ **FLOATING
C7871 S.n7163 VSUBS 2.67fF $ **FLOATING
C7872 S.t2096 VSUBS 0.02fF
C7873 S.n7164 VSUBS 0.24fF $ **FLOATING
C7874 S.n7165 VSUBS 0.36fF $ **FLOATING
C7875 S.n7166 VSUBS 0.61fF $ **FLOATING
C7876 S.n7167 VSUBS 0.12fF $ **FLOATING
C7877 S.t2290 VSUBS 0.02fF
C7878 S.n7168 VSUBS 0.14fF $ **FLOATING
C7879 S.n7170 VSUBS 1.88fF $ **FLOATING
C7880 S.n7171 VSUBS 2.68fF $ **FLOATING
C7881 S.t2125 VSUBS 0.02fF
C7882 S.n7172 VSUBS 0.24fF $ **FLOATING
C7883 S.n7173 VSUBS 0.36fF $ **FLOATING
C7884 S.n7174 VSUBS 0.61fF $ **FLOATING
C7885 S.t2464 VSUBS 0.02fF
C7886 S.n7175 VSUBS 1.22fF $ **FLOATING
C7887 S.n7176 VSUBS 0.36fF $ **FLOATING
C7888 S.n7177 VSUBS 1.22fF $ **FLOATING
C7889 S.n7178 VSUBS 0.61fF $ **FLOATING
C7890 S.n7179 VSUBS 0.35fF $ **FLOATING
C7891 S.n7180 VSUBS 0.63fF $ **FLOATING
C7892 S.n7181 VSUBS 1.15fF $ **FLOATING
C7893 S.n7182 VSUBS 3.00fF $ **FLOATING
C7894 S.n7183 VSUBS 0.59fF $ **FLOATING
C7895 S.n7184 VSUBS 0.01fF $ **FLOATING
C7896 S.n7185 VSUBS 0.97fF $ **FLOATING
C7897 S.t235 VSUBS 21.42fF
C7898 S.n7186 VSUBS 20.29fF $ **FLOATING
C7899 S.n7188 VSUBS 0.38fF $ **FLOATING
C7900 S.n7189 VSUBS 0.23fF $ **FLOATING
C7901 S.n7190 VSUBS 2.79fF $ **FLOATING
C7902 S.n7191 VSUBS 2.46fF $ **FLOATING
C7903 S.n7192 VSUBS 4.00fF $ **FLOATING
C7904 S.n7193 VSUBS 0.25fF $ **FLOATING
C7905 S.n7194 VSUBS 0.01fF $ **FLOATING
C7906 S.t1649 VSUBS 0.02fF
C7907 S.n7195 VSUBS 0.26fF $ **FLOATING
C7908 S.t242 VSUBS 0.02fF
C7909 S.n7196 VSUBS 0.95fF $ **FLOATING
C7910 S.n7197 VSUBS 0.71fF $ **FLOATING
C7911 S.n7198 VSUBS 1.89fF $ **FLOATING
C7912 S.n7199 VSUBS 1.88fF $ **FLOATING
C7913 S.t722 VSUBS 0.02fF
C7914 S.n7200 VSUBS 0.24fF $ **FLOATING
C7915 S.n7201 VSUBS 0.36fF $ **FLOATING
C7916 S.n7202 VSUBS 0.61fF $ **FLOATING
C7917 S.n7203 VSUBS 0.12fF $ **FLOATING
C7918 S.t2432 VSUBS 0.02fF
C7919 S.n7204 VSUBS 0.14fF $ **FLOATING
C7920 S.n7206 VSUBS 1.16fF $ **FLOATING
C7921 S.n7207 VSUBS 0.22fF $ **FLOATING
C7922 S.n7208 VSUBS 0.25fF $ **FLOATING
C7923 S.n7209 VSUBS 0.09fF $ **FLOATING
C7924 S.n7210 VSUBS 1.88fF $ **FLOATING
C7925 S.t1027 VSUBS 0.02fF
C7926 S.n7211 VSUBS 0.24fF $ **FLOATING
C7927 S.n7212 VSUBS 0.91fF $ **FLOATING
C7928 S.n7213 VSUBS 0.05fF $ **FLOATING
C7929 S.t779 VSUBS 0.02fF
C7930 S.n7214 VSUBS 0.12fF $ **FLOATING
C7931 S.n7215 VSUBS 0.14fF $ **FLOATING
C7932 S.n7217 VSUBS 0.78fF $ **FLOATING
C7933 S.n7218 VSUBS 1.94fF $ **FLOATING
C7934 S.n7219 VSUBS 1.88fF $ **FLOATING
C7935 S.n7220 VSUBS 0.12fF $ **FLOATING
C7936 S.t830 VSUBS 0.02fF
C7937 S.n7221 VSUBS 0.14fF $ **FLOATING
C7938 S.t1515 VSUBS 0.02fF
C7939 S.n7223 VSUBS 0.24fF $ **FLOATING
C7940 S.n7224 VSUBS 0.36fF $ **FLOATING
C7941 S.n7225 VSUBS 0.61fF $ **FLOATING
C7942 S.n7226 VSUBS 1.84fF $ **FLOATING
C7943 S.n7227 VSUBS 2.99fF $ **FLOATING
C7944 S.t1808 VSUBS 0.02fF
C7945 S.n7228 VSUBS 0.24fF $ **FLOATING
C7946 S.n7229 VSUBS 0.91fF $ **FLOATING
C7947 S.n7230 VSUBS 0.05fF $ **FLOATING
C7948 S.t1563 VSUBS 0.02fF
C7949 S.n7231 VSUBS 0.12fF $ **FLOATING
C7950 S.n7232 VSUBS 0.14fF $ **FLOATING
C7951 S.n7234 VSUBS 1.89fF $ **FLOATING
C7952 S.n7235 VSUBS 1.88fF $ **FLOATING
C7953 S.t2429 VSUBS 0.02fF
C7954 S.n7236 VSUBS 0.24fF $ **FLOATING
C7955 S.n7237 VSUBS 0.36fF $ **FLOATING
C7956 S.n7238 VSUBS 0.61fF $ **FLOATING
C7957 S.n7239 VSUBS 0.12fF $ **FLOATING
C7958 S.t1612 VSUBS 0.02fF
C7959 S.n7240 VSUBS 0.14fF $ **FLOATING
C7960 S.n7242 VSUBS 1.16fF $ **FLOATING
C7961 S.n7243 VSUBS 0.22fF $ **FLOATING
C7962 S.n7244 VSUBS 0.25fF $ **FLOATING
C7963 S.n7245 VSUBS 0.09fF $ **FLOATING
C7964 S.n7246 VSUBS 1.88fF $ **FLOATING
C7965 S.t200 VSUBS 0.02fF
C7966 S.n7247 VSUBS 0.24fF $ **FLOATING
C7967 S.n7248 VSUBS 0.91fF $ **FLOATING
C7968 S.n7249 VSUBS 0.05fF $ **FLOATING
C7969 S.t2484 VSUBS 0.02fF
C7970 S.n7250 VSUBS 0.12fF $ **FLOATING
C7971 S.n7251 VSUBS 0.14fF $ **FLOATING
C7972 S.n7253 VSUBS 0.78fF $ **FLOATING
C7973 S.n7254 VSUBS 1.94fF $ **FLOATING
C7974 S.n7255 VSUBS 1.88fF $ **FLOATING
C7975 S.n7256 VSUBS 0.12fF $ **FLOATING
C7976 S.t1237 VSUBS 0.02fF
C7977 S.n7257 VSUBS 0.14fF $ **FLOATING
C7978 S.t2054 VSUBS 0.02fF
C7979 S.n7259 VSUBS 0.24fF $ **FLOATING
C7980 S.n7260 VSUBS 0.36fF $ **FLOATING
C7981 S.n7261 VSUBS 0.61fF $ **FLOATING
C7982 S.n7262 VSUBS 1.84fF $ **FLOATING
C7983 S.n7263 VSUBS 2.99fF $ **FLOATING
C7984 S.t2326 VSUBS 0.02fF
C7985 S.n7264 VSUBS 0.24fF $ **FLOATING
C7986 S.n7265 VSUBS 0.91fF $ **FLOATING
C7987 S.n7266 VSUBS 0.05fF $ **FLOATING
C7988 S.t2102 VSUBS 0.02fF
C7989 S.n7267 VSUBS 0.12fF $ **FLOATING
C7990 S.n7268 VSUBS 0.14fF $ **FLOATING
C7991 S.n7270 VSUBS 1.89fF $ **FLOATING
C7992 S.n7271 VSUBS 1.75fF $ **FLOATING
C7993 S.t318 VSUBS 0.02fF
C7994 S.n7272 VSUBS 0.24fF $ **FLOATING
C7995 S.n7273 VSUBS 0.36fF $ **FLOATING
C7996 S.n7274 VSUBS 0.61fF $ **FLOATING
C7997 S.n7275 VSUBS 0.12fF $ **FLOATING
C7998 S.t2020 VSUBS 0.02fF
C7999 S.n7276 VSUBS 0.14fF $ **FLOATING
C8000 S.n7278 VSUBS 1.16fF $ **FLOATING
C8001 S.n7279 VSUBS 0.22fF $ **FLOATING
C8002 S.n7280 VSUBS 0.25fF $ **FLOATING
C8003 S.n7281 VSUBS 0.09fF $ **FLOATING
C8004 S.n7282 VSUBS 2.44fF $ **FLOATING
C8005 S.t590 VSUBS 0.02fF
C8006 S.n7283 VSUBS 0.24fF $ **FLOATING
C8007 S.n7284 VSUBS 0.91fF $ **FLOATING
C8008 S.n7285 VSUBS 0.05fF $ **FLOATING
C8009 S.t372 VSUBS 0.02fF
C8010 S.n7286 VSUBS 0.12fF $ **FLOATING
C8011 S.n7287 VSUBS 0.14fF $ **FLOATING
C8012 S.n7289 VSUBS 1.88fF $ **FLOATING
C8013 S.n7290 VSUBS 0.48fF $ **FLOATING
C8014 S.n7291 VSUBS 0.09fF $ **FLOATING
C8015 S.n7292 VSUBS 0.33fF $ **FLOATING
C8016 S.n7293 VSUBS 0.30fF $ **FLOATING
C8017 S.n7294 VSUBS 0.77fF $ **FLOATING
C8018 S.n7295 VSUBS 0.59fF $ **FLOATING
C8019 S.t1109 VSUBS 0.02fF
C8020 S.n7296 VSUBS 0.24fF $ **FLOATING
C8021 S.n7297 VSUBS 0.36fF $ **FLOATING
C8022 S.n7298 VSUBS 0.61fF $ **FLOATING
C8023 S.n7299 VSUBS 0.12fF $ **FLOATING
C8024 S.t294 VSUBS 0.02fF
C8025 S.n7300 VSUBS 0.14fF $ **FLOATING
C8026 S.n7302 VSUBS 2.61fF $ **FLOATING
C8027 S.n7303 VSUBS 2.15fF $ **FLOATING
C8028 S.t1384 VSUBS 0.02fF
C8029 S.n7304 VSUBS 0.24fF $ **FLOATING
C8030 S.n7305 VSUBS 0.91fF $ **FLOATING
C8031 S.n7306 VSUBS 0.05fF $ **FLOATING
C8032 S.t1161 VSUBS 0.02fF
C8033 S.n7307 VSUBS 0.12fF $ **FLOATING
C8034 S.n7308 VSUBS 0.14fF $ **FLOATING
C8035 S.n7310 VSUBS 0.78fF $ **FLOATING
C8036 S.n7311 VSUBS 2.30fF $ **FLOATING
C8037 S.n7312 VSUBS 1.88fF $ **FLOATING
C8038 S.n7313 VSUBS 0.12fF $ **FLOATING
C8039 S.t1206 VSUBS 0.02fF
C8040 S.n7314 VSUBS 0.14fF $ **FLOATING
C8041 S.t1888 VSUBS 0.02fF
C8042 S.n7316 VSUBS 0.24fF $ **FLOATING
C8043 S.n7317 VSUBS 0.36fF $ **FLOATING
C8044 S.n7318 VSUBS 0.61fF $ **FLOATING
C8045 S.n7319 VSUBS 1.39fF $ **FLOATING
C8046 S.n7320 VSUBS 0.71fF $ **FLOATING
C8047 S.n7321 VSUBS 1.14fF $ **FLOATING
C8048 S.n7322 VSUBS 0.35fF $ **FLOATING
C8049 S.n7323 VSUBS 2.02fF $ **FLOATING
C8050 S.t2169 VSUBS 0.02fF
C8051 S.n7324 VSUBS 0.24fF $ **FLOATING
C8052 S.n7325 VSUBS 0.91fF $ **FLOATING
C8053 S.n7326 VSUBS 0.05fF $ **FLOATING
C8054 S.t1945 VSUBS 0.02fF
C8055 S.n7327 VSUBS 0.12fF $ **FLOATING
C8056 S.n7328 VSUBS 0.14fF $ **FLOATING
C8057 S.n7330 VSUBS 1.89fF $ **FLOATING
C8058 S.n7331 VSUBS 1.88fF $ **FLOATING
C8059 S.t1613 VSUBS 0.02fF
C8060 S.n7332 VSUBS 0.24fF $ **FLOATING
C8061 S.n7333 VSUBS 0.36fF $ **FLOATING
C8062 S.n7334 VSUBS 0.61fF $ **FLOATING
C8063 S.n7335 VSUBS 0.12fF $ **FLOATING
C8064 S.t796 VSUBS 0.02fF
C8065 S.n7336 VSUBS 0.14fF $ **FLOATING
C8066 S.n7338 VSUBS 1.16fF $ **FLOATING
C8067 S.n7339 VSUBS 0.22fF $ **FLOATING
C8068 S.n7340 VSUBS 0.25fF $ **FLOATING
C8069 S.n7341 VSUBS 0.09fF $ **FLOATING
C8070 S.n7342 VSUBS 1.88fF $ **FLOATING
C8071 S.t1915 VSUBS 0.02fF
C8072 S.n7343 VSUBS 0.24fF $ **FLOATING
C8073 S.n7344 VSUBS 0.91fF $ **FLOATING
C8074 S.n7345 VSUBS 0.05fF $ **FLOATING
C8075 S.t336 VSUBS 0.02fF
C8076 S.n7346 VSUBS 0.12fF $ **FLOATING
C8077 S.n7347 VSUBS 0.14fF $ **FLOATING
C8078 S.n7349 VSUBS 20.78fF $ **FLOATING
C8079 S.n7350 VSUBS 1.88fF $ **FLOATING
C8080 S.n7351 VSUBS 2.67fF $ **FLOATING
C8081 S.t1452 VSUBS 0.02fF
C8082 S.n7352 VSUBS 0.24fF $ **FLOATING
C8083 S.n7353 VSUBS 0.36fF $ **FLOATING
C8084 S.n7354 VSUBS 0.61fF $ **FLOATING
C8085 S.n7355 VSUBS 0.12fF $ **FLOATING
C8086 S.t636 VSUBS 0.02fF
C8087 S.n7356 VSUBS 0.14fF $ **FLOATING
C8088 S.n7358 VSUBS 2.80fF $ **FLOATING
C8089 S.n7359 VSUBS 2.30fF $ **FLOATING
C8090 S.t1503 VSUBS 0.02fF
C8091 S.n7360 VSUBS 0.12fF $ **FLOATING
C8092 S.n7361 VSUBS 0.14fF $ **FLOATING
C8093 S.t1737 VSUBS 0.02fF
C8094 S.n7363 VSUBS 0.24fF $ **FLOATING
C8095 S.n7364 VSUBS 0.91fF $ **FLOATING
C8096 S.n7365 VSUBS 0.05fF $ **FLOATING
C8097 S.n7366 VSUBS 2.80fF $ **FLOATING
C8098 S.n7367 VSUBS 1.88fF $ **FLOATING
C8099 S.n7368 VSUBS 0.12fF $ **FLOATING
C8100 S.t1547 VSUBS 0.02fF
C8101 S.n7369 VSUBS 0.14fF $ **FLOATING
C8102 S.t2240 VSUBS 0.02fF
C8103 S.n7371 VSUBS 0.24fF $ **FLOATING
C8104 S.n7372 VSUBS 0.36fF $ **FLOATING
C8105 S.n7373 VSUBS 0.61fF $ **FLOATING
C8106 S.n7374 VSUBS 2.67fF $ **FLOATING
C8107 S.n7375 VSUBS 2.30fF $ **FLOATING
C8108 S.t2289 VSUBS 0.02fF
C8109 S.n7376 VSUBS 0.12fF $ **FLOATING
C8110 S.n7377 VSUBS 0.14fF $ **FLOATING
C8111 S.t2521 VSUBS 0.02fF
C8112 S.n7379 VSUBS 0.24fF $ **FLOATING
C8113 S.n7380 VSUBS 0.91fF $ **FLOATING
C8114 S.n7381 VSUBS 0.05fF $ **FLOATING
C8115 S.n7382 VSUBS 1.88fF $ **FLOATING
C8116 S.n7383 VSUBS 2.67fF $ **FLOATING
C8117 S.t2278 VSUBS 0.02fF
C8118 S.n7384 VSUBS 0.24fF $ **FLOATING
C8119 S.n7385 VSUBS 0.36fF $ **FLOATING
C8120 S.n7386 VSUBS 0.61fF $ **FLOATING
C8121 S.n7387 VSUBS 0.12fF $ **FLOATING
C8122 S.t2481 VSUBS 0.02fF
C8123 S.n7388 VSUBS 0.14fF $ **FLOATING
C8124 S.n7390 VSUBS 2.80fF $ **FLOATING
C8125 S.n7391 VSUBS 2.30fF $ **FLOATING
C8126 S.t825 VSUBS 0.02fF
C8127 S.n7392 VSUBS 0.12fF $ **FLOATING
C8128 S.n7393 VSUBS 0.14fF $ **FLOATING
C8129 S.t597 VSUBS 0.02fF
C8130 S.n7395 VSUBS 0.24fF $ **FLOATING
C8131 S.n7396 VSUBS 0.91fF $ **FLOATING
C8132 S.n7397 VSUBS 0.05fF $ **FLOATING
C8133 S.n7398 VSUBS 1.88fF $ **FLOATING
C8134 S.n7399 VSUBS 2.67fF $ **FLOATING
C8135 S.t549 VSUBS 0.02fF
C8136 S.n7400 VSUBS 0.24fF $ **FLOATING
C8137 S.n7401 VSUBS 0.36fF $ **FLOATING
C8138 S.n7402 VSUBS 0.61fF $ **FLOATING
C8139 S.n7403 VSUBS 0.12fF $ **FLOATING
C8140 S.t738 VSUBS 0.02fF
C8141 S.n7404 VSUBS 0.14fF $ **FLOATING
C8142 S.n7406 VSUBS 2.80fF $ **FLOATING
C8143 S.n7407 VSUBS 2.30fF $ **FLOATING
C8144 S.t1609 VSUBS 0.02fF
C8145 S.n7408 VSUBS 0.12fF $ **FLOATING
C8146 S.n7409 VSUBS 0.14fF $ **FLOATING
C8147 S.t1390 VSUBS 0.02fF
C8148 S.n7411 VSUBS 0.24fF $ **FLOATING
C8149 S.n7412 VSUBS 0.91fF $ **FLOATING
C8150 S.n7413 VSUBS 0.05fF $ **FLOATING
C8151 S.n7414 VSUBS 1.88fF $ **FLOATING
C8152 S.n7415 VSUBS 2.67fF $ **FLOATING
C8153 S.t1339 VSUBS 0.02fF
C8154 S.n7416 VSUBS 0.24fF $ **FLOATING
C8155 S.n7417 VSUBS 0.36fF $ **FLOATING
C8156 S.n7418 VSUBS 0.61fF $ **FLOATING
C8157 S.n7419 VSUBS 0.12fF $ **FLOATING
C8158 S.t1530 VSUBS 0.02fF
C8159 S.n7420 VSUBS 0.14fF $ **FLOATING
C8160 S.n7422 VSUBS 2.80fF $ **FLOATING
C8161 S.n7423 VSUBS 2.30fF $ **FLOATING
C8162 S.t2397 VSUBS 0.02fF
C8163 S.n7424 VSUBS 0.12fF $ **FLOATING
C8164 S.n7425 VSUBS 0.14fF $ **FLOATING
C8165 S.t2179 VSUBS 0.02fF
C8166 S.n7427 VSUBS 0.24fF $ **FLOATING
C8167 S.n7428 VSUBS 0.91fF $ **FLOATING
C8168 S.n7429 VSUBS 0.05fF $ **FLOATING
C8169 S.n7430 VSUBS 2.73fF $ **FLOATING
C8170 S.n7431 VSUBS 1.59fF $ **FLOATING
C8171 S.n7432 VSUBS 0.12fF $ **FLOATING
C8172 S.t103 VSUBS 0.02fF
C8173 S.n7433 VSUBS 0.14fF $ **FLOATING
C8174 S.t1329 VSUBS 0.02fF
C8175 S.n7435 VSUBS 0.24fF $ **FLOATING
C8176 S.n7436 VSUBS 0.36fF $ **FLOATING
C8177 S.n7437 VSUBS 0.61fF $ **FLOATING
C8178 S.n7438 VSUBS 0.07fF $ **FLOATING
C8179 S.n7439 VSUBS 0.01fF $ **FLOATING
C8180 S.n7440 VSUBS 0.24fF $ **FLOATING
C8181 S.n7441 VSUBS 1.16fF $ **FLOATING
C8182 S.n7442 VSUBS 1.35fF $ **FLOATING
C8183 S.n7443 VSUBS 2.30fF $ **FLOATING
C8184 S.t1449 VSUBS 0.02fF
C8185 S.n7444 VSUBS 0.12fF $ **FLOATING
C8186 S.n7445 VSUBS 0.14fF $ **FLOATING
C8187 S.t206 VSUBS 0.02fF
C8188 S.n7447 VSUBS 0.24fF $ **FLOATING
C8189 S.n7448 VSUBS 0.91fF $ **FLOATING
C8190 S.n7449 VSUBS 0.05fF $ **FLOATING
C8191 S.t102 VSUBS 48.27fF
C8192 S.t443 VSUBS 0.02fF
C8193 S.n7450 VSUBS 0.24fF $ **FLOATING
C8194 S.n7451 VSUBS 0.91fF $ **FLOATING
C8195 S.n7452 VSUBS 0.05fF $ **FLOATING
C8196 S.t660 VSUBS 0.02fF
C8197 S.n7453 VSUBS 0.12fF $ **FLOATING
C8198 S.n7454 VSUBS 0.14fF $ **FLOATING
C8199 S.n7456 VSUBS 0.12fF $ **FLOATING
C8200 S.t2315 VSUBS 0.02fF
C8201 S.n7457 VSUBS 0.14fF $ **FLOATING
C8202 S.n7459 VSUBS 5.17fF $ **FLOATING
C8203 S.n7460 VSUBS 5.44fF $ **FLOATING
C8204 S.t637 VSUBS 0.02fF
C8205 S.n7461 VSUBS 0.12fF $ **FLOATING
C8206 S.n7462 VSUBS 0.14fF $ **FLOATING
C8207 S.t420 VSUBS 0.02fF
C8208 S.n7464 VSUBS 0.24fF $ **FLOATING
C8209 S.n7465 VSUBS 0.91fF $ **FLOATING
C8210 S.n7466 VSUBS 0.05fF $ **FLOATING
C8211 S.t130 VSUBS 47.89fF
C8212 S.t1488 VSUBS 0.02fF
C8213 S.n7467 VSUBS 0.01fF $ **FLOATING
C8214 S.n7468 VSUBS 0.26fF $ **FLOATING
C8215 S.t536 VSUBS 0.02fF
C8216 S.n7470 VSUBS 1.19fF $ **FLOATING
C8217 S.n7471 VSUBS 0.05fF $ **FLOATING
C8218 S.t258 VSUBS 0.02fF
C8219 S.n7472 VSUBS 0.64fF $ **FLOATING
C8220 S.n7473 VSUBS 0.61fF $ **FLOATING
C8221 S.n7474 VSUBS 8.97fF $ **FLOATING
C8222 S.n7475 VSUBS 8.97fF $ **FLOATING
C8223 S.n7476 VSUBS 0.60fF $ **FLOATING
C8224 S.n7477 VSUBS 0.22fF $ **FLOATING
C8225 S.n7478 VSUBS 0.59fF $ **FLOATING
C8226 S.n7479 VSUBS 3.39fF $ **FLOATING
C8227 S.n7480 VSUBS 0.29fF $ **FLOATING
C8228 S.t42 VSUBS 21.42fF
C8229 S.n7481 VSUBS 21.71fF $ **FLOATING
C8230 S.n7482 VSUBS 0.77fF $ **FLOATING
C8231 S.n7483 VSUBS 0.28fF $ **FLOATING
C8232 S.n7484 VSUBS 4.00fF $ **FLOATING
C8233 S.n7485 VSUBS 1.35fF $ **FLOATING
C8234 S.n7486 VSUBS 0.01fF $ **FLOATING
C8235 S.n7487 VSUBS 0.02fF $ **FLOATING
C8236 S.n7488 VSUBS 0.03fF $ **FLOATING
C8237 S.n7489 VSUBS 0.04fF $ **FLOATING
C8238 S.n7490 VSUBS 0.17fF $ **FLOATING
C8239 S.n7491 VSUBS 0.01fF $ **FLOATING
C8240 S.n7492 VSUBS 0.02fF $ **FLOATING
C8241 S.n7493 VSUBS 0.01fF $ **FLOATING
C8242 S.n7494 VSUBS 0.01fF $ **FLOATING
C8243 S.n7495 VSUBS 0.01fF $ **FLOATING
C8244 S.n7496 VSUBS 0.01fF $ **FLOATING
C8245 S.n7497 VSUBS 0.02fF $ **FLOATING
C8246 S.n7498 VSUBS 0.01fF $ **FLOATING
C8247 S.n7499 VSUBS 0.02fF $ **FLOATING
C8248 S.n7500 VSUBS 0.05fF $ **FLOATING
C8249 S.n7501 VSUBS 0.04fF $ **FLOATING
C8250 S.n7502 VSUBS 0.11fF $ **FLOATING
C8251 S.n7503 VSUBS 0.38fF $ **FLOATING
C8252 S.n7504 VSUBS 0.20fF $ **FLOATING
C8253 S.n7505 VSUBS 4.39fF $ **FLOATING
C8254 S.n7506 VSUBS 0.24fF $ **FLOATING
C8255 S.n7507 VSUBS 1.50fF $ **FLOATING
C8256 S.n7508 VSUBS 1.31fF $ **FLOATING
C8257 S.n7509 VSUBS 0.28fF $ **FLOATING
C8258 S.n7510 VSUBS 0.25fF $ **FLOATING
C8259 S.n7511 VSUBS 0.09fF $ **FLOATING
C8260 S.n7512 VSUBS 0.21fF $ **FLOATING
C8261 S.n7513 VSUBS 0.92fF $ **FLOATING
C8262 S.n7514 VSUBS 0.44fF $ **FLOATING
C8263 S.n7515 VSUBS 1.88fF $ **FLOATING
C8264 S.n7516 VSUBS 0.12fF $ **FLOATING
C8265 S.t1290 VSUBS 0.02fF
C8266 S.n7517 VSUBS 0.14fF $ **FLOATING
C8267 S.t2108 VSUBS 0.02fF
C8268 S.n7519 VSUBS 0.24fF $ **FLOATING
C8269 S.n7520 VSUBS 0.36fF $ **FLOATING
C8270 S.n7521 VSUBS 0.61fF $ **FLOATING
C8271 S.n7522 VSUBS 0.02fF $ **FLOATING
C8272 S.n7523 VSUBS 0.01fF $ **FLOATING
C8273 S.n7524 VSUBS 0.02fF $ **FLOATING
C8274 S.n7525 VSUBS 0.08fF $ **FLOATING
C8275 S.n7526 VSUBS 0.06fF $ **FLOATING
C8276 S.n7527 VSUBS 0.03fF $ **FLOATING
C8277 S.n7528 VSUBS 0.04fF $ **FLOATING
C8278 S.n7529 VSUBS 1.00fF $ **FLOATING
C8279 S.n7530 VSUBS 0.36fF $ **FLOATING
C8280 S.n7531 VSUBS 1.87fF $ **FLOATING
C8281 S.n7532 VSUBS 1.99fF $ **FLOATING
C8282 S.t2382 VSUBS 0.02fF
C8283 S.n7533 VSUBS 0.24fF $ **FLOATING
C8284 S.n7534 VSUBS 0.91fF $ **FLOATING
C8285 S.n7535 VSUBS 0.05fF $ **FLOATING
C8286 S.t2158 VSUBS 0.02fF
C8287 S.n7536 VSUBS 0.12fF $ **FLOATING
C8288 S.n7537 VSUBS 0.14fF $ **FLOATING
C8289 S.n7539 VSUBS 1.89fF $ **FLOATING
C8290 S.n7540 VSUBS 0.06fF $ **FLOATING
C8291 S.n7541 VSUBS 0.03fF $ **FLOATING
C8292 S.n7542 VSUBS 0.04fF $ **FLOATING
C8293 S.n7543 VSUBS 0.99fF $ **FLOATING
C8294 S.n7544 VSUBS 0.02fF $ **FLOATING
C8295 S.n7545 VSUBS 0.01fF $ **FLOATING
C8296 S.n7546 VSUBS 0.02fF $ **FLOATING
C8297 S.n7547 VSUBS 0.08fF $ **FLOATING
C8298 S.n7548 VSUBS 0.36fF $ **FLOATING
C8299 S.n7549 VSUBS 1.85fF $ **FLOATING
C8300 S.t500 VSUBS 0.02fF
C8301 S.n7550 VSUBS 0.24fF $ **FLOATING
C8302 S.n7551 VSUBS 0.36fF $ **FLOATING
C8303 S.n7552 VSUBS 0.61fF $ **FLOATING
C8304 S.n7553 VSUBS 0.12fF $ **FLOATING
C8305 S.t2203 VSUBS 0.02fF
C8306 S.n7554 VSUBS 0.14fF $ **FLOATING
C8307 S.n7556 VSUBS 0.70fF $ **FLOATING
C8308 S.n7557 VSUBS 0.23fF $ **FLOATING
C8309 S.n7558 VSUBS 0.23fF $ **FLOATING
C8310 S.n7559 VSUBS 0.70fF $ **FLOATING
C8311 S.n7560 VSUBS 1.16fF $ **FLOATING
C8312 S.n7561 VSUBS 0.22fF $ **FLOATING
C8313 S.n7562 VSUBS 0.25fF $ **FLOATING
C8314 S.n7563 VSUBS 0.09fF $ **FLOATING
C8315 S.n7564 VSUBS 1.88fF $ **FLOATING
C8316 S.t775 VSUBS 0.02fF
C8317 S.n7565 VSUBS 0.24fF $ **FLOATING
C8318 S.n7566 VSUBS 0.91fF $ **FLOATING
C8319 S.n7567 VSUBS 0.05fF $ **FLOATING
C8320 S.t551 VSUBS 0.02fF
C8321 S.n7568 VSUBS 0.12fF $ **FLOATING
C8322 S.n7569 VSUBS 0.14fF $ **FLOATING
C8323 S.n7571 VSUBS 0.25fF $ **FLOATING
C8324 S.n7572 VSUBS 0.09fF $ **FLOATING
C8325 S.n7573 VSUBS 0.21fF $ **FLOATING
C8326 S.n7574 VSUBS 0.92fF $ **FLOATING
C8327 S.n7575 VSUBS 0.44fF $ **FLOATING
C8328 S.n7576 VSUBS 1.88fF $ **FLOATING
C8329 S.n7577 VSUBS 0.12fF $ **FLOATING
C8330 S.t1813 VSUBS 0.02fF
C8331 S.n7578 VSUBS 0.14fF $ **FLOATING
C8332 S.t80 VSUBS 0.02fF
C8333 S.n7580 VSUBS 0.24fF $ **FLOATING
C8334 S.n7581 VSUBS 0.36fF $ **FLOATING
C8335 S.n7582 VSUBS 0.61fF $ **FLOATING
C8336 S.n7583 VSUBS 0.02fF $ **FLOATING
C8337 S.n7584 VSUBS 0.01fF $ **FLOATING
C8338 S.n7585 VSUBS 0.02fF $ **FLOATING
C8339 S.n7586 VSUBS 0.08fF $ **FLOATING
C8340 S.n7587 VSUBS 0.06fF $ **FLOATING
C8341 S.n7588 VSUBS 0.03fF $ **FLOATING
C8342 S.n7589 VSUBS 0.04fF $ **FLOATING
C8343 S.n7590 VSUBS 1.00fF $ **FLOATING
C8344 S.n7591 VSUBS 0.36fF $ **FLOATING
C8345 S.n7592 VSUBS 1.87fF $ **FLOATING
C8346 S.n7593 VSUBS 1.99fF $ **FLOATING
C8347 S.t399 VSUBS 0.02fF
C8348 S.n7594 VSUBS 0.24fF $ **FLOATING
C8349 S.n7595 VSUBS 0.91fF $ **FLOATING
C8350 S.n7596 VSUBS 0.05fF $ **FLOATING
C8351 S.t1337 VSUBS 0.02fF
C8352 S.n7597 VSUBS 0.12fF $ **FLOATING
C8353 S.n7598 VSUBS 0.14fF $ **FLOATING
C8354 S.n7600 VSUBS 1.89fF $ **FLOATING
C8355 S.n7601 VSUBS 0.07fF $ **FLOATING
C8356 S.n7602 VSUBS 0.04fF $ **FLOATING
C8357 S.n7603 VSUBS 0.05fF $ **FLOATING
C8358 S.n7604 VSUBS 0.87fF $ **FLOATING
C8359 S.n7605 VSUBS 0.01fF $ **FLOATING
C8360 S.n7606 VSUBS 0.01fF $ **FLOATING
C8361 S.n7607 VSUBS 0.01fF $ **FLOATING
C8362 S.n7608 VSUBS 0.07fF $ **FLOATING
C8363 S.n7609 VSUBS 0.68fF $ **FLOATING
C8364 S.n7610 VSUBS 0.72fF $ **FLOATING
C8365 S.t892 VSUBS 0.02fF
C8366 S.n7611 VSUBS 0.24fF $ **FLOATING
C8367 S.n7612 VSUBS 0.36fF $ **FLOATING
C8368 S.n7613 VSUBS 0.61fF $ **FLOATING
C8369 S.n7614 VSUBS 0.12fF $ **FLOATING
C8370 S.t28 VSUBS 0.02fF
C8371 S.n7615 VSUBS 0.14fF $ **FLOATING
C8372 S.n7617 VSUBS 0.70fF $ **FLOATING
C8373 S.n7618 VSUBS 0.23fF $ **FLOATING
C8374 S.n7619 VSUBS 0.23fF $ **FLOATING
C8375 S.n7620 VSUBS 0.70fF $ **FLOATING
C8376 S.n7621 VSUBS 1.16fF $ **FLOATING
C8377 S.n7622 VSUBS 0.22fF $ **FLOATING
C8378 S.n7623 VSUBS 0.25fF $ **FLOATING
C8379 S.n7624 VSUBS 0.09fF $ **FLOATING
C8380 S.n7625 VSUBS 2.31fF $ **FLOATING
C8381 S.t1190 VSUBS 0.02fF
C8382 S.n7626 VSUBS 0.24fF $ **FLOATING
C8383 S.n7627 VSUBS 0.91fF $ **FLOATING
C8384 S.n7628 VSUBS 0.05fF $ **FLOATING
C8385 S.t945 VSUBS 0.02fF
C8386 S.n7629 VSUBS 0.12fF $ **FLOATING
C8387 S.n7630 VSUBS 0.14fF $ **FLOATING
C8388 S.n7632 VSUBS 1.88fF $ **FLOATING
C8389 S.n7633 VSUBS 0.46fF $ **FLOATING
C8390 S.n7634 VSUBS 0.22fF $ **FLOATING
C8391 S.n7635 VSUBS 0.38fF $ **FLOATING
C8392 S.n7636 VSUBS 0.16fF $ **FLOATING
C8393 S.n7637 VSUBS 0.28fF $ **FLOATING
C8394 S.n7638 VSUBS 0.21fF $ **FLOATING
C8395 S.n7639 VSUBS 0.30fF $ **FLOATING
C8396 S.n7640 VSUBS 0.42fF $ **FLOATING
C8397 S.n7641 VSUBS 0.21fF $ **FLOATING
C8398 S.t1672 VSUBS 0.02fF
C8399 S.n7642 VSUBS 0.24fF $ **FLOATING
C8400 S.n7643 VSUBS 0.36fF $ **FLOATING
C8401 S.n7644 VSUBS 0.61fF $ **FLOATING
C8402 S.n7645 VSUBS 0.12fF $ **FLOATING
C8403 S.t861 VSUBS 0.02fF
C8404 S.n7646 VSUBS 0.14fF $ **FLOATING
C8405 S.n7648 VSUBS 0.04fF $ **FLOATING
C8406 S.n7649 VSUBS 0.03fF $ **FLOATING
C8407 S.n7650 VSUBS 0.03fF $ **FLOATING
C8408 S.n7651 VSUBS 0.10fF $ **FLOATING
C8409 S.n7652 VSUBS 0.36fF $ **FLOATING
C8410 S.n7653 VSUBS 0.38fF $ **FLOATING
C8411 S.n7654 VSUBS 0.11fF $ **FLOATING
C8412 S.n7655 VSUBS 0.12fF $ **FLOATING
C8413 S.n7656 VSUBS 0.07fF $ **FLOATING
C8414 S.n7657 VSUBS 0.12fF $ **FLOATING
C8415 S.n7658 VSUBS 0.18fF $ **FLOATING
C8416 S.n7659 VSUBS 3.99fF $ **FLOATING
C8417 S.t1971 VSUBS 0.02fF
C8418 S.n7660 VSUBS 0.24fF $ **FLOATING
C8419 S.n7661 VSUBS 0.91fF $ **FLOATING
C8420 S.n7662 VSUBS 0.05fF $ **FLOATING
C8421 S.t1727 VSUBS 0.02fF
C8422 S.n7663 VSUBS 0.12fF $ **FLOATING
C8423 S.n7664 VSUBS 0.14fF $ **FLOATING
C8424 S.n7666 VSUBS 0.25fF $ **FLOATING
C8425 S.n7667 VSUBS 0.09fF $ **FLOATING
C8426 S.n7668 VSUBS 0.21fF $ **FLOATING
C8427 S.n7669 VSUBS 1.28fF $ **FLOATING
C8428 S.n7670 VSUBS 0.53fF $ **FLOATING
C8429 S.n7671 VSUBS 1.88fF $ **FLOATING
C8430 S.n7672 VSUBS 0.12fF $ **FLOATING
C8431 S.t1645 VSUBS 0.02fF
C8432 S.n7673 VSUBS 0.14fF $ **FLOATING
C8433 S.t2461 VSUBS 0.02fF
C8434 S.n7675 VSUBS 0.24fF $ **FLOATING
C8435 S.n7676 VSUBS 0.36fF $ **FLOATING
C8436 S.n7677 VSUBS 0.61fF $ **FLOATING
C8437 S.n7678 VSUBS 1.58fF $ **FLOATING
C8438 S.n7679 VSUBS 2.45fF $ **FLOATING
C8439 S.t236 VSUBS 0.02fF
C8440 S.n7680 VSUBS 0.24fF $ **FLOATING
C8441 S.n7681 VSUBS 0.91fF $ **FLOATING
C8442 S.n7682 VSUBS 0.05fF $ **FLOATING
C8443 S.t2516 VSUBS 0.02fF
C8444 S.n7683 VSUBS 0.12fF $ **FLOATING
C8445 S.n7684 VSUBS 0.14fF $ **FLOATING
C8446 S.n7686 VSUBS 1.89fF $ **FLOATING
C8447 S.n7687 VSUBS 0.06fF $ **FLOATING
C8448 S.n7688 VSUBS 0.03fF $ **FLOATING
C8449 S.n7689 VSUBS 0.04fF $ **FLOATING
C8450 S.n7690 VSUBS 0.99fF $ **FLOATING
C8451 S.n7691 VSUBS 0.02fF $ **FLOATING
C8452 S.n7692 VSUBS 0.01fF $ **FLOATING
C8453 S.n7693 VSUBS 0.02fF $ **FLOATING
C8454 S.n7694 VSUBS 0.08fF $ **FLOATING
C8455 S.n7695 VSUBS 0.36fF $ **FLOATING
C8456 S.n7696 VSUBS 1.85fF $ **FLOATING
C8457 S.t850 VSUBS 0.02fF
C8458 S.n7697 VSUBS 0.24fF $ **FLOATING
C8459 S.n7698 VSUBS 0.36fF $ **FLOATING
C8460 S.n7699 VSUBS 0.61fF $ **FLOATING
C8461 S.n7700 VSUBS 0.12fF $ **FLOATING
C8462 S.t2553 VSUBS 0.02fF
C8463 S.n7701 VSUBS 0.14fF $ **FLOATING
C8464 S.n7703 VSUBS 0.70fF $ **FLOATING
C8465 S.n7704 VSUBS 0.23fF $ **FLOATING
C8466 S.n7705 VSUBS 0.23fF $ **FLOATING
C8467 S.n7706 VSUBS 0.70fF $ **FLOATING
C8468 S.n7707 VSUBS 1.16fF $ **FLOATING
C8469 S.n7708 VSUBS 0.22fF $ **FLOATING
C8470 S.n7709 VSUBS 0.25fF $ **FLOATING
C8471 S.n7710 VSUBS 0.09fF $ **FLOATING
C8472 S.n7711 VSUBS 1.88fF $ **FLOATING
C8473 S.t1153 VSUBS 0.02fF
C8474 S.n7712 VSUBS 0.24fF $ **FLOATING
C8475 S.n7713 VSUBS 0.91fF $ **FLOATING
C8476 S.n7714 VSUBS 0.05fF $ **FLOATING
C8477 S.t906 VSUBS 0.02fF
C8478 S.n7715 VSUBS 0.12fF $ **FLOATING
C8479 S.n7716 VSUBS 0.14fF $ **FLOATING
C8480 S.n7718 VSUBS 20.78fF $ **FLOATING
C8481 S.n7719 VSUBS 1.72fF $ **FLOATING
C8482 S.n7720 VSUBS 3.05fF $ **FLOATING
C8483 S.t1322 VSUBS 0.02fF
C8484 S.n7721 VSUBS 0.24fF $ **FLOATING
C8485 S.n7722 VSUBS 0.36fF $ **FLOATING
C8486 S.n7723 VSUBS 0.61fF $ **FLOATING
C8487 S.n7724 VSUBS 0.12fF $ **FLOATING
C8488 S.t508 VSUBS 0.02fF
C8489 S.n7725 VSUBS 0.14fF $ **FLOATING
C8490 S.n7727 VSUBS 0.31fF $ **FLOATING
C8491 S.n7728 VSUBS 0.23fF $ **FLOATING
C8492 S.n7729 VSUBS 0.66fF $ **FLOATING
C8493 S.n7730 VSUBS 0.95fF $ **FLOATING
C8494 S.n7731 VSUBS 0.23fF $ **FLOATING
C8495 S.n7732 VSUBS 0.21fF $ **FLOATING
C8496 S.n7733 VSUBS 0.20fF $ **FLOATING
C8497 S.n7734 VSUBS 0.06fF $ **FLOATING
C8498 S.n7735 VSUBS 0.09fF $ **FLOATING
C8499 S.n7736 VSUBS 0.10fF $ **FLOATING
C8500 S.n7737 VSUBS 1.99fF $ **FLOATING
C8501 S.t1374 VSUBS 0.02fF
C8502 S.n7738 VSUBS 0.12fF $ **FLOATING
C8503 S.n7739 VSUBS 0.14fF $ **FLOATING
C8504 S.t1592 VSUBS 0.02fF
C8505 S.n7741 VSUBS 0.24fF $ **FLOATING
C8506 S.n7742 VSUBS 0.91fF $ **FLOATING
C8507 S.n7743 VSUBS 0.05fF $ **FLOATING
C8508 S.n7744 VSUBS 1.88fF $ **FLOATING
C8509 S.n7745 VSUBS 0.12fF $ **FLOATING
C8510 S.t238 VSUBS 0.02fF
C8511 S.n7746 VSUBS 0.14fF $ **FLOATING
C8512 S.t1908 VSUBS 0.02fF
C8513 S.n7748 VSUBS 1.22fF $ **FLOATING
C8514 S.n7749 VSUBS 0.61fF $ **FLOATING
C8515 S.n7750 VSUBS 0.35fF $ **FLOATING
C8516 S.n7751 VSUBS 0.63fF $ **FLOATING
C8517 S.n7752 VSUBS 1.15fF $ **FLOATING
C8518 S.n7753 VSUBS 3.00fF $ **FLOATING
C8519 S.n7754 VSUBS 0.59fF $ **FLOATING
C8520 S.n7755 VSUBS 0.01fF $ **FLOATING
C8521 S.n7756 VSUBS 0.97fF $ **FLOATING
C8522 S.t63 VSUBS 21.42fF
C8523 S.n7757 VSUBS 20.29fF $ **FLOATING
C8524 S.n7759 VSUBS 0.38fF $ **FLOATING
C8525 S.n7760 VSUBS 0.23fF $ **FLOATING
C8526 S.n7761 VSUBS 2.90fF $ **FLOATING
C8527 S.n7762 VSUBS 2.46fF $ **FLOATING
C8528 S.n7763 VSUBS 1.96fF $ **FLOATING
C8529 S.n7764 VSUBS 3.94fF $ **FLOATING
C8530 S.n7765 VSUBS 0.25fF $ **FLOATING
C8531 S.n7766 VSUBS 0.01fF $ **FLOATING
C8532 S.t1097 VSUBS 0.02fF
C8533 S.n7767 VSUBS 0.26fF $ **FLOATING
C8534 S.t2190 VSUBS 0.02fF
C8535 S.n7768 VSUBS 0.95fF $ **FLOATING
C8536 S.n7769 VSUBS 0.71fF $ **FLOATING
C8537 S.n7770 VSUBS 0.78fF $ **FLOATING
C8538 S.n7771 VSUBS 1.93fF $ **FLOATING
C8539 S.n7772 VSUBS 1.88fF $ **FLOATING
C8540 S.n7773 VSUBS 0.12fF $ **FLOATING
C8541 S.t1878 VSUBS 0.02fF
C8542 S.n7774 VSUBS 0.14fF $ **FLOATING
C8543 S.t163 VSUBS 0.02fF
C8544 S.n7776 VSUBS 0.24fF $ **FLOATING
C8545 S.n7777 VSUBS 0.36fF $ **FLOATING
C8546 S.n7778 VSUBS 0.61fF $ **FLOATING
C8547 S.n7779 VSUBS 1.52fF $ **FLOATING
C8548 S.n7780 VSUBS 2.99fF $ **FLOATING
C8549 S.t456 VSUBS 0.02fF
C8550 S.n7781 VSUBS 0.24fF $ **FLOATING
C8551 S.n7782 VSUBS 0.91fF $ **FLOATING
C8552 S.n7783 VSUBS 0.05fF $ **FLOATING
C8553 S.t222 VSUBS 0.02fF
C8554 S.n7784 VSUBS 0.12fF $ **FLOATING
C8555 S.n7785 VSUBS 0.14fF $ **FLOATING
C8556 S.n7787 VSUBS 1.89fF $ **FLOATING
C8557 S.n7788 VSUBS 1.88fF $ **FLOATING
C8558 S.t951 VSUBS 0.02fF
C8559 S.n7789 VSUBS 0.24fF $ **FLOATING
C8560 S.n7790 VSUBS 0.36fF $ **FLOATING
C8561 S.n7791 VSUBS 0.61fF $ **FLOATING
C8562 S.n7792 VSUBS 0.12fF $ **FLOATING
C8563 S.t274 VSUBS 0.02fF
C8564 S.n7793 VSUBS 0.14fF $ **FLOATING
C8565 S.n7795 VSUBS 1.16fF $ **FLOATING
C8566 S.n7796 VSUBS 0.22fF $ **FLOATING
C8567 S.n7797 VSUBS 0.25fF $ **FLOATING
C8568 S.n7798 VSUBS 0.09fF $ **FLOATING
C8569 S.n7799 VSUBS 1.88fF $ **FLOATING
C8570 S.t1244 VSUBS 0.02fF
C8571 S.n7800 VSUBS 0.24fF $ **FLOATING
C8572 S.n7801 VSUBS 0.91fF $ **FLOATING
C8573 S.n7802 VSUBS 0.05fF $ **FLOATING
C8574 S.t1009 VSUBS 0.02fF
C8575 S.n7803 VSUBS 0.12fF $ **FLOATING
C8576 S.n7804 VSUBS 0.14fF $ **FLOATING
C8577 S.n7806 VSUBS 0.78fF $ **FLOATING
C8578 S.n7807 VSUBS 1.94fF $ **FLOATING
C8579 S.n7808 VSUBS 1.88fF $ **FLOATING
C8580 S.n7809 VSUBS 0.12fF $ **FLOATING
C8581 S.t1052 VSUBS 0.02fF
C8582 S.n7810 VSUBS 0.14fF $ **FLOATING
C8583 S.t1865 VSUBS 0.02fF
C8584 S.n7812 VSUBS 0.24fF $ **FLOATING
C8585 S.n7813 VSUBS 0.36fF $ **FLOATING
C8586 S.n7814 VSUBS 0.61fF $ **FLOATING
C8587 S.n7815 VSUBS 1.84fF $ **FLOATING
C8588 S.n7816 VSUBS 2.99fF $ **FLOATING
C8589 S.t2152 VSUBS 0.02fF
C8590 S.n7817 VSUBS 0.24fF $ **FLOATING
C8591 S.n7818 VSUBS 0.91fF $ **FLOATING
C8592 S.n7819 VSUBS 0.05fF $ **FLOATING
C8593 S.t1923 VSUBS 0.02fF
C8594 S.n7820 VSUBS 0.12fF $ **FLOATING
C8595 S.n7821 VSUBS 0.14fF $ **FLOATING
C8596 S.n7823 VSUBS 1.89fF $ **FLOATING
C8597 S.n7824 VSUBS 1.75fF $ **FLOATING
C8598 S.t1470 VSUBS 0.02fF
C8599 S.n7825 VSUBS 0.24fF $ **FLOATING
C8600 S.n7826 VSUBS 0.36fF $ **FLOATING
C8601 S.n7827 VSUBS 0.61fF $ **FLOATING
C8602 S.n7828 VSUBS 0.12fF $ **FLOATING
C8603 S.t651 VSUBS 0.02fF
C8604 S.n7829 VSUBS 0.14fF $ **FLOATING
C8605 S.n7831 VSUBS 1.16fF $ **FLOATING
C8606 S.n7832 VSUBS 0.22fF $ **FLOATING
C8607 S.n7833 VSUBS 0.25fF $ **FLOATING
C8608 S.n7834 VSUBS 0.09fF $ **FLOATING
C8609 S.n7835 VSUBS 2.44fF $ **FLOATING
C8610 S.t1761 VSUBS 0.02fF
C8611 S.n7836 VSUBS 0.24fF $ **FLOATING
C8612 S.n7837 VSUBS 0.91fF $ **FLOATING
C8613 S.n7838 VSUBS 0.05fF $ **FLOATING
C8614 S.t1518 VSUBS 0.02fF
C8615 S.n7839 VSUBS 0.12fF $ **FLOATING
C8616 S.n7840 VSUBS 0.14fF $ **FLOATING
C8617 S.n7842 VSUBS 1.88fF $ **FLOATING
C8618 S.n7843 VSUBS 0.48fF $ **FLOATING
C8619 S.n7844 VSUBS 0.09fF $ **FLOATING
C8620 S.n7845 VSUBS 0.33fF $ **FLOATING
C8621 S.n7846 VSUBS 0.30fF $ **FLOATING
C8622 S.n7847 VSUBS 0.77fF $ **FLOATING
C8623 S.n7848 VSUBS 0.59fF $ **FLOATING
C8624 S.t2257 VSUBS 0.02fF
C8625 S.n7849 VSUBS 0.24fF $ **FLOATING
C8626 S.n7850 VSUBS 0.36fF $ **FLOATING
C8627 S.n7851 VSUBS 0.61fF $ **FLOATING
C8628 S.n7852 VSUBS 0.12fF $ **FLOATING
C8629 S.t1439 VSUBS 0.02fF
C8630 S.n7853 VSUBS 0.14fF $ **FLOATING
C8631 S.n7855 VSUBS 2.61fF $ **FLOATING
C8632 S.n7856 VSUBS 2.15fF $ **FLOATING
C8633 S.t2542 VSUBS 0.02fF
C8634 S.n7857 VSUBS 0.24fF $ **FLOATING
C8635 S.n7858 VSUBS 0.91fF $ **FLOATING
C8636 S.n7859 VSUBS 0.05fF $ **FLOATING
C8637 S.t2308 VSUBS 0.02fF
C8638 S.n7860 VSUBS 0.12fF $ **FLOATING
C8639 S.n7861 VSUBS 0.14fF $ **FLOATING
C8640 S.n7863 VSUBS 0.78fF $ **FLOATING
C8641 S.n7864 VSUBS 2.30fF $ **FLOATING
C8642 S.n7865 VSUBS 1.88fF $ **FLOATING
C8643 S.n7866 VSUBS 0.12fF $ **FLOATING
C8644 S.t2231 VSUBS 0.02fF
C8645 S.n7867 VSUBS 0.14fF $ **FLOATING
C8646 S.t527 VSUBS 0.02fF
C8647 S.n7869 VSUBS 0.24fF $ **FLOATING
C8648 S.n7870 VSUBS 0.36fF $ **FLOATING
C8649 S.n7871 VSUBS 0.61fF $ **FLOATING
C8650 S.n7872 VSUBS 1.39fF $ **FLOATING
C8651 S.n7873 VSUBS 0.71fF $ **FLOATING
C8652 S.n7874 VSUBS 1.14fF $ **FLOATING
C8653 S.n7875 VSUBS 0.35fF $ **FLOATING
C8654 S.n7876 VSUBS 2.02fF $ **FLOATING
C8655 S.t806 VSUBS 0.02fF
C8656 S.n7877 VSUBS 0.24fF $ **FLOATING
C8657 S.n7878 VSUBS 0.91fF $ **FLOATING
C8658 S.n7879 VSUBS 0.05fF $ **FLOATING
C8659 S.t576 VSUBS 0.02fF
C8660 S.n7880 VSUBS 0.12fF $ **FLOATING
C8661 S.n7881 VSUBS 0.14fF $ **FLOATING
C8662 S.n7883 VSUBS 1.89fF $ **FLOATING
C8663 S.n7884 VSUBS 1.88fF $ **FLOATING
C8664 S.t1313 VSUBS 0.02fF
C8665 S.n7885 VSUBS 0.24fF $ **FLOATING
C8666 S.n7886 VSUBS 0.36fF $ **FLOATING
C8667 S.n7887 VSUBS 0.61fF $ **FLOATING
C8668 S.n7888 VSUBS 0.12fF $ **FLOATING
C8669 S.t619 VSUBS 0.02fF
C8670 S.n7889 VSUBS 0.14fF $ **FLOATING
C8671 S.n7891 VSUBS 1.16fF $ **FLOATING
C8672 S.n7892 VSUBS 0.22fF $ **FLOATING
C8673 S.n7893 VSUBS 0.25fF $ **FLOATING
C8674 S.n7894 VSUBS 0.09fF $ **FLOATING
C8675 S.n7895 VSUBS 1.88fF $ **FLOATING
C8676 S.t1587 VSUBS 0.02fF
C8677 S.n7896 VSUBS 0.24fF $ **FLOATING
C8678 S.n7897 VSUBS 0.91fF $ **FLOATING
C8679 S.n7898 VSUBS 0.05fF $ **FLOATING
C8680 S.t1367 VSUBS 0.02fF
C8681 S.n7899 VSUBS 0.12fF $ **FLOATING
C8682 S.n7900 VSUBS 0.14fF $ **FLOATING
C8683 S.n7902 VSUBS 20.78fF $ **FLOATING
C8684 S.n7903 VSUBS 1.88fF $ **FLOATING
C8685 S.n7904 VSUBS 2.67fF $ **FLOATING
C8686 S.t64 VSUBS 0.02fF
C8687 S.n7905 VSUBS 0.24fF $ **FLOATING
C8688 S.n7906 VSUBS 0.36fF $ **FLOATING
C8689 S.n7907 VSUBS 0.61fF $ **FLOATING
C8690 S.n7908 VSUBS 0.12fF $ **FLOATING
C8691 S.t1802 VSUBS 0.02fF
C8692 S.n7909 VSUBS 0.14fF $ **FLOATING
C8693 S.n7911 VSUBS 2.80fF $ **FLOATING
C8694 S.n7912 VSUBS 2.30fF $ **FLOATING
C8695 S.t140 VSUBS 0.02fF
C8696 S.n7913 VSUBS 0.12fF $ **FLOATING
C8697 S.n7914 VSUBS 0.14fF $ **FLOATING
C8698 S.t391 VSUBS 0.02fF
C8699 S.n7916 VSUBS 0.24fF $ **FLOATING
C8700 S.n7917 VSUBS 0.91fF $ **FLOATING
C8701 S.n7918 VSUBS 0.05fF $ **FLOATING
C8702 S.n7919 VSUBS 2.80fF $ **FLOATING
C8703 S.n7920 VSUBS 1.88fF $ **FLOATING
C8704 S.n7921 VSUBS 0.12fF $ **FLOATING
C8705 S.t12 VSUBS 0.02fF
C8706 S.n7922 VSUBS 0.14fF $ **FLOATING
C8707 S.t881 VSUBS 0.02fF
C8708 S.n7924 VSUBS 0.24fF $ **FLOATING
C8709 S.n7925 VSUBS 0.36fF $ **FLOATING
C8710 S.n7926 VSUBS 0.61fF $ **FLOATING
C8711 S.n7927 VSUBS 2.67fF $ **FLOATING
C8712 S.n7928 VSUBS 2.30fF $ **FLOATING
C8713 S.t937 VSUBS 0.02fF
C8714 S.n7929 VSUBS 0.12fF $ **FLOATING
C8715 S.n7930 VSUBS 0.14fF $ **FLOATING
C8716 S.t1183 VSUBS 0.02fF
C8717 S.n7932 VSUBS 0.24fF $ **FLOATING
C8718 S.n7933 VSUBS 0.91fF $ **FLOATING
C8719 S.n7934 VSUBS 0.05fF $ **FLOATING
C8720 S.n7935 VSUBS 1.88fF $ **FLOATING
C8721 S.n7936 VSUBS 2.67fF $ **FLOATING
C8722 S.t1662 VSUBS 0.02fF
C8723 S.n7937 VSUBS 0.24fF $ **FLOATING
C8724 S.n7938 VSUBS 0.36fF $ **FLOATING
C8725 S.n7939 VSUBS 0.61fF $ **FLOATING
C8726 S.n7940 VSUBS 0.12fF $ **FLOATING
C8727 S.t986 VSUBS 0.02fF
C8728 S.n7941 VSUBS 0.14fF $ **FLOATING
C8729 S.n7943 VSUBS 2.80fF $ **FLOATING
C8730 S.n7944 VSUBS 2.30fF $ **FLOATING
C8731 S.t1718 VSUBS 0.02fF
C8732 S.n7945 VSUBS 0.12fF $ **FLOATING
C8733 S.n7946 VSUBS 0.14fF $ **FLOATING
C8734 S.t1966 VSUBS 0.02fF
C8735 S.n7948 VSUBS 0.24fF $ **FLOATING
C8736 S.n7949 VSUBS 0.91fF $ **FLOATING
C8737 S.n7950 VSUBS 0.05fF $ **FLOATING
C8738 S.n7951 VSUBS 1.88fF $ **FLOATING
C8739 S.n7952 VSUBS 2.67fF $ **FLOATING
C8740 S.t594 VSUBS 0.02fF
C8741 S.n7953 VSUBS 0.24fF $ **FLOATING
C8742 S.n7954 VSUBS 0.36fF $ **FLOATING
C8743 S.n7955 VSUBS 0.61fF $ **FLOATING
C8744 S.n7956 VSUBS 0.12fF $ **FLOATING
C8745 S.t790 VSUBS 0.02fF
C8746 S.n7957 VSUBS 0.14fF $ **FLOATING
C8747 S.n7959 VSUBS 2.80fF $ **FLOATING
C8748 S.n7960 VSUBS 2.30fF $ **FLOATING
C8749 S.t1658 VSUBS 0.02fF
C8750 S.n7961 VSUBS 0.12fF $ **FLOATING
C8751 S.n7962 VSUBS 0.14fF $ **FLOATING
C8752 S.t1435 VSUBS 0.02fF
C8753 S.n7964 VSUBS 0.24fF $ **FLOATING
C8754 S.n7965 VSUBS 0.91fF $ **FLOATING
C8755 S.n7966 VSUBS 0.05fF $ **FLOATING
C8756 S.n7967 VSUBS 1.88fF $ **FLOATING
C8757 S.n7968 VSUBS 2.67fF $ **FLOATING
C8758 S.t1387 VSUBS 0.02fF
C8759 S.n7969 VSUBS 0.24fF $ **FLOATING
C8760 S.n7970 VSUBS 0.36fF $ **FLOATING
C8761 S.n7971 VSUBS 0.61fF $ **FLOATING
C8762 S.n7972 VSUBS 0.12fF $ **FLOATING
C8763 S.t1571 VSUBS 0.02fF
C8764 S.n7973 VSUBS 0.14fF $ **FLOATING
C8765 S.n7975 VSUBS 2.80fF $ **FLOATING
C8766 S.n7976 VSUBS 2.30fF $ **FLOATING
C8767 S.t2446 VSUBS 0.02fF
C8768 S.n7977 VSUBS 0.12fF $ **FLOATING
C8769 S.n7978 VSUBS 0.14fF $ **FLOATING
C8770 S.t2227 VSUBS 0.02fF
C8771 S.n7980 VSUBS 0.24fF $ **FLOATING
C8772 S.n7981 VSUBS 0.91fF $ **FLOATING
C8773 S.n7982 VSUBS 0.05fF $ **FLOATING
C8774 S.n7983 VSUBS 1.88fF $ **FLOATING
C8775 S.n7984 VSUBS 2.67fF $ **FLOATING
C8776 S.t2172 VSUBS 0.02fF
C8777 S.n7985 VSUBS 0.24fF $ **FLOATING
C8778 S.n7986 VSUBS 0.36fF $ **FLOATING
C8779 S.n7987 VSUBS 0.61fF $ **FLOATING
C8780 S.n7988 VSUBS 0.12fF $ **FLOATING
C8781 S.t2364 VSUBS 0.02fF
C8782 S.n7989 VSUBS 0.14fF $ **FLOATING
C8783 S.n7991 VSUBS 2.80fF $ **FLOATING
C8784 S.n7992 VSUBS 2.30fF $ **FLOATING
C8785 S.t703 VSUBS 0.02fF
C8786 S.n7993 VSUBS 0.12fF $ **FLOATING
C8787 S.n7994 VSUBS 0.14fF $ **FLOATING
C8788 S.t494 VSUBS 0.02fF
C8789 S.n7996 VSUBS 0.24fF $ **FLOATING
C8790 S.n7997 VSUBS 0.91fF $ **FLOATING
C8791 S.n7998 VSUBS 0.05fF $ **FLOATING
C8792 S.n7999 VSUBS 1.88fF $ **FLOATING
C8793 S.n8000 VSUBS 2.68fF $ **FLOATING
C8794 S.t437 VSUBS 0.02fF
C8795 S.n8001 VSUBS 0.24fF $ **FLOATING
C8796 S.n8002 VSUBS 0.36fF $ **FLOATING
C8797 S.n8003 VSUBS 0.61fF $ **FLOATING
C8798 S.n8004 VSUBS 0.12fF $ **FLOATING
C8799 S.t632 VSUBS 0.02fF
C8800 S.n8005 VSUBS 0.14fF $ **FLOATING
C8801 S.n8007 VSUBS 5.17fF $ **FLOATING
C8802 S.t1499 VSUBS 0.02fF
C8803 S.n8008 VSUBS 0.12fF $ **FLOATING
C8804 S.n8009 VSUBS 0.14fF $ **FLOATING
C8805 S.t1283 VSUBS 0.02fF
C8806 S.n8011 VSUBS 0.24fF $ **FLOATING
C8807 S.n8012 VSUBS 0.91fF $ **FLOATING
C8808 S.n8013 VSUBS 0.05fF $ **FLOATING
C8809 S.n8014 VSUBS 2.73fF $ **FLOATING
C8810 S.n8015 VSUBS 1.59fF $ **FLOATING
C8811 S.n8016 VSUBS 0.12fF $ **FLOATING
C8812 S.t2427 VSUBS 0.02fF
C8813 S.n8017 VSUBS 0.14fF $ **FLOATING
C8814 S.t1055 VSUBS 0.02fF
C8815 S.n8019 VSUBS 0.24fF $ **FLOATING
C8816 S.n8020 VSUBS 0.36fF $ **FLOATING
C8817 S.n8021 VSUBS 0.61fF $ **FLOATING
C8818 S.n8022 VSUBS 0.07fF $ **FLOATING
C8819 S.n8023 VSUBS 0.01fF $ **FLOATING
C8820 S.n8024 VSUBS 0.24fF $ **FLOATING
C8821 S.n8025 VSUBS 1.16fF $ **FLOATING
C8822 S.n8026 VSUBS 1.35fF $ **FLOATING
C8823 S.n8027 VSUBS 2.30fF $ **FLOATING
C8824 S.t2285 VSUBS 0.02fF
C8825 S.n8028 VSUBS 0.12fF $ **FLOATING
C8826 S.n8029 VSUBS 0.14fF $ **FLOATING
C8827 S.t2437 VSUBS 0.02fF
C8828 S.n8031 VSUBS 0.24fF $ **FLOATING
C8829 S.n8032 VSUBS 0.91fF $ **FLOATING
C8830 S.n8033 VSUBS 0.05fF $ **FLOATING
C8831 S.t11 VSUBS 48.27fF
C8832 S.t2271 VSUBS 0.02fF
C8833 S.n8034 VSUBS 0.12fF $ **FLOATING
C8834 S.n8035 VSUBS 0.14fF $ **FLOATING
C8835 S.t1338 VSUBS 0.02fF
C8836 S.n8037 VSUBS 0.24fF $ **FLOATING
C8837 S.n8038 VSUBS 0.91fF $ **FLOATING
C8838 S.n8039 VSUBS 0.05fF $ **FLOATING
C8839 S.t1053 VSUBS 0.02fF
C8840 S.n8040 VSUBS 0.24fF $ **FLOATING
C8841 S.n8041 VSUBS 0.36fF $ **FLOATING
C8842 S.n8042 VSUBS 0.61fF $ **FLOATING
C8843 S.n8043 VSUBS 0.32fF $ **FLOATING
C8844 S.n8044 VSUBS 1.09fF $ **FLOATING
C8845 S.n8045 VSUBS 0.15fF $ **FLOATING
C8846 S.n8046 VSUBS 2.10fF $ **FLOATING
C8847 S.n8047 VSUBS 2.94fF $ **FLOATING
C8848 S.n8048 VSUBS 1.88fF $ **FLOATING
C8849 S.n8049 VSUBS 0.12fF $ **FLOATING
C8850 S.t2174 VSUBS 0.02fF
C8851 S.n8050 VSUBS 0.14fF $ **FLOATING
C8852 S.t470 VSUBS 0.02fF
C8853 S.n8052 VSUBS 0.24fF $ **FLOATING
C8854 S.n8053 VSUBS 0.36fF $ **FLOATING
C8855 S.n8054 VSUBS 0.61fF $ **FLOATING
C8856 S.n8055 VSUBS 0.92fF $ **FLOATING
C8857 S.n8056 VSUBS 0.32fF $ **FLOATING
C8858 S.n8057 VSUBS 0.92fF $ **FLOATING
C8859 S.n8058 VSUBS 1.09fF $ **FLOATING
C8860 S.n8059 VSUBS 0.15fF $ **FLOATING
C8861 S.n8060 VSUBS 4.96fF $ **FLOATING
C8862 S.t519 VSUBS 0.02fF
C8863 S.n8061 VSUBS 0.12fF $ **FLOATING
C8864 S.n8062 VSUBS 0.14fF $ **FLOATING
C8865 S.t739 VSUBS 0.02fF
C8866 S.n8064 VSUBS 0.24fF $ **FLOATING
C8867 S.n8065 VSUBS 0.91fF $ **FLOATING
C8868 S.n8066 VSUBS 0.05fF $ **FLOATING
C8869 S.n8067 VSUBS 1.88fF $ **FLOATING
C8870 S.n8068 VSUBS 2.67fF $ **FLOATING
C8871 S.t1256 VSUBS 0.02fF
C8872 S.n8069 VSUBS 0.24fF $ **FLOATING
C8873 S.n8070 VSUBS 0.36fF $ **FLOATING
C8874 S.n8071 VSUBS 0.61fF $ **FLOATING
C8875 S.n8072 VSUBS 0.12fF $ **FLOATING
C8876 S.t439 VSUBS 0.02fF
C8877 S.n8073 VSUBS 0.14fF $ **FLOATING
C8878 S.n8075 VSUBS 1.88fF $ **FLOATING
C8879 S.n8076 VSUBS 2.67fF $ **FLOATING
C8880 S.t1837 VSUBS 0.02fF
C8881 S.n8077 VSUBS 0.24fF $ **FLOATING
C8882 S.n8078 VSUBS 0.36fF $ **FLOATING
C8883 S.n8079 VSUBS 0.61fF $ **FLOATING
C8884 S.t2123 VSUBS 0.02fF
C8885 S.n8080 VSUBS 0.24fF $ **FLOATING
C8886 S.n8081 VSUBS 0.91fF $ **FLOATING
C8887 S.n8082 VSUBS 0.05fF $ **FLOATING
C8888 S.t1891 VSUBS 0.02fF
C8889 S.n8083 VSUBS 0.12fF $ **FLOATING
C8890 S.n8084 VSUBS 0.14fF $ **FLOATING
C8891 S.n8086 VSUBS 0.12fF $ **FLOATING
C8892 S.t1023 VSUBS 0.02fF
C8893 S.n8087 VSUBS 0.14fF $ **FLOATING
C8894 S.n8089 VSUBS 2.30fF $ **FLOATING
C8895 S.n8090 VSUBS 2.94fF $ **FLOATING
C8896 S.n8091 VSUBS 5.16fF $ **FLOATING
C8897 S.t1306 VSUBS 0.02fF
C8898 S.n8092 VSUBS 0.12fF $ **FLOATING
C8899 S.n8093 VSUBS 0.14fF $ **FLOATING
C8900 S.t1531 VSUBS 0.02fF
C8901 S.n8095 VSUBS 0.24fF $ **FLOATING
C8902 S.n8096 VSUBS 0.91fF $ **FLOATING
C8903 S.n8097 VSUBS 0.05fF $ **FLOATING
C8904 S.n8098 VSUBS 1.88fF $ **FLOATING
C8905 S.n8099 VSUBS 2.67fF $ **FLOATING
C8906 S.t2044 VSUBS 0.02fF
C8907 S.n8100 VSUBS 0.24fF $ **FLOATING
C8908 S.n8101 VSUBS 0.36fF $ **FLOATING
C8909 S.n8102 VSUBS 0.61fF $ **FLOATING
C8910 S.n8103 VSUBS 0.12fF $ **FLOATING
C8911 S.t1232 VSUBS 0.02fF
C8912 S.n8104 VSUBS 0.14fF $ **FLOATING
C8913 S.n8106 VSUBS 5.17fF $ **FLOATING
C8914 S.t2093 VSUBS 0.02fF
C8915 S.n8107 VSUBS 0.12fF $ **FLOATING
C8916 S.n8108 VSUBS 0.14fF $ **FLOATING
C8917 S.t2317 VSUBS 0.02fF
C8918 S.n8110 VSUBS 0.24fF $ **FLOATING
C8919 S.n8111 VSUBS 0.91fF $ **FLOATING
C8920 S.n8112 VSUBS 0.05fF $ **FLOATING
C8921 S.n8113 VSUBS 1.88fF $ **FLOATING
C8922 S.n8114 VSUBS 0.12fF $ **FLOATING
C8923 S.t2013 VSUBS 0.02fF
C8924 S.n8115 VSUBS 0.14fF $ **FLOATING
C8925 S.t312 VSUBS 0.02fF
C8926 S.n8117 VSUBS 0.24fF $ **FLOATING
C8927 S.n8118 VSUBS 0.36fF $ **FLOATING
C8928 S.n8119 VSUBS 0.61fF $ **FLOATING
C8929 S.n8120 VSUBS 2.67fF $ **FLOATING
C8930 S.n8121 VSUBS 5.17fF $ **FLOATING
C8931 S.t365 VSUBS 0.02fF
C8932 S.n8122 VSUBS 0.12fF $ **FLOATING
C8933 S.n8123 VSUBS 0.14fF $ **FLOATING
C8934 S.t583 VSUBS 0.02fF
C8935 S.n8125 VSUBS 0.24fF $ **FLOATING
C8936 S.n8126 VSUBS 0.91fF $ **FLOATING
C8937 S.n8127 VSUBS 0.05fF $ **FLOATING
C8938 S.n8128 VSUBS 1.88fF $ **FLOATING
C8939 S.n8129 VSUBS 2.67fF $ **FLOATING
C8940 S.t2303 VSUBS 0.02fF
C8941 S.n8130 VSUBS 0.24fF $ **FLOATING
C8942 S.n8131 VSUBS 0.36fF $ **FLOATING
C8943 S.n8132 VSUBS 0.61fF $ **FLOATING
C8944 S.n8133 VSUBS 0.12fF $ **FLOATING
C8945 S.t2505 VSUBS 0.02fF
C8946 S.n8134 VSUBS 0.14fF $ **FLOATING
C8947 S.n8136 VSUBS 5.17fF $ **FLOATING
C8948 S.t1272 VSUBS 0.02fF
C8949 S.n8137 VSUBS 0.12fF $ **FLOATING
C8950 S.n8138 VSUBS 0.14fF $ **FLOATING
C8951 S.t625 VSUBS 0.02fF
C8952 S.n8140 VSUBS 0.24fF $ **FLOATING
C8953 S.n8141 VSUBS 0.91fF $ **FLOATING
C8954 S.n8142 VSUBS 0.05fF $ **FLOATING
C8955 S.n8143 VSUBS 1.88fF $ **FLOATING
C8956 S.n8144 VSUBS 2.67fF $ **FLOATING
C8957 S.t573 VSUBS 0.02fF
C8958 S.n8145 VSUBS 0.24fF $ **FLOATING
C8959 S.n8146 VSUBS 0.36fF $ **FLOATING
C8960 S.n8147 VSUBS 0.61fF $ **FLOATING
C8961 S.n8148 VSUBS 0.12fF $ **FLOATING
C8962 S.t763 VSUBS 0.02fF
C8963 S.n8149 VSUBS 0.14fF $ **FLOATING
C8964 S.n8151 VSUBS 5.17fF $ **FLOATING
C8965 S.t1634 VSUBS 0.02fF
C8966 S.n8152 VSUBS 0.12fF $ **FLOATING
C8967 S.n8153 VSUBS 0.14fF $ **FLOATING
C8968 S.t1414 VSUBS 0.02fF
C8969 S.n8155 VSUBS 0.24fF $ **FLOATING
C8970 S.n8156 VSUBS 0.91fF $ **FLOATING
C8971 S.n8157 VSUBS 0.05fF $ **FLOATING
C8972 S.n8158 VSUBS 1.88fF $ **FLOATING
C8973 S.n8159 VSUBS 2.67fF $ **FLOATING
C8974 S.t1362 VSUBS 0.02fF
C8975 S.n8160 VSUBS 0.24fF $ **FLOATING
C8976 S.n8161 VSUBS 0.36fF $ **FLOATING
C8977 S.n8162 VSUBS 0.61fF $ **FLOATING
C8978 S.n8163 VSUBS 0.12fF $ **FLOATING
C8979 S.t1551 VSUBS 0.02fF
C8980 S.n8164 VSUBS 0.14fF $ **FLOATING
C8981 S.n8166 VSUBS 5.17fF $ **FLOATING
C8982 S.t2419 VSUBS 0.02fF
C8983 S.n8167 VSUBS 0.12fF $ **FLOATING
C8984 S.n8168 VSUBS 0.14fF $ **FLOATING
C8985 S.t2204 VSUBS 0.02fF
C8986 S.n8170 VSUBS 0.24fF $ **FLOATING
C8987 S.n8171 VSUBS 0.91fF $ **FLOATING
C8988 S.n8172 VSUBS 0.05fF $ **FLOATING
C8989 S.n8173 VSUBS 1.88fF $ **FLOATING
C8990 S.n8174 VSUBS 2.67fF $ **FLOATING
C8991 S.t2148 VSUBS 0.02fF
C8992 S.n8175 VSUBS 0.24fF $ **FLOATING
C8993 S.n8176 VSUBS 0.36fF $ **FLOATING
C8994 S.n8177 VSUBS 0.61fF $ **FLOATING
C8995 S.n8178 VSUBS 0.12fF $ **FLOATING
C8996 S.t2341 VSUBS 0.02fF
C8997 S.n8179 VSUBS 0.14fF $ **FLOATING
C8998 S.n8181 VSUBS 4.89fF $ **FLOATING
C8999 S.t683 VSUBS 0.02fF
C9000 S.n8182 VSUBS 0.12fF $ **FLOATING
C9001 S.n8183 VSUBS 0.14fF $ **FLOATING
C9002 S.t471 VSUBS 0.02fF
C9003 S.n8185 VSUBS 0.24fF $ **FLOATING
C9004 S.n8186 VSUBS 0.91fF $ **FLOATING
C9005 S.n8187 VSUBS 0.05fF $ **FLOATING
C9006 S.n8188 VSUBS 1.88fF $ **FLOATING
C9007 S.n8189 VSUBS 2.67fF $ **FLOATING
C9008 S.t417 VSUBS 0.02fF
C9009 S.n8190 VSUBS 0.24fF $ **FLOATING
C9010 S.n8191 VSUBS 0.36fF $ **FLOATING
C9011 S.n8192 VSUBS 0.61fF $ **FLOATING
C9012 S.n8193 VSUBS 0.12fF $ **FLOATING
C9013 S.t606 VSUBS 0.02fF
C9014 S.n8194 VSUBS 0.14fF $ **FLOATING
C9015 S.n8196 VSUBS 5.44fF $ **FLOATING
C9016 S.t1474 VSUBS 0.02fF
C9017 S.n8197 VSUBS 0.12fF $ **FLOATING
C9018 S.n8198 VSUBS 0.14fF $ **FLOATING
C9019 S.t1257 VSUBS 0.02fF
C9020 S.n8200 VSUBS 0.24fF $ **FLOATING
C9021 S.n8201 VSUBS 0.91fF $ **FLOATING
C9022 S.n8202 VSUBS 0.05fF $ **FLOATING
C9023 S.t27 VSUBS 47.89fF
C9024 S.t1282 VSUBS 0.02fF
C9025 S.n8203 VSUBS 0.01fF $ **FLOATING
C9026 S.n8204 VSUBS 0.26fF $ **FLOATING
C9027 S.t2480 VSUBS 0.02fF
C9028 S.n8206 VSUBS 1.19fF $ **FLOATING
C9029 S.n8207 VSUBS 0.05fF $ **FLOATING
C9030 S.t2201 VSUBS 0.02fF
C9031 S.n8208 VSUBS 0.64fF $ **FLOATING
C9032 S.n8209 VSUBS 0.61fF $ **FLOATING
C9033 S.n8210 VSUBS 8.97fF $ **FLOATING
C9034 S.n8211 VSUBS 8.97fF $ **FLOATING
C9035 S.n8212 VSUBS 0.60fF $ **FLOATING
C9036 S.n8213 VSUBS 0.22fF $ **FLOATING
C9037 S.n8214 VSUBS 0.59fF $ **FLOATING
C9038 S.n8215 VSUBS 3.39fF $ **FLOATING
C9039 S.n8216 VSUBS 0.29fF $ **FLOATING
C9040 S.t79 VSUBS 21.42fF
C9041 S.n8217 VSUBS 21.71fF $ **FLOATING
C9042 S.n8218 VSUBS 0.77fF $ **FLOATING
C9043 S.n8219 VSUBS 0.28fF $ **FLOATING
C9044 S.n8220 VSUBS 4.00fF $ **FLOATING
C9045 S.n8221 VSUBS 1.35fF $ **FLOATING
C9046 S.n8222 VSUBS 0.01fF $ **FLOATING
C9047 S.n8223 VSUBS 0.02fF $ **FLOATING
C9048 S.n8224 VSUBS 0.03fF $ **FLOATING
C9049 S.n8225 VSUBS 0.04fF $ **FLOATING
C9050 S.n8226 VSUBS 0.17fF $ **FLOATING
C9051 S.n8227 VSUBS 0.01fF $ **FLOATING
C9052 S.n8228 VSUBS 0.02fF $ **FLOATING
C9053 S.n8229 VSUBS 0.01fF $ **FLOATING
C9054 S.n8230 VSUBS 0.01fF $ **FLOATING
C9055 S.n8231 VSUBS 0.01fF $ **FLOATING
C9056 S.n8232 VSUBS 0.01fF $ **FLOATING
C9057 S.n8233 VSUBS 0.02fF $ **FLOATING
C9058 S.n8234 VSUBS 0.01fF $ **FLOATING
C9059 S.n8235 VSUBS 0.02fF $ **FLOATING
C9060 S.n8236 VSUBS 0.05fF $ **FLOATING
C9061 S.n8237 VSUBS 0.04fF $ **FLOATING
C9062 S.n8238 VSUBS 0.11fF $ **FLOATING
C9063 S.n8239 VSUBS 0.38fF $ **FLOATING
C9064 S.n8240 VSUBS 0.20fF $ **FLOATING
C9065 S.n8241 VSUBS 4.39fF $ **FLOATING
C9066 S.n8242 VSUBS 0.24fF $ **FLOATING
C9067 S.n8243 VSUBS 1.50fF $ **FLOATING
C9068 S.n8244 VSUBS 1.31fF $ **FLOATING
C9069 S.n8245 VSUBS 0.28fF $ **FLOATING
C9070 S.n8246 VSUBS 1.89fF $ **FLOATING
C9071 S.n8247 VSUBS 0.06fF $ **FLOATING
C9072 S.n8248 VSUBS 0.03fF $ **FLOATING
C9073 S.n8249 VSUBS 0.04fF $ **FLOATING
C9074 S.n8250 VSUBS 0.99fF $ **FLOATING
C9075 S.n8251 VSUBS 0.02fF $ **FLOATING
C9076 S.n8252 VSUBS 0.01fF $ **FLOATING
C9077 S.n8253 VSUBS 0.02fF $ **FLOATING
C9078 S.n8254 VSUBS 0.08fF $ **FLOATING
C9079 S.n8255 VSUBS 0.36fF $ **FLOATING
C9080 S.n8256 VSUBS 1.85fF $ **FLOATING
C9081 S.t1528 VSUBS 0.02fF
C9082 S.n8257 VSUBS 0.24fF $ **FLOATING
C9083 S.n8258 VSUBS 0.36fF $ **FLOATING
C9084 S.n8259 VSUBS 0.61fF $ **FLOATING
C9085 S.n8260 VSUBS 0.12fF $ **FLOATING
C9086 S.t705 VSUBS 0.02fF
C9087 S.n8261 VSUBS 0.14fF $ **FLOATING
C9088 S.n8263 VSUBS 0.70fF $ **FLOATING
C9089 S.n8264 VSUBS 0.23fF $ **FLOATING
C9090 S.n8265 VSUBS 0.23fF $ **FLOATING
C9091 S.n8266 VSUBS 0.70fF $ **FLOATING
C9092 S.n8267 VSUBS 1.16fF $ **FLOATING
C9093 S.n8268 VSUBS 0.22fF $ **FLOATING
C9094 S.n8269 VSUBS 0.25fF $ **FLOATING
C9095 S.n8270 VSUBS 0.09fF $ **FLOATING
C9096 S.n8271 VSUBS 1.88fF $ **FLOATING
C9097 S.t1822 VSUBS 0.02fF
C9098 S.n8272 VSUBS 0.24fF $ **FLOATING
C9099 S.n8273 VSUBS 0.91fF $ **FLOATING
C9100 S.n8274 VSUBS 0.05fF $ **FLOATING
C9101 S.t1573 VSUBS 0.02fF
C9102 S.n8275 VSUBS 0.12fF $ **FLOATING
C9103 S.n8276 VSUBS 0.14fF $ **FLOATING
C9104 S.n8278 VSUBS 0.25fF $ **FLOATING
C9105 S.n8279 VSUBS 0.09fF $ **FLOATING
C9106 S.n8280 VSUBS 0.21fF $ **FLOATING
C9107 S.n8281 VSUBS 0.92fF $ **FLOATING
C9108 S.n8282 VSUBS 0.44fF $ **FLOATING
C9109 S.n8283 VSUBS 1.88fF $ **FLOATING
C9110 S.n8284 VSUBS 0.12fF $ **FLOATING
C9111 S.t1621 VSUBS 0.02fF
C9112 S.n8285 VSUBS 0.14fF $ **FLOATING
C9113 S.t2434 VSUBS 0.02fF
C9114 S.n8287 VSUBS 0.24fF $ **FLOATING
C9115 S.n8288 VSUBS 0.36fF $ **FLOATING
C9116 S.n8289 VSUBS 0.61fF $ **FLOATING
C9117 S.n8290 VSUBS 0.02fF $ **FLOATING
C9118 S.n8291 VSUBS 0.01fF $ **FLOATING
C9119 S.n8292 VSUBS 0.02fF $ **FLOATING
C9120 S.n8293 VSUBS 0.08fF $ **FLOATING
C9121 S.n8294 VSUBS 0.06fF $ **FLOATING
C9122 S.n8295 VSUBS 0.03fF $ **FLOATING
C9123 S.n8296 VSUBS 0.04fF $ **FLOATING
C9124 S.n8297 VSUBS 1.00fF $ **FLOATING
C9125 S.n8298 VSUBS 0.36fF $ **FLOATING
C9126 S.n8299 VSUBS 1.87fF $ **FLOATING
C9127 S.n8300 VSUBS 1.99fF $ **FLOATING
C9128 S.t211 VSUBS 0.02fF
C9129 S.n8301 VSUBS 0.24fF $ **FLOATING
C9130 S.n8302 VSUBS 0.91fF $ **FLOATING
C9131 S.n8303 VSUBS 0.05fF $ **FLOATING
C9132 S.t2492 VSUBS 0.02fF
C9133 S.n8304 VSUBS 0.12fF $ **FLOATING
C9134 S.n8305 VSUBS 0.14fF $ **FLOATING
C9135 S.n8307 VSUBS 1.89fF $ **FLOATING
C9136 S.n8308 VSUBS 0.07fF $ **FLOATING
C9137 S.n8309 VSUBS 0.04fF $ **FLOATING
C9138 S.n8310 VSUBS 0.05fF $ **FLOATING
C9139 S.n8311 VSUBS 0.87fF $ **FLOATING
C9140 S.n8312 VSUBS 0.01fF $ **FLOATING
C9141 S.n8313 VSUBS 0.01fF $ **FLOATING
C9142 S.n8314 VSUBS 0.01fF $ **FLOATING
C9143 S.n8315 VSUBS 0.07fF $ **FLOATING
C9144 S.n8316 VSUBS 0.68fF $ **FLOATING
C9145 S.n8317 VSUBS 0.72fF $ **FLOATING
C9146 S.t2063 VSUBS 0.02fF
C9147 S.n8318 VSUBS 0.24fF $ **FLOATING
C9148 S.n8319 VSUBS 0.36fF $ **FLOATING
C9149 S.n8320 VSUBS 0.61fF $ **FLOATING
C9150 S.n8321 VSUBS 0.12fF $ **FLOATING
C9151 S.t1245 VSUBS 0.02fF
C9152 S.n8322 VSUBS 0.14fF $ **FLOATING
C9153 S.n8324 VSUBS 0.70fF $ **FLOATING
C9154 S.n8325 VSUBS 0.23fF $ **FLOATING
C9155 S.n8326 VSUBS 0.23fF $ **FLOATING
C9156 S.n8327 VSUBS 0.70fF $ **FLOATING
C9157 S.n8328 VSUBS 1.16fF $ **FLOATING
C9158 S.n8329 VSUBS 0.22fF $ **FLOATING
C9159 S.n8330 VSUBS 0.25fF $ **FLOATING
C9160 S.n8331 VSUBS 0.09fF $ **FLOATING
C9161 S.n8332 VSUBS 2.31fF $ **FLOATING
C9162 S.t2337 VSUBS 0.02fF
C9163 S.n8333 VSUBS 0.24fF $ **FLOATING
C9164 S.n8334 VSUBS 0.91fF $ **FLOATING
C9165 S.n8335 VSUBS 0.05fF $ **FLOATING
C9166 S.t749 VSUBS 0.02fF
C9167 S.n8336 VSUBS 0.12fF $ **FLOATING
C9168 S.n8337 VSUBS 0.14fF $ **FLOATING
C9169 S.n8339 VSUBS 1.88fF $ **FLOATING
C9170 S.n8340 VSUBS 0.46fF $ **FLOATING
C9171 S.n8341 VSUBS 0.22fF $ **FLOATING
C9172 S.n8342 VSUBS 0.38fF $ **FLOATING
C9173 S.n8343 VSUBS 0.16fF $ **FLOATING
C9174 S.n8344 VSUBS 0.28fF $ **FLOATING
C9175 S.n8345 VSUBS 0.21fF $ **FLOATING
C9176 S.n8346 VSUBS 0.30fF $ **FLOATING
C9177 S.n8347 VSUBS 0.42fF $ **FLOATING
C9178 S.n8348 VSUBS 0.21fF $ **FLOATING
C9179 S.t328 VSUBS 0.02fF
C9180 S.n8349 VSUBS 0.24fF $ **FLOATING
C9181 S.n8350 VSUBS 0.36fF $ **FLOATING
C9182 S.n8351 VSUBS 0.61fF $ **FLOATING
C9183 S.n8352 VSUBS 0.12fF $ **FLOATING
C9184 S.t2030 VSUBS 0.02fF
C9185 S.n8353 VSUBS 0.14fF $ **FLOATING
C9186 S.n8355 VSUBS 0.04fF $ **FLOATING
C9187 S.n8356 VSUBS 0.03fF $ **FLOATING
C9188 S.n8357 VSUBS 0.03fF $ **FLOATING
C9189 S.n8358 VSUBS 0.10fF $ **FLOATING
C9190 S.n8359 VSUBS 0.36fF $ **FLOATING
C9191 S.n8360 VSUBS 0.38fF $ **FLOATING
C9192 S.n8361 VSUBS 0.11fF $ **FLOATING
C9193 S.n8362 VSUBS 0.12fF $ **FLOATING
C9194 S.n8363 VSUBS 0.07fF $ **FLOATING
C9195 S.n8364 VSUBS 0.12fF $ **FLOATING
C9196 S.n8365 VSUBS 0.18fF $ **FLOATING
C9197 S.n8366 VSUBS 3.99fF $ **FLOATING
C9198 S.t601 VSUBS 0.02fF
C9199 S.n8367 VSUBS 0.24fF $ **FLOATING
C9200 S.n8368 VSUBS 0.91fF $ **FLOATING
C9201 S.n8369 VSUBS 0.05fF $ **FLOATING
C9202 S.t380 VSUBS 0.02fF
C9203 S.n8370 VSUBS 0.12fF $ **FLOATING
C9204 S.n8371 VSUBS 0.14fF $ **FLOATING
C9205 S.n8373 VSUBS 0.25fF $ **FLOATING
C9206 S.n8374 VSUBS 0.09fF $ **FLOATING
C9207 S.n8375 VSUBS 0.21fF $ **FLOATING
C9208 S.n8376 VSUBS 1.28fF $ **FLOATING
C9209 S.n8377 VSUBS 0.53fF $ **FLOATING
C9210 S.n8378 VSUBS 1.88fF $ **FLOATING
C9211 S.n8379 VSUBS 0.12fF $ **FLOATING
C9212 S.t301 VSUBS 0.02fF
C9213 S.n8380 VSUBS 0.14fF $ **FLOATING
C9214 S.t1118 VSUBS 0.02fF
C9215 S.n8382 VSUBS 0.24fF $ **FLOATING
C9216 S.n8383 VSUBS 0.36fF $ **FLOATING
C9217 S.n8384 VSUBS 0.61fF $ **FLOATING
C9218 S.n8385 VSUBS 1.58fF $ **FLOATING
C9219 S.n8386 VSUBS 2.45fF $ **FLOATING
C9220 S.t1394 VSUBS 0.02fF
C9221 S.n8387 VSUBS 0.24fF $ **FLOATING
C9222 S.n8388 VSUBS 0.91fF $ **FLOATING
C9223 S.n8389 VSUBS 0.05fF $ **FLOATING
C9224 S.t1166 VSUBS 0.02fF
C9225 S.n8390 VSUBS 0.12fF $ **FLOATING
C9226 S.n8391 VSUBS 0.14fF $ **FLOATING
C9227 S.n8393 VSUBS 1.89fF $ **FLOATING
C9228 S.n8394 VSUBS 0.06fF $ **FLOATING
C9229 S.n8395 VSUBS 0.03fF $ **FLOATING
C9230 S.n8396 VSUBS 0.04fF $ **FLOATING
C9231 S.n8397 VSUBS 0.99fF $ **FLOATING
C9232 S.n8398 VSUBS 0.02fF $ **FLOATING
C9233 S.n8399 VSUBS 0.01fF $ **FLOATING
C9234 S.n8400 VSUBS 0.02fF $ **FLOATING
C9235 S.n8401 VSUBS 0.08fF $ **FLOATING
C9236 S.n8402 VSUBS 0.36fF $ **FLOATING
C9237 S.n8403 VSUBS 1.85fF $ **FLOATING
C9238 S.t1899 VSUBS 0.02fF
C9239 S.n8404 VSUBS 0.24fF $ **FLOATING
C9240 S.n8405 VSUBS 0.36fF $ **FLOATING
C9241 S.n8406 VSUBS 0.61fF $ **FLOATING
C9242 S.n8407 VSUBS 0.12fF $ **FLOATING
C9243 S.t1085 VSUBS 0.02fF
C9244 S.n8408 VSUBS 0.14fF $ **FLOATING
C9245 S.n8410 VSUBS 0.70fF $ **FLOATING
C9246 S.n8411 VSUBS 0.23fF $ **FLOATING
C9247 S.n8412 VSUBS 0.23fF $ **FLOATING
C9248 S.n8413 VSUBS 0.70fF $ **FLOATING
C9249 S.n8414 VSUBS 1.16fF $ **FLOATING
C9250 S.n8415 VSUBS 0.22fF $ **FLOATING
C9251 S.n8416 VSUBS 0.25fF $ **FLOATING
C9252 S.n8417 VSUBS 0.09fF $ **FLOATING
C9253 S.n8418 VSUBS 1.88fF $ **FLOATING
C9254 S.t2182 VSUBS 0.02fF
C9255 S.n8419 VSUBS 0.24fF $ **FLOATING
C9256 S.n8420 VSUBS 0.91fF $ **FLOATING
C9257 S.n8421 VSUBS 0.05fF $ **FLOATING
C9258 S.t1953 VSUBS 0.02fF
C9259 S.n8422 VSUBS 0.12fF $ **FLOATING
C9260 S.n8423 VSUBS 0.14fF $ **FLOATING
C9261 S.n8425 VSUBS 20.78fF $ **FLOATING
C9262 S.n8426 VSUBS 0.06fF $ **FLOATING
C9263 S.n8427 VSUBS 0.20fF $ **FLOATING
C9264 S.n8428 VSUBS 0.09fF $ **FLOATING
C9265 S.n8429 VSUBS 0.21fF $ **FLOATING
C9266 S.n8430 VSUBS 0.10fF $ **FLOATING
C9267 S.n8431 VSUBS 0.30fF $ **FLOATING
C9268 S.n8432 VSUBS 0.69fF $ **FLOATING
C9269 S.n8433 VSUBS 0.45fF $ **FLOATING
C9270 S.n8434 VSUBS 2.33fF $ **FLOATING
C9271 S.n8435 VSUBS 0.12fF $ **FLOATING
C9272 S.t2442 VSUBS 0.02fF
C9273 S.n8436 VSUBS 0.14fF $ **FLOATING
C9274 S.t735 VSUBS 0.02fF
C9275 S.n8438 VSUBS 0.24fF $ **FLOATING
C9276 S.n8439 VSUBS 0.36fF $ **FLOATING
C9277 S.n8440 VSUBS 0.61fF $ **FLOATING
C9278 S.n8441 VSUBS 1.90fF $ **FLOATING
C9279 S.n8442 VSUBS 0.17fF $ **FLOATING
C9280 S.n8443 VSUBS 0.76fF $ **FLOATING
C9281 S.n8444 VSUBS 0.25fF $ **FLOATING
C9282 S.n8445 VSUBS 0.30fF $ **FLOATING
C9283 S.n8446 VSUBS 0.32fF $ **FLOATING
C9284 S.n8447 VSUBS 0.47fF $ **FLOATING
C9285 S.n8448 VSUBS 0.16fF $ **FLOATING
C9286 S.n8449 VSUBS 1.93fF $ **FLOATING
C9287 S.t787 VSUBS 0.02fF
C9288 S.n8450 VSUBS 0.12fF $ **FLOATING
C9289 S.n8451 VSUBS 0.14fF $ **FLOATING
C9290 S.t1041 VSUBS 0.02fF
C9291 S.n8453 VSUBS 0.24fF $ **FLOATING
C9292 S.n8454 VSUBS 0.91fF $ **FLOATING
C9293 S.n8455 VSUBS 0.05fF $ **FLOATING
C9294 S.n8456 VSUBS 1.88fF $ **FLOATING
C9295 S.n8457 VSUBS 0.12fF $ **FLOATING
C9296 S.t2568 VSUBS 0.02fF
C9297 S.n8458 VSUBS 0.14fF $ **FLOATING
C9298 S.t1333 VSUBS 0.02fF
C9299 S.n8460 VSUBS 1.22fF $ **FLOATING
C9300 S.n8461 VSUBS 0.36fF $ **FLOATING
C9301 S.n8462 VSUBS 1.22fF $ **FLOATING
C9302 S.n8463 VSUBS 0.61fF $ **FLOATING
C9303 S.n8464 VSUBS 0.35fF $ **FLOATING
C9304 S.n8465 VSUBS 0.63fF $ **FLOATING
C9305 S.n8466 VSUBS 1.15fF $ **FLOATING
C9306 S.n8467 VSUBS 3.00fF $ **FLOATING
C9307 S.n8468 VSUBS 0.59fF $ **FLOATING
C9308 S.n8469 VSUBS 0.01fF $ **FLOATING
C9309 S.n8470 VSUBS 0.97fF $ **FLOATING
C9310 S.t320 VSUBS 21.42fF
C9311 S.n8471 VSUBS 20.29fF $ **FLOATING
C9312 S.n8473 VSUBS 0.38fF $ **FLOATING
C9313 S.n8474 VSUBS 0.23fF $ **FLOATING
C9314 S.n8475 VSUBS 2.79fF $ **FLOATING
C9315 S.n8476 VSUBS 2.46fF $ **FLOATING
C9316 S.n8477 VSUBS 4.00fF $ **FLOATING
C9317 S.n8478 VSUBS 0.25fF $ **FLOATING
C9318 S.n8479 VSUBS 0.01fF $ **FLOATING
C9319 S.t515 VSUBS 0.02fF
C9320 S.n8480 VSUBS 0.26fF $ **FLOATING
C9321 S.t1607 VSUBS 0.02fF
C9322 S.n8481 VSUBS 0.95fF $ **FLOATING
C9323 S.n8482 VSUBS 0.71fF $ **FLOATING
C9324 S.n8483 VSUBS 1.89fF $ **FLOATING
C9325 S.n8484 VSUBS 1.88fF $ **FLOATING
C9326 S.t2118 VSUBS 0.02fF
C9327 S.n8485 VSUBS 0.24fF $ **FLOATING
C9328 S.n8486 VSUBS 0.36fF $ **FLOATING
C9329 S.n8487 VSUBS 0.61fF $ **FLOATING
C9330 S.n8488 VSUBS 0.12fF $ **FLOATING
C9331 S.t1302 VSUBS 0.02fF
C9332 S.n8489 VSUBS 0.14fF $ **FLOATING
C9333 S.n8491 VSUBS 1.16fF $ **FLOATING
C9334 S.n8492 VSUBS 0.22fF $ **FLOATING
C9335 S.n8493 VSUBS 0.25fF $ **FLOATING
C9336 S.n8494 VSUBS 0.09fF $ **FLOATING
C9337 S.n8495 VSUBS 1.88fF $ **FLOATING
C9338 S.t2396 VSUBS 0.02fF
C9339 S.n8496 VSUBS 0.24fF $ **FLOATING
C9340 S.n8497 VSUBS 0.91fF $ **FLOATING
C9341 S.n8498 VSUBS 0.05fF $ **FLOATING
C9342 S.t2168 VSUBS 0.02fF
C9343 S.n8499 VSUBS 0.12fF $ **FLOATING
C9344 S.n8500 VSUBS 0.14fF $ **FLOATING
C9345 S.n8502 VSUBS 0.78fF $ **FLOATING
C9346 S.n8503 VSUBS 1.94fF $ **FLOATING
C9347 S.n8504 VSUBS 1.88fF $ **FLOATING
C9348 S.n8505 VSUBS 0.12fF $ **FLOATING
C9349 S.t2212 VSUBS 0.02fF
C9350 S.n8506 VSUBS 0.14fF $ **FLOATING
C9351 S.t387 VSUBS 0.02fF
C9352 S.n8508 VSUBS 0.24fF $ **FLOATING
C9353 S.n8509 VSUBS 0.36fF $ **FLOATING
C9354 S.n8510 VSUBS 0.61fF $ **FLOATING
C9355 S.n8511 VSUBS 1.84fF $ **FLOATING
C9356 S.n8512 VSUBS 2.99fF $ **FLOATING
C9357 S.t658 VSUBS 0.02fF
C9358 S.n8513 VSUBS 0.24fF $ **FLOATING
C9359 S.n8514 VSUBS 0.91fF $ **FLOATING
C9360 S.n8515 VSUBS 0.05fF $ **FLOATING
C9361 S.t436 VSUBS 0.02fF
C9362 S.n8516 VSUBS 0.12fF $ **FLOATING
C9363 S.n8517 VSUBS 0.14fF $ **FLOATING
C9364 S.n8519 VSUBS 1.89fF $ **FLOATING
C9365 S.n8520 VSUBS 1.75fF $ **FLOATING
C9366 S.t1293 VSUBS 0.02fF
C9367 S.n8521 VSUBS 0.24fF $ **FLOATING
C9368 S.n8522 VSUBS 0.36fF $ **FLOATING
C9369 S.n8523 VSUBS 0.61fF $ **FLOATING
C9370 S.n8524 VSUBS 0.12fF $ **FLOATING
C9371 S.t480 VSUBS 0.02fF
C9372 S.n8525 VSUBS 0.14fF $ **FLOATING
C9373 S.n8527 VSUBS 1.16fF $ **FLOATING
C9374 S.n8528 VSUBS 0.22fF $ **FLOATING
C9375 S.n8529 VSUBS 0.25fF $ **FLOATING
C9376 S.n8530 VSUBS 0.09fF $ **FLOATING
C9377 S.n8531 VSUBS 2.44fF $ **FLOATING
C9378 S.t1565 VSUBS 0.02fF
C9379 S.n8532 VSUBS 0.24fF $ **FLOATING
C9380 S.n8533 VSUBS 0.91fF $ **FLOATING
C9381 S.n8534 VSUBS 0.05fF $ **FLOATING
C9382 S.t1347 VSUBS 0.02fF
C9383 S.n8535 VSUBS 0.12fF $ **FLOATING
C9384 S.n8536 VSUBS 0.14fF $ **FLOATING
C9385 S.n8538 VSUBS 1.88fF $ **FLOATING
C9386 S.n8539 VSUBS 0.48fF $ **FLOATING
C9387 S.n8540 VSUBS 0.09fF $ **FLOATING
C9388 S.n8541 VSUBS 0.33fF $ **FLOATING
C9389 S.n8542 VSUBS 0.30fF $ **FLOATING
C9390 S.n8543 VSUBS 0.77fF $ **FLOATING
C9391 S.n8544 VSUBS 0.59fF $ **FLOATING
C9392 S.t902 VSUBS 0.02fF
C9393 S.n8545 VSUBS 0.24fF $ **FLOATING
C9394 S.n8546 VSUBS 0.36fF $ **FLOATING
C9395 S.n8547 VSUBS 0.61fF $ **FLOATING
C9396 S.n8548 VSUBS 0.12fF $ **FLOATING
C9397 S.t41 VSUBS 0.02fF
C9398 S.n8549 VSUBS 0.14fF $ **FLOATING
C9399 S.n8551 VSUBS 2.61fF $ **FLOATING
C9400 S.n8552 VSUBS 2.15fF $ **FLOATING
C9401 S.t1201 VSUBS 0.02fF
C9402 S.n8553 VSUBS 0.24fF $ **FLOATING
C9403 S.n8554 VSUBS 0.91fF $ **FLOATING
C9404 S.n8555 VSUBS 0.05fF $ **FLOATING
C9405 S.t953 VSUBS 0.02fF
C9406 S.n8556 VSUBS 0.12fF $ **FLOATING
C9407 S.n8557 VSUBS 0.14fF $ **FLOATING
C9408 S.n8559 VSUBS 0.78fF $ **FLOATING
C9409 S.n8560 VSUBS 2.30fF $ **FLOATING
C9410 S.n8561 VSUBS 1.88fF $ **FLOATING
C9411 S.n8562 VSUBS 0.12fF $ **FLOATING
C9412 S.t867 VSUBS 0.02fF
C9413 S.n8563 VSUBS 0.14fF $ **FLOATING
C9414 S.t1681 VSUBS 0.02fF
C9415 S.n8565 VSUBS 0.24fF $ **FLOATING
C9416 S.n8566 VSUBS 0.36fF $ **FLOATING
C9417 S.n8567 VSUBS 0.61fF $ **FLOATING
C9418 S.n8568 VSUBS 1.39fF $ **FLOATING
C9419 S.n8569 VSUBS 0.71fF $ **FLOATING
C9420 S.n8570 VSUBS 1.14fF $ **FLOATING
C9421 S.n8571 VSUBS 0.35fF $ **FLOATING
C9422 S.n8572 VSUBS 2.02fF $ **FLOATING
C9423 S.t1981 VSUBS 0.02fF
C9424 S.n8573 VSUBS 0.24fF $ **FLOATING
C9425 S.n8574 VSUBS 0.91fF $ **FLOATING
C9426 S.n8575 VSUBS 0.05fF $ **FLOATING
C9427 S.t1736 VSUBS 0.02fF
C9428 S.n8576 VSUBS 0.12fF $ **FLOATING
C9429 S.n8577 VSUBS 0.14fF $ **FLOATING
C9430 S.n8579 VSUBS 1.89fF $ **FLOATING
C9431 S.n8580 VSUBS 1.88fF $ **FLOATING
C9432 S.t2470 VSUBS 0.02fF
C9433 S.n8581 VSUBS 0.24fF $ **FLOATING
C9434 S.n8582 VSUBS 0.36fF $ **FLOATING
C9435 S.n8583 VSUBS 0.61fF $ **FLOATING
C9436 S.n8584 VSUBS 0.12fF $ **FLOATING
C9437 S.t1651 VSUBS 0.02fF
C9438 S.n8585 VSUBS 0.14fF $ **FLOATING
C9439 S.n8587 VSUBS 1.16fF $ **FLOATING
C9440 S.n8588 VSUBS 0.22fF $ **FLOATING
C9441 S.n8589 VSUBS 0.25fF $ **FLOATING
C9442 S.n8590 VSUBS 0.09fF $ **FLOATING
C9443 S.n8591 VSUBS 1.88fF $ **FLOATING
C9444 S.t249 VSUBS 0.02fF
C9445 S.n8592 VSUBS 0.24fF $ **FLOATING
C9446 S.n8593 VSUBS 0.91fF $ **FLOATING
C9447 S.n8594 VSUBS 0.05fF $ **FLOATING
C9448 S.t2520 VSUBS 0.02fF
C9449 S.n8595 VSUBS 0.12fF $ **FLOATING
C9450 S.n8596 VSUBS 0.14fF $ **FLOATING
C9451 S.n8598 VSUBS 20.78fF $ **FLOATING
C9452 S.n8599 VSUBS 1.88fF $ **FLOATING
C9453 S.n8600 VSUBS 2.67fF $ **FLOATING
C9454 S.t1267 VSUBS 0.02fF
C9455 S.n8601 VSUBS 0.24fF $ **FLOATING
C9456 S.n8602 VSUBS 0.36fF $ **FLOATING
C9457 S.n8603 VSUBS 0.61fF $ **FLOATING
C9458 S.n8604 VSUBS 0.12fF $ **FLOATING
C9459 S.t449 VSUBS 0.02fF
C9460 S.n8605 VSUBS 0.14fF $ **FLOATING
C9461 S.n8607 VSUBS 2.80fF $ **FLOATING
C9462 S.n8608 VSUBS 2.30fF $ **FLOATING
C9463 S.t1316 VSUBS 0.02fF
C9464 S.n8609 VSUBS 0.12fF $ **FLOATING
C9465 S.n8610 VSUBS 0.14fF $ **FLOATING
C9466 S.t1540 VSUBS 0.02fF
C9467 S.n8612 VSUBS 0.24fF $ **FLOATING
C9468 S.n8613 VSUBS 0.91fF $ **FLOATING
C9469 S.n8614 VSUBS 0.05fF $ **FLOATING
C9470 S.n8615 VSUBS 2.80fF $ **FLOATING
C9471 S.n8616 VSUBS 1.88fF $ **FLOATING
C9472 S.n8617 VSUBS 0.12fF $ **FLOATING
C9473 S.t1239 VSUBS 0.02fF
C9474 S.n8618 VSUBS 0.14fF $ **FLOATING
C9475 S.t2057 VSUBS 0.02fF
C9476 S.n8620 VSUBS 0.24fF $ **FLOATING
C9477 S.n8621 VSUBS 0.36fF $ **FLOATING
C9478 S.n8622 VSUBS 0.61fF $ **FLOATING
C9479 S.n8623 VSUBS 2.67fF $ **FLOATING
C9480 S.n8624 VSUBS 2.30fF $ **FLOATING
C9481 S.t2104 VSUBS 0.02fF
C9482 S.n8625 VSUBS 0.12fF $ **FLOATING
C9483 S.n8626 VSUBS 0.14fF $ **FLOATING
C9484 S.t2328 VSUBS 0.02fF
C9485 S.n8628 VSUBS 0.24fF $ **FLOATING
C9486 S.n8629 VSUBS 0.91fF $ **FLOATING
C9487 S.n8630 VSUBS 0.05fF $ **FLOATING
C9488 S.n8631 VSUBS 1.88fF $ **FLOATING
C9489 S.n8632 VSUBS 2.67fF $ **FLOATING
C9490 S.t321 VSUBS 0.02fF
C9491 S.n8633 VSUBS 0.24fF $ **FLOATING
C9492 S.n8634 VSUBS 0.36fF $ **FLOATING
C9493 S.n8635 VSUBS 0.61fF $ **FLOATING
C9494 S.n8636 VSUBS 0.12fF $ **FLOATING
C9495 S.t2023 VSUBS 0.02fF
C9496 S.n8637 VSUBS 0.14fF $ **FLOATING
C9497 S.n8639 VSUBS 2.80fF $ **FLOATING
C9498 S.n8640 VSUBS 2.30fF $ **FLOATING
C9499 S.t374 VSUBS 0.02fF
C9500 S.n8641 VSUBS 0.12fF $ **FLOATING
C9501 S.n8642 VSUBS 0.14fF $ **FLOATING
C9502 S.t592 VSUBS 0.02fF
C9503 S.n8644 VSUBS 0.24fF $ **FLOATING
C9504 S.n8645 VSUBS 0.91fF $ **FLOATING
C9505 S.n8646 VSUBS 0.05fF $ **FLOATING
C9506 S.n8647 VSUBS 1.88fF $ **FLOATING
C9507 S.n8648 VSUBS 2.67fF $ **FLOATING
C9508 S.t1111 VSUBS 0.02fF
C9509 S.n8649 VSUBS 0.24fF $ **FLOATING
C9510 S.n8650 VSUBS 0.36fF $ **FLOATING
C9511 S.n8651 VSUBS 0.61fF $ **FLOATING
C9512 S.n8652 VSUBS 0.12fF $ **FLOATING
C9513 S.t416 VSUBS 0.02fF
C9514 S.n8653 VSUBS 0.14fF $ **FLOATING
C9515 S.n8655 VSUBS 2.80fF $ **FLOATING
C9516 S.n8656 VSUBS 2.30fF $ **FLOATING
C9517 S.t1162 VSUBS 0.02fF
C9518 S.n8657 VSUBS 0.12fF $ **FLOATING
C9519 S.n8658 VSUBS 0.14fF $ **FLOATING
C9520 S.t1386 VSUBS 0.02fF
C9521 S.n8660 VSUBS 0.24fF $ **FLOATING
C9522 S.n8661 VSUBS 0.91fF $ **FLOATING
C9523 S.n8662 VSUBS 0.05fF $ **FLOATING
C9524 S.n8663 VSUBS 1.88fF $ **FLOATING
C9525 S.n8664 VSUBS 2.67fF $ **FLOATING
C9526 S.t1432 VSUBS 0.02fF
C9527 S.n8665 VSUBS 0.24fF $ **FLOATING
C9528 S.n8666 VSUBS 0.36fF $ **FLOATING
C9529 S.n8667 VSUBS 0.61fF $ **FLOATING
C9530 S.n8668 VSUBS 0.12fF $ **FLOATING
C9531 S.t1629 VSUBS 0.02fF
C9532 S.n8669 VSUBS 0.14fF $ **FLOATING
C9533 S.n8671 VSUBS 2.80fF $ **FLOATING
C9534 S.n8672 VSUBS 2.30fF $ **FLOATING
C9535 S.t2500 VSUBS 0.02fF
C9536 S.n8673 VSUBS 0.12fF $ **FLOATING
C9537 S.n8674 VSUBS 0.14fF $ **FLOATING
C9538 S.t2274 VSUBS 0.02fF
C9539 S.n8676 VSUBS 0.24fF $ **FLOATING
C9540 S.n8677 VSUBS 0.91fF $ **FLOATING
C9541 S.n8678 VSUBS 0.05fF $ **FLOATING
C9542 S.n8679 VSUBS 1.88fF $ **FLOATING
C9543 S.n8680 VSUBS 2.67fF $ **FLOATING
C9544 S.t2223 VSUBS 0.02fF
C9545 S.n8681 VSUBS 0.24fF $ **FLOATING
C9546 S.n8682 VSUBS 0.36fF $ **FLOATING
C9547 S.n8683 VSUBS 0.61fF $ **FLOATING
C9548 S.n8684 VSUBS 0.12fF $ **FLOATING
C9549 S.t2415 VSUBS 0.02fF
C9550 S.n8685 VSUBS 0.14fF $ **FLOATING
C9551 S.n8687 VSUBS 2.80fF $ **FLOATING
C9552 S.n8688 VSUBS 2.30fF $ **FLOATING
C9553 S.t758 VSUBS 0.02fF
C9554 S.n8689 VSUBS 0.12fF $ **FLOATING
C9555 S.n8690 VSUBS 0.14fF $ **FLOATING
C9556 S.t546 VSUBS 0.02fF
C9557 S.n8692 VSUBS 0.24fF $ **FLOATING
C9558 S.n8693 VSUBS 0.91fF $ **FLOATING
C9559 S.n8694 VSUBS 0.05fF $ **FLOATING
C9560 S.n8695 VSUBS 1.88fF $ **FLOATING
C9561 S.n8696 VSUBS 2.67fF $ **FLOATING
C9562 S.t489 VSUBS 0.02fF
C9563 S.n8697 VSUBS 0.24fF $ **FLOATING
C9564 S.n8698 VSUBS 0.36fF $ **FLOATING
C9565 S.n8699 VSUBS 0.61fF $ **FLOATING
C9566 S.n8700 VSUBS 0.12fF $ **FLOATING
C9567 S.t679 VSUBS 0.02fF
C9568 S.n8701 VSUBS 0.14fF $ **FLOATING
C9569 S.n8703 VSUBS 2.80fF $ **FLOATING
C9570 S.n8704 VSUBS 2.30fF $ **FLOATING
C9571 S.t1548 VSUBS 0.02fF
C9572 S.n8705 VSUBS 0.12fF $ **FLOATING
C9573 S.n8706 VSUBS 0.14fF $ **FLOATING
C9574 S.t1334 VSUBS 0.02fF
C9575 S.n8708 VSUBS 0.24fF $ **FLOATING
C9576 S.n8709 VSUBS 0.91fF $ **FLOATING
C9577 S.n8710 VSUBS 0.05fF $ **FLOATING
C9578 S.n8711 VSUBS 1.88fF $ **FLOATING
C9579 S.n8712 VSUBS 2.68fF $ **FLOATING
C9580 S.t1275 VSUBS 0.02fF
C9581 S.n8713 VSUBS 0.24fF $ **FLOATING
C9582 S.n8714 VSUBS 0.36fF $ **FLOATING
C9583 S.n8715 VSUBS 0.61fF $ **FLOATING
C9584 S.n8716 VSUBS 0.12fF $ **FLOATING
C9585 S.t1469 VSUBS 0.02fF
C9586 S.n8717 VSUBS 0.14fF $ **FLOATING
C9587 S.n8719 VSUBS 5.17fF $ **FLOATING
C9588 S.t2336 VSUBS 0.02fF
C9589 S.n8720 VSUBS 0.12fF $ **FLOATING
C9590 S.n8721 VSUBS 0.14fF $ **FLOATING
C9591 S.t2121 VSUBS 0.02fF
C9592 S.n8723 VSUBS 0.24fF $ **FLOATING
C9593 S.n8724 VSUBS 0.91fF $ **FLOATING
C9594 S.n8725 VSUBS 0.05fF $ **FLOATING
C9595 S.n8726 VSUBS 2.73fF $ **FLOATING
C9596 S.n8727 VSUBS 1.59fF $ **FLOATING
C9597 S.n8728 VSUBS 0.12fF $ **FLOATING
C9598 S.t2220 VSUBS 0.02fF
C9599 S.n8729 VSUBS 0.14fF $ **FLOATING
C9600 S.t760 VSUBS 0.02fF
C9601 S.n8731 VSUBS 0.24fF $ **FLOATING
C9602 S.n8732 VSUBS 0.36fF $ **FLOATING
C9603 S.n8733 VSUBS 0.61fF $ **FLOATING
C9604 S.n8734 VSUBS 0.07fF $ **FLOATING
C9605 S.n8735 VSUBS 0.01fF $ **FLOATING
C9606 S.n8736 VSUBS 0.24fF $ **FLOATING
C9607 S.n8737 VSUBS 1.16fF $ **FLOATING
C9608 S.n8738 VSUBS 1.35fF $ **FLOATING
C9609 S.n8739 VSUBS 2.30fF $ **FLOATING
C9610 S.t599 VSUBS 0.02fF
C9611 S.n8740 VSUBS 0.12fF $ **FLOATING
C9612 S.n8741 VSUBS 0.14fF $ **FLOATING
C9613 S.t2171 VSUBS 0.02fF
C9614 S.n8743 VSUBS 0.24fF $ **FLOATING
C9615 S.n8744 VSUBS 0.91fF $ **FLOATING
C9616 S.n8745 VSUBS 0.05fF $ **FLOATING
C9617 S.t40 VSUBS 48.27fF
C9618 S.t782 VSUBS 0.02fF
C9619 S.n8746 VSUBS 0.12fF $ **FLOATING
C9620 S.n8747 VSUBS 0.14fF $ **FLOATING
C9621 S.t1029 VSUBS 0.02fF
C9622 S.n8749 VSUBS 0.24fF $ **FLOATING
C9623 S.n8750 VSUBS 0.91fF $ **FLOATING
C9624 S.n8751 VSUBS 0.05fF $ **FLOATING
C9625 S.t725 VSUBS 0.02fF
C9626 S.n8752 VSUBS 0.24fF $ **FLOATING
C9627 S.n8753 VSUBS 0.36fF $ **FLOATING
C9628 S.n8754 VSUBS 0.61fF $ **FLOATING
C9629 S.n8755 VSUBS 0.32fF $ **FLOATING
C9630 S.n8756 VSUBS 1.09fF $ **FLOATING
C9631 S.n8757 VSUBS 0.15fF $ **FLOATING
C9632 S.n8758 VSUBS 2.10fF $ **FLOATING
C9633 S.n8759 VSUBS 2.94fF $ **FLOATING
C9634 S.n8760 VSUBS 1.88fF $ **FLOATING
C9635 S.n8761 VSUBS 0.12fF $ **FLOATING
C9636 S.t1996 VSUBS 0.02fF
C9637 S.n8762 VSUBS 0.14fF $ **FLOATING
C9638 S.t295 VSUBS 0.02fF
C9639 S.n8764 VSUBS 0.24fF $ **FLOATING
C9640 S.n8765 VSUBS 0.36fF $ **FLOATING
C9641 S.n8766 VSUBS 0.61fF $ **FLOATING
C9642 S.n8767 VSUBS 0.92fF $ **FLOATING
C9643 S.n8768 VSUBS 0.32fF $ **FLOATING
C9644 S.n8769 VSUBS 0.92fF $ **FLOATING
C9645 S.n8770 VSUBS 1.09fF $ **FLOATING
C9646 S.n8771 VSUBS 0.15fF $ **FLOATING
C9647 S.n8772 VSUBS 4.96fF $ **FLOATING
C9648 S.t348 VSUBS 0.02fF
C9649 S.n8773 VSUBS 0.12fF $ **FLOATING
C9650 S.n8774 VSUBS 0.14fF $ **FLOATING
C9651 S.t569 VSUBS 0.02fF
C9652 S.n8776 VSUBS 0.24fF $ **FLOATING
C9653 S.n8777 VSUBS 0.91fF $ **FLOATING
C9654 S.n8778 VSUBS 0.05fF $ **FLOATING
C9655 S.n8779 VSUBS 1.88fF $ **FLOATING
C9656 S.n8780 VSUBS 2.67fF $ **FLOATING
C9657 S.t2407 VSUBS 0.02fF
C9658 S.n8781 VSUBS 0.24fF $ **FLOATING
C9659 S.n8782 VSUBS 0.36fF $ **FLOATING
C9660 S.n8783 VSUBS 0.61fF $ **FLOATING
C9661 S.n8784 VSUBS 0.12fF $ **FLOATING
C9662 S.t1589 VSUBS 0.02fF
C9663 S.n8785 VSUBS 0.14fF $ **FLOATING
C9664 S.n8787 VSUBS 1.88fF $ **FLOATING
C9665 S.n8788 VSUBS 2.67fF $ **FLOATING
C9666 S.t479 VSUBS 0.02fF
C9667 S.n8789 VSUBS 0.24fF $ **FLOATING
C9668 S.n8790 VSUBS 0.36fF $ **FLOATING
C9669 S.n8791 VSUBS 0.61fF $ **FLOATING
C9670 S.t748 VSUBS 0.02fF
C9671 S.n8792 VSUBS 0.24fF $ **FLOATING
C9672 S.n8793 VSUBS 0.91fF $ **FLOATING
C9673 S.n8794 VSUBS 0.05fF $ **FLOATING
C9674 S.t1698 VSUBS 0.02fF
C9675 S.n8795 VSUBS 0.12fF $ **FLOATING
C9676 S.n8796 VSUBS 0.14fF $ **FLOATING
C9677 S.n8798 VSUBS 0.12fF $ **FLOATING
C9678 S.t2184 VSUBS 0.02fF
C9679 S.n8799 VSUBS 0.14fF $ **FLOATING
C9680 S.n8801 VSUBS 2.30fF $ **FLOATING
C9681 S.n8802 VSUBS 2.94fF $ **FLOATING
C9682 S.n8803 VSUBS 5.16fF $ **FLOATING
C9683 S.t2462 VSUBS 0.02fF
C9684 S.n8804 VSUBS 0.12fF $ **FLOATING
C9685 S.n8805 VSUBS 0.14fF $ **FLOATING
C9686 S.t179 VSUBS 0.02fF
C9687 S.n8807 VSUBS 0.24fF $ **FLOATING
C9688 S.n8808 VSUBS 0.91fF $ **FLOATING
C9689 S.n8809 VSUBS 0.05fF $ **FLOATING
C9690 S.n8810 VSUBS 1.88fF $ **FLOATING
C9691 S.n8811 VSUBS 2.67fF $ **FLOATING
C9692 S.t671 VSUBS 0.02fF
C9693 S.n8812 VSUBS 0.24fF $ **FLOATING
C9694 S.n8813 VSUBS 0.36fF $ **FLOATING
C9695 S.n8814 VSUBS 0.61fF $ **FLOATING
C9696 S.n8815 VSUBS 0.12fF $ **FLOATING
C9697 S.t2380 VSUBS 0.02fF
C9698 S.n8816 VSUBS 0.14fF $ **FLOATING
C9699 S.n8818 VSUBS 5.17fF $ **FLOATING
C9700 S.t720 VSUBS 0.02fF
C9701 S.n8819 VSUBS 0.12fF $ **FLOATING
C9702 S.n8820 VSUBS 0.14fF $ **FLOATING
C9703 S.t966 VSUBS 0.02fF
C9704 S.n8822 VSUBS 0.24fF $ **FLOATING
C9705 S.n8823 VSUBS 0.91fF $ **FLOATING
C9706 S.n8824 VSUBS 0.05fF $ **FLOATING
C9707 S.n8825 VSUBS 1.88fF $ **FLOATING
C9708 S.n8826 VSUBS 0.12fF $ **FLOATING
C9709 S.t645 VSUBS 0.02fF
C9710 S.n8827 VSUBS 0.14fF $ **FLOATING
C9711 S.t1458 VSUBS 0.02fF
C9712 S.n8829 VSUBS 0.24fF $ **FLOATING
C9713 S.n8830 VSUBS 0.36fF $ **FLOATING
C9714 S.n8831 VSUBS 0.61fF $ **FLOATING
C9715 S.n8832 VSUBS 2.67fF $ **FLOATING
C9716 S.n8833 VSUBS 5.17fF $ **FLOATING
C9717 S.t1512 VSUBS 0.02fF
C9718 S.n8834 VSUBS 0.12fF $ **FLOATING
C9719 S.n8835 VSUBS 0.14fF $ **FLOATING
C9720 S.t1748 VSUBS 0.02fF
C9721 S.n8837 VSUBS 0.24fF $ **FLOATING
C9722 S.n8838 VSUBS 0.91fF $ **FLOATING
C9723 S.n8839 VSUBS 0.05fF $ **FLOATING
C9724 S.n8840 VSUBS 1.88fF $ **FLOATING
C9725 S.n8841 VSUBS 2.67fF $ **FLOATING
C9726 S.t2249 VSUBS 0.02fF
C9727 S.n8842 VSUBS 0.24fF $ **FLOATING
C9728 S.n8843 VSUBS 0.36fF $ **FLOATING
C9729 S.n8844 VSUBS 0.61fF $ **FLOATING
C9730 S.n8845 VSUBS 0.12fF $ **FLOATING
C9731 S.t1433 VSUBS 0.02fF
C9732 S.n8846 VSUBS 0.14fF $ **FLOATING
C9733 S.n8848 VSUBS 5.17fF $ **FLOATING
C9734 S.t2301 VSUBS 0.02fF
C9735 S.n8849 VSUBS 0.12fF $ **FLOATING
C9736 S.n8850 VSUBS 0.14fF $ **FLOATING
C9737 S.t2531 VSUBS 0.02fF
C9738 S.n8852 VSUBS 0.24fF $ **FLOATING
C9739 S.n8853 VSUBS 0.91fF $ **FLOATING
C9740 S.n8854 VSUBS 0.05fF $ **FLOATING
C9741 S.n8855 VSUBS 1.88fF $ **FLOATING
C9742 S.n8856 VSUBS 2.67fF $ **FLOATING
C9743 S.t621 VSUBS 0.02fF
C9744 S.n8857 VSUBS 0.24fF $ **FLOATING
C9745 S.n8858 VSUBS 0.36fF $ **FLOATING
C9746 S.n8859 VSUBS 0.61fF $ **FLOATING
C9747 S.n8860 VSUBS 0.12fF $ **FLOATING
C9748 S.t820 VSUBS 0.02fF
C9749 S.n8861 VSUBS 0.14fF $ **FLOATING
C9750 S.n8863 VSUBS 5.17fF $ **FLOATING
C9751 S.t689 VSUBS 0.02fF
C9752 S.n8864 VSUBS 0.12fF $ **FLOATING
C9753 S.n8865 VSUBS 0.14fF $ **FLOATING
C9754 S.t1460 VSUBS 0.02fF
C9755 S.n8867 VSUBS 0.24fF $ **FLOATING
C9756 S.n8868 VSUBS 0.91fF $ **FLOATING
C9757 S.n8869 VSUBS 0.05fF $ **FLOATING
C9758 S.n8870 VSUBS 1.88fF $ **FLOATING
C9759 S.n8871 VSUBS 2.67fF $ **FLOATING
C9760 S.t1411 VSUBS 0.02fF
C9761 S.n8872 VSUBS 0.24fF $ **FLOATING
C9762 S.n8873 VSUBS 0.36fF $ **FLOATING
C9763 S.n8874 VSUBS 0.61fF $ **FLOATING
C9764 S.n8875 VSUBS 0.12fF $ **FLOATING
C9765 S.t1602 VSUBS 0.02fF
C9766 S.n8876 VSUBS 0.14fF $ **FLOATING
C9767 S.n8878 VSUBS 5.17fF $ **FLOATING
C9768 S.t2473 VSUBS 0.02fF
C9769 S.n8879 VSUBS 0.12fF $ **FLOATING
C9770 S.n8880 VSUBS 0.14fF $ **FLOATING
C9771 S.t2250 VSUBS 0.02fF
C9772 S.n8882 VSUBS 0.24fF $ **FLOATING
C9773 S.n8883 VSUBS 0.91fF $ **FLOATING
C9774 S.n8884 VSUBS 0.05fF $ **FLOATING
C9775 S.n8885 VSUBS 1.88fF $ **FLOATING
C9776 S.n8886 VSUBS 2.67fF $ **FLOATING
C9777 S.t2200 VSUBS 0.02fF
C9778 S.n8887 VSUBS 0.24fF $ **FLOATING
C9779 S.n8888 VSUBS 0.36fF $ **FLOATING
C9780 S.n8889 VSUBS 0.61fF $ **FLOATING
C9781 S.n8890 VSUBS 0.12fF $ **FLOATING
C9782 S.t2390 VSUBS 0.02fF
C9783 S.n8891 VSUBS 0.14fF $ **FLOATING
C9784 S.n8893 VSUBS 5.17fF $ **FLOATING
C9785 S.t731 VSUBS 0.02fF
C9786 S.n8894 VSUBS 0.12fF $ **FLOATING
C9787 S.n8895 VSUBS 0.14fF $ **FLOATING
C9788 S.t518 VSUBS 0.02fF
C9789 S.n8897 VSUBS 0.24fF $ **FLOATING
C9790 S.n8898 VSUBS 0.91fF $ **FLOATING
C9791 S.n8899 VSUBS 0.05fF $ **FLOATING
C9792 S.n8900 VSUBS 1.88fF $ **FLOATING
C9793 S.n8901 VSUBS 2.67fF $ **FLOATING
C9794 S.t467 VSUBS 0.02fF
C9795 S.n8902 VSUBS 0.24fF $ **FLOATING
C9796 S.n8903 VSUBS 0.36fF $ **FLOATING
C9797 S.n8904 VSUBS 0.61fF $ **FLOATING
C9798 S.n8905 VSUBS 0.12fF $ **FLOATING
C9799 S.t654 VSUBS 0.02fF
C9800 S.n8906 VSUBS 0.14fF $ **FLOATING
C9801 S.n8908 VSUBS 4.89fF $ **FLOATING
C9802 S.t1524 VSUBS 0.02fF
C9803 S.n8909 VSUBS 0.12fF $ **FLOATING
C9804 S.n8910 VSUBS 0.14fF $ **FLOATING
C9805 S.t1304 VSUBS 0.02fF
C9806 S.n8912 VSUBS 0.24fF $ **FLOATING
C9807 S.n8913 VSUBS 0.91fF $ **FLOATING
C9808 S.n8914 VSUBS 0.05fF $ **FLOATING
C9809 S.n8915 VSUBS 1.88fF $ **FLOATING
C9810 S.n8916 VSUBS 2.67fF $ **FLOATING
C9811 S.t1254 VSUBS 0.02fF
C9812 S.n8917 VSUBS 0.24fF $ **FLOATING
C9813 S.n8918 VSUBS 0.36fF $ **FLOATING
C9814 S.n8919 VSUBS 0.61fF $ **FLOATING
C9815 S.n8920 VSUBS 0.12fF $ **FLOATING
C9816 S.t1444 VSUBS 0.02fF
C9817 S.n8921 VSUBS 0.14fF $ **FLOATING
C9818 S.n8923 VSUBS 5.44fF $ **FLOATING
C9819 S.t2312 VSUBS 0.02fF
C9820 S.n8924 VSUBS 0.12fF $ **FLOATING
C9821 S.n8925 VSUBS 0.14fF $ **FLOATING
C9822 S.t2091 VSUBS 0.02fF
C9823 S.n8927 VSUBS 0.24fF $ **FLOATING
C9824 S.n8928 VSUBS 0.91fF $ **FLOATING
C9825 S.n8929 VSUBS 0.05fF $ **FLOATING
C9826 S.t300 VSUBS 47.89fF
C9827 S.t1073 VSUBS 0.02fF
C9828 S.n8930 VSUBS 0.01fF $ **FLOATING
C9829 S.n8931 VSUBS 0.26fF $ **FLOATING
C9830 S.t1922 VSUBS 0.02fF
C9831 S.n8933 VSUBS 1.19fF $ **FLOATING
C9832 S.n8934 VSUBS 0.05fF $ **FLOATING
C9833 S.t1620 VSUBS 0.02fF
C9834 S.n8935 VSUBS 0.64fF $ **FLOATING
C9835 S.n8936 VSUBS 0.61fF $ **FLOATING
C9836 S.n8937 VSUBS 8.97fF $ **FLOATING
C9837 S.n8938 VSUBS 8.97fF $ **FLOATING
C9838 S.n8939 VSUBS 0.60fF $ **FLOATING
C9839 S.n8940 VSUBS 0.22fF $ **FLOATING
C9840 S.n8941 VSUBS 0.59fF $ **FLOATING
C9841 S.n8942 VSUBS 3.39fF $ **FLOATING
C9842 S.n8943 VSUBS 0.29fF $ **FLOATING
C9843 S.t248 VSUBS 21.42fF
C9844 S.n8944 VSUBS 21.71fF $ **FLOATING
C9845 S.n8945 VSUBS 0.77fF $ **FLOATING
C9846 S.n8946 VSUBS 0.28fF $ **FLOATING
C9847 S.n8947 VSUBS 4.00fF $ **FLOATING
C9848 S.n8948 VSUBS 1.35fF $ **FLOATING
C9849 S.n8949 VSUBS 0.01fF $ **FLOATING
C9850 S.n8950 VSUBS 0.02fF $ **FLOATING
C9851 S.n8951 VSUBS 0.03fF $ **FLOATING
C9852 S.n8952 VSUBS 0.04fF $ **FLOATING
C9853 S.n8953 VSUBS 0.17fF $ **FLOATING
C9854 S.n8954 VSUBS 0.01fF $ **FLOATING
C9855 S.n8955 VSUBS 0.02fF $ **FLOATING
C9856 S.n8956 VSUBS 0.01fF $ **FLOATING
C9857 S.n8957 VSUBS 0.01fF $ **FLOATING
C9858 S.n8958 VSUBS 0.01fF $ **FLOATING
C9859 S.n8959 VSUBS 0.01fF $ **FLOATING
C9860 S.n8960 VSUBS 0.02fF $ **FLOATING
C9861 S.n8961 VSUBS 0.01fF $ **FLOATING
C9862 S.n8962 VSUBS 0.02fF $ **FLOATING
C9863 S.n8963 VSUBS 0.05fF $ **FLOATING
C9864 S.n8964 VSUBS 0.04fF $ **FLOATING
C9865 S.n8965 VSUBS 0.11fF $ **FLOATING
C9866 S.n8966 VSUBS 0.38fF $ **FLOATING
C9867 S.n8967 VSUBS 0.20fF $ **FLOATING
C9868 S.n8968 VSUBS 4.39fF $ **FLOATING
C9869 S.n8969 VSUBS 0.24fF $ **FLOATING
C9870 S.n8970 VSUBS 1.50fF $ **FLOATING
C9871 S.n8971 VSUBS 1.31fF $ **FLOATING
C9872 S.n8972 VSUBS 0.28fF $ **FLOATING
C9873 S.n8973 VSUBS 0.25fF $ **FLOATING
C9874 S.n8974 VSUBS 0.09fF $ **FLOATING
C9875 S.n8975 VSUBS 0.21fF $ **FLOATING
C9876 S.n8976 VSUBS 0.92fF $ **FLOATING
C9877 S.n8977 VSUBS 0.44fF $ **FLOATING
C9878 S.n8978 VSUBS 1.88fF $ **FLOATING
C9879 S.n8979 VSUBS 0.12fF $ **FLOATING
C9880 S.t136 VSUBS 0.02fF
C9881 S.n8980 VSUBS 0.14fF $ **FLOATING
C9882 S.t961 VSUBS 0.02fF
C9883 S.n8982 VSUBS 0.24fF $ **FLOATING
C9884 S.n8983 VSUBS 0.36fF $ **FLOATING
C9885 S.n8984 VSUBS 0.61fF $ **FLOATING
C9886 S.n8985 VSUBS 0.02fF $ **FLOATING
C9887 S.n8986 VSUBS 0.01fF $ **FLOATING
C9888 S.n8987 VSUBS 0.02fF $ **FLOATING
C9889 S.n8988 VSUBS 0.08fF $ **FLOATING
C9890 S.n8989 VSUBS 0.06fF $ **FLOATING
C9891 S.n8990 VSUBS 0.03fF $ **FLOATING
C9892 S.n8991 VSUBS 0.04fF $ **FLOATING
C9893 S.n8992 VSUBS 1.00fF $ **FLOATING
C9894 S.n8993 VSUBS 0.36fF $ **FLOATING
C9895 S.n8994 VSUBS 1.87fF $ **FLOATING
C9896 S.n8995 VSUBS 1.99fF $ **FLOATING
C9897 S.t1253 VSUBS 0.02fF
C9898 S.n8996 VSUBS 0.24fF $ **FLOATING
C9899 S.n8997 VSUBS 0.91fF $ **FLOATING
C9900 S.n8998 VSUBS 0.05fF $ **FLOATING
C9901 S.t1020 VSUBS 0.02fF
C9902 S.n8999 VSUBS 0.12fF $ **FLOATING
C9903 S.n9000 VSUBS 0.14fF $ **FLOATING
C9904 S.n9002 VSUBS 1.89fF $ **FLOATING
C9905 S.n9003 VSUBS 0.07fF $ **FLOATING
C9906 S.n9004 VSUBS 0.04fF $ **FLOATING
C9907 S.n9005 VSUBS 0.05fF $ **FLOATING
C9908 S.n9006 VSUBS 0.87fF $ **FLOATING
C9909 S.n9007 VSUBS 0.01fF $ **FLOATING
C9910 S.n9008 VSUBS 0.01fF $ **FLOATING
C9911 S.n9009 VSUBS 0.01fF $ **FLOATING
C9912 S.n9010 VSUBS 0.07fF $ **FLOATING
C9913 S.n9011 VSUBS 0.68fF $ **FLOATING
C9914 S.n9012 VSUBS 0.72fF $ **FLOATING
C9915 S.t1880 VSUBS 0.02fF
C9916 S.n9013 VSUBS 0.24fF $ **FLOATING
C9917 S.n9014 VSUBS 0.36fF $ **FLOATING
C9918 S.n9015 VSUBS 0.61fF $ **FLOATING
C9919 S.n9016 VSUBS 0.12fF $ **FLOATING
C9920 S.t1065 VSUBS 0.02fF
C9921 S.n9017 VSUBS 0.14fF $ **FLOATING
C9922 S.n9019 VSUBS 0.70fF $ **FLOATING
C9923 S.n9020 VSUBS 0.23fF $ **FLOATING
C9924 S.n9021 VSUBS 0.23fF $ **FLOATING
C9925 S.n9022 VSUBS 0.70fF $ **FLOATING
C9926 S.n9023 VSUBS 1.16fF $ **FLOATING
C9927 S.n9024 VSUBS 0.22fF $ **FLOATING
C9928 S.n9025 VSUBS 0.25fF $ **FLOATING
C9929 S.n9026 VSUBS 0.09fF $ **FLOATING
C9930 S.n9027 VSUBS 2.31fF $ **FLOATING
C9931 S.t2161 VSUBS 0.02fF
C9932 S.n9028 VSUBS 0.24fF $ **FLOATING
C9933 S.n9029 VSUBS 0.91fF $ **FLOATING
C9934 S.n9030 VSUBS 0.05fF $ **FLOATING
C9935 S.t1934 VSUBS 0.02fF
C9936 S.n9031 VSUBS 0.12fF $ **FLOATING
C9937 S.n9032 VSUBS 0.14fF $ **FLOATING
C9938 S.n9034 VSUBS 1.88fF $ **FLOATING
C9939 S.n9035 VSUBS 0.46fF $ **FLOATING
C9940 S.n9036 VSUBS 0.22fF $ **FLOATING
C9941 S.n9037 VSUBS 0.38fF $ **FLOATING
C9942 S.n9038 VSUBS 0.16fF $ **FLOATING
C9943 S.n9039 VSUBS 0.28fF $ **FLOATING
C9944 S.n9040 VSUBS 0.21fF $ **FLOATING
C9945 S.n9041 VSUBS 0.30fF $ **FLOATING
C9946 S.n9042 VSUBS 0.42fF $ **FLOATING
C9947 S.n9043 VSUBS 0.21fF $ **FLOATING
C9948 S.t1482 VSUBS 0.02fF
C9949 S.n9044 VSUBS 0.24fF $ **FLOATING
C9950 S.n9045 VSUBS 0.36fF $ **FLOATING
C9951 S.n9046 VSUBS 0.61fF $ **FLOATING
C9952 S.n9047 VSUBS 0.12fF $ **FLOATING
C9953 S.t661 VSUBS 0.02fF
C9954 S.n9048 VSUBS 0.14fF $ **FLOATING
C9955 S.n9050 VSUBS 0.04fF $ **FLOATING
C9956 S.n9051 VSUBS 0.03fF $ **FLOATING
C9957 S.n9052 VSUBS 0.03fF $ **FLOATING
C9958 S.n9053 VSUBS 0.10fF $ **FLOATING
C9959 S.n9054 VSUBS 0.36fF $ **FLOATING
C9960 S.n9055 VSUBS 0.38fF $ **FLOATING
C9961 S.n9056 VSUBS 0.11fF $ **FLOATING
C9962 S.n9057 VSUBS 0.12fF $ **FLOATING
C9963 S.n9058 VSUBS 0.07fF $ **FLOATING
C9964 S.n9059 VSUBS 0.12fF $ **FLOATING
C9965 S.n9060 VSUBS 0.18fF $ **FLOATING
C9966 S.n9061 VSUBS 3.99fF $ **FLOATING
C9967 S.t1771 VSUBS 0.02fF
C9968 S.n9062 VSUBS 0.24fF $ **FLOATING
C9969 S.n9063 VSUBS 0.91fF $ **FLOATING
C9970 S.n9064 VSUBS 0.05fF $ **FLOATING
C9971 S.t191 VSUBS 0.02fF
C9972 S.n9065 VSUBS 0.12fF $ **FLOATING
C9973 S.n9066 VSUBS 0.14fF $ **FLOATING
C9974 S.n9068 VSUBS 0.25fF $ **FLOATING
C9975 S.n9069 VSUBS 0.09fF $ **FLOATING
C9976 S.n9070 VSUBS 0.21fF $ **FLOATING
C9977 S.n9071 VSUBS 1.28fF $ **FLOATING
C9978 S.n9072 VSUBS 0.53fF $ **FLOATING
C9979 S.n9073 VSUBS 1.88fF $ **FLOATING
C9980 S.n9074 VSUBS 0.12fF $ **FLOATING
C9981 S.t1451 VSUBS 0.02fF
C9982 S.n9075 VSUBS 0.14fF $ **FLOATING
C9983 S.t2265 VSUBS 0.02fF
C9984 S.n9077 VSUBS 0.24fF $ **FLOATING
C9985 S.n9078 VSUBS 0.36fF $ **FLOATING
C9986 S.n9079 VSUBS 0.61fF $ **FLOATING
C9987 S.n9080 VSUBS 1.58fF $ **FLOATING
C9988 S.n9081 VSUBS 2.45fF $ **FLOATING
C9989 S.t2548 VSUBS 0.02fF
C9990 S.n9082 VSUBS 0.24fF $ **FLOATING
C9991 S.n9083 VSUBS 0.91fF $ **FLOATING
C9992 S.n9084 VSUBS 0.05fF $ **FLOATING
C9993 S.t2316 VSUBS 0.02fF
C9994 S.n9085 VSUBS 0.12fF $ **FLOATING
C9995 S.n9086 VSUBS 0.14fF $ **FLOATING
C9996 S.n9088 VSUBS 1.89fF $ **FLOATING
C9997 S.n9089 VSUBS 0.06fF $ **FLOATING
C9998 S.n9090 VSUBS 0.03fF $ **FLOATING
C9999 S.n9091 VSUBS 0.04fF $ **FLOATING
C10000 S.n9092 VSUBS 0.99fF $ **FLOATING
C10001 S.n9093 VSUBS 0.02fF $ **FLOATING
C10002 S.n9094 VSUBS 0.01fF $ **FLOATING
C10003 S.n9095 VSUBS 0.02fF $ **FLOATING
C10004 S.n9096 VSUBS 0.08fF $ **FLOATING
C10005 S.n9097 VSUBS 0.36fF $ **FLOATING
C10006 S.n9098 VSUBS 1.85fF $ **FLOATING
C10007 S.t538 VSUBS 0.02fF
C10008 S.n9099 VSUBS 0.24fF $ **FLOATING
C10009 S.n9100 VSUBS 0.36fF $ **FLOATING
C10010 S.n9101 VSUBS 0.61fF $ **FLOATING
C10011 S.n9102 VSUBS 0.12fF $ **FLOATING
C10012 S.t2241 VSUBS 0.02fF
C10013 S.n9103 VSUBS 0.14fF $ **FLOATING
C10014 S.n9105 VSUBS 0.70fF $ **FLOATING
C10015 S.n9106 VSUBS 0.23fF $ **FLOATING
C10016 S.n9107 VSUBS 0.23fF $ **FLOATING
C10017 S.n9108 VSUBS 0.70fF $ **FLOATING
C10018 S.n9109 VSUBS 1.16fF $ **FLOATING
C10019 S.n9110 VSUBS 0.22fF $ **FLOATING
C10020 S.n9111 VSUBS 0.25fF $ **FLOATING
C10021 S.n9112 VSUBS 0.09fF $ **FLOATING
C10022 S.n9113 VSUBS 1.88fF $ **FLOATING
C10023 S.t816 VSUBS 0.02fF
C10024 S.n9114 VSUBS 0.24fF $ **FLOATING
C10025 S.n9115 VSUBS 0.91fF $ **FLOATING
C10026 S.n9116 VSUBS 0.05fF $ **FLOATING
C10027 S.t582 VSUBS 0.02fF
C10028 S.n9117 VSUBS 0.12fF $ **FLOATING
C10029 S.n9118 VSUBS 0.14fF $ **FLOATING
C10030 S.n9120 VSUBS 20.78fF $ **FLOATING
C10031 S.n9121 VSUBS 1.72fF $ **FLOATING
C10032 S.n9122 VSUBS 3.05fF $ **FLOATING
C10033 S.t177 VSUBS 0.02fF
C10034 S.n9123 VSUBS 0.24fF $ **FLOATING
C10035 S.n9124 VSUBS 0.36fF $ **FLOATING
C10036 S.n9125 VSUBS 0.61fF $ **FLOATING
C10037 S.n9126 VSUBS 0.12fF $ **FLOATING
C10038 S.t1887 VSUBS 0.02fF
C10039 S.n9127 VSUBS 0.14fF $ **FLOATING
C10040 S.n9129 VSUBS 0.31fF $ **FLOATING
C10041 S.n9130 VSUBS 0.23fF $ **FLOATING
C10042 S.n9131 VSUBS 0.66fF $ **FLOATING
C10043 S.n9132 VSUBS 0.95fF $ **FLOATING
C10044 S.n9133 VSUBS 0.23fF $ **FLOATING
C10045 S.n9134 VSUBS 0.21fF $ **FLOATING
C10046 S.n9135 VSUBS 0.20fF $ **FLOATING
C10047 S.n9136 VSUBS 0.06fF $ **FLOATING
C10048 S.n9137 VSUBS 0.09fF $ **FLOATING
C10049 S.n9138 VSUBS 0.10fF $ **FLOATING
C10050 S.n9139 VSUBS 1.99fF $ **FLOATING
C10051 S.t233 VSUBS 0.02fF
C10052 S.n9140 VSUBS 0.12fF $ **FLOATING
C10053 S.n9141 VSUBS 0.14fF $ **FLOATING
C10054 S.t466 VSUBS 0.02fF
C10055 S.n9143 VSUBS 0.24fF $ **FLOATING
C10056 S.n9144 VSUBS 0.91fF $ **FLOATING
C10057 S.n9145 VSUBS 0.05fF $ **FLOATING
C10058 S.n9146 VSUBS 1.88fF $ **FLOATING
C10059 S.n9147 VSUBS 0.12fF $ **FLOATING
C10060 S.t1100 VSUBS 0.02fF
C10061 S.n9148 VSUBS 0.14fF $ **FLOATING
C10062 S.t1965 VSUBS 0.02fF
C10063 S.n9150 VSUBS 0.12fF $ **FLOATING
C10064 S.n9151 VSUBS 0.14fF $ **FLOATING
C10065 S.t2193 VSUBS 0.02fF
C10066 S.n9153 VSUBS 0.24fF $ **FLOATING
C10067 S.n9154 VSUBS 0.91fF $ **FLOATING
C10068 S.n9155 VSUBS 0.05fF $ **FLOATING
C10069 S.t1913 VSUBS 0.02fF
C10070 S.n9156 VSUBS 0.24fF $ **FLOATING
C10071 S.n9157 VSUBS 0.36fF $ **FLOATING
C10072 S.n9158 VSUBS 0.61fF $ **FLOATING
C10073 S.n9159 VSUBS 0.32fF $ **FLOATING
C10074 S.n9160 VSUBS 1.09fF $ **FLOATING
C10075 S.n9161 VSUBS 0.15fF $ **FLOATING
C10076 S.n9162 VSUBS 2.10fF $ **FLOATING
C10077 S.n9163 VSUBS 2.94fF $ **FLOATING
C10078 S.n9164 VSUBS 1.88fF $ **FLOATING
C10079 S.n9165 VSUBS 0.12fF $ **FLOATING
C10080 S.t510 VSUBS 0.02fF
C10081 S.n9166 VSUBS 0.14fF $ **FLOATING
C10082 S.t1325 VSUBS 0.02fF
C10083 S.n9168 VSUBS 0.24fF $ **FLOATING
C10084 S.n9169 VSUBS 0.36fF $ **FLOATING
C10085 S.n9170 VSUBS 0.61fF $ **FLOATING
C10086 S.n9171 VSUBS 0.92fF $ **FLOATING
C10087 S.n9172 VSUBS 0.32fF $ **FLOATING
C10088 S.n9173 VSUBS 0.92fF $ **FLOATING
C10089 S.n9174 VSUBS 1.09fF $ **FLOATING
C10090 S.n9175 VSUBS 0.15fF $ **FLOATING
C10091 S.n9176 VSUBS 4.96fF $ **FLOATING
C10092 S.t1376 VSUBS 0.02fF
C10093 S.n9177 VSUBS 0.12fF $ **FLOATING
C10094 S.n9178 VSUBS 0.14fF $ **FLOATING
C10095 S.t1597 VSUBS 0.02fF
C10096 S.n9180 VSUBS 0.24fF $ **FLOATING
C10097 S.n9181 VSUBS 0.91fF $ **FLOATING
C10098 S.n9182 VSUBS 0.05fF $ **FLOATING
C10099 S.n9183 VSUBS 1.88fF $ **FLOATING
C10100 S.n9184 VSUBS 2.67fF $ **FLOATING
C10101 S.t2233 VSUBS 0.02fF
C10102 S.n9185 VSUBS 0.24fF $ **FLOATING
C10103 S.n9186 VSUBS 0.36fF $ **FLOATING
C10104 S.n9187 VSUBS 0.61fF $ **FLOATING
C10105 S.n9188 VSUBS 0.12fF $ **FLOATING
C10106 S.t1417 VSUBS 0.02fF
C10107 S.n9189 VSUBS 0.14fF $ **FLOATING
C10108 S.n9191 VSUBS 1.88fF $ **FLOATING
C10109 S.n9192 VSUBS 2.67fF $ **FLOATING
C10110 S.t167 VSUBS 0.02fF
C10111 S.n9193 VSUBS 0.24fF $ **FLOATING
C10112 S.n9194 VSUBS 0.36fF $ **FLOATING
C10113 S.n9195 VSUBS 0.61fF $ **FLOATING
C10114 S.t458 VSUBS 0.02fF
C10115 S.n9196 VSUBS 0.24fF $ **FLOATING
C10116 S.n9197 VSUBS 0.91fF $ **FLOATING
C10117 S.n9198 VSUBS 0.05fF $ **FLOATING
C10118 S.t226 VSUBS 0.02fF
C10119 S.n9199 VSUBS 0.12fF $ **FLOATING
C10120 S.n9200 VSUBS 0.14fF $ **FLOATING
C10121 S.n9202 VSUBS 0.12fF $ **FLOATING
C10122 S.t2003 VSUBS 0.02fF
C10123 S.n9203 VSUBS 0.14fF $ **FLOATING
C10124 S.n9205 VSUBS 2.30fF $ **FLOATING
C10125 S.n9206 VSUBS 2.94fF $ **FLOATING
C10126 S.n9207 VSUBS 5.16fF $ **FLOATING
C10127 S.t2279 VSUBS 0.02fF
C10128 S.n9208 VSUBS 0.12fF $ **FLOATING
C10129 S.n9209 VSUBS 0.14fF $ **FLOATING
C10130 S.t2517 VSUBS 0.02fF
C10131 S.n9211 VSUBS 0.24fF $ **FLOATING
C10132 S.n9212 VSUBS 0.91fF $ **FLOATING
C10133 S.n9213 VSUBS 0.05fF $ **FLOATING
C10134 S.n9214 VSUBS 1.88fF $ **FLOATING
C10135 S.n9215 VSUBS 2.67fF $ **FLOATING
C10136 S.t1850 VSUBS 0.02fF
C10137 S.n9216 VSUBS 0.24fF $ **FLOATING
C10138 S.n9217 VSUBS 0.36fF $ **FLOATING
C10139 S.n9218 VSUBS 0.61fF $ **FLOATING
C10140 S.n9219 VSUBS 0.12fF $ **FLOATING
C10141 S.t1034 VSUBS 0.02fF
C10142 S.n9220 VSUBS 0.14fF $ **FLOATING
C10143 S.n9222 VSUBS 5.17fF $ **FLOATING
C10144 S.t1902 VSUBS 0.02fF
C10145 S.n9223 VSUBS 0.12fF $ **FLOATING
C10146 S.n9224 VSUBS 0.14fF $ **FLOATING
C10147 S.t2133 VSUBS 0.02fF
C10148 S.n9226 VSUBS 0.24fF $ **FLOATING
C10149 S.n9227 VSUBS 0.91fF $ **FLOATING
C10150 S.n9228 VSUBS 0.05fF $ **FLOATING
C10151 S.n9229 VSUBS 1.88fF $ **FLOATING
C10152 S.n9230 VSUBS 0.12fF $ **FLOATING
C10153 S.t1816 VSUBS 0.02fF
C10154 S.n9231 VSUBS 0.14fF $ **FLOATING
C10155 S.t82 VSUBS 0.02fF
C10156 S.n9233 VSUBS 0.24fF $ **FLOATING
C10157 S.n9234 VSUBS 0.36fF $ **FLOATING
C10158 S.n9235 VSUBS 0.61fF $ **FLOATING
C10159 S.n9236 VSUBS 2.67fF $ **FLOATING
C10160 S.n9237 VSUBS 5.17fF $ **FLOATING
C10161 S.t153 VSUBS 0.02fF
C10162 S.n9238 VSUBS 0.12fF $ **FLOATING
C10163 S.n9239 VSUBS 0.14fF $ **FLOATING
C10164 S.t402 VSUBS 0.02fF
C10165 S.n9241 VSUBS 0.24fF $ **FLOATING
C10166 S.n9242 VSUBS 0.91fF $ **FLOATING
C10167 S.n9243 VSUBS 0.05fF $ **FLOATING
C10168 S.n9244 VSUBS 1.88fF $ **FLOATING
C10169 S.n9245 VSUBS 2.67fF $ **FLOATING
C10170 S.t894 VSUBS 0.02fF
C10171 S.n9246 VSUBS 0.24fF $ **FLOATING
C10172 S.n9247 VSUBS 0.36fF $ **FLOATING
C10173 S.n9248 VSUBS 0.61fF $ **FLOATING
C10174 S.n9249 VSUBS 0.12fF $ **FLOATING
C10175 S.t32 VSUBS 0.02fF
C10176 S.n9250 VSUBS 0.14fF $ **FLOATING
C10177 S.n9252 VSUBS 5.17fF $ **FLOATING
C10178 S.t947 VSUBS 0.02fF
C10179 S.n9253 VSUBS 0.12fF $ **FLOATING
C10180 S.n9254 VSUBS 0.14fF $ **FLOATING
C10181 S.t1192 VSUBS 0.02fF
C10182 S.n9256 VSUBS 0.24fF $ **FLOATING
C10183 S.n9257 VSUBS 0.91fF $ **FLOATING
C10184 S.n9258 VSUBS 0.05fF $ **FLOATING
C10185 S.n9259 VSUBS 1.88fF $ **FLOATING
C10186 S.n9260 VSUBS 2.67fF $ **FLOATING
C10187 S.t1675 VSUBS 0.02fF
C10188 S.n9261 VSUBS 0.24fF $ **FLOATING
C10189 S.n9262 VSUBS 0.36fF $ **FLOATING
C10190 S.n9263 VSUBS 0.61fF $ **FLOATING
C10191 S.n9264 VSUBS 0.12fF $ **FLOATING
C10192 S.t863 VSUBS 0.02fF
C10193 S.n9265 VSUBS 0.14fF $ **FLOATING
C10194 S.n9267 VSUBS 5.17fF $ **FLOATING
C10195 S.t1730 VSUBS 0.02fF
C10196 S.n9268 VSUBS 0.12fF $ **FLOATING
C10197 S.n9269 VSUBS 0.14fF $ **FLOATING
C10198 S.t1972 VSUBS 0.02fF
C10199 S.n9271 VSUBS 0.24fF $ **FLOATING
C10200 S.n9272 VSUBS 0.91fF $ **FLOATING
C10201 S.n9273 VSUBS 0.05fF $ **FLOATING
C10202 S.n9274 VSUBS 1.88fF $ **FLOATING
C10203 S.n9275 VSUBS 2.67fF $ **FLOATING
C10204 S.t1455 VSUBS 0.02fF
C10205 S.n9276 VSUBS 0.24fF $ **FLOATING
C10206 S.n9277 VSUBS 0.36fF $ **FLOATING
C10207 S.n9278 VSUBS 0.61fF $ **FLOATING
C10208 S.n9279 VSUBS 0.12fF $ **FLOATING
C10209 S.t1654 VSUBS 0.02fF
C10210 S.n9280 VSUBS 0.14fF $ **FLOATING
C10211 S.n9282 VSUBS 5.17fF $ **FLOATING
C10212 S.t101 VSUBS 0.02fF
C10213 S.n9283 VSUBS 0.12fF $ **FLOATING
C10214 S.n9284 VSUBS 0.14fF $ **FLOATING
C10215 S.t2300 VSUBS 0.02fF
C10216 S.n9286 VSUBS 0.24fF $ **FLOATING
C10217 S.n9287 VSUBS 0.91fF $ **FLOATING
C10218 S.n9288 VSUBS 0.05fF $ **FLOATING
C10219 S.n9289 VSUBS 1.88fF $ **FLOATING
C10220 S.n9290 VSUBS 2.67fF $ **FLOATING
C10221 S.t2245 VSUBS 0.02fF
C10222 S.n9291 VSUBS 0.24fF $ **FLOATING
C10223 S.n9292 VSUBS 0.36fF $ **FLOATING
C10224 S.n9293 VSUBS 0.61fF $ **FLOATING
C10225 S.n9294 VSUBS 0.12fF $ **FLOATING
C10226 S.t2436 VSUBS 0.02fF
C10227 S.n9295 VSUBS 0.14fF $ **FLOATING
C10228 S.n9297 VSUBS 5.17fF $ **FLOATING
C10229 S.t784 VSUBS 0.02fF
C10230 S.n9298 VSUBS 0.12fF $ **FLOATING
C10231 S.n9299 VSUBS 0.14fF $ **FLOATING
C10232 S.t570 VSUBS 0.02fF
C10233 S.n9301 VSUBS 0.24fF $ **FLOATING
C10234 S.n9302 VSUBS 0.91fF $ **FLOATING
C10235 S.n9303 VSUBS 0.05fF $ **FLOATING
C10236 S.n9304 VSUBS 1.88fF $ **FLOATING
C10237 S.n9305 VSUBS 2.67fF $ **FLOATING
C10238 S.t514 VSUBS 0.02fF
C10239 S.n9306 VSUBS 0.24fF $ **FLOATING
C10240 S.n9307 VSUBS 0.36fF $ **FLOATING
C10241 S.n9308 VSUBS 0.61fF $ **FLOATING
C10242 S.n9309 VSUBS 0.12fF $ **FLOATING
C10243 S.t701 VSUBS 0.02fF
C10244 S.n9310 VSUBS 0.14fF $ **FLOATING
C10245 S.n9312 VSUBS 5.17fF $ **FLOATING
C10246 S.t1566 VSUBS 0.02fF
C10247 S.n9313 VSUBS 0.12fF $ **FLOATING
C10248 S.n9314 VSUBS 0.14fF $ **FLOATING
C10249 S.t1357 VSUBS 0.02fF
C10250 S.n9316 VSUBS 0.24fF $ **FLOATING
C10251 S.n9317 VSUBS 0.91fF $ **FLOATING
C10252 S.n9318 VSUBS 0.05fF $ **FLOATING
C10253 S.n9319 VSUBS 1.88fF $ **FLOATING
C10254 S.n9320 VSUBS 2.67fF $ **FLOATING
C10255 S.t1301 VSUBS 0.02fF
C10256 S.n9321 VSUBS 0.24fF $ **FLOATING
C10257 S.n9322 VSUBS 0.36fF $ **FLOATING
C10258 S.n9323 VSUBS 0.61fF $ **FLOATING
C10259 S.n9324 VSUBS 0.12fF $ **FLOATING
C10260 S.t1496 VSUBS 0.02fF
C10261 S.n9325 VSUBS 0.14fF $ **FLOATING
C10262 S.n9327 VSUBS 4.89fF $ **FLOATING
C10263 S.t2359 VSUBS 0.02fF
C10264 S.n9328 VSUBS 0.12fF $ **FLOATING
C10265 S.n9329 VSUBS 0.14fF $ **FLOATING
C10266 S.t2142 VSUBS 0.02fF
C10267 S.n9331 VSUBS 0.24fF $ **FLOATING
C10268 S.n9332 VSUBS 0.91fF $ **FLOATING
C10269 S.n9333 VSUBS 0.05fF $ **FLOATING
C10270 S.n9334 VSUBS 1.88fF $ **FLOATING
C10271 S.n9335 VSUBS 2.67fF $ **FLOATING
C10272 S.t2090 VSUBS 0.02fF
C10273 S.n9336 VSUBS 0.24fF $ **FLOATING
C10274 S.n9337 VSUBS 0.36fF $ **FLOATING
C10275 S.n9338 VSUBS 0.61fF $ **FLOATING
C10276 S.n9339 VSUBS 0.12fF $ **FLOATING
C10277 S.t2280 VSUBS 0.02fF
C10278 S.n9340 VSUBS 0.14fF $ **FLOATING
C10279 S.n9342 VSUBS 1.88fF $ **FLOATING
C10280 S.n9343 VSUBS 2.68fF $ **FLOATING
C10281 S.t2115 VSUBS 0.02fF
C10282 S.n9344 VSUBS 0.24fF $ **FLOATING
C10283 S.n9345 VSUBS 0.36fF $ **FLOATING
C10284 S.n9346 VSUBS 0.61fF $ **FLOATING
C10285 S.t747 VSUBS 0.02fF
C10286 S.n9347 VSUBS 1.22fF $ **FLOATING
C10287 S.n9348 VSUBS 0.61fF $ **FLOATING
C10288 S.n9349 VSUBS 0.35fF $ **FLOATING
C10289 S.n9350 VSUBS 0.63fF $ **FLOATING
C10290 S.n9351 VSUBS 1.15fF $ **FLOATING
C10291 S.n9352 VSUBS 3.00fF $ **FLOATING
C10292 S.n9353 VSUBS 0.59fF $ **FLOATING
C10293 S.n9354 VSUBS 0.01fF $ **FLOATING
C10294 S.n9355 VSUBS 0.97fF $ **FLOATING
C10295 S.t166 VSUBS 21.42fF
C10296 S.n9356 VSUBS 20.29fF $ **FLOATING
C10297 S.n9358 VSUBS 0.38fF $ **FLOATING
C10298 S.n9359 VSUBS 0.23fF $ **FLOATING
C10299 S.n9360 VSUBS 2.90fF $ **FLOATING
C10300 S.n9361 VSUBS 2.46fF $ **FLOATING
C10301 S.n9362 VSUBS 1.96fF $ **FLOATING
C10302 S.n9363 VSUBS 3.94fF $ **FLOATING
C10303 S.n9364 VSUBS 0.25fF $ **FLOATING
C10304 S.n9365 VSUBS 0.01fF $ **FLOATING
C10305 S.t2460 VSUBS 0.02fF
C10306 S.n9366 VSUBS 0.26fF $ **FLOATING
C10307 S.t1051 VSUBS 0.02fF
C10308 S.n9367 VSUBS 0.95fF $ **FLOATING
C10309 S.n9368 VSUBS 0.71fF $ **FLOATING
C10310 S.n9369 VSUBS 0.78fF $ **FLOATING
C10311 S.n9370 VSUBS 1.93fF $ **FLOATING
C10312 S.n9371 VSUBS 1.88fF $ **FLOATING
C10313 S.n9372 VSUBS 0.12fF $ **FLOATING
C10314 S.t718 VSUBS 0.02fF
C10315 S.n9373 VSUBS 0.14fF $ **FLOATING
C10316 S.t1539 VSUBS 0.02fF
C10317 S.n9375 VSUBS 0.24fF $ **FLOATING
C10318 S.n9376 VSUBS 0.36fF $ **FLOATING
C10319 S.n9377 VSUBS 0.61fF $ **FLOATING
C10320 S.n9378 VSUBS 1.52fF $ **FLOATING
C10321 S.n9379 VSUBS 2.99fF $ **FLOATING
C10322 S.t1834 VSUBS 0.02fF
C10323 S.n9380 VSUBS 0.24fF $ **FLOATING
C10324 S.n9381 VSUBS 0.91fF $ **FLOATING
C10325 S.n9382 VSUBS 0.05fF $ **FLOATING
C10326 S.t1586 VSUBS 0.02fF
C10327 S.n9383 VSUBS 0.12fF $ **FLOATING
C10328 S.n9384 VSUBS 0.14fF $ **FLOATING
C10329 S.n9386 VSUBS 1.89fF $ **FLOATING
C10330 S.n9387 VSUBS 1.75fF $ **FLOATING
C10331 S.t2324 VSUBS 0.02fF
C10332 S.n9388 VSUBS 0.24fF $ **FLOATING
C10333 S.n9389 VSUBS 0.36fF $ **FLOATING
C10334 S.n9390 VSUBS 0.61fF $ **FLOATING
C10335 S.n9391 VSUBS 0.12fF $ **FLOATING
C10336 S.t1632 VSUBS 0.02fF
C10337 S.n9392 VSUBS 0.14fF $ **FLOATING
C10338 S.n9394 VSUBS 1.16fF $ **FLOATING
C10339 S.n9395 VSUBS 0.22fF $ **FLOATING
C10340 S.n9396 VSUBS 0.25fF $ **FLOATING
C10341 S.n9397 VSUBS 0.09fF $ **FLOATING
C10342 S.n9398 VSUBS 2.44fF $ **FLOATING
C10343 S.t56 VSUBS 0.02fF
C10344 S.n9399 VSUBS 0.24fF $ **FLOATING
C10345 S.n9400 VSUBS 0.91fF $ **FLOATING
C10346 S.n9401 VSUBS 0.05fF $ **FLOATING
C10347 S.t2376 VSUBS 0.02fF
C10348 S.n9402 VSUBS 0.12fF $ **FLOATING
C10349 S.n9403 VSUBS 0.14fF $ **FLOATING
C10350 S.n9405 VSUBS 1.88fF $ **FLOATING
C10351 S.n9406 VSUBS 0.48fF $ **FLOATING
C10352 S.n9407 VSUBS 0.09fF $ **FLOATING
C10353 S.n9408 VSUBS 0.33fF $ **FLOATING
C10354 S.n9409 VSUBS 0.30fF $ **FLOATING
C10355 S.n9410 VSUBS 0.77fF $ **FLOATING
C10356 S.n9411 VSUBS 0.59fF $ **FLOATING
C10357 S.t706 VSUBS 0.02fF
C10358 S.n9412 VSUBS 0.24fF $ **FLOATING
C10359 S.n9413 VSUBS 0.36fF $ **FLOATING
C10360 S.n9414 VSUBS 0.61fF $ **FLOATING
C10361 S.n9415 VSUBS 0.12fF $ **FLOATING
C10362 S.t2416 VSUBS 0.02fF
C10363 S.n9416 VSUBS 0.14fF $ **FLOATING
C10364 S.n9418 VSUBS 2.61fF $ **FLOATING
C10365 S.n9419 VSUBS 2.15fF $ **FLOATING
C10366 S.t1012 VSUBS 0.02fF
C10367 S.n9420 VSUBS 0.24fF $ **FLOATING
C10368 S.n9421 VSUBS 0.91fF $ **FLOATING
C10369 S.n9422 VSUBS 0.05fF $ **FLOATING
C10370 S.t761 VSUBS 0.02fF
C10371 S.n9423 VSUBS 0.12fF $ **FLOATING
C10372 S.n9424 VSUBS 0.14fF $ **FLOATING
C10373 S.n9426 VSUBS 0.78fF $ **FLOATING
C10374 S.n9427 VSUBS 2.30fF $ **FLOATING
C10375 S.n9428 VSUBS 1.88fF $ **FLOATING
C10376 S.n9429 VSUBS 0.12fF $ **FLOATING
C10377 S.t2043 VSUBS 0.02fF
C10378 S.n9430 VSUBS 0.14fF $ **FLOATING
C10379 S.t343 VSUBS 0.02fF
C10380 S.n9432 VSUBS 0.24fF $ **FLOATING
C10381 S.n9433 VSUBS 0.36fF $ **FLOATING
C10382 S.n9434 VSUBS 0.61fF $ **FLOATING
C10383 S.n9435 VSUBS 1.39fF $ **FLOATING
C10384 S.n9436 VSUBS 0.71fF $ **FLOATING
C10385 S.n9437 VSUBS 1.14fF $ **FLOATING
C10386 S.n9438 VSUBS 0.35fF $ **FLOATING
C10387 S.n9439 VSUBS 2.02fF $ **FLOATING
C10388 S.t613 VSUBS 0.02fF
C10389 S.n9440 VSUBS 0.24fF $ **FLOATING
C10390 S.n9441 VSUBS 0.91fF $ **FLOATING
C10391 S.n9442 VSUBS 0.05fF $ **FLOATING
C10392 S.t390 VSUBS 0.02fF
C10393 S.n9443 VSUBS 0.12fF $ **FLOATING
C10394 S.n9444 VSUBS 0.14fF $ **FLOATING
C10395 S.n9446 VSUBS 1.89fF $ **FLOATING
C10396 S.n9447 VSUBS 1.88fF $ **FLOATING
C10397 S.t1131 VSUBS 0.02fF
C10398 S.n9448 VSUBS 0.24fF $ **FLOATING
C10399 S.n9449 VSUBS 0.36fF $ **FLOATING
C10400 S.n9450 VSUBS 0.61fF $ **FLOATING
C10401 S.n9451 VSUBS 0.12fF $ **FLOATING
C10402 S.t311 VSUBS 0.02fF
C10403 S.n9452 VSUBS 0.14fF $ **FLOATING
C10404 S.n9454 VSUBS 1.16fF $ **FLOATING
C10405 S.n9455 VSUBS 0.22fF $ **FLOATING
C10406 S.n9456 VSUBS 0.25fF $ **FLOATING
C10407 S.n9457 VSUBS 0.09fF $ **FLOATING
C10408 S.n9458 VSUBS 1.88fF $ **FLOATING
C10409 S.t1403 VSUBS 0.02fF
C10410 S.n9459 VSUBS 0.24fF $ **FLOATING
C10411 S.n9460 VSUBS 0.91fF $ **FLOATING
C10412 S.n9461 VSUBS 0.05fF $ **FLOATING
C10413 S.t1182 VSUBS 0.02fF
C10414 S.n9462 VSUBS 0.12fF $ **FLOATING
C10415 S.n9463 VSUBS 0.14fF $ **FLOATING
C10416 S.n9465 VSUBS 20.78fF $ **FLOATING
C10417 S.n9466 VSUBS 1.88fF $ **FLOATING
C10418 S.n9467 VSUBS 2.67fF $ **FLOATING
C10419 S.t2417 VSUBS 0.02fF
C10420 S.n9468 VSUBS 0.24fF $ **FLOATING
C10421 S.n9469 VSUBS 0.36fF $ **FLOATING
C10422 S.n9470 VSUBS 0.61fF $ **FLOATING
C10423 S.n9471 VSUBS 0.12fF $ **FLOATING
C10424 S.t1600 VSUBS 0.02fF
C10425 S.n9472 VSUBS 0.14fF $ **FLOATING
C10426 S.n9474 VSUBS 2.80fF $ **FLOATING
C10427 S.n9475 VSUBS 2.30fF $ **FLOATING
C10428 S.t1143 VSUBS 0.02fF
C10429 S.n9476 VSUBS 0.12fF $ **FLOATING
C10430 S.n9477 VSUBS 0.14fF $ **FLOATING
C10431 S.t192 VSUBS 0.02fF
C10432 S.n9479 VSUBS 0.24fF $ **FLOATING
C10433 S.n9480 VSUBS 0.91fF $ **FLOATING
C10434 S.n9481 VSUBS 0.05fF $ **FLOATING
C10435 S.n9482 VSUBS 2.80fF $ **FLOATING
C10436 S.n9483 VSUBS 1.88fF $ **FLOATING
C10437 S.n9484 VSUBS 0.12fF $ **FLOATING
C10438 S.t2388 VSUBS 0.02fF
C10439 S.n9485 VSUBS 0.14fF $ **FLOATING
C10440 S.t680 VSUBS 0.02fF
C10441 S.n9487 VSUBS 0.24fF $ **FLOATING
C10442 S.n9488 VSUBS 0.36fF $ **FLOATING
C10443 S.n9489 VSUBS 0.61fF $ **FLOATING
C10444 S.n9490 VSUBS 2.67fF $ **FLOATING
C10445 S.n9491 VSUBS 2.30fF $ **FLOATING
C10446 S.t729 VSUBS 0.02fF
C10447 S.n9492 VSUBS 0.12fF $ **FLOATING
C10448 S.n9493 VSUBS 0.14fF $ **FLOATING
C10449 S.t979 VSUBS 0.02fF
C10450 S.n9495 VSUBS 0.24fF $ **FLOATING
C10451 S.n9496 VSUBS 0.91fF $ **FLOATING
C10452 S.n9497 VSUBS 0.05fF $ **FLOATING
C10453 S.n9498 VSUBS 1.88fF $ **FLOATING
C10454 S.n9499 VSUBS 2.67fF $ **FLOATING
C10455 S.t1471 VSUBS 0.02fF
C10456 S.n9500 VSUBS 0.24fF $ **FLOATING
C10457 S.n9501 VSUBS 0.36fF $ **FLOATING
C10458 S.n9502 VSUBS 0.61fF $ **FLOATING
C10459 S.n9503 VSUBS 0.12fF $ **FLOATING
C10460 S.t653 VSUBS 0.02fF
C10461 S.n9504 VSUBS 0.14fF $ **FLOATING
C10462 S.n9506 VSUBS 2.80fF $ **FLOATING
C10463 S.n9507 VSUBS 2.30fF $ **FLOATING
C10464 S.t1520 VSUBS 0.02fF
C10465 S.n9508 VSUBS 0.12fF $ **FLOATING
C10466 S.n9509 VSUBS 0.14fF $ **FLOATING
C10467 S.t1763 VSUBS 0.02fF
C10468 S.n9511 VSUBS 0.24fF $ **FLOATING
C10469 S.n9512 VSUBS 0.91fF $ **FLOATING
C10470 S.n9513 VSUBS 0.05fF $ **FLOATING
C10471 S.n9514 VSUBS 1.88fF $ **FLOATING
C10472 S.n9515 VSUBS 2.67fF $ **FLOATING
C10473 S.t2260 VSUBS 0.02fF
C10474 S.n9516 VSUBS 0.24fF $ **FLOATING
C10475 S.n9517 VSUBS 0.36fF $ **FLOATING
C10476 S.n9518 VSUBS 0.61fF $ **FLOATING
C10477 S.n9519 VSUBS 0.12fF $ **FLOATING
C10478 S.t1443 VSUBS 0.02fF
C10479 S.n9520 VSUBS 0.14fF $ **FLOATING
C10480 S.n9522 VSUBS 2.80fF $ **FLOATING
C10481 S.n9523 VSUBS 2.30fF $ **FLOATING
C10482 S.t2311 VSUBS 0.02fF
C10483 S.n9524 VSUBS 0.12fF $ **FLOATING
C10484 S.n9525 VSUBS 0.14fF $ **FLOATING
C10485 S.t2543 VSUBS 0.02fF
C10486 S.n9527 VSUBS 0.24fF $ **FLOATING
C10487 S.n9528 VSUBS 0.91fF $ **FLOATING
C10488 S.n9529 VSUBS 0.05fF $ **FLOATING
C10489 S.n9530 VSUBS 1.88fF $ **FLOATING
C10490 S.n9531 VSUBS 2.67fF $ **FLOATING
C10491 S.t529 VSUBS 0.02fF
C10492 S.n9532 VSUBS 0.24fF $ **FLOATING
C10493 S.n9533 VSUBS 0.36fF $ **FLOATING
C10494 S.n9534 VSUBS 0.61fF $ **FLOATING
C10495 S.n9535 VSUBS 0.12fF $ **FLOATING
C10496 S.t2354 VSUBS 0.02fF
C10497 S.n9536 VSUBS 0.14fF $ **FLOATING
C10498 S.n9538 VSUBS 2.80fF $ **FLOATING
C10499 S.n9539 VSUBS 2.30fF $ **FLOATING
C10500 S.t579 VSUBS 0.02fF
C10501 S.n9540 VSUBS 0.12fF $ **FLOATING
C10502 S.n9541 VSUBS 0.14fF $ **FLOATING
C10503 S.t810 VSUBS 0.02fF
C10504 S.n9543 VSUBS 0.24fF $ **FLOATING
C10505 S.n9544 VSUBS 0.91fF $ **FLOATING
C10506 S.n9545 VSUBS 0.05fF $ **FLOATING
C10507 S.n9546 VSUBS 1.88fF $ **FLOATING
C10508 S.n9547 VSUBS 2.67fF $ **FLOATING
C10509 S.t2269 VSUBS 0.02fF
C10510 S.n9548 VSUBS 0.24fF $ **FLOATING
C10511 S.n9549 VSUBS 0.36fF $ **FLOATING
C10512 S.n9550 VSUBS 0.61fF $ **FLOATING
C10513 S.n9551 VSUBS 0.12fF $ **FLOATING
C10514 S.t2468 VSUBS 0.02fF
C10515 S.n9552 VSUBS 0.14fF $ **FLOATING
C10516 S.n9554 VSUBS 2.80fF $ **FLOATING
C10517 S.n9555 VSUBS 2.30fF $ **FLOATING
C10518 S.t814 VSUBS 0.02fF
C10519 S.n9556 VSUBS 0.12fF $ **FLOATING
C10520 S.n9557 VSUBS 0.14fF $ **FLOATING
C10521 S.t588 VSUBS 0.02fF
C10522 S.n9559 VSUBS 0.24fF $ **FLOATING
C10523 S.n9560 VSUBS 0.91fF $ **FLOATING
C10524 S.n9561 VSUBS 0.05fF $ **FLOATING
C10525 S.n9562 VSUBS 1.88fF $ **FLOATING
C10526 S.n9563 VSUBS 2.67fF $ **FLOATING
C10527 S.t541 VSUBS 0.02fF
C10528 S.n9564 VSUBS 0.24fF $ **FLOATING
C10529 S.n9565 VSUBS 0.36fF $ **FLOATING
C10530 S.n9566 VSUBS 0.61fF $ **FLOATING
C10531 S.n9567 VSUBS 0.12fF $ **FLOATING
C10532 S.t726 VSUBS 0.02fF
C10533 S.n9568 VSUBS 0.14fF $ **FLOATING
C10534 S.n9570 VSUBS 2.80fF $ **FLOATING
C10535 S.n9571 VSUBS 2.30fF $ **FLOATING
C10536 S.t1595 VSUBS 0.02fF
C10537 S.n9572 VSUBS 0.12fF $ **FLOATING
C10538 S.n9573 VSUBS 0.14fF $ **FLOATING
C10539 S.t1381 VSUBS 0.02fF
C10540 S.n9575 VSUBS 0.24fF $ **FLOATING
C10541 S.n9576 VSUBS 0.91fF $ **FLOATING
C10542 S.n9577 VSUBS 0.05fF $ **FLOATING
C10543 S.n9578 VSUBS 1.88fF $ **FLOATING
C10544 S.n9579 VSUBS 2.67fF $ **FLOATING
C10545 S.t1327 VSUBS 0.02fF
C10546 S.n9580 VSUBS 0.24fF $ **FLOATING
C10547 S.n9581 VSUBS 0.36fF $ **FLOATING
C10548 S.n9582 VSUBS 0.61fF $ **FLOATING
C10549 S.n9583 VSUBS 0.12fF $ **FLOATING
C10550 S.t1517 VSUBS 0.02fF
C10551 S.n9584 VSUBS 0.14fF $ **FLOATING
C10552 S.n9586 VSUBS 2.80fF $ **FLOATING
C10553 S.n9587 VSUBS 2.30fF $ **FLOATING
C10554 S.t2386 VSUBS 0.02fF
C10555 S.n9588 VSUBS 0.12fF $ **FLOATING
C10556 S.n9589 VSUBS 0.14fF $ **FLOATING
C10557 S.t2167 VSUBS 0.02fF
C10558 S.n9591 VSUBS 0.24fF $ **FLOATING
C10559 S.n9592 VSUBS 0.91fF $ **FLOATING
C10560 S.n9593 VSUBS 0.05fF $ **FLOATING
C10561 S.n9594 VSUBS 2.73fF $ **FLOATING
C10562 S.n9595 VSUBS 1.59fF $ **FLOATING
C10563 S.n9596 VSUBS 0.12fF $ **FLOATING
C10564 S.t2010 VSUBS 0.02fF
C10565 S.n9597 VSUBS 0.14fF $ **FLOATING
C10566 S.t499 VSUBS 0.02fF
C10567 S.n9599 VSUBS 0.24fF $ **FLOATING
C10568 S.n9600 VSUBS 0.36fF $ **FLOATING
C10569 S.n9601 VSUBS 0.61fF $ **FLOATING
C10570 S.n9602 VSUBS 0.07fF $ **FLOATING
C10571 S.n9603 VSUBS 0.01fF $ **FLOATING
C10572 S.n9604 VSUBS 0.24fF $ **FLOATING
C10573 S.n9605 VSUBS 1.16fF $ **FLOATING
C10574 S.n9606 VSUBS 1.35fF $ **FLOATING
C10575 S.n9607 VSUBS 2.30fF $ **FLOATING
C10576 S.t1437 VSUBS 0.02fF
C10577 S.n9608 VSUBS 0.12fF $ **FLOATING
C10578 S.n9609 VSUBS 0.14fF $ **FLOATING
C10579 S.t1900 VSUBS 0.02fF
C10580 S.n9611 VSUBS 0.24fF $ **FLOATING
C10581 S.n9612 VSUBS 0.91fF $ **FLOATING
C10582 S.n9613 VSUBS 0.05fF $ **FLOATING
C10583 S.t225 VSUBS 48.27fF
C10584 S.t434 VSUBS 0.02fF
C10585 S.n9614 VSUBS 0.24fF $ **FLOATING
C10586 S.n9615 VSUBS 0.91fF $ **FLOATING
C10587 S.n9616 VSUBS 0.05fF $ **FLOATING
C10588 S.t649 VSUBS 0.02fF
C10589 S.n9617 VSUBS 0.12fF $ **FLOATING
C10590 S.n9618 VSUBS 0.14fF $ **FLOATING
C10591 S.n9620 VSUBS 0.12fF $ **FLOATING
C10592 S.t2305 VSUBS 0.02fF
C10593 S.n9621 VSUBS 0.14fF $ **FLOATING
C10594 S.n9623 VSUBS 5.17fF $ **FLOATING
C10595 S.n9624 VSUBS 5.44fF $ **FLOATING
C10596 S.t626 VSUBS 0.02fF
C10597 S.n9625 VSUBS 0.12fF $ **FLOATING
C10598 S.n9626 VSUBS 0.14fF $ **FLOATING
C10599 S.t410 VSUBS 0.02fF
C10600 S.n9628 VSUBS 0.24fF $ **FLOATING
C10601 S.n9629 VSUBS 0.91fF $ **FLOATING
C10602 S.n9630 VSUBS 0.05fF $ **FLOATING
C10603 S.t31 VSUBS 47.89fF
C10604 S.t846 VSUBS 0.02fF
C10605 S.n9631 VSUBS 0.01fF $ **FLOATING
C10606 S.n9632 VSUBS 0.26fF $ **FLOATING
C10607 S.t1345 VSUBS 0.02fF
C10608 S.n9634 VSUBS 1.19fF $ **FLOATING
C10609 S.n9635 VSUBS 0.05fF $ **FLOATING
C10610 S.t1061 VSUBS 0.02fF
C10611 S.n9636 VSUBS 0.64fF $ **FLOATING
C10612 S.n9637 VSUBS 0.61fF $ **FLOATING
C10613 S.n9638 VSUBS 8.97fF $ **FLOATING
C10614 S.n9639 VSUBS 8.97fF $ **FLOATING
C10615 S.n9640 VSUBS 0.60fF $ **FLOATING
C10616 S.n9641 VSUBS 0.22fF $ **FLOATING
C10617 S.n9642 VSUBS 0.59fF $ **FLOATING
C10618 S.n9643 VSUBS 3.39fF $ **FLOATING
C10619 S.n9644 VSUBS 0.29fF $ **FLOATING
C10620 S.t55 VSUBS 21.42fF
C10621 S.n9645 VSUBS 21.71fF $ **FLOATING
C10622 S.n9646 VSUBS 0.77fF $ **FLOATING
C10623 S.n9647 VSUBS 0.28fF $ **FLOATING
C10624 S.n9648 VSUBS 4.00fF $ **FLOATING
C10625 S.n9649 VSUBS 1.35fF $ **FLOATING
C10626 S.n9650 VSUBS 0.01fF $ **FLOATING
C10627 S.n9651 VSUBS 0.02fF $ **FLOATING
C10628 S.n9652 VSUBS 0.03fF $ **FLOATING
C10629 S.n9653 VSUBS 0.04fF $ **FLOATING
C10630 S.n9654 VSUBS 0.17fF $ **FLOATING
C10631 S.n9655 VSUBS 0.01fF $ **FLOATING
C10632 S.n9656 VSUBS 0.02fF $ **FLOATING
C10633 S.n9657 VSUBS 0.01fF $ **FLOATING
C10634 S.n9658 VSUBS 0.01fF $ **FLOATING
C10635 S.n9659 VSUBS 0.01fF $ **FLOATING
C10636 S.n9660 VSUBS 0.01fF $ **FLOATING
C10637 S.n9661 VSUBS 0.02fF $ **FLOATING
C10638 S.n9662 VSUBS 0.01fF $ **FLOATING
C10639 S.n9663 VSUBS 0.02fF $ **FLOATING
C10640 S.n9664 VSUBS 0.05fF $ **FLOATING
C10641 S.n9665 VSUBS 0.04fF $ **FLOATING
C10642 S.n9666 VSUBS 0.11fF $ **FLOATING
C10643 S.n9667 VSUBS 0.38fF $ **FLOATING
C10644 S.n9668 VSUBS 0.20fF $ **FLOATING
C10645 S.n9669 VSUBS 4.39fF $ **FLOATING
C10646 S.n9670 VSUBS 0.24fF $ **FLOATING
C10647 S.n9671 VSUBS 1.50fF $ **FLOATING
C10648 S.n9672 VSUBS 1.31fF $ **FLOATING
C10649 S.n9673 VSUBS 0.28fF $ **FLOATING
C10650 S.n9674 VSUBS 1.89fF $ **FLOATING
C10651 S.n9675 VSUBS 0.07fF $ **FLOATING
C10652 S.n9676 VSUBS 0.04fF $ **FLOATING
C10653 S.n9677 VSUBS 0.05fF $ **FLOATING
C10654 S.n9678 VSUBS 0.87fF $ **FLOATING
C10655 S.n9679 VSUBS 0.01fF $ **FLOATING
C10656 S.n9680 VSUBS 0.01fF $ **FLOATING
C10657 S.n9681 VSUBS 0.01fF $ **FLOATING
C10658 S.n9682 VSUBS 0.07fF $ **FLOATING
C10659 S.n9683 VSUBS 0.68fF $ **FLOATING
C10660 S.n9684 VSUBS 0.72fF $ **FLOATING
C10661 S.t593 VSUBS 0.02fF
C10662 S.n9685 VSUBS 0.24fF $ **FLOATING
C10663 S.n9686 VSUBS 0.36fF $ **FLOATING
C10664 S.n9687 VSUBS 0.61fF $ **FLOATING
C10665 S.n9688 VSUBS 0.12fF $ **FLOATING
C10666 S.t2099 VSUBS 0.02fF
C10667 S.n9689 VSUBS 0.14fF $ **FLOATING
C10668 S.n9691 VSUBS 0.70fF $ **FLOATING
C10669 S.n9692 VSUBS 0.23fF $ **FLOATING
C10670 S.n9693 VSUBS 0.23fF $ **FLOATING
C10671 S.n9694 VSUBS 0.70fF $ **FLOATING
C10672 S.n9695 VSUBS 1.16fF $ **FLOATING
C10673 S.n9696 VSUBS 0.22fF $ **FLOATING
C10674 S.n9697 VSUBS 0.25fF $ **FLOATING
C10675 S.n9698 VSUBS 0.09fF $ **FLOATING
C10676 S.n9699 VSUBS 2.31fF $ **FLOATING
C10677 S.t667 VSUBS 0.02fF
C10678 S.n9700 VSUBS 0.24fF $ **FLOATING
C10679 S.n9701 VSUBS 0.91fF $ **FLOATING
C10680 S.n9702 VSUBS 0.05fF $ **FLOATING
C10681 S.t446 VSUBS 0.02fF
C10682 S.n9703 VSUBS 0.12fF $ **FLOATING
C10683 S.n9704 VSUBS 0.14fF $ **FLOATING
C10684 S.n9706 VSUBS 1.88fF $ **FLOATING
C10685 S.n9707 VSUBS 0.46fF $ **FLOATING
C10686 S.n9708 VSUBS 0.22fF $ **FLOATING
C10687 S.n9709 VSUBS 0.38fF $ **FLOATING
C10688 S.n9710 VSUBS 0.16fF $ **FLOATING
C10689 S.n9711 VSUBS 0.28fF $ **FLOATING
C10690 S.n9712 VSUBS 0.21fF $ **FLOATING
C10691 S.n9713 VSUBS 0.30fF $ **FLOATING
C10692 S.n9714 VSUBS 0.42fF $ **FLOATING
C10693 S.n9715 VSUBS 0.21fF $ **FLOATING
C10694 S.t1506 VSUBS 0.02fF
C10695 S.n9716 VSUBS 0.24fF $ **FLOATING
C10696 S.n9717 VSUBS 0.36fF $ **FLOATING
C10697 S.n9718 VSUBS 0.61fF $ **FLOATING
C10698 S.n9719 VSUBS 0.12fF $ **FLOATING
C10699 S.t488 VSUBS 0.02fF
C10700 S.n9720 VSUBS 0.14fF $ **FLOATING
C10701 S.n9722 VSUBS 0.04fF $ **FLOATING
C10702 S.n9723 VSUBS 0.03fF $ **FLOATING
C10703 S.n9724 VSUBS 0.03fF $ **FLOATING
C10704 S.n9725 VSUBS 0.10fF $ **FLOATING
C10705 S.n9726 VSUBS 0.36fF $ **FLOATING
C10706 S.n9727 VSUBS 0.38fF $ **FLOATING
C10707 S.n9728 VSUBS 0.11fF $ **FLOATING
C10708 S.n9729 VSUBS 0.12fF $ **FLOATING
C10709 S.n9730 VSUBS 0.07fF $ **FLOATING
C10710 S.n9731 VSUBS 0.12fF $ **FLOATING
C10711 S.n9732 VSUBS 0.18fF $ **FLOATING
C10712 S.n9733 VSUBS 3.99fF $ **FLOATING
C10713 S.t1574 VSUBS 0.02fF
C10714 S.n9734 VSUBS 0.24fF $ **FLOATING
C10715 S.n9735 VSUBS 0.91fF $ **FLOATING
C10716 S.n9736 VSUBS 0.05fF $ **FLOATING
C10717 S.t1356 VSUBS 0.02fF
C10718 S.n9737 VSUBS 0.12fF $ **FLOATING
C10719 S.n9738 VSUBS 0.14fF $ **FLOATING
C10720 S.n9740 VSUBS 0.25fF $ **FLOATING
C10721 S.n9741 VSUBS 0.09fF $ **FLOATING
C10722 S.n9742 VSUBS 0.21fF $ **FLOATING
C10723 S.n9743 VSUBS 1.28fF $ **FLOATING
C10724 S.n9744 VSUBS 0.53fF $ **FLOATING
C10725 S.n9745 VSUBS 1.88fF $ **FLOATING
C10726 S.n9746 VSUBS 0.12fF $ **FLOATING
C10727 S.t62 VSUBS 0.02fF
C10728 S.n9747 VSUBS 0.14fF $ **FLOATING
C10729 S.t1136 VSUBS 0.02fF
C10730 S.n9749 VSUBS 0.24fF $ **FLOATING
C10731 S.n9750 VSUBS 0.36fF $ **FLOATING
C10732 S.n9751 VSUBS 0.61fF $ **FLOATING
C10733 S.n9752 VSUBS 1.58fF $ **FLOATING
C10734 S.n9753 VSUBS 2.45fF $ **FLOATING
C10735 S.t1213 VSUBS 0.02fF
C10736 S.n9754 VSUBS 0.24fF $ **FLOATING
C10737 S.n9755 VSUBS 0.91fF $ **FLOATING
C10738 S.n9756 VSUBS 0.05fF $ **FLOATING
C10739 S.t2141 VSUBS 0.02fF
C10740 S.n9757 VSUBS 0.12fF $ **FLOATING
C10741 S.n9758 VSUBS 0.14fF $ **FLOATING
C10742 S.n9760 VSUBS 1.89fF $ **FLOATING
C10743 S.n9761 VSUBS 0.06fF $ **FLOATING
C10744 S.n9762 VSUBS 0.03fF $ **FLOATING
C10745 S.n9763 VSUBS 0.04fF $ **FLOATING
C10746 S.n9764 VSUBS 0.99fF $ **FLOATING
C10747 S.n9765 VSUBS 0.02fF $ **FLOATING
C10748 S.n9766 VSUBS 0.01fF $ **FLOATING
C10749 S.n9767 VSUBS 0.02fF $ **FLOATING
C10750 S.n9768 VSUBS 0.08fF $ **FLOATING
C10751 S.n9769 VSUBS 0.36fF $ **FLOATING
C10752 S.n9770 VSUBS 1.85fF $ **FLOATING
C10753 S.t1918 VSUBS 0.02fF
C10754 S.n9771 VSUBS 0.24fF $ **FLOATING
C10755 S.n9772 VSUBS 0.36fF $ **FLOATING
C10756 S.n9773 VSUBS 0.61fF $ **FLOATING
C10757 S.n9774 VSUBS 0.12fF $ **FLOATING
C10758 S.t880 VSUBS 0.02fF
C10759 S.n9775 VSUBS 0.14fF $ **FLOATING
C10760 S.n9777 VSUBS 0.70fF $ **FLOATING
C10761 S.n9778 VSUBS 0.23fF $ **FLOATING
C10762 S.n9779 VSUBS 0.23fF $ **FLOATING
C10763 S.n9780 VSUBS 0.70fF $ **FLOATING
C10764 S.n9781 VSUBS 1.16fF $ **FLOATING
C10765 S.n9782 VSUBS 0.22fF $ **FLOATING
C10766 S.n9783 VSUBS 0.25fF $ **FLOATING
C10767 S.n9784 VSUBS 0.09fF $ **FLOATING
C10768 S.n9785 VSUBS 1.88fF $ **FLOATING
C10769 S.t1991 VSUBS 0.02fF
C10770 S.n9786 VSUBS 0.24fF $ **FLOATING
C10771 S.n9787 VSUBS 0.91fF $ **FLOATING
C10772 S.n9788 VSUBS 0.05fF $ **FLOATING
C10773 S.t1747 VSUBS 0.02fF
C10774 S.n9789 VSUBS 0.12fF $ **FLOATING
C10775 S.n9790 VSUBS 0.14fF $ **FLOATING
C10776 S.n9792 VSUBS 20.78fF $ **FLOATING
C10777 S.n9793 VSUBS 0.06fF $ **FLOATING
C10778 S.n9794 VSUBS 0.20fF $ **FLOATING
C10779 S.n9795 VSUBS 0.09fF $ **FLOATING
C10780 S.n9796 VSUBS 0.21fF $ **FLOATING
C10781 S.n9797 VSUBS 0.10fF $ **FLOATING
C10782 S.n9798 VSUBS 0.30fF $ **FLOATING
C10783 S.n9799 VSUBS 0.69fF $ **FLOATING
C10784 S.n9800 VSUBS 0.45fF $ **FLOATING
C10785 S.n9801 VSUBS 2.33fF $ **FLOATING
C10786 S.n9802 VSUBS 0.12fF $ **FLOATING
C10787 S.t1312 VSUBS 0.02fF
C10788 S.n9803 VSUBS 0.14fF $ **FLOATING
C10789 S.t2329 VSUBS 0.02fF
C10790 S.n9805 VSUBS 0.24fF $ **FLOATING
C10791 S.n9806 VSUBS 0.36fF $ **FLOATING
C10792 S.n9807 VSUBS 0.61fF $ **FLOATING
C10793 S.n9808 VSUBS 1.90fF $ **FLOATING
C10794 S.n9809 VSUBS 0.17fF $ **FLOATING
C10795 S.n9810 VSUBS 0.76fF $ **FLOATING
C10796 S.n9811 VSUBS 0.32fF $ **FLOATING
C10797 S.n9812 VSUBS 0.25fF $ **FLOATING
C10798 S.n9813 VSUBS 0.30fF $ **FLOATING
C10799 S.n9814 VSUBS 0.47fF $ **FLOATING
C10800 S.n9815 VSUBS 0.16fF $ **FLOATING
C10801 S.n9816 VSUBS 1.93fF $ **FLOATING
C10802 S.t2180 VSUBS 0.02fF
C10803 S.n9817 VSUBS 0.12fF $ **FLOATING
C10804 S.n9818 VSUBS 0.14fF $ **FLOATING
C10805 S.t2406 VSUBS 0.02fF
C10806 S.n9820 VSUBS 0.24fF $ **FLOATING
C10807 S.n9821 VSUBS 0.91fF $ **FLOATING
C10808 S.n9822 VSUBS 0.05fF $ **FLOATING
C10809 S.n9823 VSUBS 1.88fF $ **FLOATING
C10810 S.n9824 VSUBS 0.12fF $ **FLOATING
C10811 S.t2456 VSUBS 0.02fF
C10812 S.n9825 VSUBS 0.14fF $ **FLOATING
C10813 S.t801 VSUBS 0.02fF
C10814 S.n9827 VSUBS 0.12fF $ **FLOATING
C10815 S.n9828 VSUBS 0.14fF $ **FLOATING
C10816 S.t1047 VSUBS 0.02fF
C10817 S.n9830 VSUBS 0.24fF $ **FLOATING
C10818 S.n9831 VSUBS 0.91fF $ **FLOATING
C10819 S.n9832 VSUBS 0.05fF $ **FLOATING
C10820 S.t742 VSUBS 0.02fF
C10821 S.n9833 VSUBS 0.24fF $ **FLOATING
C10822 S.n9834 VSUBS 0.36fF $ **FLOATING
C10823 S.n9835 VSUBS 0.61fF $ **FLOATING
C10824 S.n9836 VSUBS 0.32fF $ **FLOATING
C10825 S.n9837 VSUBS 1.09fF $ **FLOATING
C10826 S.n9838 VSUBS 0.15fF $ **FLOATING
C10827 S.n9839 VSUBS 2.10fF $ **FLOATING
C10828 S.n9840 VSUBS 2.94fF $ **FLOATING
C10829 S.n9841 VSUBS 1.88fF $ **FLOATING
C10830 S.n9842 VSUBS 0.12fF $ **FLOATING
C10831 S.t1661 VSUBS 0.02fF
C10832 S.n9843 VSUBS 0.14fF $ **FLOATING
C10833 S.t171 VSUBS 0.02fF
C10834 S.n9845 VSUBS 0.24fF $ **FLOATING
C10835 S.n9846 VSUBS 0.36fF $ **FLOATING
C10836 S.n9847 VSUBS 0.61fF $ **FLOATING
C10837 S.n9848 VSUBS 0.92fF $ **FLOATING
C10838 S.n9849 VSUBS 0.32fF $ **FLOATING
C10839 S.n9850 VSUBS 0.92fF $ **FLOATING
C10840 S.n9851 VSUBS 1.09fF $ **FLOATING
C10841 S.n9852 VSUBS 0.15fF $ **FLOATING
C10842 S.n9853 VSUBS 4.96fF $ **FLOATING
C10843 S.t2530 VSUBS 0.02fF
C10844 S.n9854 VSUBS 0.12fF $ **FLOATING
C10845 S.n9855 VSUBS 0.14fF $ **FLOATING
C10846 S.t262 VSUBS 0.02fF
C10847 S.n9857 VSUBS 0.24fF $ **FLOATING
C10848 S.n9858 VSUBS 0.91fF $ **FLOATING
C10849 S.n9859 VSUBS 0.05fF $ **FLOATING
C10850 S.n9860 VSUBS 1.88fF $ **FLOATING
C10851 S.n9861 VSUBS 2.67fF $ **FLOATING
C10852 S.t959 VSUBS 0.02fF
C10853 S.n9862 VSUBS 0.24fF $ **FLOATING
C10854 S.n9863 VSUBS 0.36fF $ **FLOATING
C10855 S.n9864 VSUBS 0.61fF $ **FLOATING
C10856 S.n9865 VSUBS 0.12fF $ **FLOATING
C10857 S.t2448 VSUBS 0.02fF
C10858 S.n9866 VSUBS 0.14fF $ **FLOATING
C10859 S.n9868 VSUBS 1.88fF $ **FLOATING
C10860 S.n9869 VSUBS 2.67fF $ **FLOATING
C10861 S.t1533 VSUBS 0.02fF
C10862 S.n9870 VSUBS 0.24fF $ **FLOATING
C10863 S.n9871 VSUBS 0.36fF $ **FLOATING
C10864 S.n9872 VSUBS 0.61fF $ **FLOATING
C10865 S.t1827 VSUBS 0.02fF
C10866 S.n9873 VSUBS 0.24fF $ **FLOATING
C10867 S.n9874 VSUBS 0.91fF $ **FLOATING
C10868 S.n9875 VSUBS 0.05fF $ **FLOATING
C10869 S.t1581 VSUBS 0.02fF
C10870 S.n9876 VSUBS 0.12fF $ **FLOATING
C10871 S.n9877 VSUBS 0.14fF $ **FLOATING
C10872 S.n9879 VSUBS 0.12fF $ **FLOATING
C10873 S.t713 VSUBS 0.02fF
C10874 S.n9880 VSUBS 0.14fF $ **FLOATING
C10875 S.n9882 VSUBS 2.30fF $ **FLOATING
C10876 S.n9883 VSUBS 2.94fF $ **FLOATING
C10877 S.n9884 VSUBS 5.16fF $ **FLOATING
C10878 S.t793 VSUBS 0.02fF
C10879 S.n9885 VSUBS 0.12fF $ **FLOATING
C10880 S.n9886 VSUBS 0.14fF $ **FLOATING
C10881 S.t1045 VSUBS 0.02fF
C10882 S.n9888 VSUBS 0.24fF $ **FLOATING
C10883 S.n9889 VSUBS 0.91fF $ **FLOATING
C10884 S.n9890 VSUBS 0.05fF $ **FLOATING
C10885 S.n9891 VSUBS 1.88fF $ **FLOATING
C10886 S.n9892 VSUBS 2.67fF $ **FLOATING
C10887 S.t1873 VSUBS 0.02fF
C10888 S.n9893 VSUBS 0.24fF $ **FLOATING
C10889 S.n9894 VSUBS 0.36fF $ **FLOATING
C10890 S.n9895 VSUBS 0.61fF $ **FLOATING
C10891 S.n9896 VSUBS 0.12fF $ **FLOATING
C10892 S.t840 VSUBS 0.02fF
C10893 S.n9897 VSUBS 0.14fF $ **FLOATING
C10894 S.n9899 VSUBS 5.17fF $ **FLOATING
C10895 S.t1708 VSUBS 0.02fF
C10896 S.n9900 VSUBS 0.12fF $ **FLOATING
C10897 S.n9901 VSUBS 0.14fF $ **FLOATING
C10898 S.t1954 VSUBS 0.02fF
C10899 S.n9903 VSUBS 0.24fF $ **FLOATING
C10900 S.n9904 VSUBS 0.91fF $ **FLOATING
C10901 S.n9905 VSUBS 0.05fF $ **FLOATING
C10902 S.n9906 VSUBS 1.88fF $ **FLOATING
C10903 S.n9907 VSUBS 0.12fF $ **FLOATING
C10904 S.t462 VSUBS 0.02fF
C10905 S.n9908 VSUBS 0.14fF $ **FLOATING
C10906 S.t1478 VSUBS 0.02fF
C10907 S.n9910 VSUBS 0.24fF $ **FLOATING
C10908 S.n9911 VSUBS 0.36fF $ **FLOATING
C10909 S.n9912 VSUBS 0.61fF $ **FLOATING
C10910 S.n9913 VSUBS 2.67fF $ **FLOATING
C10911 S.n9914 VSUBS 5.17fF $ **FLOATING
C10912 S.t1328 VSUBS 0.02fF
C10913 S.n9915 VSUBS 0.12fF $ **FLOATING
C10914 S.n9916 VSUBS 0.14fF $ **FLOATING
C10915 S.t1550 VSUBS 0.02fF
C10916 S.n9918 VSUBS 0.24fF $ **FLOATING
C10917 S.n9919 VSUBS 0.91fF $ **FLOATING
C10918 S.n9920 VSUBS 0.05fF $ **FLOATING
C10919 S.n9921 VSUBS 1.88fF $ **FLOATING
C10920 S.n9922 VSUBS 2.67fF $ **FLOATING
C10921 S.t2262 VSUBS 0.02fF
C10922 S.n9923 VSUBS 0.24fF $ **FLOATING
C10923 S.n9924 VSUBS 0.36fF $ **FLOATING
C10924 S.n9925 VSUBS 0.61fF $ **FLOATING
C10925 S.n9926 VSUBS 0.12fF $ **FLOATING
C10926 S.t1247 VSUBS 0.02fF
C10927 S.n9927 VSUBS 0.14fF $ **FLOATING
C10928 S.n9929 VSUBS 5.17fF $ **FLOATING
C10929 S.t2114 VSUBS 0.02fF
C10930 S.n9930 VSUBS 0.12fF $ **FLOATING
C10931 S.n9931 VSUBS 0.14fF $ **FLOATING
C10932 S.t2338 VSUBS 0.02fF
C10933 S.n9933 VSUBS 0.24fF $ **FLOATING
C10934 S.n9934 VSUBS 0.91fF $ **FLOATING
C10935 S.n9935 VSUBS 0.05fF $ **FLOATING
C10936 S.n9936 VSUBS 1.88fF $ **FLOATING
C10937 S.n9937 VSUBS 2.67fF $ **FLOATING
C10938 S.t535 VSUBS 0.02fF
C10939 S.n9938 VSUBS 0.24fF $ **FLOATING
C10940 S.n9939 VSUBS 0.36fF $ **FLOATING
C10941 S.n9940 VSUBS 0.61fF $ **FLOATING
C10942 S.n9941 VSUBS 0.12fF $ **FLOATING
C10943 S.t2033 VSUBS 0.02fF
C10944 S.n9942 VSUBS 0.14fF $ **FLOATING
C10945 S.n9944 VSUBS 5.17fF $ **FLOATING
C10946 S.t382 VSUBS 0.02fF
C10947 S.n9945 VSUBS 0.12fF $ **FLOATING
C10948 S.n9946 VSUBS 0.14fF $ **FLOATING
C10949 S.t603 VSUBS 0.02fF
C10950 S.n9948 VSUBS 0.24fF $ **FLOATING
C10951 S.n9949 VSUBS 0.91fF $ **FLOATING
C10952 S.n9950 VSUBS 0.05fF $ **FLOATING
C10953 S.n9951 VSUBS 1.88fF $ **FLOATING
C10954 S.n9952 VSUBS 2.67fF $ **FLOATING
C10955 S.t1320 VSUBS 0.02fF
C10956 S.n9953 VSUBS 0.24fF $ **FLOATING
C10957 S.n9954 VSUBS 0.36fF $ **FLOATING
C10958 S.n9955 VSUBS 0.61fF $ **FLOATING
C10959 S.n9956 VSUBS 0.12fF $ **FLOATING
C10960 S.t303 VSUBS 0.02fF
C10961 S.n9957 VSUBS 0.14fF $ **FLOATING
C10962 S.n9959 VSUBS 5.17fF $ **FLOATING
C10963 S.t1170 VSUBS 0.02fF
C10964 S.n9960 VSUBS 0.12fF $ **FLOATING
C10965 S.n9961 VSUBS 0.14fF $ **FLOATING
C10966 S.t1395 VSUBS 0.02fF
C10967 S.n9963 VSUBS 0.24fF $ **FLOATING
C10968 S.n9964 VSUBS 0.91fF $ **FLOATING
C10969 S.n9965 VSUBS 0.05fF $ **FLOATING
C10970 S.n9966 VSUBS 1.88fF $ **FLOATING
C10971 S.n9967 VSUBS 2.67fF $ **FLOATING
C10972 S.t149 VSUBS 0.02fF
C10973 S.n9968 VSUBS 0.24fF $ **FLOATING
C10974 S.n9969 VSUBS 0.36fF $ **FLOATING
C10975 S.n9970 VSUBS 0.61fF $ **FLOATING
C10976 S.n9971 VSUBS 0.12fF $ **FLOATING
C10977 S.t2494 VSUBS 0.02fF
C10978 S.n9972 VSUBS 0.14fF $ **FLOATING
C10979 S.n9974 VSUBS 5.17fF $ **FLOATING
C10980 S.t2078 VSUBS 0.02fF
C10981 S.n9975 VSUBS 0.12fF $ **FLOATING
C10982 S.n9976 VSUBS 0.14fF $ **FLOATING
C10983 S.t617 VSUBS 0.02fF
C10984 S.n9978 VSUBS 0.24fF $ **FLOATING
C10985 S.n9979 VSUBS 0.91fF $ **FLOATING
C10986 S.n9980 VSUBS 0.05fF $ **FLOATING
C10987 S.n9981 VSUBS 1.88fF $ **FLOATING
C10988 S.n9982 VSUBS 2.67fF $ **FLOATING
C10989 S.t942 VSUBS 0.02fF
C10990 S.n9983 VSUBS 0.24fF $ **FLOATING
C10991 S.n9984 VSUBS 0.36fF $ **FLOATING
C10992 S.n9985 VSUBS 0.61fF $ **FLOATING
C10993 S.n9986 VSUBS 0.12fF $ **FLOATING
C10994 S.t750 VSUBS 0.02fF
C10995 S.n9987 VSUBS 0.14fF $ **FLOATING
C10996 S.n9989 VSUBS 5.17fF $ **FLOATING
C10997 S.t1622 VSUBS 0.02fF
C10998 S.n9990 VSUBS 0.12fF $ **FLOATING
C10999 S.n9991 VSUBS 0.14fF $ **FLOATING
C11000 S.t1408 VSUBS 0.02fF
C11001 S.n9993 VSUBS 0.24fF $ **FLOATING
C11002 S.n9994 VSUBS 0.91fF $ **FLOATING
C11003 S.n9995 VSUBS 0.05fF $ **FLOATING
C11004 S.n9996 VSUBS 1.88fF $ **FLOATING
C11005 S.n9997 VSUBS 2.67fF $ **FLOATING
C11006 S.t1724 VSUBS 0.02fF
C11007 S.n9998 VSUBS 0.24fF $ **FLOATING
C11008 S.n9999 VSUBS 0.36fF $ **FLOATING
C11009 S.n10000 VSUBS 0.61fF $ **FLOATING
C11010 S.n10001 VSUBS 0.12fF $ **FLOATING
C11011 S.t1544 VSUBS 0.02fF
C11012 S.n10002 VSUBS 0.14fF $ **FLOATING
C11013 S.n10004 VSUBS 5.17fF $ **FLOATING
C11014 S.t2409 VSUBS 0.02fF
C11015 S.n10005 VSUBS 0.12fF $ **FLOATING
C11016 S.n10006 VSUBS 0.14fF $ **FLOATING
C11017 S.t2196 VSUBS 0.02fF
C11018 S.n10008 VSUBS 0.24fF $ **FLOATING
C11019 S.n10009 VSUBS 0.91fF $ **FLOATING
C11020 S.n10010 VSUBS 0.05fF $ **FLOATING
C11021 S.n10011 VSUBS 1.88fF $ **FLOATING
C11022 S.n10012 VSUBS 2.67fF $ **FLOATING
C11023 S.t2512 VSUBS 0.02fF
C11024 S.n10013 VSUBS 0.24fF $ **FLOATING
C11025 S.n10014 VSUBS 0.36fF $ **FLOATING
C11026 S.n10015 VSUBS 0.61fF $ **FLOATING
C11027 S.n10016 VSUBS 0.12fF $ **FLOATING
C11028 S.t2331 VSUBS 0.02fF
C11029 S.n10017 VSUBS 0.14fF $ **FLOATING
C11030 S.n10019 VSUBS 4.89fF $ **FLOATING
C11031 S.t675 VSUBS 0.02fF
C11032 S.n10020 VSUBS 0.12fF $ **FLOATING
C11033 S.n10021 VSUBS 0.14fF $ **FLOATING
C11034 S.t461 VSUBS 0.02fF
C11035 S.n10023 VSUBS 0.24fF $ **FLOATING
C11036 S.n10024 VSUBS 0.91fF $ **FLOATING
C11037 S.n10025 VSUBS 0.05fF $ **FLOATING
C11038 S.n10026 VSUBS 1.88fF $ **FLOATING
C11039 S.n10027 VSUBS 2.67fF $ **FLOATING
C11040 S.t773 VSUBS 0.02fF
C11041 S.n10028 VSUBS 0.24fF $ **FLOATING
C11042 S.n10029 VSUBS 0.36fF $ **FLOATING
C11043 S.n10030 VSUBS 0.61fF $ **FLOATING
C11044 S.n10031 VSUBS 0.12fF $ **FLOATING
C11045 S.t595 VSUBS 0.02fF
C11046 S.n10032 VSUBS 0.14fF $ **FLOATING
C11047 S.n10034 VSUBS 1.88fF $ **FLOATING
C11048 S.n10035 VSUBS 2.68fF $ **FLOATING
C11049 S.t798 VSUBS 0.02fF
C11050 S.n10036 VSUBS 0.24fF $ **FLOATING
C11051 S.n10037 VSUBS 0.36fF $ **FLOATING
C11052 S.n10038 VSUBS 0.61fF $ **FLOATING
C11053 S.t401 VSUBS 0.02fF
C11054 S.n10039 VSUBS 1.22fF $ **FLOATING
C11055 S.n10040 VSUBS 0.36fF $ **FLOATING
C11056 S.n10041 VSUBS 1.22fF $ **FLOATING
C11057 S.n10042 VSUBS 0.61fF $ **FLOATING
C11058 S.n10043 VSUBS 0.35fF $ **FLOATING
C11059 S.n10044 VSUBS 0.63fF $ **FLOATING
C11060 S.n10045 VSUBS 1.15fF $ **FLOATING
C11061 S.n10046 VSUBS 3.00fF $ **FLOATING
C11062 S.n10047 VSUBS 0.59fF $ **FLOATING
C11063 S.n10048 VSUBS 0.01fF $ **FLOATING
C11064 S.n10049 VSUBS 0.97fF $ **FLOATING
C11065 S.t67 VSUBS 21.42fF
C11066 S.n10050 VSUBS 20.29fF $ **FLOATING
C11067 S.n10052 VSUBS 0.38fF $ **FLOATING
C11068 S.n10053 VSUBS 0.23fF $ **FLOATING
C11069 S.n10054 VSUBS 2.79fF $ **FLOATING
C11070 S.n10055 VSUBS 2.46fF $ **FLOATING
C11071 S.n10056 VSUBS 4.00fF $ **FLOATING
C11072 S.n10057 VSUBS 0.25fF $ **FLOATING
C11073 S.n10058 VSUBS 0.01fF $ **FLOATING
C11074 S.t2103 VSUBS 0.02fF
C11075 S.n10059 VSUBS 0.26fF $ **FLOATING
C11076 S.t672 VSUBS 0.02fF
C11077 S.n10060 VSUBS 0.95fF $ **FLOATING
C11078 S.n10061 VSUBS 0.71fF $ **FLOATING
C11079 S.n10062 VSUBS 1.89fF $ **FLOATING
C11080 S.n10063 VSUBS 1.73fF $ **FLOATING
C11081 S.t1193 VSUBS 0.02fF
C11082 S.n10064 VSUBS 0.24fF $ **FLOATING
C11083 S.n10065 VSUBS 0.36fF $ **FLOATING
C11084 S.n10066 VSUBS 0.61fF $ **FLOATING
C11085 S.n10067 VSUBS 0.12fF $ **FLOATING
C11086 S.t376 VSUBS 0.02fF
C11087 S.n10068 VSUBS 0.14fF $ **FLOATING
C11088 S.n10070 VSUBS 1.16fF $ **FLOATING
C11089 S.n10071 VSUBS 0.22fF $ **FLOATING
C11090 S.n10072 VSUBS 0.25fF $ **FLOATING
C11091 S.n10073 VSUBS 0.09fF $ **FLOATING
C11092 S.n10074 VSUBS 2.44fF $ **FLOATING
C11093 S.t1459 VSUBS 0.02fF
C11094 S.n10075 VSUBS 0.24fF $ **FLOATING
C11095 S.n10076 VSUBS 0.91fF $ **FLOATING
C11096 S.n10077 VSUBS 0.05fF $ **FLOATING
C11097 S.t1241 VSUBS 0.02fF
C11098 S.n10078 VSUBS 0.12fF $ **FLOATING
C11099 S.n10079 VSUBS 0.14fF $ **FLOATING
C11100 S.n10081 VSUBS 1.88fF $ **FLOATING
C11101 S.n10082 VSUBS 0.48fF $ **FLOATING
C11102 S.n10083 VSUBS 0.09fF $ **FLOATING
C11103 S.n10084 VSUBS 0.33fF $ **FLOATING
C11104 S.n10085 VSUBS 0.30fF $ **FLOATING
C11105 S.n10086 VSUBS 0.77fF $ **FLOATING
C11106 S.n10087 VSUBS 0.59fF $ **FLOATING
C11107 S.t1974 VSUBS 0.02fF
C11108 S.n10088 VSUBS 0.24fF $ **FLOATING
C11109 S.n10089 VSUBS 0.36fF $ **FLOATING
C11110 S.n10090 VSUBS 0.61fF $ **FLOATING
C11111 S.n10091 VSUBS 0.12fF $ **FLOATING
C11112 S.t1281 VSUBS 0.02fF
C11113 S.n10092 VSUBS 0.14fF $ **FLOATING
C11114 S.n10094 VSUBS 2.61fF $ **FLOATING
C11115 S.n10095 VSUBS 2.15fF $ **FLOATING
C11116 S.t2248 VSUBS 0.02fF
C11117 S.n10096 VSUBS 0.24fF $ **FLOATING
C11118 S.n10097 VSUBS 0.91fF $ **FLOATING
C11119 S.n10098 VSUBS 0.05fF $ **FLOATING
C11120 S.t2024 VSUBS 0.02fF
C11121 S.n10099 VSUBS 0.12fF $ **FLOATING
C11122 S.n10100 VSUBS 0.14fF $ **FLOATING
C11123 S.n10102 VSUBS 0.78fF $ **FLOATING
C11124 S.n10103 VSUBS 2.30fF $ **FLOATING
C11125 S.n10104 VSUBS 1.88fF $ **FLOATING
C11126 S.n10105 VSUBS 0.12fF $ **FLOATING
C11127 S.t2071 VSUBS 0.02fF
C11128 S.n10106 VSUBS 0.14fF $ **FLOATING
C11129 S.t368 VSUBS 0.02fF
C11130 S.n10108 VSUBS 0.24fF $ **FLOATING
C11131 S.n10109 VSUBS 0.36fF $ **FLOATING
C11132 S.n10110 VSUBS 0.61fF $ **FLOATING
C11133 S.n10111 VSUBS 1.39fF $ **FLOATING
C11134 S.n10112 VSUBS 0.71fF $ **FLOATING
C11135 S.n10113 VSUBS 1.14fF $ **FLOATING
C11136 S.n10114 VSUBS 0.35fF $ **FLOATING
C11137 S.n10115 VSUBS 2.02fF $ **FLOATING
C11138 S.t640 VSUBS 0.02fF
C11139 S.n10116 VSUBS 0.24fF $ **FLOATING
C11140 S.n10117 VSUBS 0.91fF $ **FLOATING
C11141 S.n10118 VSUBS 0.05fF $ **FLOATING
C11142 S.t418 VSUBS 0.02fF
C11143 S.n10119 VSUBS 0.12fF $ **FLOATING
C11144 S.n10120 VSUBS 0.14fF $ **FLOATING
C11145 S.n10122 VSUBS 1.89fF $ **FLOATING
C11146 S.n10123 VSUBS 1.88fF $ **FLOATING
C11147 S.t2487 VSUBS 0.02fF
C11148 S.n10124 VSUBS 0.24fF $ **FLOATING
C11149 S.n10125 VSUBS 0.36fF $ **FLOATING
C11150 S.n10126 VSUBS 0.61fF $ **FLOATING
C11151 S.n10127 VSUBS 0.12fF $ **FLOATING
C11152 S.t1667 VSUBS 0.02fF
C11153 S.n10128 VSUBS 0.14fF $ **FLOATING
C11154 S.n10130 VSUBS 1.16fF $ **FLOATING
C11155 S.n10131 VSUBS 0.22fF $ **FLOATING
C11156 S.n10132 VSUBS 0.25fF $ **FLOATING
C11157 S.n10133 VSUBS 0.09fF $ **FLOATING
C11158 S.n10134 VSUBS 1.88fF $ **FLOATING
C11159 S.t267 VSUBS 0.02fF
C11160 S.n10135 VSUBS 0.24fF $ **FLOATING
C11161 S.n10136 VSUBS 0.91fF $ **FLOATING
C11162 S.n10137 VSUBS 0.05fF $ **FLOATING
C11163 S.t2537 VSUBS 0.02fF
C11164 S.n10138 VSUBS 0.12fF $ **FLOATING
C11165 S.n10139 VSUBS 0.14fF $ **FLOATING
C11166 S.n10141 VSUBS 20.78fF $ **FLOATING
C11167 S.n10142 VSUBS 1.88fF $ **FLOATING
C11168 S.n10143 VSUBS 2.67fF $ **FLOATING
C11169 S.t2319 VSUBS 0.02fF
C11170 S.n10144 VSUBS 0.24fF $ **FLOATING
C11171 S.n10145 VSUBS 0.36fF $ **FLOATING
C11172 S.n10146 VSUBS 0.61fF $ **FLOATING
C11173 S.n10147 VSUBS 0.12fF $ **FLOATING
C11174 S.t1628 VSUBS 0.02fF
C11175 S.n10148 VSUBS 0.14fF $ **FLOATING
C11176 S.n10150 VSUBS 2.80fF $ **FLOATING
C11177 S.n10151 VSUBS 2.30fF $ **FLOATING
C11178 S.t2372 VSUBS 0.02fF
C11179 S.n10152 VSUBS 0.12fF $ **FLOATING
C11180 S.n10153 VSUBS 0.14fF $ **FLOATING
C11181 S.t49 VSUBS 0.02fF
C11182 S.n10155 VSUBS 0.24fF $ **FLOATING
C11183 S.n10156 VSUBS 0.91fF $ **FLOATING
C11184 S.n10157 VSUBS 0.05fF $ **FLOATING
C11185 S.n10158 VSUBS 2.80fF $ **FLOATING
C11186 S.n10159 VSUBS 1.88fF $ **FLOATING
C11187 S.n10160 VSUBS 0.12fF $ **FLOATING
C11188 S.t1255 VSUBS 0.02fF
C11189 S.n10161 VSUBS 0.14fF $ **FLOATING
C11190 S.t2070 VSUBS 0.02fF
C11191 S.n10163 VSUBS 0.24fF $ **FLOATING
C11192 S.n10164 VSUBS 0.36fF $ **FLOATING
C11193 S.n10165 VSUBS 0.61fF $ **FLOATING
C11194 S.n10166 VSUBS 2.67fF $ **FLOATING
C11195 S.n10167 VSUBS 2.30fF $ **FLOATING
C11196 S.t757 VSUBS 0.02fF
C11197 S.n10168 VSUBS 0.12fF $ **FLOATING
C11198 S.n10169 VSUBS 0.14fF $ **FLOATING
C11199 S.t2346 VSUBS 0.02fF
C11200 S.n10171 VSUBS 0.24fF $ **FLOATING
C11201 S.n10172 VSUBS 0.91fF $ **FLOATING
C11202 S.n10173 VSUBS 0.05fF $ **FLOATING
C11203 S.n10174 VSUBS 1.88fF $ **FLOATING
C11204 S.n10175 VSUBS 2.67fF $ **FLOATING
C11205 S.t339 VSUBS 0.02fF
C11206 S.n10176 VSUBS 0.24fF $ **FLOATING
C11207 S.n10177 VSUBS 0.36fF $ **FLOATING
C11208 S.n10178 VSUBS 0.61fF $ **FLOATING
C11209 S.n10179 VSUBS 0.12fF $ **FLOATING
C11210 S.t2038 VSUBS 0.02fF
C11211 S.n10180 VSUBS 0.14fF $ **FLOATING
C11212 S.n10182 VSUBS 2.80fF $ **FLOATING
C11213 S.n10183 VSUBS 2.30fF $ **FLOATING
C11214 S.t388 VSUBS 0.02fF
C11215 S.n10184 VSUBS 0.12fF $ **FLOATING
C11216 S.n10185 VSUBS 0.14fF $ **FLOATING
C11217 S.t609 VSUBS 0.02fF
C11218 S.n10187 VSUBS 0.24fF $ **FLOATING
C11219 S.n10188 VSUBS 0.91fF $ **FLOATING
C11220 S.n10189 VSUBS 0.05fF $ **FLOATING
C11221 S.n10190 VSUBS 1.88fF $ **FLOATING
C11222 S.n10191 VSUBS 2.67fF $ **FLOATING
C11223 S.t1125 VSUBS 0.02fF
C11224 S.n10192 VSUBS 0.24fF $ **FLOATING
C11225 S.n10193 VSUBS 0.36fF $ **FLOATING
C11226 S.n10194 VSUBS 0.61fF $ **FLOATING
C11227 S.n10195 VSUBS 0.12fF $ **FLOATING
C11228 S.t307 VSUBS 0.02fF
C11229 S.n10196 VSUBS 0.14fF $ **FLOATING
C11230 S.n10198 VSUBS 2.80fF $ **FLOATING
C11231 S.n10199 VSUBS 2.30fF $ **FLOATING
C11232 S.t1176 VSUBS 0.02fF
C11233 S.n10200 VSUBS 0.12fF $ **FLOATING
C11234 S.n10201 VSUBS 0.14fF $ **FLOATING
C11235 S.t1399 VSUBS 0.02fF
C11236 S.n10203 VSUBS 0.24fF $ **FLOATING
C11237 S.n10204 VSUBS 0.91fF $ **FLOATING
C11238 S.n10205 VSUBS 0.05fF $ **FLOATING
C11239 S.n10206 VSUBS 1.88fF $ **FLOATING
C11240 S.n10207 VSUBS 2.67fF $ **FLOATING
C11241 S.t1909 VSUBS 0.02fF
C11242 S.n10208 VSUBS 0.24fF $ **FLOATING
C11243 S.n10209 VSUBS 0.36fF $ **FLOATING
C11244 S.n10210 VSUBS 0.61fF $ **FLOATING
C11245 S.n10211 VSUBS 0.12fF $ **FLOATING
C11246 S.t1093 VSUBS 0.02fF
C11247 S.n10212 VSUBS 0.14fF $ **FLOATING
C11248 S.n10214 VSUBS 2.80fF $ **FLOATING
C11249 S.n10215 VSUBS 2.30fF $ **FLOATING
C11250 S.t1961 VSUBS 0.02fF
C11251 S.n10216 VSUBS 0.12fF $ **FLOATING
C11252 S.n10217 VSUBS 0.14fF $ **FLOATING
C11253 S.t2189 VSUBS 0.02fF
C11254 S.n10219 VSUBS 0.24fF $ **FLOATING
C11255 S.n10220 VSUBS 0.91fF $ **FLOATING
C11256 S.n10221 VSUBS 0.05fF $ **FLOATING
C11257 S.n10222 VSUBS 1.88fF $ **FLOATING
C11258 S.n10223 VSUBS 2.67fF $ **FLOATING
C11259 S.t162 VSUBS 0.02fF
C11260 S.n10224 VSUBS 0.24fF $ **FLOATING
C11261 S.n10225 VSUBS 0.36fF $ **FLOATING
C11262 S.n10226 VSUBS 0.61fF $ **FLOATING
C11263 S.n10227 VSUBS 0.12fF $ **FLOATING
C11264 S.t2001 VSUBS 0.02fF
C11265 S.n10228 VSUBS 0.14fF $ **FLOATING
C11266 S.n10230 VSUBS 2.80fF $ **FLOATING
C11267 S.n10231 VSUBS 2.30fF $ **FLOATING
C11268 S.t218 VSUBS 0.02fF
C11269 S.n10232 VSUBS 0.12fF $ **FLOATING
C11270 S.n10233 VSUBS 0.14fF $ **FLOATING
C11271 S.t455 VSUBS 0.02fF
C11272 S.n10235 VSUBS 0.24fF $ **FLOATING
C11273 S.n10236 VSUBS 0.91fF $ **FLOATING
C11274 S.n10237 VSUBS 0.05fF $ **FLOATING
C11275 S.n10238 VSUBS 1.88fF $ **FLOATING
C11276 S.n10239 VSUBS 2.67fF $ **FLOATING
C11277 S.t969 VSUBS 0.02fF
C11278 S.n10240 VSUBS 0.24fF $ **FLOATING
C11279 S.n10241 VSUBS 0.36fF $ **FLOATING
C11280 S.n10242 VSUBS 0.61fF $ **FLOATING
C11281 S.n10243 VSUBS 0.12fF $ **FLOATING
C11282 S.t1178 VSUBS 0.02fF
C11283 S.n10244 VSUBS 0.14fF $ **FLOATING
C11284 S.n10246 VSUBS 2.80fF $ **FLOATING
C11285 S.n10247 VSUBS 2.30fF $ **FLOATING
C11286 S.t2041 VSUBS 0.02fF
C11287 S.n10248 VSUBS 0.12fF $ **FLOATING
C11288 S.n10249 VSUBS 0.14fF $ **FLOATING
C11289 S.t1809 VSUBS 0.02fF
C11290 S.n10251 VSUBS 0.24fF $ **FLOATING
C11291 S.n10252 VSUBS 0.91fF $ **FLOATING
C11292 S.n10253 VSUBS 0.05fF $ **FLOATING
C11293 S.n10254 VSUBS 1.88fF $ **FLOATING
C11294 S.n10255 VSUBS 2.67fF $ **FLOATING
C11295 S.t1752 VSUBS 0.02fF
C11296 S.n10256 VSUBS 0.24fF $ **FLOATING
C11297 S.n10257 VSUBS 0.36fF $ **FLOATING
C11298 S.n10258 VSUBS 0.61fF $ **FLOATING
C11299 S.n10259 VSUBS 0.12fF $ **FLOATING
C11300 S.t1964 VSUBS 0.02fF
C11301 S.n10260 VSUBS 0.14fF $ **FLOATING
C11302 S.n10262 VSUBS 2.80fF $ **FLOATING
C11303 S.n10263 VSUBS 2.30fF $ **FLOATING
C11304 S.t309 VSUBS 0.02fF
C11305 S.n10264 VSUBS 0.12fF $ **FLOATING
C11306 S.n10265 VSUBS 0.14fF $ **FLOATING
C11307 S.t24 VSUBS 0.02fF
C11308 S.n10267 VSUBS 0.24fF $ **FLOATING
C11309 S.n10268 VSUBS 0.91fF $ **FLOATING
C11310 S.n10269 VSUBS 0.05fF $ **FLOATING
C11311 S.n10270 VSUBS 1.88fF $ **FLOATING
C11312 S.n10271 VSUBS 2.67fF $ **FLOATING
C11313 S.t2533 VSUBS 0.02fF
C11314 S.n10272 VSUBS 0.24fF $ **FLOATING
C11315 S.n10273 VSUBS 0.36fF $ **FLOATING
C11316 S.n10274 VSUBS 0.61fF $ **FLOATING
C11317 S.n10275 VSUBS 0.12fF $ **FLOATING
C11318 S.t224 VSUBS 0.02fF
C11319 S.n10276 VSUBS 0.14fF $ **FLOATING
C11320 S.n10278 VSUBS 2.80fF $ **FLOATING
C11321 S.n10279 VSUBS 2.30fF $ **FLOATING
C11322 S.t1099 VSUBS 0.02fF
C11323 S.n10280 VSUBS 0.12fF $ **FLOATING
C11324 S.n10281 VSUBS 0.14fF $ **FLOATING
C11325 S.t859 VSUBS 0.02fF
C11326 S.n10283 VSUBS 0.24fF $ **FLOATING
C11327 S.n10284 VSUBS 0.91fF $ **FLOATING
C11328 S.n10285 VSUBS 0.05fF $ **FLOATING
C11329 S.n10286 VSUBS 2.73fF $ **FLOATING
C11330 S.n10287 VSUBS 1.59fF $ **FLOATING
C11331 S.n10288 VSUBS 0.12fF $ **FLOATING
C11332 S.t1106 VSUBS 0.02fF
C11333 S.n10289 VSUBS 0.14fF $ **FLOATING
C11334 S.t1095 VSUBS 0.02fF
C11335 S.n10291 VSUBS 0.24fF $ **FLOATING
C11336 S.n10292 VSUBS 0.36fF $ **FLOATING
C11337 S.n10293 VSUBS 0.61fF $ **FLOATING
C11338 S.n10294 VSUBS 0.07fF $ **FLOATING
C11339 S.n10295 VSUBS 0.01fF $ **FLOATING
C11340 S.n10296 VSUBS 0.24fF $ **FLOATING
C11341 S.n10297 VSUBS 1.16fF $ **FLOATING
C11342 S.n10298 VSUBS 1.35fF $ **FLOATING
C11343 S.n10299 VSUBS 2.30fF $ **FLOATING
C11344 S.t125 VSUBS 0.02fF
C11345 S.n10300 VSUBS 0.12fF $ **FLOATING
C11346 S.n10301 VSUBS 0.14fF $ **FLOATING
C11347 S.t2483 VSUBS 0.02fF
C11348 S.n10303 VSUBS 0.24fF $ **FLOATING
C11349 S.n10304 VSUBS 0.91fF $ **FLOATING
C11350 S.n10305 VSUBS 0.05fF $ **FLOATING
C11351 S.t124 VSUBS 48.27fF
C11352 S.t1643 VSUBS 0.02fF
C11353 S.n10306 VSUBS 0.24fF $ **FLOATING
C11354 S.n10307 VSUBS 0.91fF $ **FLOATING
C11355 S.n10308 VSUBS 0.05fF $ **FLOATING
C11356 S.t1879 VSUBS 0.02fF
C11357 S.n10309 VSUBS 0.12fF $ **FLOATING
C11358 S.n10310 VSUBS 0.14fF $ **FLOATING
C11359 S.n10312 VSUBS 0.12fF $ **FLOATING
C11360 S.t1011 VSUBS 0.02fF
C11361 S.n10313 VSUBS 0.14fF $ **FLOATING
C11362 S.n10315 VSUBS 5.17fF $ **FLOATING
C11363 S.n10316 VSUBS 5.44fF $ **FLOATING
C11364 S.t1462 VSUBS 0.02fF
C11365 S.n10317 VSUBS 0.12fF $ **FLOATING
C11366 S.n10318 VSUBS 0.14fF $ **FLOATING
C11367 S.t1248 VSUBS 0.02fF
C11368 S.n10320 VSUBS 0.24fF $ **FLOATING
C11369 S.n10321 VSUBS 0.91fF $ **FLOATING
C11370 S.n10322 VSUBS 0.05fF $ **FLOATING
C11371 S.t61 VSUBS 47.89fF
C11372 S.t634 VSUBS 0.02fF
C11373 S.n10323 VSUBS 0.01fF $ **FLOATING
C11374 S.n10324 VSUBS 0.26fF $ **FLOATING
C11375 S.t755 VSUBS 0.02fF
C11376 S.n10326 VSUBS 1.19fF $ **FLOATING
C11377 S.n10327 VSUBS 0.05fF $ **FLOATING
C11378 S.t681 VSUBS 0.02fF
C11379 S.n10328 VSUBS 0.64fF $ **FLOATING
C11380 S.n10329 VSUBS 0.61fF $ **FLOATING
C11381 S.n10330 VSUBS 8.97fF $ **FLOATING
C11382 S.n10331 VSUBS 8.97fF $ **FLOATING
C11383 S.n10332 VSUBS 0.60fF $ **FLOATING
C11384 S.n10333 VSUBS 0.22fF $ **FLOATING
C11385 S.n10334 VSUBS 0.59fF $ **FLOATING
C11386 S.n10335 VSUBS 3.39fF $ **FLOATING
C11387 S.n10336 VSUBS 0.29fF $ **FLOATING
C11388 S.t23 VSUBS 21.42fF
C11389 S.n10337 VSUBS 21.71fF $ **FLOATING
C11390 S.n10338 VSUBS 0.77fF $ **FLOATING
C11391 S.n10339 VSUBS 0.28fF $ **FLOATING
C11392 S.n10340 VSUBS 4.00fF $ **FLOATING
C11393 S.n10341 VSUBS 1.35fF $ **FLOATING
C11394 S.n10342 VSUBS 0.01fF $ **FLOATING
C11395 S.n10343 VSUBS 0.02fF $ **FLOATING
C11396 S.n10344 VSUBS 0.03fF $ **FLOATING
C11397 S.n10345 VSUBS 0.04fF $ **FLOATING
C11398 S.n10346 VSUBS 0.17fF $ **FLOATING
C11399 S.n10347 VSUBS 0.01fF $ **FLOATING
C11400 S.n10348 VSUBS 0.02fF $ **FLOATING
C11401 S.n10349 VSUBS 0.01fF $ **FLOATING
C11402 S.n10350 VSUBS 0.01fF $ **FLOATING
C11403 S.n10351 VSUBS 0.01fF $ **FLOATING
C11404 S.n10352 VSUBS 0.01fF $ **FLOATING
C11405 S.n10353 VSUBS 0.02fF $ **FLOATING
C11406 S.n10354 VSUBS 0.01fF $ **FLOATING
C11407 S.n10355 VSUBS 0.02fF $ **FLOATING
C11408 S.n10356 VSUBS 0.05fF $ **FLOATING
C11409 S.n10357 VSUBS 0.04fF $ **FLOATING
C11410 S.n10358 VSUBS 0.11fF $ **FLOATING
C11411 S.n10359 VSUBS 0.38fF $ **FLOATING
C11412 S.n10360 VSUBS 0.20fF $ **FLOATING
C11413 S.n10361 VSUBS 4.39fF $ **FLOATING
C11414 S.n10362 VSUBS 0.24fF $ **FLOATING
C11415 S.n10363 VSUBS 1.50fF $ **FLOATING
C11416 S.n10364 VSUBS 1.31fF $ **FLOATING
C11417 S.n10365 VSUBS 0.28fF $ **FLOATING
C11418 S.n10366 VSUBS 1.88fF $ **FLOATING
C11419 S.n10367 VSUBS 0.46fF $ **FLOATING
C11420 S.n10368 VSUBS 0.22fF $ **FLOATING
C11421 S.n10369 VSUBS 0.38fF $ **FLOATING
C11422 S.n10370 VSUBS 0.16fF $ **FLOATING
C11423 S.n10371 VSUBS 0.28fF $ **FLOATING
C11424 S.n10372 VSUBS 0.21fF $ **FLOATING
C11425 S.n10373 VSUBS 0.30fF $ **FLOATING
C11426 S.n10374 VSUBS 0.42fF $ **FLOATING
C11427 S.n10375 VSUBS 0.21fF $ **FLOATING
C11428 S.t2544 VSUBS 0.02fF
C11429 S.n10376 VSUBS 0.24fF $ **FLOATING
C11430 S.n10377 VSUBS 0.36fF $ **FLOATING
C11431 S.n10378 VSUBS 0.61fF $ **FLOATING
C11432 S.n10379 VSUBS 0.12fF $ **FLOATING
C11433 S.t1732 VSUBS 0.02fF
C11434 S.n10380 VSUBS 0.14fF $ **FLOATING
C11435 S.n10382 VSUBS 0.04fF $ **FLOATING
C11436 S.n10383 VSUBS 0.03fF $ **FLOATING
C11437 S.n10384 VSUBS 0.03fF $ **FLOATING
C11438 S.n10385 VSUBS 0.10fF $ **FLOATING
C11439 S.n10386 VSUBS 0.36fF $ **FLOATING
C11440 S.n10387 VSUBS 0.38fF $ **FLOATING
C11441 S.n10388 VSUBS 0.11fF $ **FLOATING
C11442 S.n10389 VSUBS 0.12fF $ **FLOATING
C11443 S.n10390 VSUBS 0.07fF $ **FLOATING
C11444 S.n10391 VSUBS 0.12fF $ **FLOATING
C11445 S.n10392 VSUBS 0.18fF $ **FLOATING
C11446 S.n10393 VSUBS 3.99fF $ **FLOATING
C11447 S.t323 VSUBS 0.02fF
C11448 S.n10394 VSUBS 0.24fF $ **FLOATING
C11449 S.n10395 VSUBS 0.91fF $ **FLOATING
C11450 S.n10396 VSUBS 0.05fF $ **FLOATING
C11451 S.t36 VSUBS 0.02fF
C11452 S.n10397 VSUBS 0.12fF $ **FLOATING
C11453 S.n10398 VSUBS 0.14fF $ **FLOATING
C11454 S.n10400 VSUBS 0.25fF $ **FLOATING
C11455 S.n10401 VSUBS 0.09fF $ **FLOATING
C11456 S.n10402 VSUBS 0.21fF $ **FLOATING
C11457 S.n10403 VSUBS 1.28fF $ **FLOATING
C11458 S.n10404 VSUBS 0.53fF $ **FLOATING
C11459 S.n10405 VSUBS 1.88fF $ **FLOATING
C11460 S.n10406 VSUBS 0.12fF $ **FLOATING
C11461 S.t100 VSUBS 0.02fF
C11462 S.n10407 VSUBS 0.14fF $ **FLOATING
C11463 S.t940 VSUBS 0.02fF
C11464 S.n10409 VSUBS 0.24fF $ **FLOATING
C11465 S.n10410 VSUBS 0.36fF $ **FLOATING
C11466 S.n10411 VSUBS 0.61fF $ **FLOATING
C11467 S.n10412 VSUBS 1.58fF $ **FLOATING
C11468 S.n10413 VSUBS 2.45fF $ **FLOATING
C11469 S.t1234 VSUBS 0.02fF
C11470 S.n10414 VSUBS 0.24fF $ **FLOATING
C11471 S.n10415 VSUBS 0.91fF $ **FLOATING
C11472 S.n10416 VSUBS 0.05fF $ **FLOATING
C11473 S.t997 VSUBS 0.02fF
C11474 S.n10417 VSUBS 0.12fF $ **FLOATING
C11475 S.n10418 VSUBS 0.14fF $ **FLOATING
C11476 S.n10420 VSUBS 1.89fF $ **FLOATING
C11477 S.n10421 VSUBS 0.06fF $ **FLOATING
C11478 S.n10422 VSUBS 0.03fF $ **FLOATING
C11479 S.n10423 VSUBS 0.04fF $ **FLOATING
C11480 S.n10424 VSUBS 0.99fF $ **FLOATING
C11481 S.n10425 VSUBS 0.02fF $ **FLOATING
C11482 S.n10426 VSUBS 0.01fF $ **FLOATING
C11483 S.n10427 VSUBS 0.02fF $ **FLOATING
C11484 S.n10428 VSUBS 0.08fF $ **FLOATING
C11485 S.n10429 VSUBS 0.36fF $ **FLOATING
C11486 S.n10430 VSUBS 1.85fF $ **FLOATING
C11487 S.t553 VSUBS 0.02fF
C11488 S.n10431 VSUBS 0.24fF $ **FLOATING
C11489 S.n10432 VSUBS 0.36fF $ **FLOATING
C11490 S.n10433 VSUBS 0.61fF $ **FLOATING
C11491 S.n10434 VSUBS 0.12fF $ **FLOATING
C11492 S.t2253 VSUBS 0.02fF
C11493 S.n10435 VSUBS 0.14fF $ **FLOATING
C11494 S.n10437 VSUBS 0.70fF $ **FLOATING
C11495 S.n10438 VSUBS 0.23fF $ **FLOATING
C11496 S.n10439 VSUBS 0.23fF $ **FLOATING
C11497 S.n10440 VSUBS 0.70fF $ **FLOATING
C11498 S.n10441 VSUBS 1.16fF $ **FLOATING
C11499 S.n10442 VSUBS 0.22fF $ **FLOATING
C11500 S.n10443 VSUBS 0.25fF $ **FLOATING
C11501 S.n10444 VSUBS 0.09fF $ **FLOATING
C11502 S.n10445 VSUBS 1.88fF $ **FLOATING
C11503 S.t833 VSUBS 0.02fF
C11504 S.n10446 VSUBS 0.24fF $ **FLOATING
C11505 S.n10447 VSUBS 0.91fF $ **FLOATING
C11506 S.n10448 VSUBS 0.05fF $ **FLOATING
C11507 S.t1780 VSUBS 0.02fF
C11508 S.n10449 VSUBS 0.12fF $ **FLOATING
C11509 S.n10450 VSUBS 0.14fF $ **FLOATING
C11510 S.n10452 VSUBS 20.78fF $ **FLOATING
C11511 S.n10453 VSUBS 1.72fF $ **FLOATING
C11512 S.n10454 VSUBS 0.66fF $ **FLOATING
C11513 S.n10455 VSUBS 0.69fF $ **FLOATING
C11514 S.n10456 VSUBS 0.72fF $ **FLOATING
C11515 S.n10457 VSUBS 0.36fF $ **FLOATING
C11516 S.t1762 VSUBS 0.02fF
C11517 S.n10458 VSUBS 0.24fF $ **FLOATING
C11518 S.n10459 VSUBS 0.36fF $ **FLOATING
C11519 S.n10460 VSUBS 0.61fF $ **FLOATING
C11520 S.n10461 VSUBS 0.12fF $ **FLOATING
C11521 S.t946 VSUBS 0.02fF
C11522 S.n10462 VSUBS 0.14fF $ **FLOATING
C11523 S.n10464 VSUBS 0.31fF $ **FLOATING
C11524 S.n10465 VSUBS 0.23fF $ **FLOATING
C11525 S.n10466 VSUBS 0.66fF $ **FLOATING
C11526 S.n10467 VSUBS 0.95fF $ **FLOATING
C11527 S.n10468 VSUBS 0.23fF $ **FLOATING
C11528 S.n10469 VSUBS 0.21fF $ **FLOATING
C11529 S.n10470 VSUBS 0.20fF $ **FLOATING
C11530 S.n10471 VSUBS 0.06fF $ **FLOATING
C11531 S.n10472 VSUBS 0.09fF $ **FLOATING
C11532 S.n10473 VSUBS 0.10fF $ **FLOATING
C11533 S.n10474 VSUBS 1.67fF $ **FLOATING
C11534 S.t1815 VSUBS 0.02fF
C11535 S.n10475 VSUBS 0.12fF $ **FLOATING
C11536 S.n10476 VSUBS 0.14fF $ **FLOATING
C11537 S.t2056 VSUBS 0.02fF
C11538 S.n10478 VSUBS 0.24fF $ **FLOATING
C11539 S.n10479 VSUBS 0.91fF $ **FLOATING
C11540 S.n10480 VSUBS 0.05fF $ **FLOATING
C11541 S.n10481 VSUBS 1.88fF $ **FLOATING
C11542 S.n10482 VSUBS 0.12fF $ **FLOATING
C11543 S.t1114 VSUBS 0.02fF
C11544 S.n10483 VSUBS 0.14fF $ **FLOATING
C11545 S.t1978 VSUBS 0.02fF
C11546 S.n10485 VSUBS 0.12fF $ **FLOATING
C11547 S.n10486 VSUBS 0.14fF $ **FLOATING
C11548 S.t2205 VSUBS 0.02fF
C11549 S.n10488 VSUBS 0.24fF $ **FLOATING
C11550 S.n10489 VSUBS 0.91fF $ **FLOATING
C11551 S.n10490 VSUBS 0.05fF $ **FLOATING
C11552 S.t1925 VSUBS 0.02fF
C11553 S.n10491 VSUBS 0.24fF $ **FLOATING
C11554 S.n10492 VSUBS 0.36fF $ **FLOATING
C11555 S.n10493 VSUBS 0.61fF $ **FLOATING
C11556 S.n10494 VSUBS 0.32fF $ **FLOATING
C11557 S.n10495 VSUBS 1.09fF $ **FLOATING
C11558 S.n10496 VSUBS 0.15fF $ **FLOATING
C11559 S.n10497 VSUBS 2.10fF $ **FLOATING
C11560 S.n10498 VSUBS 2.94fF $ **FLOATING
C11561 S.n10499 VSUBS 1.88fF $ **FLOATING
C11562 S.n10500 VSUBS 0.12fF $ **FLOATING
C11563 S.t521 VSUBS 0.02fF
C11564 S.n10501 VSUBS 0.14fF $ **FLOATING
C11565 S.t1340 VSUBS 0.02fF
C11566 S.n10503 VSUBS 0.24fF $ **FLOATING
C11567 S.n10504 VSUBS 0.36fF $ **FLOATING
C11568 S.n10505 VSUBS 0.61fF $ **FLOATING
C11569 S.n10506 VSUBS 0.92fF $ **FLOATING
C11570 S.n10507 VSUBS 0.32fF $ **FLOATING
C11571 S.n10508 VSUBS 0.92fF $ **FLOATING
C11572 S.n10509 VSUBS 1.09fF $ **FLOATING
C11573 S.n10510 VSUBS 0.15fF $ **FLOATING
C11574 S.n10511 VSUBS 4.96fF $ **FLOATING
C11575 S.t1389 VSUBS 0.02fF
C11576 S.n10512 VSUBS 0.12fF $ **FLOATING
C11577 S.n10513 VSUBS 0.14fF $ **FLOATING
C11578 S.t1615 VSUBS 0.02fF
C11579 S.n10515 VSUBS 0.24fF $ **FLOATING
C11580 S.n10516 VSUBS 0.91fF $ **FLOATING
C11581 S.n10517 VSUBS 0.05fF $ **FLOATING
C11582 S.n10518 VSUBS 1.88fF $ **FLOATING
C11583 S.n10519 VSUBS 2.67fF $ **FLOATING
C11584 S.t2128 VSUBS 0.02fF
C11585 S.n10520 VSUBS 0.24fF $ **FLOATING
C11586 S.n10521 VSUBS 0.36fF $ **FLOATING
C11587 S.n10522 VSUBS 0.61fF $ **FLOATING
C11588 S.n10523 VSUBS 0.12fF $ **FLOATING
C11589 S.t1308 VSUBS 0.02fF
C11590 S.n10524 VSUBS 0.14fF $ **FLOATING
C11591 S.n10526 VSUBS 1.88fF $ **FLOATING
C11592 S.n10527 VSUBS 2.67fF $ **FLOATING
C11593 S.t180 VSUBS 0.02fF
C11594 S.n10528 VSUBS 0.24fF $ **FLOATING
C11595 S.n10529 VSUBS 0.36fF $ **FLOATING
C11596 S.n10530 VSUBS 0.61fF $ **FLOATING
C11597 S.t473 VSUBS 0.02fF
C11598 S.n10531 VSUBS 0.24fF $ **FLOATING
C11599 S.n10532 VSUBS 0.91fF $ **FLOATING
C11600 S.n10533 VSUBS 0.05fF $ **FLOATING
C11601 S.t241 VSUBS 0.02fF
C11602 S.n10534 VSUBS 0.12fF $ **FLOATING
C11603 S.n10535 VSUBS 0.14fF $ **FLOATING
C11604 S.n10537 VSUBS 0.12fF $ **FLOATING
C11605 S.t1894 VSUBS 0.02fF
C11606 S.n10538 VSUBS 0.14fF $ **FLOATING
C11607 S.n10540 VSUBS 2.30fF $ **FLOATING
C11608 S.n10541 VSUBS 2.94fF $ **FLOATING
C11609 S.n10542 VSUBS 5.16fF $ **FLOATING
C11610 S.t2176 VSUBS 0.02fF
C11611 S.n10543 VSUBS 0.12fF $ **FLOATING
C11612 S.n10544 VSUBS 0.14fF $ **FLOATING
C11613 S.t2401 VSUBS 0.02fF
C11614 S.n10546 VSUBS 0.24fF $ **FLOATING
C11615 S.n10547 VSUBS 0.91fF $ **FLOATING
C11616 S.n10548 VSUBS 0.05fF $ **FLOATING
C11617 S.n10549 VSUBS 1.88fF $ **FLOATING
C11618 S.n10550 VSUBS 2.67fF $ **FLOATING
C11619 S.t394 VSUBS 0.02fF
C11620 S.n10551 VSUBS 0.24fF $ **FLOATING
C11621 S.n10552 VSUBS 0.36fF $ **FLOATING
C11622 S.n10553 VSUBS 0.61fF $ **FLOATING
C11623 S.n10554 VSUBS 0.12fF $ **FLOATING
C11624 S.t2095 VSUBS 0.02fF
C11625 S.n10555 VSUBS 0.14fF $ **FLOATING
C11626 S.n10557 VSUBS 5.17fF $ **FLOATING
C11627 S.t441 VSUBS 0.02fF
C11628 S.n10558 VSUBS 0.12fF $ **FLOATING
C11629 S.n10559 VSUBS 0.14fF $ **FLOATING
C11630 S.t664 VSUBS 0.02fF
C11631 S.n10561 VSUBS 0.24fF $ **FLOATING
C11632 S.n10562 VSUBS 0.91fF $ **FLOATING
C11633 S.n10563 VSUBS 0.05fF $ **FLOATING
C11634 S.n10564 VSUBS 1.88fF $ **FLOATING
C11635 S.n10565 VSUBS 0.12fF $ **FLOATING
C11636 S.t486 VSUBS 0.02fF
C11637 S.n10566 VSUBS 0.14fF $ **FLOATING
C11638 S.t1300 VSUBS 0.02fF
C11639 S.n10568 VSUBS 0.24fF $ **FLOATING
C11640 S.n10569 VSUBS 0.36fF $ **FLOATING
C11641 S.n10570 VSUBS 0.61fF $ **FLOATING
C11642 S.n10571 VSUBS 2.67fF $ **FLOATING
C11643 S.n10572 VSUBS 5.17fF $ **FLOATING
C11644 S.t1353 VSUBS 0.02fF
C11645 S.n10573 VSUBS 0.12fF $ **FLOATING
C11646 S.n10574 VSUBS 0.14fF $ **FLOATING
C11647 S.t1569 VSUBS 0.02fF
C11648 S.n10576 VSUBS 0.24fF $ **FLOATING
C11649 S.n10577 VSUBS 0.91fF $ **FLOATING
C11650 S.n10578 VSUBS 0.05fF $ **FLOATING
C11651 S.n10579 VSUBS 1.88fF $ **FLOATING
C11652 S.n10580 VSUBS 2.67fF $ **FLOATING
C11653 S.t909 VSUBS 0.02fF
C11654 S.n10581 VSUBS 0.24fF $ **FLOATING
C11655 S.n10582 VSUBS 0.36fF $ **FLOATING
C11656 S.n10583 VSUBS 0.61fF $ **FLOATING
C11657 S.n10584 VSUBS 0.12fF $ **FLOATING
C11658 S.t57 VSUBS 0.02fF
C11659 S.n10585 VSUBS 0.14fF $ **FLOATING
C11660 S.n10587 VSUBS 5.17fF $ **FLOATING
C11661 S.t963 VSUBS 0.02fF
C11662 S.n10588 VSUBS 0.12fF $ **FLOATING
C11663 S.n10589 VSUBS 0.14fF $ **FLOATING
C11664 S.t1210 VSUBS 0.02fF
C11665 S.n10591 VSUBS 0.24fF $ **FLOATING
C11666 S.n10592 VSUBS 0.91fF $ **FLOATING
C11667 S.n10593 VSUBS 0.05fF $ **FLOATING
C11668 S.n10594 VSUBS 1.88fF $ **FLOATING
C11669 S.n10595 VSUBS 2.67fF $ **FLOATING
C11670 S.t1690 VSUBS 0.02fF
C11671 S.n10596 VSUBS 0.24fF $ **FLOATING
C11672 S.n10597 VSUBS 0.36fF $ **FLOATING
C11673 S.n10598 VSUBS 0.61fF $ **FLOATING
C11674 S.n10599 VSUBS 0.12fF $ **FLOATING
C11675 S.t875 VSUBS 0.02fF
C11676 S.n10600 VSUBS 0.14fF $ **FLOATING
C11677 S.n10602 VSUBS 5.17fF $ **FLOATING
C11678 S.t1744 VSUBS 0.02fF
C11679 S.n10603 VSUBS 0.12fF $ **FLOATING
C11680 S.n10604 VSUBS 0.14fF $ **FLOATING
C11681 S.t1987 VSUBS 0.02fF
C11682 S.n10606 VSUBS 0.24fF $ **FLOATING
C11683 S.n10607 VSUBS 0.91fF $ **FLOATING
C11684 S.n10608 VSUBS 0.05fF $ **FLOATING
C11685 S.n10609 VSUBS 1.88fF $ **FLOATING
C11686 S.n10610 VSUBS 2.67fF $ **FLOATING
C11687 S.t2476 VSUBS 0.02fF
C11688 S.n10611 VSUBS 0.24fF $ **FLOATING
C11689 S.n10612 VSUBS 0.36fF $ **FLOATING
C11690 S.n10613 VSUBS 0.61fF $ **FLOATING
C11691 S.n10614 VSUBS 0.12fF $ **FLOATING
C11692 S.t1656 VSUBS 0.02fF
C11693 S.n10615 VSUBS 0.14fF $ **FLOATING
C11694 S.n10617 VSUBS 5.17fF $ **FLOATING
C11695 S.t2525 VSUBS 0.02fF
C11696 S.n10618 VSUBS 0.12fF $ **FLOATING
C11697 S.n10619 VSUBS 0.14fF $ **FLOATING
C11698 S.t255 VSUBS 0.02fF
C11699 S.n10621 VSUBS 0.24fF $ **FLOATING
C11700 S.n10622 VSUBS 0.91fF $ **FLOATING
C11701 S.n10623 VSUBS 0.05fF $ **FLOATING
C11702 S.n10624 VSUBS 1.88fF $ **FLOATING
C11703 S.n10625 VSUBS 2.67fF $ **FLOATING
C11704 S.t736 VSUBS 0.02fF
C11705 S.n10626 VSUBS 0.24fF $ **FLOATING
C11706 S.n10627 VSUBS 0.36fF $ **FLOATING
C11707 S.n10628 VSUBS 0.61fF $ **FLOATING
C11708 S.n10629 VSUBS 0.12fF $ **FLOATING
C11709 S.t2445 VSUBS 0.02fF
C11710 S.n10630 VSUBS 0.14fF $ **FLOATING
C11711 S.n10632 VSUBS 5.17fF $ **FLOATING
C11712 S.t789 VSUBS 0.02fF
C11713 S.n10633 VSUBS 0.12fF $ **FLOATING
C11714 S.n10634 VSUBS 0.14fF $ **FLOATING
C11715 S.t1040 VSUBS 0.02fF
C11716 S.n10636 VSUBS 0.24fF $ **FLOATING
C11717 S.n10637 VSUBS 0.91fF $ **FLOATING
C11718 S.n10638 VSUBS 0.05fF $ **FLOATING
C11719 S.n10639 VSUBS 1.88fF $ **FLOATING
C11720 S.n10640 VSUBS 2.67fF $ **FLOATING
C11721 S.t998 VSUBS 0.02fF
C11722 S.n10641 VSUBS 0.24fF $ **FLOATING
C11723 S.n10642 VSUBS 0.36fF $ **FLOATING
C11724 S.n10643 VSUBS 0.61fF $ **FLOATING
C11725 S.n10644 VSUBS 0.12fF $ **FLOATING
C11726 S.t1209 VSUBS 0.02fF
C11727 S.n10645 VSUBS 0.14fF $ **FLOATING
C11728 S.n10647 VSUBS 5.17fF $ **FLOATING
C11729 S.t1705 VSUBS 0.02fF
C11730 S.n10648 VSUBS 0.12fF $ **FLOATING
C11731 S.n10649 VSUBS 0.14fF $ **FLOATING
C11732 S.t1839 VSUBS 0.02fF
C11733 S.n10651 VSUBS 0.24fF $ **FLOATING
C11734 S.n10652 VSUBS 0.91fF $ **FLOATING
C11735 S.n10653 VSUBS 0.05fF $ **FLOATING
C11736 S.n10654 VSUBS 1.88fF $ **FLOATING
C11737 S.n10655 VSUBS 2.67fF $ **FLOATING
C11738 S.t1781 VSUBS 0.02fF
C11739 S.n10656 VSUBS 0.24fF $ **FLOATING
C11740 S.n10657 VSUBS 0.36fF $ **FLOATING
C11741 S.n10658 VSUBS 0.61fF $ **FLOATING
C11742 S.n10659 VSUBS 0.12fF $ **FLOATING
C11743 S.t1986 VSUBS 0.02fF
C11744 S.n10660 VSUBS 0.14fF $ **FLOATING
C11745 S.n10662 VSUBS 5.17fF $ **FLOATING
C11746 S.t337 VSUBS 0.02fF
C11747 S.n10663 VSUBS 0.12fF $ **FLOATING
C11748 S.n10664 VSUBS 0.14fF $ **FLOATING
C11749 S.t68 VSUBS 0.02fF
C11750 S.n10666 VSUBS 0.24fF $ **FLOATING
C11751 S.n10667 VSUBS 0.91fF $ **FLOATING
C11752 S.n10668 VSUBS 0.05fF $ **FLOATING
C11753 S.n10669 VSUBS 1.88fF $ **FLOATING
C11754 S.n10670 VSUBS 2.67fF $ **FLOATING
C11755 S.t2561 VSUBS 0.02fF
C11756 S.n10671 VSUBS 0.24fF $ **FLOATING
C11757 S.n10672 VSUBS 0.36fF $ **FLOATING
C11758 S.n10673 VSUBS 0.61fF $ **FLOATING
C11759 S.n10674 VSUBS 0.12fF $ **FLOATING
C11760 S.t253 VSUBS 0.02fF
C11761 S.n10675 VSUBS 0.14fF $ **FLOATING
C11762 S.n10677 VSUBS 5.17fF $ **FLOATING
C11763 S.t1123 VSUBS 0.02fF
C11764 S.n10678 VSUBS 0.12fF $ **FLOATING
C11765 S.n10679 VSUBS 0.14fF $ **FLOATING
C11766 S.t884 VSUBS 0.02fF
C11767 S.n10681 VSUBS 0.24fF $ **FLOATING
C11768 S.n10682 VSUBS 0.91fF $ **FLOATING
C11769 S.n10683 VSUBS 0.05fF $ **FLOATING
C11770 S.n10684 VSUBS 1.88fF $ **FLOATING
C11771 S.n10685 VSUBS 2.67fF $ **FLOATING
C11772 S.t827 VSUBS 0.02fF
C11773 S.n10686 VSUBS 0.24fF $ **FLOATING
C11774 S.n10687 VSUBS 0.36fF $ **FLOATING
C11775 S.n10688 VSUBS 0.61fF $ **FLOATING
C11776 S.n10689 VSUBS 0.12fF $ **FLOATING
C11777 S.t1037 VSUBS 0.02fF
C11778 S.n10690 VSUBS 0.14fF $ **FLOATING
C11779 S.n10692 VSUBS 4.89fF $ **FLOATING
C11780 S.t1905 VSUBS 0.02fF
C11781 S.n10693 VSUBS 0.12fF $ **FLOATING
C11782 S.n10694 VSUBS 0.14fF $ **FLOATING
C11783 S.t1666 VSUBS 0.02fF
C11784 S.n10696 VSUBS 0.24fF $ **FLOATING
C11785 S.n10697 VSUBS 0.91fF $ **FLOATING
C11786 S.n10698 VSUBS 0.05fF $ **FLOATING
C11787 S.n10699 VSUBS 1.88fF $ **FLOATING
C11788 S.n10700 VSUBS 2.67fF $ **FLOATING
C11789 S.t1610 VSUBS 0.02fF
C11790 S.n10701 VSUBS 0.24fF $ **FLOATING
C11791 S.n10702 VSUBS 0.36fF $ **FLOATING
C11792 S.n10703 VSUBS 0.61fF $ **FLOATING
C11793 S.n10704 VSUBS 0.12fF $ **FLOATING
C11794 S.t1818 VSUBS 0.02fF
C11795 S.n10705 VSUBS 0.14fF $ **FLOATING
C11796 S.n10707 VSUBS 1.88fF $ **FLOATING
C11797 S.n10708 VSUBS 2.68fF $ **FLOATING
C11798 S.t1635 VSUBS 0.02fF
C11799 S.n10709 VSUBS 0.24fF $ **FLOATING
C11800 S.n10710 VSUBS 0.36fF $ **FLOATING
C11801 S.n10711 VSUBS 0.61fF $ **FLOATING
C11802 S.t2339 VSUBS 0.02fF
C11803 S.n10712 VSUBS 1.22fF $ **FLOATING
C11804 S.n10713 VSUBS 0.61fF $ **FLOATING
C11805 S.n10714 VSUBS 1.15fF $ **FLOATING
C11806 S.n10715 VSUBS 3.00fF $ **FLOATING
C11807 S.n10716 VSUBS 0.01fF $ **FLOATING
C11808 S.n10717 VSUBS 0.97fF $ **FLOATING
C11809 S.t15 VSUBS 21.42fF
C11810 S.n10718 VSUBS 20.29fF $ **FLOATING
C11811 S.n10720 VSUBS 0.38fF $ **FLOATING
C11812 S.n10721 VSUBS 0.23fF $ **FLOATING
C11813 S.n10722 VSUBS 2.89fF $ **FLOATING
C11814 S.n10723 VSUBS 2.46fF $ **FLOATING
C11815 S.n10724 VSUBS 2.53fF $ **FLOATING
C11816 S.n10725 VSUBS 3.94fF $ **FLOATING
C11817 S.n10726 VSUBS 0.25fF $ **FLOATING
C11818 S.n10727 VSUBS 0.01fF $ **FLOATING
C11819 S.t1522 VSUBS 0.02fF
C11820 S.n10728 VSUBS 0.26fF $ **FLOATING
C11821 S.t81 VSUBS 0.02fF
C11822 S.n10729 VSUBS 0.95fF $ **FLOATING
C11823 S.n10730 VSUBS 0.71fF $ **FLOATING
C11824 S.n10731 VSUBS 1.88fF $ **FLOATING
C11825 S.n10732 VSUBS 0.48fF $ **FLOATING
C11826 S.n10733 VSUBS 0.09fF $ **FLOATING
C11827 S.n10734 VSUBS 0.33fF $ **FLOATING
C11828 S.n10735 VSUBS 0.30fF $ **FLOATING
C11829 S.n10736 VSUBS 0.77fF $ **FLOATING
C11830 S.n10737 VSUBS 0.59fF $ **FLOATING
C11831 S.t602 VSUBS 0.02fF
C11832 S.n10738 VSUBS 0.24fF $ **FLOATING
C11833 S.n10739 VSUBS 0.36fF $ **FLOATING
C11834 S.n10740 VSUBS 0.61fF $ **FLOATING
C11835 S.n10741 VSUBS 0.12fF $ **FLOATING
C11836 S.t2310 VSUBS 0.02fF
C11837 S.n10742 VSUBS 0.14fF $ **FLOATING
C11838 S.n10744 VSUBS 1.44fF $ **FLOATING
C11839 S.n10745 VSUBS 2.15fF $ **FLOATING
C11840 S.t893 VSUBS 0.02fF
C11841 S.n10746 VSUBS 0.24fF $ **FLOATING
C11842 S.n10747 VSUBS 0.91fF $ **FLOATING
C11843 S.n10748 VSUBS 0.05fF $ **FLOATING
C11844 S.t652 VSUBS 0.02fF
C11845 S.n10749 VSUBS 0.12fF $ **FLOATING
C11846 S.n10750 VSUBS 0.14fF $ **FLOATING
C11847 S.n10752 VSUBS 0.78fF $ **FLOATING
C11848 S.n10753 VSUBS 2.30fF $ **FLOATING
C11849 S.n10754 VSUBS 1.88fF $ **FLOATING
C11850 S.n10755 VSUBS 0.12fF $ **FLOATING
C11851 S.t696 VSUBS 0.02fF
C11852 S.n10756 VSUBS 0.14fF $ **FLOATING
C11853 S.t1396 VSUBS 0.02fF
C11854 S.n10758 VSUBS 0.24fF $ **FLOATING
C11855 S.n10759 VSUBS 0.36fF $ **FLOATING
C11856 S.n10760 VSUBS 0.61fF $ **FLOATING
C11857 S.n10761 VSUBS 1.39fF $ **FLOATING
C11858 S.n10762 VSUBS 0.71fF $ **FLOATING
C11859 S.n10763 VSUBS 1.14fF $ **FLOATING
C11860 S.n10764 VSUBS 0.35fF $ **FLOATING
C11861 S.n10765 VSUBS 2.02fF $ **FLOATING
C11862 S.t1676 VSUBS 0.02fF
C11863 S.n10766 VSUBS 0.24fF $ **FLOATING
C11864 S.n10767 VSUBS 0.91fF $ **FLOATING
C11865 S.n10768 VSUBS 0.05fF $ **FLOATING
C11866 S.t1445 VSUBS 0.02fF
C11867 S.n10769 VSUBS 0.12fF $ **FLOATING
C11868 S.n10770 VSUBS 0.14fF $ **FLOATING
C11869 S.n10772 VSUBS 1.89fF $ **FLOATING
C11870 S.n10773 VSUBS 1.88fF $ **FLOATING
C11871 S.t2302 VSUBS 0.02fF
C11872 S.n10774 VSUBS 0.24fF $ **FLOATING
C11873 S.n10775 VSUBS 0.36fF $ **FLOATING
C11874 S.n10776 VSUBS 0.61fF $ **FLOATING
C11875 S.n10777 VSUBS 0.12fF $ **FLOATING
C11876 S.t1489 VSUBS 0.02fF
C11877 S.n10778 VSUBS 0.14fF $ **FLOATING
C11878 S.n10780 VSUBS 1.16fF $ **FLOATING
C11879 S.n10781 VSUBS 0.22fF $ **FLOATING
C11880 S.n10782 VSUBS 0.25fF $ **FLOATING
C11881 S.n10783 VSUBS 0.09fF $ **FLOATING
C11882 S.n10784 VSUBS 1.88fF $ **FLOATING
C11883 S.t18 VSUBS 0.02fF
C11884 S.n10785 VSUBS 0.24fF $ **FLOATING
C11885 S.n10786 VSUBS 0.91fF $ **FLOATING
C11886 S.n10787 VSUBS 0.05fF $ **FLOATING
C11887 S.t2353 VSUBS 0.02fF
C11888 S.n10788 VSUBS 0.12fF $ **FLOATING
C11889 S.n10789 VSUBS 0.14fF $ **FLOATING
C11890 S.n10791 VSUBS 20.78fF $ **FLOATING
C11891 S.n10792 VSUBS 1.88fF $ **FLOATING
C11892 S.n10793 VSUBS 2.67fF $ **FLOATING
C11893 S.t971 VSUBS 0.02fF
C11894 S.n10794 VSUBS 0.24fF $ **FLOATING
C11895 S.n10795 VSUBS 0.36fF $ **FLOATING
C11896 S.n10796 VSUBS 0.61fF $ **FLOATING
C11897 S.n10797 VSUBS 0.12fF $ **FLOATING
C11898 S.t145 VSUBS 0.02fF
C11899 S.n10798 VSUBS 0.14fF $ **FLOATING
C11900 S.n10800 VSUBS 2.80fF $ **FLOATING
C11901 S.n10801 VSUBS 2.30fF $ **FLOATING
C11902 S.t1026 VSUBS 0.02fF
C11903 S.n10802 VSUBS 0.12fF $ **FLOATING
C11904 S.n10803 VSUBS 0.14fF $ **FLOATING
C11905 S.t1260 VSUBS 0.02fF
C11906 S.n10805 VSUBS 0.24fF $ **FLOATING
C11907 S.n10806 VSUBS 0.91fF $ **FLOATING
C11908 S.n10807 VSUBS 0.05fF $ **FLOATING
C11909 S.n10808 VSUBS 2.80fF $ **FLOATING
C11910 S.n10809 VSUBS 1.88fF $ **FLOATING
C11911 S.n10810 VSUBS 0.12fF $ **FLOATING
C11912 S.t1072 VSUBS 0.02fF
C11913 S.n10811 VSUBS 0.14fF $ **FLOATING
C11914 S.t1751 VSUBS 0.02fF
C11915 S.n10813 VSUBS 0.24fF $ **FLOATING
C11916 S.n10814 VSUBS 0.36fF $ **FLOATING
C11917 S.n10815 VSUBS 0.61fF $ **FLOATING
C11918 S.n10816 VSUBS 2.67fF $ **FLOATING
C11919 S.n10817 VSUBS 2.30fF $ **FLOATING
C11920 S.t1807 VSUBS 0.02fF
C11921 S.n10818 VSUBS 0.12fF $ **FLOATING
C11922 S.n10819 VSUBS 0.14fF $ **FLOATING
C11923 S.t2047 VSUBS 0.02fF
C11924 S.n10821 VSUBS 0.24fF $ **FLOATING
C11925 S.n10822 VSUBS 0.91fF $ **FLOATING
C11926 S.n10823 VSUBS 0.05fF $ **FLOATING
C11927 S.n10824 VSUBS 1.88fF $ **FLOATING
C11928 S.n10825 VSUBS 2.67fF $ **FLOATING
C11929 S.t1490 VSUBS 0.02fF
C11930 S.n10826 VSUBS 0.24fF $ **FLOATING
C11931 S.n10827 VSUBS 0.36fF $ **FLOATING
C11932 S.n10828 VSUBS 0.61fF $ **FLOATING
C11933 S.n10829 VSUBS 0.12fF $ **FLOATING
C11934 S.t669 VSUBS 0.02fF
C11935 S.n10830 VSUBS 0.14fF $ **FLOATING
C11936 S.n10832 VSUBS 2.80fF $ **FLOATING
C11937 S.n10833 VSUBS 2.30fF $ **FLOATING
C11938 S.t199 VSUBS 0.02fF
C11939 S.n10834 VSUBS 0.12fF $ **FLOATING
C11940 S.n10835 VSUBS 0.14fF $ **FLOATING
C11941 S.t1778 VSUBS 0.02fF
C11942 S.n10837 VSUBS 0.24fF $ **FLOATING
C11943 S.n10838 VSUBS 0.91fF $ **FLOATING
C11944 S.n10839 VSUBS 0.05fF $ **FLOATING
C11945 S.n10840 VSUBS 1.88fF $ **FLOATING
C11946 S.n10841 VSUBS 2.67fF $ **FLOATING
C11947 S.t2272 VSUBS 0.02fF
C11948 S.n10842 VSUBS 0.24fF $ **FLOATING
C11949 S.n10843 VSUBS 0.36fF $ **FLOATING
C11950 S.n10844 VSUBS 0.61fF $ **FLOATING
C11951 S.n10845 VSUBS 0.12fF $ **FLOATING
C11952 S.t1456 VSUBS 0.02fF
C11953 S.n10846 VSUBS 0.14fF $ **FLOATING
C11954 S.n10848 VSUBS 2.80fF $ **FLOATING
C11955 S.n10849 VSUBS 2.30fF $ **FLOATING
C11956 S.t2325 VSUBS 0.02fF
C11957 S.n10850 VSUBS 0.12fF $ **FLOATING
C11958 S.n10851 VSUBS 0.14fF $ **FLOATING
C11959 S.t2559 VSUBS 0.02fF
C11960 S.n10853 VSUBS 0.24fF $ **FLOATING
C11961 S.n10854 VSUBS 0.91fF $ **FLOATING
C11962 S.n10855 VSUBS 0.05fF $ **FLOATING
C11963 S.n10856 VSUBS 1.88fF $ **FLOATING
C11964 S.n10857 VSUBS 2.67fF $ **FLOATING
C11965 S.t545 VSUBS 0.02fF
C11966 S.n10858 VSUBS 0.24fF $ **FLOATING
C11967 S.n10859 VSUBS 0.36fF $ **FLOATING
C11968 S.n10860 VSUBS 0.61fF $ **FLOATING
C11969 S.n10861 VSUBS 0.12fF $ **FLOATING
C11970 S.t2244 VSUBS 0.02fF
C11971 S.n10862 VSUBS 0.14fF $ **FLOATING
C11972 S.n10864 VSUBS 2.80fF $ **FLOATING
C11973 S.n10865 VSUBS 2.30fF $ **FLOATING
C11974 S.t589 VSUBS 0.02fF
C11975 S.n10866 VSUBS 0.12fF $ **FLOATING
C11976 S.n10867 VSUBS 0.14fF $ **FLOATING
C11977 S.t823 VSUBS 0.02fF
C11978 S.n10869 VSUBS 0.24fF $ **FLOATING
C11979 S.n10870 VSUBS 0.91fF $ **FLOATING
C11980 S.n10871 VSUBS 0.05fF $ **FLOATING
C11981 S.n10872 VSUBS 1.88fF $ **FLOATING
C11982 S.n10873 VSUBS 2.67fF $ **FLOATING
C11983 S.t1331 VSUBS 0.02fF
C11984 S.n10874 VSUBS 0.24fF $ **FLOATING
C11985 S.n10875 VSUBS 0.36fF $ **FLOATING
C11986 S.n10876 VSUBS 0.61fF $ **FLOATING
C11987 S.n10877 VSUBS 0.12fF $ **FLOATING
C11988 S.t513 VSUBS 0.02fF
C11989 S.n10878 VSUBS 0.14fF $ **FLOATING
C11990 S.n10880 VSUBS 2.80fF $ **FLOATING
C11991 S.n10881 VSUBS 2.30fF $ **FLOATING
C11992 S.t1380 VSUBS 0.02fF
C11993 S.n10882 VSUBS 0.12fF $ **FLOATING
C11994 S.n10883 VSUBS 0.14fF $ **FLOATING
C11995 S.t1605 VSUBS 0.02fF
C11996 S.n10885 VSUBS 0.24fF $ **FLOATING
C11997 S.n10886 VSUBS 0.91fF $ **FLOATING
C11998 S.n10887 VSUBS 0.05fF $ **FLOATING
C11999 S.n10888 VSUBS 1.88fF $ **FLOATING
C12000 S.n10889 VSUBS 2.67fF $ **FLOATING
C12001 S.t2120 VSUBS 0.02fF
C12002 S.n10890 VSUBS 0.24fF $ **FLOATING
C12003 S.n10891 VSUBS 0.36fF $ **FLOATING
C12004 S.n10892 VSUBS 0.61fF $ **FLOATING
C12005 S.n10893 VSUBS 0.12fF $ **FLOATING
C12006 S.t1423 VSUBS 0.02fF
C12007 S.n10894 VSUBS 0.14fF $ **FLOATING
C12008 S.n10896 VSUBS 2.80fF $ **FLOATING
C12009 S.n10897 VSUBS 2.30fF $ **FLOATING
C12010 S.t2166 VSUBS 0.02fF
C12011 S.n10898 VSUBS 0.12fF $ **FLOATING
C12012 S.n10899 VSUBS 0.14fF $ **FLOATING
C12013 S.t2395 VSUBS 0.02fF
C12014 S.n10901 VSUBS 0.24fF $ **FLOATING
C12015 S.n10902 VSUBS 0.91fF $ **FLOATING
C12016 S.n10903 VSUBS 0.05fF $ **FLOATING
C12017 S.n10904 VSUBS 1.88fF $ **FLOATING
C12018 S.n10905 VSUBS 2.67fF $ **FLOATING
C12019 S.t1804 VSUBS 0.02fF
C12020 S.n10906 VSUBS 0.24fF $ **FLOATING
C12021 S.n10907 VSUBS 0.36fF $ **FLOATING
C12022 S.n10908 VSUBS 0.61fF $ **FLOATING
C12023 S.n10909 VSUBS 0.12fF $ **FLOATING
C12024 S.t2009 VSUBS 0.02fF
C12025 S.n10910 VSUBS 0.14fF $ **FLOATING
C12026 S.n10912 VSUBS 2.80fF $ **FLOATING
C12027 S.n10913 VSUBS 2.30fF $ **FLOATING
C12028 S.t363 VSUBS 0.02fF
C12029 S.n10914 VSUBS 0.12fF $ **FLOATING
C12030 S.n10915 VSUBS 0.14fF $ **FLOATING
C12031 S.t105 VSUBS 0.02fF
C12032 S.n10917 VSUBS 0.24fF $ **FLOATING
C12033 S.n10918 VSUBS 0.91fF $ **FLOATING
C12034 S.n10919 VSUBS 0.05fF $ **FLOATING
C12035 S.n10920 VSUBS 1.88fF $ **FLOATING
C12036 S.n10921 VSUBS 2.67fF $ **FLOATING
C12037 S.t16 VSUBS 0.02fF
C12038 S.n10922 VSUBS 0.24fF $ **FLOATING
C12039 S.n10923 VSUBS 0.36fF $ **FLOATING
C12040 S.n10924 VSUBS 0.61fF $ **FLOATING
C12041 S.n10925 VSUBS 0.12fF $ **FLOATING
C12042 S.t283 VSUBS 0.02fF
C12043 S.n10926 VSUBS 0.14fF $ **FLOATING
C12044 S.n10928 VSUBS 2.80fF $ **FLOATING
C12045 S.n10929 VSUBS 2.30fF $ **FLOATING
C12046 S.t1149 VSUBS 0.02fF
C12047 S.n10930 VSUBS 0.12fF $ **FLOATING
C12048 S.n10931 VSUBS 0.14fF $ **FLOATING
C12049 S.t912 VSUBS 0.02fF
C12050 S.n10933 VSUBS 0.24fF $ **FLOATING
C12051 S.n10934 VSUBS 0.91fF $ **FLOATING
C12052 S.n10935 VSUBS 0.05fF $ **FLOATING
C12053 S.n10936 VSUBS 1.88fF $ **FLOATING
C12054 S.n10937 VSUBS 2.67fF $ **FLOATING
C12055 S.t854 VSUBS 0.02fF
C12056 S.n10938 VSUBS 0.24fF $ **FLOATING
C12057 S.n10939 VSUBS 0.36fF $ **FLOATING
C12058 S.n10940 VSUBS 0.61fF $ **FLOATING
C12059 S.n10941 VSUBS 0.12fF $ **FLOATING
C12060 S.t1064 VSUBS 0.02fF
C12061 S.n10942 VSUBS 0.14fF $ **FLOATING
C12062 S.n10944 VSUBS 2.80fF $ **FLOATING
C12063 S.n10945 VSUBS 2.30fF $ **FLOATING
C12064 S.t1932 VSUBS 0.02fF
C12065 S.n10946 VSUBS 0.12fF $ **FLOATING
C12066 S.n10947 VSUBS 0.14fF $ **FLOATING
C12067 S.t1692 VSUBS 0.02fF
C12068 S.n10949 VSUBS 0.24fF $ **FLOATING
C12069 S.n10950 VSUBS 0.91fF $ **FLOATING
C12070 S.n10951 VSUBS 0.05fF $ **FLOATING
C12071 S.n10952 VSUBS 2.73fF $ **FLOATING
C12072 S.n10953 VSUBS 1.59fF $ **FLOATING
C12073 S.n10954 VSUBS 0.12fF $ **FLOATING
C12074 S.t874 VSUBS 0.02fF
C12075 S.n10955 VSUBS 0.14fF $ **FLOATING
C12076 S.t800 VSUBS 0.02fF
C12077 S.n10957 VSUBS 0.24fF $ **FLOATING
C12078 S.n10958 VSUBS 0.36fF $ **FLOATING
C12079 S.n10959 VSUBS 0.61fF $ **FLOATING
C12080 S.n10960 VSUBS 0.07fF $ **FLOATING
C12081 S.n10961 VSUBS 0.01fF $ **FLOATING
C12082 S.n10962 VSUBS 0.24fF $ **FLOATING
C12083 S.n10963 VSUBS 1.16fF $ **FLOATING
C12084 S.n10964 VSUBS 1.35fF $ **FLOATING
C12085 S.n10965 VSUBS 2.30fF $ **FLOATING
C12086 S.t978 VSUBS 0.02fF
C12087 S.n10966 VSUBS 0.12fF $ **FLOATING
C12088 S.n10967 VSUBS 0.14fF $ **FLOATING
C12089 S.t2210 VSUBS 0.02fF
C12090 S.n10969 VSUBS 0.24fF $ **FLOATING
C12091 S.n10970 VSUBS 0.91fF $ **FLOATING
C12092 S.n10971 VSUBS 0.05fF $ **FLOATING
C12093 S.t144 VSUBS 48.27fF
C12094 S.t2482 VSUBS 0.02fF
C12095 S.n10972 VSUBS 0.24fF $ **FLOATING
C12096 S.n10973 VSUBS 0.91fF $ **FLOATING
C12097 S.n10974 VSUBS 0.05fF $ **FLOATING
C12098 S.t190 VSUBS 0.02fF
C12099 S.n10975 VSUBS 0.12fF $ **FLOATING
C12100 S.n10976 VSUBS 0.14fF $ **FLOATING
C12101 S.n10978 VSUBS 0.12fF $ **FLOATING
C12102 S.t1849 VSUBS 0.02fF
C12103 S.n10979 VSUBS 0.14fF $ **FLOATING
C12104 S.n10981 VSUBS 5.17fF $ **FLOATING
C12105 S.n10982 VSUBS 5.44fF $ **FLOATING
C12106 S.t156 VSUBS 0.02fF
C12107 S.n10983 VSUBS 0.12fF $ **FLOATING
C12108 S.n10984 VSUBS 0.14fF $ **FLOATING
C12109 S.t2454 VSUBS 0.02fF
C12110 S.n10986 VSUBS 0.24fF $ **FLOATING
C12111 S.n10987 VSUBS 0.91fF $ **FLOATING
C12112 S.n10988 VSUBS 0.05fF $ **FLOATING
C12113 S.t35 VSUBS 47.89fF
C12114 S.t2243 VSUBS 0.02fF
C12115 S.n10989 VSUBS 0.01fF $ **FLOATING
C12116 S.n10990 VSUBS 0.26fF $ **FLOATING
C12117 S.t409 VSUBS 0.02fF
C12118 S.n10992 VSUBS 1.19fF $ **FLOATING
C12119 S.n10993 VSUBS 0.05fF $ **FLOATING
C12120 S.t92 VSUBS 0.02fF
C12121 S.n10994 VSUBS 0.64fF $ **FLOATING
C12122 S.n10995 VSUBS 0.61fF $ **FLOATING
C12123 S.n10996 VSUBS 0.60fF $ **FLOATING
C12124 S.n10997 VSUBS 0.22fF $ **FLOATING
C12125 S.n10998 VSUBS 0.59fF $ **FLOATING
C12126 S.n10999 VSUBS 3.39fF $ **FLOATING
C12127 S.n11000 VSUBS 0.29fF $ **FLOATING
C12128 S.t17 VSUBS 21.42fF
C12129 S.n11001 VSUBS 21.71fF $ **FLOATING
C12130 S.n11002 VSUBS 0.77fF $ **FLOATING
C12131 S.n11003 VSUBS 0.28fF $ **FLOATING
C12132 S.n11004 VSUBS 4.00fF $ **FLOATING
C12133 S.n11005 VSUBS 1.35fF $ **FLOATING
C12134 S.n11006 VSUBS 0.01fF $ **FLOATING
C12135 S.n11007 VSUBS 0.02fF $ **FLOATING
C12136 S.n11008 VSUBS 0.03fF $ **FLOATING
C12137 S.n11009 VSUBS 0.04fF $ **FLOATING
C12138 S.n11010 VSUBS 0.17fF $ **FLOATING
C12139 S.n11011 VSUBS 0.01fF $ **FLOATING
C12140 S.n11012 VSUBS 0.02fF $ **FLOATING
C12141 S.n11013 VSUBS 0.01fF $ **FLOATING
C12142 S.n11014 VSUBS 0.01fF $ **FLOATING
C12143 S.n11015 VSUBS 0.01fF $ **FLOATING
C12144 S.n11016 VSUBS 0.01fF $ **FLOATING
C12145 S.n11017 VSUBS 0.02fF $ **FLOATING
C12146 S.n11018 VSUBS 0.01fF $ **FLOATING
C12147 S.n11019 VSUBS 0.02fF $ **FLOATING
C12148 S.n11020 VSUBS 0.05fF $ **FLOATING
C12149 S.n11021 VSUBS 0.04fF $ **FLOATING
C12150 S.n11022 VSUBS 0.11fF $ **FLOATING
C12151 S.n11023 VSUBS 0.38fF $ **FLOATING
C12152 S.n11024 VSUBS 0.20fF $ **FLOATING
C12153 S.n11025 VSUBS 4.39fF $ **FLOATING
C12154 S.n11026 VSUBS 0.24fF $ **FLOATING
C12155 S.n11027 VSUBS 1.50fF $ **FLOATING
C12156 S.n11028 VSUBS 1.26fF $ **FLOATING
C12157 S.n11029 VSUBS 0.28fF $ **FLOATING
C12158 S.n11030 VSUBS 0.25fF $ **FLOATING
C12159 S.n11031 VSUBS 0.09fF $ **FLOATING
C12160 S.n11032 VSUBS 0.21fF $ **FLOATING
C12161 S.n11033 VSUBS 1.28fF $ **FLOATING
C12162 S.n11034 VSUBS 0.53fF $ **FLOATING
C12163 S.n11035 VSUBS 1.88fF $ **FLOATING
C12164 S.n11036 VSUBS 0.12fF $ **FLOATING
C12165 S.t1169 VSUBS 0.02fF
C12166 S.n11037 VSUBS 0.14fF $ **FLOATING
C12167 S.t1983 VSUBS 0.02fF
C12168 S.n11039 VSUBS 0.24fF $ **FLOATING
C12169 S.n11040 VSUBS 0.36fF $ **FLOATING
C12170 S.n11041 VSUBS 0.61fF $ **FLOATING
C12171 S.n11042 VSUBS 1.58fF $ **FLOATING
C12172 S.n11043 VSUBS 2.45fF $ **FLOATING
C12173 S.t2259 VSUBS 0.02fF
C12174 S.n11044 VSUBS 0.24fF $ **FLOATING
C12175 S.n11045 VSUBS 0.91fF $ **FLOATING
C12176 S.n11046 VSUBS 0.05fF $ **FLOATING
C12177 S.t2032 VSUBS 0.02fF
C12178 S.n11047 VSUBS 0.12fF $ **FLOATING
C12179 S.n11048 VSUBS 0.14fF $ **FLOATING
C12180 S.n11050 VSUBS 1.89fF $ **FLOATING
C12181 S.n11051 VSUBS 0.06fF $ **FLOATING
C12182 S.n11052 VSUBS 0.03fF $ **FLOATING
C12183 S.n11053 VSUBS 0.04fF $ **FLOATING
C12184 S.n11054 VSUBS 0.99fF $ **FLOATING
C12185 S.n11055 VSUBS 0.02fF $ **FLOATING
C12186 S.n11056 VSUBS 0.01fF $ **FLOATING
C12187 S.n11057 VSUBS 0.02fF $ **FLOATING
C12188 S.n11058 VSUBS 0.08fF $ **FLOATING
C12189 S.n11059 VSUBS 0.36fF $ **FLOATING
C12190 S.n11060 VSUBS 1.85fF $ **FLOATING
C12191 S.t377 VSUBS 0.02fF
C12192 S.n11061 VSUBS 0.24fF $ **FLOATING
C12193 S.n11062 VSUBS 0.36fF $ **FLOATING
C12194 S.n11063 VSUBS 0.61fF $ **FLOATING
C12195 S.n11064 VSUBS 0.12fF $ **FLOATING
C12196 S.t2080 VSUBS 0.02fF
C12197 S.n11065 VSUBS 0.14fF $ **FLOATING
C12198 S.n11067 VSUBS 0.70fF $ **FLOATING
C12199 S.n11068 VSUBS 0.23fF $ **FLOATING
C12200 S.n11069 VSUBS 0.23fF $ **FLOATING
C12201 S.n11070 VSUBS 0.70fF $ **FLOATING
C12202 S.n11071 VSUBS 1.16fF $ **FLOATING
C12203 S.n11072 VSUBS 0.22fF $ **FLOATING
C12204 S.n11073 VSUBS 0.25fF $ **FLOATING
C12205 S.n11074 VSUBS 0.09fF $ **FLOATING
C12206 S.n11075 VSUBS 1.88fF $ **FLOATING
C12207 S.t646 VSUBS 0.02fF
C12208 S.n11076 VSUBS 0.24fF $ **FLOATING
C12209 S.n11077 VSUBS 0.91fF $ **FLOATING
C12210 S.n11078 VSUBS 0.05fF $ **FLOATING
C12211 S.t426 VSUBS 0.02fF
C12212 S.n11079 VSUBS 0.12fF $ **FLOATING
C12213 S.n11080 VSUBS 0.14fF $ **FLOATING
C12214 S.n11082 VSUBS 20.78fF $ **FLOATING
C12215 S.n11083 VSUBS 2.39fF $ **FLOATING
C12216 S.n11084 VSUBS 0.46fF $ **FLOATING
C12217 S.n11085 VSUBS 0.22fF $ **FLOATING
C12218 S.n11086 VSUBS 0.38fF $ **FLOATING
C12219 S.n11087 VSUBS 0.16fF $ **FLOATING
C12220 S.n11088 VSUBS 0.28fF $ **FLOATING
C12221 S.n11089 VSUBS 0.21fF $ **FLOATING
C12222 S.n11090 VSUBS 0.30fF $ **FLOATING
C12223 S.n11091 VSUBS 0.21fF $ **FLOATING
C12224 S.t1203 VSUBS 0.02fF
C12225 S.n11092 VSUBS 0.24fF $ **FLOATING
C12226 S.n11093 VSUBS 0.36fF $ **FLOATING
C12227 S.n11094 VSUBS 0.61fF $ **FLOATING
C12228 S.n11095 VSUBS 0.12fF $ **FLOATING
C12229 S.t383 VSUBS 0.02fF
C12230 S.n11096 VSUBS 0.14fF $ **FLOATING
C12231 S.n11098 VSUBS 0.19fF $ **FLOATING
C12232 S.n11099 VSUBS 1.57fF $ **FLOATING
C12233 S.n11100 VSUBS 2.21fF $ **FLOATING
C12234 S.n11101 VSUBS 0.32fF $ **FLOATING
C12235 S.n11102 VSUBS 2.39fF $ **FLOATING
C12236 S.t1249 VSUBS 0.02fF
C12237 S.n11103 VSUBS 0.12fF $ **FLOATING
C12238 S.n11104 VSUBS 0.14fF $ **FLOATING
C12239 S.t1472 VSUBS 0.02fF
C12240 S.n11106 VSUBS 0.24fF $ **FLOATING
C12241 S.n11107 VSUBS 0.91fF $ **FLOATING
C12242 S.n11108 VSUBS 0.05fF $ **FLOATING
C12243 S.n11109 VSUBS 1.88fF $ **FLOATING
C12244 S.n11110 VSUBS 0.12fF $ **FLOATING
C12245 S.t922 VSUBS 0.02fF
C12246 S.n11111 VSUBS 0.14fF $ **FLOATING
C12247 S.t1788 VSUBS 0.02fF
C12248 S.n11113 VSUBS 0.12fF $ **FLOATING
C12249 S.n11114 VSUBS 0.14fF $ **FLOATING
C12250 S.t2026 VSUBS 0.02fF
C12251 S.n11116 VSUBS 0.24fF $ **FLOATING
C12252 S.n11117 VSUBS 0.91fF $ **FLOATING
C12253 S.n11118 VSUBS 0.05fF $ **FLOATING
C12254 S.t1733 VSUBS 0.02fF
C12255 S.n11119 VSUBS 0.24fF $ **FLOATING
C12256 S.n11120 VSUBS 0.36fF $ **FLOATING
C12257 S.n11121 VSUBS 0.61fF $ **FLOATING
C12258 S.n11122 VSUBS 0.32fF $ **FLOATING
C12259 S.n11123 VSUBS 1.09fF $ **FLOATING
C12260 S.n11124 VSUBS 0.15fF $ **FLOATING
C12261 S.n11125 VSUBS 2.10fF $ **FLOATING
C12262 S.n11126 VSUBS 2.94fF $ **FLOATING
C12263 S.n11127 VSUBS 1.88fF $ **FLOATING
C12264 S.n11128 VSUBS 0.12fF $ **FLOATING
C12265 S.t1678 VSUBS 0.02fF
C12266 S.n11129 VSUBS 0.14fF $ **FLOATING
C12267 S.t2495 VSUBS 0.02fF
C12268 S.n11131 VSUBS 0.24fF $ **FLOATING
C12269 S.n11132 VSUBS 0.36fF $ **FLOATING
C12270 S.n11133 VSUBS 0.61fF $ **FLOATING
C12271 S.n11134 VSUBS 0.92fF $ **FLOATING
C12272 S.n11135 VSUBS 0.32fF $ **FLOATING
C12273 S.n11136 VSUBS 0.92fF $ **FLOATING
C12274 S.n11137 VSUBS 1.09fF $ **FLOATING
C12275 S.n11138 VSUBS 0.15fF $ **FLOATING
C12276 S.n11139 VSUBS 4.96fF $ **FLOATING
C12277 S.t1221 VSUBS 0.02fF
C12278 S.n11140 VSUBS 0.12fF $ **FLOATING
C12279 S.n11141 VSUBS 0.14fF $ **FLOATING
C12280 S.t276 VSUBS 0.02fF
C12281 S.n11143 VSUBS 0.24fF $ **FLOATING
C12282 S.n11144 VSUBS 0.91fF $ **FLOATING
C12283 S.n11145 VSUBS 0.05fF $ **FLOATING
C12284 S.n11146 VSUBS 1.88fF $ **FLOATING
C12285 S.n11147 VSUBS 2.67fF $ **FLOATING
C12286 S.t751 VSUBS 0.02fF
C12287 S.n11148 VSUBS 0.24fF $ **FLOATING
C12288 S.n11149 VSUBS 0.36fF $ **FLOATING
C12289 S.n11150 VSUBS 0.61fF $ **FLOATING
C12290 S.n11151 VSUBS 0.12fF $ **FLOATING
C12291 S.t2463 VSUBS 0.02fF
C12292 S.n11152 VSUBS 0.14fF $ **FLOATING
C12293 S.n11154 VSUBS 1.88fF $ **FLOATING
C12294 S.n11155 VSUBS 2.67fF $ **FLOATING
C12295 S.t1349 VSUBS 0.02fF
C12296 S.n11156 VSUBS 0.24fF $ **FLOATING
C12297 S.n11157 VSUBS 0.36fF $ **FLOATING
C12298 S.n11158 VSUBS 0.61fF $ **FLOATING
C12299 S.t1623 VSUBS 0.02fF
C12300 S.n11159 VSUBS 0.24fF $ **FLOATING
C12301 S.n11160 VSUBS 0.91fF $ **FLOATING
C12302 S.n11161 VSUBS 0.05fF $ **FLOATING
C12303 S.t1401 VSUBS 0.02fF
C12304 S.n11162 VSUBS 0.12fF $ **FLOATING
C12305 S.n11163 VSUBS 0.14fF $ **FLOATING
C12306 S.n11165 VSUBS 0.12fF $ **FLOATING
C12307 S.t534 VSUBS 0.02fF
C12308 S.n11166 VSUBS 0.14fF $ **FLOATING
C12309 S.n11168 VSUBS 2.30fF $ **FLOATING
C12310 S.n11169 VSUBS 2.94fF $ **FLOATING
C12311 S.n11170 VSUBS 5.16fF $ **FLOATING
C12312 S.t811 VSUBS 0.02fF
C12313 S.n11171 VSUBS 0.12fF $ **FLOATING
C12314 S.n11172 VSUBS 0.14fF $ **FLOATING
C12315 S.t1056 VSUBS 0.02fF
C12316 S.n11174 VSUBS 0.24fF $ **FLOATING
C12317 S.n11175 VSUBS 0.91fF $ **FLOATING
C12318 S.n11176 VSUBS 0.05fF $ **FLOATING
C12319 S.n11177 VSUBS 1.88fF $ **FLOATING
C12320 S.n11178 VSUBS 2.67fF $ **FLOATING
C12321 S.t1541 VSUBS 0.02fF
C12322 S.n11179 VSUBS 0.24fF $ **FLOATING
C12323 S.n11180 VSUBS 0.36fF $ **FLOATING
C12324 S.n11181 VSUBS 0.61fF $ **FLOATING
C12325 S.n11182 VSUBS 0.12fF $ **FLOATING
C12326 S.t721 VSUBS 0.02fF
C12327 S.n11183 VSUBS 0.14fF $ **FLOATING
C12328 S.n11185 VSUBS 5.17fF $ **FLOATING
C12329 S.t1590 VSUBS 0.02fF
C12330 S.n11186 VSUBS 0.12fF $ **FLOATING
C12331 S.n11187 VSUBS 0.14fF $ **FLOATING
C12332 S.t1841 VSUBS 0.02fF
C12333 S.n11189 VSUBS 0.24fF $ **FLOATING
C12334 S.n11190 VSUBS 0.91fF $ **FLOATING
C12335 S.n11191 VSUBS 0.05fF $ **FLOATING
C12336 S.n11192 VSUBS 1.88fF $ **FLOATING
C12337 S.n11193 VSUBS 0.12fF $ **FLOATING
C12338 S.t1514 VSUBS 0.02fF
C12339 S.n11194 VSUBS 0.14fF $ **FLOATING
C12340 S.t2332 VSUBS 0.02fF
C12341 S.n11196 VSUBS 0.24fF $ **FLOATING
C12342 S.n11197 VSUBS 0.36fF $ **FLOATING
C12343 S.n11198 VSUBS 0.61fF $ **FLOATING
C12344 S.n11199 VSUBS 2.67fF $ **FLOATING
C12345 S.n11200 VSUBS 5.17fF $ **FLOATING
C12346 S.t2381 VSUBS 0.02fF
C12347 S.n11201 VSUBS 0.12fF $ **FLOATING
C12348 S.n11202 VSUBS 0.14fF $ **FLOATING
C12349 S.t71 VSUBS 0.02fF
C12350 S.n11204 VSUBS 0.24fF $ **FLOATING
C12351 S.n11205 VSUBS 0.91fF $ **FLOATING
C12352 S.n11206 VSUBS 0.05fF $ **FLOATING
C12353 S.n11207 VSUBS 1.88fF $ **FLOATING
C12354 S.n11208 VSUBS 2.67fF $ **FLOATING
C12355 S.t714 VSUBS 0.02fF
C12356 S.n11209 VSUBS 0.24fF $ **FLOATING
C12357 S.n11210 VSUBS 0.36fF $ **FLOATING
C12358 S.n11211 VSUBS 0.61fF $ **FLOATING
C12359 S.n11212 VSUBS 0.12fF $ **FLOATING
C12360 S.t2428 VSUBS 0.02fF
C12361 S.n11213 VSUBS 0.14fF $ **FLOATING
C12362 S.n11215 VSUBS 5.17fF $ **FLOATING
C12363 S.t770 VSUBS 0.02fF
C12364 S.n11216 VSUBS 0.12fF $ **FLOATING
C12365 S.n11217 VSUBS 0.14fF $ **FLOATING
C12366 S.t1019 VSUBS 0.02fF
C12367 S.n11219 VSUBS 0.24fF $ **FLOATING
C12368 S.n11220 VSUBS 0.91fF $ **FLOATING
C12369 S.n11221 VSUBS 0.05fF $ **FLOATING
C12370 S.n11222 VSUBS 1.88fF $ **FLOATING
C12371 S.n11223 VSUBS 2.67fF $ **FLOATING
C12372 S.t352 VSUBS 0.02fF
C12373 S.n11224 VSUBS 0.24fF $ **FLOATING
C12374 S.n11225 VSUBS 0.36fF $ **FLOATING
C12375 S.n11226 VSUBS 0.61fF $ **FLOATING
C12376 S.n11227 VSUBS 0.12fF $ **FLOATING
C12377 S.t2052 VSUBS 0.02fF
C12378 S.n11228 VSUBS 0.14fF $ **FLOATING
C12379 S.n11230 VSUBS 5.17fF $ **FLOATING
C12380 S.t397 VSUBS 0.02fF
C12381 S.n11231 VSUBS 0.12fF $ **FLOATING
C12382 S.n11232 VSUBS 0.14fF $ **FLOATING
C12383 S.t620 VSUBS 0.02fF
C12384 S.n11234 VSUBS 0.24fF $ **FLOATING
C12385 S.n11235 VSUBS 0.91fF $ **FLOATING
C12386 S.n11236 VSUBS 0.05fF $ **FLOATING
C12387 S.n11237 VSUBS 1.88fF $ **FLOATING
C12388 S.n11238 VSUBS 2.67fF $ **FLOATING
C12389 S.t1137 VSUBS 0.02fF
C12390 S.n11239 VSUBS 0.24fF $ **FLOATING
C12391 S.n11240 VSUBS 0.36fF $ **FLOATING
C12392 S.n11241 VSUBS 0.61fF $ **FLOATING
C12393 S.n11242 VSUBS 0.12fF $ **FLOATING
C12394 S.t317 VSUBS 0.02fF
C12395 S.n11243 VSUBS 0.14fF $ **FLOATING
C12396 S.n11245 VSUBS 5.17fF $ **FLOATING
C12397 S.t1188 VSUBS 0.02fF
C12398 S.n11246 VSUBS 0.12fF $ **FLOATING
C12399 S.n11247 VSUBS 0.14fF $ **FLOATING
C12400 S.t1410 VSUBS 0.02fF
C12401 S.n11249 VSUBS 0.24fF $ **FLOATING
C12402 S.n11250 VSUBS 0.91fF $ **FLOATING
C12403 S.n11251 VSUBS 0.05fF $ **FLOATING
C12404 S.n11252 VSUBS 1.88fF $ **FLOATING
C12405 S.n11253 VSUBS 2.67fF $ **FLOATING
C12406 S.t1921 VSUBS 0.02fF
C12407 S.n11254 VSUBS 0.24fF $ **FLOATING
C12408 S.n11255 VSUBS 0.36fF $ **FLOATING
C12409 S.n11256 VSUBS 0.61fF $ **FLOATING
C12410 S.n11257 VSUBS 0.12fF $ **FLOATING
C12411 S.t1107 VSUBS 0.02fF
C12412 S.n11258 VSUBS 0.14fF $ **FLOATING
C12413 S.n11260 VSUBS 5.17fF $ **FLOATING
C12414 S.t1970 VSUBS 0.02fF
C12415 S.n11261 VSUBS 0.12fF $ **FLOATING
C12416 S.n11262 VSUBS 0.14fF $ **FLOATING
C12417 S.t2198 VSUBS 0.02fF
C12418 S.n11264 VSUBS 0.24fF $ **FLOATING
C12419 S.n11265 VSUBS 0.91fF $ **FLOATING
C12420 S.n11266 VSUBS 0.05fF $ **FLOATING
C12421 S.n11267 VSUBS 1.88fF $ **FLOATING
C12422 S.n11268 VSUBS 2.67fF $ **FLOATING
C12423 S.t174 VSUBS 0.02fF
C12424 S.n11269 VSUBS 0.24fF $ **FLOATING
C12425 S.n11270 VSUBS 0.36fF $ **FLOATING
C12426 S.n11271 VSUBS 0.61fF $ **FLOATING
C12427 S.n11272 VSUBS 0.12fF $ **FLOATING
C12428 S.t1886 VSUBS 0.02fF
C12429 S.n11273 VSUBS 0.14fF $ **FLOATING
C12430 S.n11275 VSUBS 5.17fF $ **FLOATING
C12431 S.t232 VSUBS 0.02fF
C12432 S.n11276 VSUBS 0.12fF $ **FLOATING
C12433 S.n11277 VSUBS 0.14fF $ **FLOATING
C12434 S.t464 VSUBS 0.02fF
C12435 S.n11279 VSUBS 0.24fF $ **FLOATING
C12436 S.n11280 VSUBS 0.91fF $ **FLOATING
C12437 S.n11281 VSUBS 0.05fF $ **FLOATING
C12438 S.n11282 VSUBS 1.88fF $ **FLOATING
C12439 S.n11283 VSUBS 2.67fF $ **FLOATING
C12440 S.t1836 VSUBS 0.02fF
C12441 S.n11284 VSUBS 0.24fF $ **FLOATING
C12442 S.n11285 VSUBS 0.36fF $ **FLOATING
C12443 S.n11286 VSUBS 0.61fF $ **FLOATING
C12444 S.n11287 VSUBS 0.12fF $ **FLOATING
C12445 S.t2037 VSUBS 0.02fF
C12446 S.n11288 VSUBS 0.14fF $ **FLOATING
C12447 S.n11290 VSUBS 5.17fF $ **FLOATING
C12448 S.t1152 VSUBS 0.02fF
C12449 S.n11291 VSUBS 0.12fF $ **FLOATING
C12450 S.n11292 VSUBS 0.14fF $ **FLOATING
C12451 S.t142 VSUBS 0.02fF
C12452 S.n11294 VSUBS 0.24fF $ **FLOATING
C12453 S.n11295 VSUBS 0.91fF $ **FLOATING
C12454 S.n11296 VSUBS 0.05fF $ **FLOATING
C12455 S.n11297 VSUBS 1.88fF $ **FLOATING
C12456 S.n11298 VSUBS 2.67fF $ **FLOATING
C12457 S.t58 VSUBS 0.02fF
C12458 S.n11299 VSUBS 0.24fF $ **FLOATING
C12459 S.n11300 VSUBS 0.36fF $ **FLOATING
C12460 S.n11301 VSUBS 0.61fF $ **FLOATING
C12461 S.n11302 VSUBS 0.12fF $ **FLOATING
C12462 S.t306 VSUBS 0.02fF
C12463 S.n11303 VSUBS 0.14fF $ **FLOATING
C12464 S.n11305 VSUBS 5.17fF $ **FLOATING
C12465 S.t1174 VSUBS 0.02fF
C12466 S.n11306 VSUBS 0.12fF $ **FLOATING
C12467 S.n11307 VSUBS 0.14fF $ **FLOATING
C12468 S.t939 VSUBS 0.02fF
C12469 S.n11309 VSUBS 0.24fF $ **FLOATING
C12470 S.n11310 VSUBS 0.91fF $ **FLOATING
C12471 S.n11311 VSUBS 0.05fF $ **FLOATING
C12472 S.n11312 VSUBS 1.88fF $ **FLOATING
C12473 S.n11313 VSUBS 2.67fF $ **FLOATING
C12474 S.t877 VSUBS 0.02fF
C12475 S.n11314 VSUBS 0.24fF $ **FLOATING
C12476 S.n11315 VSUBS 0.36fF $ **FLOATING
C12477 S.n11316 VSUBS 0.61fF $ **FLOATING
C12478 S.n11317 VSUBS 0.12fF $ **FLOATING
C12479 S.t1089 VSUBS 0.02fF
C12480 S.n11318 VSUBS 0.14fF $ **FLOATING
C12481 S.n11320 VSUBS 5.17fF $ **FLOATING
C12482 S.t1958 VSUBS 0.02fF
C12483 S.n11321 VSUBS 0.12fF $ **FLOATING
C12484 S.n11322 VSUBS 0.14fF $ **FLOATING
C12485 S.t1720 VSUBS 0.02fF
C12486 S.n11324 VSUBS 0.24fF $ **FLOATING
C12487 S.n11325 VSUBS 0.91fF $ **FLOATING
C12488 S.n11326 VSUBS 0.05fF $ **FLOATING
C12489 S.n11327 VSUBS 1.88fF $ **FLOATING
C12490 S.n11328 VSUBS 2.67fF $ **FLOATING
C12491 S.t1659 VSUBS 0.02fF
C12492 S.n11329 VSUBS 0.24fF $ **FLOATING
C12493 S.n11330 VSUBS 0.36fF $ **FLOATING
C12494 S.n11331 VSUBS 0.61fF $ **FLOATING
C12495 S.n11332 VSUBS 0.12fF $ **FLOATING
C12496 S.t1871 VSUBS 0.02fF
C12497 S.n11333 VSUBS 0.14fF $ **FLOATING
C12498 S.n11335 VSUBS 4.89fF $ **FLOATING
C12499 S.t216 VSUBS 0.02fF
C12500 S.n11336 VSUBS 0.12fF $ **FLOATING
C12501 S.n11337 VSUBS 0.14fF $ **FLOATING
C12502 S.t2506 VSUBS 0.02fF
C12503 S.n11339 VSUBS 0.24fF $ **FLOATING
C12504 S.n11340 VSUBS 0.91fF $ **FLOATING
C12505 S.n11341 VSUBS 0.05fF $ **FLOATING
C12506 S.n11342 VSUBS 1.88fF $ **FLOATING
C12507 S.n11343 VSUBS 2.67fF $ **FLOATING
C12508 S.t2447 VSUBS 0.02fF
C12509 S.n11344 VSUBS 0.24fF $ **FLOATING
C12510 S.n11345 VSUBS 0.36fF $ **FLOATING
C12511 S.n11346 VSUBS 0.61fF $ **FLOATING
C12512 S.n11347 VSUBS 0.12fF $ **FLOATING
C12513 S.t116 VSUBS 0.02fF
C12514 S.n11348 VSUBS 0.14fF $ **FLOATING
C12515 S.n11350 VSUBS 1.88fF $ **FLOATING
C12516 S.n11351 VSUBS 2.68fF $ **FLOATING
C12517 S.t2474 VSUBS 0.02fF
C12518 S.n11352 VSUBS 0.24fF $ **FLOATING
C12519 S.n11353 VSUBS 0.36fF $ **FLOATING
C12520 S.n11354 VSUBS 0.61fF $ **FLOATING
C12521 S.t1772 VSUBS 0.02fF
C12522 S.n11355 VSUBS 1.22fF $ **FLOATING
C12523 S.n11356 VSUBS 0.42fF $ **FLOATING
C12524 S.n11357 VSUBS 0.44fF $ **FLOATING
C12525 S.n11358 VSUBS 0.36fF $ **FLOATING
C12526 S.n11359 VSUBS 0.21fF $ **FLOATING
C12527 S.n11360 VSUBS 0.25fF $ **FLOATING
C12528 S.n11361 VSUBS 1.28fF $ **FLOATING
C12529 S.n11362 VSUBS 2.00fF $ **FLOATING
C12530 S.n11363 VSUBS 4.08fF $ **FLOATING
C12531 S.n11364 VSUBS 0.25fF $ **FLOATING
C12532 S.n11365 VSUBS 0.01fF $ **FLOATING
C12533 S.t957 VSUBS 0.02fF
C12534 S.n11366 VSUBS 0.26fF $ **FLOATING
C12535 S.t2064 VSUBS 0.02fF
C12536 S.n11367 VSUBS 0.95fF $ **FLOATING
C12537 S.n11368 VSUBS 0.71fF $ **FLOATING
C12538 S.n11369 VSUBS 0.78fF $ **FLOATING
C12539 S.n11370 VSUBS 2.26fF $ **FLOATING
C12540 S.n11371 VSUBS 1.88fF $ **FLOATING
C12541 S.n11372 VSUBS 0.12fF $ **FLOATING
C12542 S.t1739 VSUBS 0.02fF
C12543 S.n11373 VSUBS 0.14fF $ **FLOATING
C12544 S.t2551 VSUBS 0.02fF
C12545 S.n11375 VSUBS 0.24fF $ **FLOATING
C12546 S.n11376 VSUBS 0.36fF $ **FLOATING
C12547 S.n11377 VSUBS 0.61fF $ **FLOATING
C12548 S.n11378 VSUBS 1.39fF $ **FLOATING
C12549 S.n11379 VSUBS 0.71fF $ **FLOATING
C12550 S.n11380 VSUBS 1.14fF $ **FLOATING
C12551 S.n11381 VSUBS 0.35fF $ **FLOATING
C12552 S.n11382 VSUBS 2.02fF $ **FLOATING
C12553 S.t330 VSUBS 0.02fF
C12554 S.n11383 VSUBS 0.24fF $ **FLOATING
C12555 S.n11384 VSUBS 0.91fF $ **FLOATING
C12556 S.n11385 VSUBS 0.05fF $ **FLOATING
C12557 S.t48 VSUBS 0.02fF
C12558 S.n11386 VSUBS 0.12fF $ **FLOATING
C12559 S.n11387 VSUBS 0.14fF $ **FLOATING
C12560 S.n11389 VSUBS 1.89fF $ **FLOATING
C12561 S.n11390 VSUBS 1.88fF $ **FLOATING
C12562 S.t817 VSUBS 0.02fF
C12563 S.n11391 VSUBS 0.24fF $ **FLOATING
C12564 S.n11392 VSUBS 0.36fF $ **FLOATING
C12565 S.n11393 VSUBS 0.61fF $ **FLOATING
C12566 S.n11394 VSUBS 0.12fF $ **FLOATING
C12567 S.t120 VSUBS 0.02fF
C12568 S.n11395 VSUBS 0.14fF $ **FLOATING
C12569 S.n11397 VSUBS 1.16fF $ **FLOATING
C12570 S.n11398 VSUBS 0.22fF $ **FLOATING
C12571 S.n11399 VSUBS 0.25fF $ **FLOATING
C12572 S.n11400 VSUBS 0.09fF $ **FLOATING
C12573 S.n11401 VSUBS 1.88fF $ **FLOATING
C12574 S.t1120 VSUBS 0.02fF
C12575 S.n11402 VSUBS 0.24fF $ **FLOATING
C12576 S.n11403 VSUBS 0.91fF $ **FLOATING
C12577 S.n11404 VSUBS 0.05fF $ **FLOATING
C12578 S.t869 VSUBS 0.02fF
C12579 S.n11405 VSUBS 0.12fF $ **FLOATING
C12580 S.n11406 VSUBS 0.14fF $ **FLOATING
C12581 S.n11408 VSUBS 1.88fF $ **FLOATING
C12582 S.n11409 VSUBS 2.67fF $ **FLOATING
C12583 S.t2135 VSUBS 0.02fF
C12584 S.n11410 VSUBS 0.24fF $ **FLOATING
C12585 S.n11411 VSUBS 0.36fF $ **FLOATING
C12586 S.n11412 VSUBS 0.61fF $ **FLOATING
C12587 S.n11413 VSUBS 0.12fF $ **FLOATING
C12588 S.t1319 VSUBS 0.02fF
C12589 S.n11414 VSUBS 0.14fF $ **FLOATING
C12590 S.n11416 VSUBS 2.80fF $ **FLOATING
C12591 S.n11417 VSUBS 2.30fF $ **FLOATING
C12592 S.t2188 VSUBS 0.02fF
C12593 S.n11418 VSUBS 0.12fF $ **FLOATING
C12594 S.n11419 VSUBS 0.14fF $ **FLOATING
C12595 S.t2410 VSUBS 0.02fF
C12596 S.n11421 VSUBS 0.24fF $ **FLOATING
C12597 S.n11422 VSUBS 0.91fF $ **FLOATING
C12598 S.n11423 VSUBS 0.05fF $ **FLOATING
C12599 S.n11424 VSUBS 2.80fF $ **FLOATING
C12600 S.n11425 VSUBS 1.88fF $ **FLOATING
C12601 S.n11426 VSUBS 0.12fF $ **FLOATING
C12602 S.t2106 VSUBS 0.02fF
C12603 S.n11427 VSUBS 0.14fF $ **FLOATING
C12604 S.t403 VSUBS 0.02fF
C12605 S.n11429 VSUBS 0.24fF $ **FLOATING
C12606 S.n11430 VSUBS 0.36fF $ **FLOATING
C12607 S.n11431 VSUBS 0.61fF $ **FLOATING
C12608 S.n11432 VSUBS 2.67fF $ **FLOATING
C12609 S.n11433 VSUBS 2.30fF $ **FLOATING
C12610 S.t452 VSUBS 0.02fF
C12611 S.n11434 VSUBS 0.12fF $ **FLOATING
C12612 S.n11435 VSUBS 0.14fF $ **FLOATING
C12613 S.t673 VSUBS 0.02fF
C12614 S.n11437 VSUBS 0.24fF $ **FLOATING
C12615 S.n11438 VSUBS 0.91fF $ **FLOATING
C12616 S.n11439 VSUBS 0.05fF $ **FLOATING
C12617 S.n11440 VSUBS 1.88fF $ **FLOATING
C12618 S.n11441 VSUBS 2.67fF $ **FLOATING
C12619 S.t1195 VSUBS 0.02fF
C12620 S.n11442 VSUBS 0.24fF $ **FLOATING
C12621 S.n11443 VSUBS 0.36fF $ **FLOATING
C12622 S.n11444 VSUBS 0.61fF $ **FLOATING
C12623 S.n11445 VSUBS 0.12fF $ **FLOATING
C12624 S.t495 VSUBS 0.02fF
C12625 S.n11446 VSUBS 0.14fF $ **FLOATING
C12626 S.n11448 VSUBS 2.80fF $ **FLOATING
C12627 S.n11449 VSUBS 2.30fF $ **FLOATING
C12628 S.t1243 VSUBS 0.02fF
C12629 S.n11450 VSUBS 0.12fF $ **FLOATING
C12630 S.n11451 VSUBS 0.14fF $ **FLOATING
C12631 S.t1461 VSUBS 0.02fF
C12632 S.n11453 VSUBS 0.24fF $ **FLOATING
C12633 S.n11454 VSUBS 0.91fF $ **FLOATING
C12634 S.n11455 VSUBS 0.05fF $ **FLOATING
C12635 S.n11456 VSUBS 1.88fF $ **FLOATING
C12636 S.n11457 VSUBS 2.67fF $ **FLOATING
C12637 S.t923 VSUBS 0.02fF
C12638 S.n11458 VSUBS 0.24fF $ **FLOATING
C12639 S.n11459 VSUBS 0.36fF $ **FLOATING
C12640 S.n11460 VSUBS 0.61fF $ **FLOATING
C12641 S.n11461 VSUBS 0.12fF $ **FLOATING
C12642 S.t75 VSUBS 0.02fF
C12643 S.n11462 VSUBS 0.14fF $ **FLOATING
C12644 S.n11464 VSUBS 2.80fF $ **FLOATING
C12645 S.n11465 VSUBS 2.30fF $ **FLOATING
C12646 S.t2149 VSUBS 0.02fF
C12647 S.n11466 VSUBS 0.12fF $ **FLOATING
C12648 S.n11467 VSUBS 0.14fF $ **FLOATING
C12649 S.t1222 VSUBS 0.02fF
C12650 S.n11469 VSUBS 0.24fF $ **FLOATING
C12651 S.n11470 VSUBS 0.91fF $ **FLOATING
C12652 S.n11471 VSUBS 0.05fF $ **FLOATING
C12653 S.n11472 VSUBS 1.88fF $ **FLOATING
C12654 S.n11473 VSUBS 2.67fF $ **FLOATING
C12655 S.t1700 VSUBS 0.02fF
C12656 S.n11474 VSUBS 0.24fF $ **FLOATING
C12657 S.n11475 VSUBS 0.36fF $ **FLOATING
C12658 S.n11476 VSUBS 0.61fF $ **FLOATING
C12659 S.n11477 VSUBS 0.12fF $ **FLOATING
C12660 S.t888 VSUBS 0.02fF
C12661 S.n11478 VSUBS 0.14fF $ **FLOATING
C12662 S.n11480 VSUBS 2.80fF $ **FLOATING
C12663 S.n11481 VSUBS 2.30fF $ **FLOATING
C12664 S.t1758 VSUBS 0.02fF
C12665 S.n11482 VSUBS 0.12fF $ **FLOATING
C12666 S.n11483 VSUBS 0.14fF $ **FLOATING
C12667 S.t1998 VSUBS 0.02fF
C12668 S.n11485 VSUBS 0.24fF $ **FLOATING
C12669 S.n11486 VSUBS 0.91fF $ **FLOATING
C12670 S.n11487 VSUBS 0.05fF $ **FLOATING
C12671 S.n11488 VSUBS 1.88fF $ **FLOATING
C12672 S.n11489 VSUBS 2.67fF $ **FLOATING
C12673 S.t2489 VSUBS 0.02fF
C12674 S.n11490 VSUBS 0.24fF $ **FLOATING
C12675 S.n11491 VSUBS 0.36fF $ **FLOATING
C12676 S.n11492 VSUBS 0.61fF $ **FLOATING
C12677 S.n11493 VSUBS 0.12fF $ **FLOATING
C12678 S.t1670 VSUBS 0.02fF
C12679 S.n11494 VSUBS 0.14fF $ **FLOATING
C12680 S.n11496 VSUBS 2.80fF $ **FLOATING
C12681 S.n11497 VSUBS 2.30fF $ **FLOATING
C12682 S.t2539 VSUBS 0.02fF
C12683 S.n11498 VSUBS 0.12fF $ **FLOATING
C12684 S.n11499 VSUBS 0.14fF $ **FLOATING
C12685 S.t270 VSUBS 0.02fF
C12686 S.n11501 VSUBS 0.24fF $ **FLOATING
C12687 S.n11502 VSUBS 0.91fF $ **FLOATING
C12688 S.n11503 VSUBS 0.05fF $ **FLOATING
C12689 S.n11504 VSUBS 1.88fF $ **FLOATING
C12690 S.n11505 VSUBS 2.67fF $ **FLOATING
C12691 S.t745 VSUBS 0.02fF
C12692 S.n11506 VSUBS 0.24fF $ **FLOATING
C12693 S.n11507 VSUBS 0.36fF $ **FLOATING
C12694 S.n11508 VSUBS 0.61fF $ **FLOATING
C12695 S.n11509 VSUBS 0.12fF $ **FLOATING
C12696 S.t2458 VSUBS 0.02fF
C12697 S.n11510 VSUBS 0.14fF $ **FLOATING
C12698 S.n11512 VSUBS 2.80fF $ **FLOATING
C12699 S.n11513 VSUBS 2.30fF $ **FLOATING
C12700 S.t804 VSUBS 0.02fF
C12701 S.n11514 VSUBS 0.12fF $ **FLOATING
C12702 S.n11515 VSUBS 0.14fF $ **FLOATING
C12703 S.t1049 VSUBS 0.02fF
C12704 S.n11517 VSUBS 0.24fF $ **FLOATING
C12705 S.n11518 VSUBS 0.91fF $ **FLOATING
C12706 S.n11519 VSUBS 0.05fF $ **FLOATING
C12707 S.n11520 VSUBS 1.88fF $ **FLOATING
C12708 S.n11521 VSUBS 2.67fF $ **FLOATING
C12709 S.t1538 VSUBS 0.02fF
C12710 S.n11522 VSUBS 0.24fF $ **FLOATING
C12711 S.n11523 VSUBS 0.36fF $ **FLOATING
C12712 S.n11524 VSUBS 0.61fF $ **FLOATING
C12713 S.n11525 VSUBS 0.12fF $ **FLOATING
C12714 S.t851 VSUBS 0.02fF
C12715 S.n11526 VSUBS 0.14fF $ **FLOATING
C12716 S.n11528 VSUBS 2.80fF $ **FLOATING
C12717 S.n11529 VSUBS 2.30fF $ **FLOATING
C12718 S.t1583 VSUBS 0.02fF
C12719 S.n11530 VSUBS 0.12fF $ **FLOATING
C12720 S.n11531 VSUBS 0.14fF $ **FLOATING
C12721 S.t1833 VSUBS 0.02fF
C12722 S.n11533 VSUBS 0.24fF $ **FLOATING
C12723 S.n11534 VSUBS 0.91fF $ **FLOATING
C12724 S.n11535 VSUBS 0.05fF $ **FLOATING
C12725 S.n11536 VSUBS 1.88fF $ **FLOATING
C12726 S.n11537 VSUBS 2.67fF $ **FLOATING
C12727 S.t96 VSUBS 0.02fF
C12728 S.n11538 VSUBS 0.24fF $ **FLOATING
C12729 S.n11539 VSUBS 0.36fF $ **FLOATING
C12730 S.n11540 VSUBS 0.61fF $ **FLOATING
C12731 S.n11541 VSUBS 0.12fF $ **FLOATING
C12732 S.t329 VSUBS 0.02fF
C12733 S.n11542 VSUBS 0.14fF $ **FLOATING
C12734 S.n11544 VSUBS 2.80fF $ **FLOATING
C12735 S.n11545 VSUBS 2.30fF $ **FLOATING
C12736 S.t1202 VSUBS 0.02fF
C12737 S.n11546 VSUBS 0.12fF $ **FLOATING
C12738 S.n11547 VSUBS 0.14fF $ **FLOATING
C12739 S.t964 VSUBS 0.02fF
C12740 S.n11549 VSUBS 0.24fF $ **FLOATING
C12741 S.n11550 VSUBS 0.91fF $ **FLOATING
C12742 S.n11551 VSUBS 0.05fF $ **FLOATING
C12743 S.n11552 VSUBS 1.88fF $ **FLOATING
C12744 S.n11553 VSUBS 2.67fF $ **FLOATING
C12745 S.t907 VSUBS 0.02fF
C12746 S.n11554 VSUBS 0.24fF $ **FLOATING
C12747 S.n11555 VSUBS 0.36fF $ **FLOATING
C12748 S.n11556 VSUBS 0.61fF $ **FLOATING
C12749 S.n11557 VSUBS 0.12fF $ **FLOATING
C12750 S.t1119 VSUBS 0.02fF
C12751 S.n11558 VSUBS 0.14fF $ **FLOATING
C12752 S.n11560 VSUBS 2.80fF $ **FLOATING
C12753 S.n11561 VSUBS 2.30fF $ **FLOATING
C12754 S.t1982 VSUBS 0.02fF
C12755 S.n11562 VSUBS 0.12fF $ **FLOATING
C12756 S.n11563 VSUBS 0.14fF $ **FLOATING
C12757 S.t1745 VSUBS 0.02fF
C12758 S.n11565 VSUBS 0.24fF $ **FLOATING
C12759 S.n11566 VSUBS 0.91fF $ **FLOATING
C12760 S.n11567 VSUBS 0.05fF $ **FLOATING
C12761 S.n11568 VSUBS 1.88fF $ **FLOATING
C12762 S.n11569 VSUBS 2.67fF $ **FLOATING
C12763 S.t1687 VSUBS 0.02fF
C12764 S.n11570 VSUBS 0.24fF $ **FLOATING
C12765 S.n11571 VSUBS 0.36fF $ **FLOATING
C12766 S.n11572 VSUBS 0.61fF $ **FLOATING
C12767 S.n11573 VSUBS 0.12fF $ **FLOATING
C12768 S.t1901 VSUBS 0.02fF
C12769 S.n11574 VSUBS 0.14fF $ **FLOATING
C12770 S.n11576 VSUBS 2.80fF $ **FLOATING
C12771 S.n11577 VSUBS 2.30fF $ **FLOATING
C12772 S.t250 VSUBS 0.02fF
C12773 S.n11578 VSUBS 0.12fF $ **FLOATING
C12774 S.n11579 VSUBS 0.14fF $ **FLOATING
C12775 S.t2527 VSUBS 0.02fF
C12776 S.n11581 VSUBS 0.24fF $ **FLOATING
C12777 S.n11582 VSUBS 0.91fF $ **FLOATING
C12778 S.n11583 VSUBS 0.05fF $ **FLOATING
C12779 S.n11584 VSUBS 0.12fF $ **FLOATING
C12780 S.t659 VSUBS 0.02fF
C12781 S.n11585 VSUBS 0.14fF $ **FLOATING
C12782 S.t531 VSUBS 0.02fF
C12783 S.n11587 VSUBS 0.24fF $ **FLOATING
C12784 S.n11588 VSUBS 0.36fF $ **FLOATING
C12785 S.n11589 VSUBS 0.61fF $ **FLOATING
C12786 S.n11590 VSUBS 1.60fF $ **FLOATING
C12787 S.n11591 VSUBS 0.03fF $ **FLOATING
C12788 S.n11592 VSUBS 0.14fF $ **FLOATING
C12789 S.n11593 VSUBS 0.58fF $ **FLOATING
C12790 S.n11594 VSUBS 0.12fF $ **FLOATING
C12791 S.n11595 VSUBS 0.53fF $ **FLOATING
C12792 S.n11596 VSUBS 0.41fF $ **FLOATING
C12793 S.n11597 VSUBS 0.25fF $ **FLOATING
C12794 S.n11598 VSUBS 0.25fF $ **FLOATING
C12795 S.n11599 VSUBS 0.68fF $ **FLOATING
C12796 S.n11600 VSUBS 1.97fF $ **FLOATING
C12797 S.t1811 VSUBS 0.02fF
C12798 S.n11601 VSUBS 0.12fF $ **FLOATING
C12799 S.n11602 VSUBS 0.14fF $ **FLOATING
C12800 S.t1941 VSUBS 0.02fF
C12801 S.n11604 VSUBS 0.24fF $ **FLOATING
C12802 S.n11605 VSUBS 0.91fF $ **FLOATING
C12803 S.n11606 VSUBS 0.05fF $ **FLOATING
C12804 S.t47 VSUBS 48.27fF
C12805 S.t791 VSUBS 0.02fF
C12806 S.n11607 VSUBS 0.24fF $ **FLOATING
C12807 S.n11608 VSUBS 0.91fF $ **FLOATING
C12808 S.n11609 VSUBS 0.05fF $ **FLOATING
C12809 S.t1032 VSUBS 0.02fF
C12810 S.n11610 VSUBS 0.12fF $ **FLOATING
C12811 S.n11611 VSUBS 0.14fF $ **FLOATING
C12812 S.n11613 VSUBS 0.12fF $ **FLOATING
C12813 S.t151 VSUBS 0.02fF
C12814 S.n11614 VSUBS 0.14fF $ **FLOATING
C12815 S.n11616 VSUBS 5.17fF $ **FLOATING
C12816 S.n11617 VSUBS 5.44fF $ **FLOATING
C12817 S.t1005 VSUBS 0.02fF
C12818 S.n11618 VSUBS 0.12fF $ **FLOATING
C12819 S.n11619 VSUBS 0.14fF $ **FLOATING
C12820 S.t764 VSUBS 0.02fF
C12821 S.n11621 VSUBS 0.24fF $ **FLOATING
C12822 S.n11622 VSUBS 0.91fF $ **FLOATING
C12823 S.n11623 VSUBS 0.05fF $ **FLOATING
C12824 S.t115 VSUBS 47.89fF
C12825 S.t2040 VSUBS 0.02fF
C12826 S.n11624 VSUBS 0.01fF $ **FLOATING
C12827 S.n11625 VSUBS 0.26fF $ **FLOATING
C12828 S.t2349 VSUBS 0.02fF
C12829 S.n11627 VSUBS 1.19fF $ **FLOATING
C12830 S.n11628 VSUBS 0.05fF $ **FLOATING
C12831 S.t2074 VSUBS 0.02fF
C12832 S.n11629 VSUBS 0.64fF $ **FLOATING
C12833 S.n11630 VSUBS 0.61fF $ **FLOATING
C12834 S.n11631 VSUBS 0.56fF $ **FLOATING
C12835 S.n11632 VSUBS 0.03fF $ **FLOATING
C12836 S.n11633 VSUBS 0.86fF $ **FLOATING
C12837 S.n11634 VSUBS 0.22fF $ **FLOATING
C12838 S.n11635 VSUBS 0.15fF $ **FLOATING
C12839 S.n11636 VSUBS 0.77fF $ **FLOATING
C12840 S.n11637 VSUBS 0.28fF $ **FLOATING
C12841 S.n11638 VSUBS 4.00fF $ **FLOATING
C12842 S.n11639 VSUBS 1.14fF $ **FLOATING
C12843 S.n11640 VSUBS 0.02fF $ **FLOATING
C12844 S.n11641 VSUBS 0.03fF $ **FLOATING
C12845 S.n11642 VSUBS 0.24fF $ **FLOATING
C12846 S.n11643 VSUBS 0.13fF $ **FLOATING
C12847 S.n11644 VSUBS 4.38fF $ **FLOATING
C12848 S.t926 VSUBS 0.02fF
C12849 S.n11645 VSUBS 1.22fF $ **FLOATING
C12850 S.n11646 VSUBS 0.36fF $ **FLOATING
C12851 S.n11647 VSUBS 0.47fF $ **FLOATING
C12852 S.n11648 VSUBS 1.14fF $ **FLOATING
C12853 S.n11649 VSUBS 1.88fF $ **FLOATING
C12854 S.n11650 VSUBS 0.12fF $ **FLOATING
C12855 S.t1025 VSUBS 0.02fF
C12856 S.n11651 VSUBS 0.14fF $ **FLOATING
C12857 S.t815 VSUBS 0.02fF
C12858 S.n11653 VSUBS 0.24fF $ **FLOATING
C12859 S.n11654 VSUBS 0.36fF $ **FLOATING
C12860 S.n11655 VSUBS 0.61fF $ **FLOATING
C12861 S.n11656 VSUBS 2.67fF $ **FLOATING
C12862 S.n11657 VSUBS 3.93fF $ **FLOATING
C12863 S.t1655 VSUBS 0.02fF
C12864 S.n11658 VSUBS 0.24fF $ **FLOATING
C12865 S.n11659 VSUBS 0.91fF $ **FLOATING
C12866 S.n11660 VSUBS 0.05fF $ **FLOATING
C12867 S.t1893 VSUBS 0.02fF
C12868 S.n11661 VSUBS 0.12fF $ **FLOATING
C12869 S.n11662 VSUBS 0.14fF $ **FLOATING
C12870 S.n11664 VSUBS 1.88fF $ **FLOATING
C12871 S.n11665 VSUBS 2.67fF $ **FLOATING
C12872 S.t2549 VSUBS 0.02fF
C12873 S.n11666 VSUBS 0.24fF $ **FLOATING
C12874 S.n11667 VSUBS 0.36fF $ **FLOATING
C12875 S.n11668 VSUBS 0.61fF $ **FLOATING
C12876 S.n11669 VSUBS 0.12fF $ **FLOATING
C12877 S.t240 VSUBS 0.02fF
C12878 S.n11670 VSUBS 0.14fF $ **FLOATING
C12879 S.n11672 VSUBS 5.17fF $ **FLOATING
C12880 S.t873 VSUBS 0.02fF
C12881 S.n11673 VSUBS 0.24fF $ **FLOATING
C12882 S.n11674 VSUBS 0.91fF $ **FLOATING
C12883 S.n11675 VSUBS 0.05fF $ **FLOATING
C12884 S.t1113 VSUBS 0.02fF
C12885 S.n11676 VSUBS 0.12fF $ **FLOATING
C12886 S.n11677 VSUBS 0.14fF $ **FLOATING
C12887 S.n11679 VSUBS 1.88fF $ **FLOATING
C12888 S.n11680 VSUBS 2.67fF $ **FLOATING
C12889 S.t1770 VSUBS 0.02fF
C12890 S.n11681 VSUBS 0.24fF $ **FLOATING
C12891 S.n11682 VSUBS 0.36fF $ **FLOATING
C12892 S.n11683 VSUBS 0.61fF $ **FLOATING
C12893 S.n11684 VSUBS 0.12fF $ **FLOATING
C12894 S.t1977 VSUBS 0.02fF
C12895 S.n11685 VSUBS 0.14fF $ **FLOATING
C12896 S.n11687 VSUBS 5.17fF $ **FLOATING
C12897 S.t50 VSUBS 0.02fF
C12898 S.n11688 VSUBS 0.24fF $ **FLOATING
C12899 S.n11689 VSUBS 0.91fF $ **FLOATING
C12900 S.n11690 VSUBS 0.05fF $ **FLOATING
C12901 S.t325 VSUBS 0.02fF
C12902 S.n11691 VSUBS 0.12fF $ **FLOATING
C12903 S.n11692 VSUBS 0.14fF $ **FLOATING
C12904 S.n11694 VSUBS 1.88fF $ **FLOATING
C12905 S.n11695 VSUBS 2.67fF $ **FLOATING
C12906 S.t988 VSUBS 0.02fF
C12907 S.n11696 VSUBS 0.24fF $ **FLOATING
C12908 S.n11697 VSUBS 0.36fF $ **FLOATING
C12909 S.n11698 VSUBS 0.61fF $ **FLOATING
C12910 S.n11699 VSUBS 0.12fF $ **FLOATING
C12911 S.t1197 VSUBS 0.02fF
C12912 S.n11700 VSUBS 0.14fF $ **FLOATING
C12913 S.n11702 VSUBS 5.17fF $ **FLOATING
C12914 S.t1830 VSUBS 0.02fF
C12915 S.n11703 VSUBS 0.24fF $ **FLOATING
C12916 S.n11704 VSUBS 0.91fF $ **FLOATING
C12917 S.n11705 VSUBS 0.05fF $ **FLOATING
C12918 S.t2515 VSUBS 0.02fF
C12919 S.n11706 VSUBS 0.12fF $ **FLOATING
C12920 S.n11707 VSUBS 0.14fF $ **FLOATING
C12921 S.n11709 VSUBS 1.88fF $ **FLOATING
C12922 S.n11710 VSUBS 2.67fF $ **FLOATING
C12923 S.t1545 VSUBS 0.02fF
C12924 S.n11711 VSUBS 0.24fF $ **FLOATING
C12925 S.n11712 VSUBS 0.36fF $ **FLOATING
C12926 S.n11713 VSUBS 0.61fF $ **FLOATING
C12927 S.n11714 VSUBS 0.12fF $ **FLOATING
C12928 S.t724 VSUBS 0.02fF
C12929 S.n11715 VSUBS 0.14fF $ **FLOATING
C12930 S.n11717 VSUBS 5.17fF $ **FLOATING
C12931 S.t1843 VSUBS 0.02fF
C12932 S.n11718 VSUBS 0.24fF $ **FLOATING
C12933 S.n11719 VSUBS 0.91fF $ **FLOATING
C12934 S.n11720 VSUBS 0.05fF $ **FLOATING
C12935 S.t1594 VSUBS 0.02fF
C12936 S.n11721 VSUBS 0.12fF $ **FLOATING
C12937 S.n11722 VSUBS 0.14fF $ **FLOATING
C12938 S.n11724 VSUBS 1.88fF $ **FLOATING
C12939 S.n11725 VSUBS 2.67fF $ **FLOATING
C12940 S.t752 VSUBS 0.02fF
C12941 S.n11726 VSUBS 0.24fF $ **FLOATING
C12942 S.n11727 VSUBS 0.36fF $ **FLOATING
C12943 S.n11728 VSUBS 0.61fF $ **FLOATING
C12944 S.n11729 VSUBS 0.12fF $ **FLOATING
C12945 S.t2465 VSUBS 0.02fF
C12946 S.n11730 VSUBS 0.14fF $ **FLOATING
C12947 S.n11732 VSUBS 5.17fF $ **FLOATING
C12948 S.t1058 VSUBS 0.02fF
C12949 S.n11733 VSUBS 0.24fF $ **FLOATING
C12950 S.n11734 VSUBS 0.91fF $ **FLOATING
C12951 S.n11735 VSUBS 0.05fF $ **FLOATING
C12952 S.t812 VSUBS 0.02fF
C12953 S.n11736 VSUBS 0.12fF $ **FLOATING
C12954 S.n11737 VSUBS 0.14fF $ **FLOATING
C12955 S.n11739 VSUBS 1.88fF $ **FLOATING
C12956 S.n11740 VSUBS 2.67fF $ **FLOATING
C12957 S.t2496 VSUBS 0.02fF
C12958 S.n11741 VSUBS 0.24fF $ **FLOATING
C12959 S.n11742 VSUBS 0.36fF $ **FLOATING
C12960 S.n11743 VSUBS 0.61fF $ **FLOATING
C12961 S.n11744 VSUBS 0.12fF $ **FLOATING
C12962 S.t1679 VSUBS 0.02fF
C12963 S.n11745 VSUBS 0.14fF $ **FLOATING
C12964 S.n11747 VSUBS 5.17fF $ **FLOATING
C12965 S.t278 VSUBS 0.02fF
C12966 S.n11748 VSUBS 0.24fF $ **FLOATING
C12967 S.n11749 VSUBS 0.91fF $ **FLOATING
C12968 S.n11750 VSUBS 0.05fF $ **FLOATING
C12969 S.t2546 VSUBS 0.02fF
C12970 S.n11751 VSUBS 0.12fF $ **FLOATING
C12971 S.n11752 VSUBS 0.14fF $ **FLOATING
C12972 S.n11754 VSUBS 1.88fF $ **FLOATING
C12973 S.n11755 VSUBS 2.67fF $ **FLOATING
C12974 S.t1709 VSUBS 0.02fF
C12975 S.n11756 VSUBS 0.24fF $ **FLOATING
C12976 S.n11757 VSUBS 0.36fF $ **FLOATING
C12977 S.n11758 VSUBS 0.61fF $ **FLOATING
C12978 S.n11759 VSUBS 0.12fF $ **FLOATING
C12979 S.t899 VSUBS 0.02fF
C12980 S.n11760 VSUBS 0.14fF $ **FLOATING
C12981 S.n11762 VSUBS 5.17fF $ **FLOATING
C12982 S.t2005 VSUBS 0.02fF
C12983 S.n11763 VSUBS 0.24fF $ **FLOATING
C12984 S.n11764 VSUBS 0.91fF $ **FLOATING
C12985 S.n11765 VSUBS 0.05fF $ **FLOATING
C12986 S.t1768 VSUBS 0.02fF
C12987 S.n11766 VSUBS 0.12fF $ **FLOATING
C12988 S.n11767 VSUBS 0.14fF $ **FLOATING
C12989 S.n11769 VSUBS 1.88fF $ **FLOATING
C12990 S.n11770 VSUBS 2.67fF $ **FLOATING
C12991 S.t2109 VSUBS 0.02fF
C12992 S.n11771 VSUBS 0.24fF $ **FLOATING
C12993 S.n11772 VSUBS 0.36fF $ **FLOATING
C12994 S.n11773 VSUBS 0.61fF $ **FLOATING
C12995 S.n11774 VSUBS 0.12fF $ **FLOATING
C12996 S.t1291 VSUBS 0.02fF
C12997 S.n11775 VSUBS 0.14fF $ **FLOATING
C12998 S.n11777 VSUBS 5.17fF $ **FLOATING
C12999 S.t2383 VSUBS 0.02fF
C13000 S.n11778 VSUBS 0.24fF $ **FLOATING
C13001 S.n11779 VSUBS 0.91fF $ **FLOATING
C13002 S.n11780 VSUBS 0.05fF $ **FLOATING
C13003 S.t2159 VSUBS 0.02fF
C13004 S.n11781 VSUBS 0.12fF $ **FLOATING
C13005 S.n11782 VSUBS 0.14fF $ **FLOATING
C13006 S.n11784 VSUBS 1.88fF $ **FLOATING
C13007 S.n11785 VSUBS 2.67fF $ **FLOATING
C13008 S.t1208 VSUBS 0.02fF
C13009 S.n11786 VSUBS 0.24fF $ **FLOATING
C13010 S.n11787 VSUBS 0.36fF $ **FLOATING
C13011 S.n11788 VSUBS 0.61fF $ **FLOATING
C13012 S.n11789 VSUBS 0.12fF $ **FLOATING
C13013 S.t385 VSUBS 0.02fF
C13014 S.n11790 VSUBS 0.14fF $ **FLOATING
C13015 S.n11792 VSUBS 5.17fF $ **FLOATING
C13016 S.t1475 VSUBS 0.02fF
C13017 S.n11793 VSUBS 0.24fF $ **FLOATING
C13018 S.n11794 VSUBS 0.91fF $ **FLOATING
C13019 S.n11795 VSUBS 0.05fF $ **FLOATING
C13020 S.t1250 VSUBS 0.02fF
C13021 S.n11796 VSUBS 0.12fF $ **FLOATING
C13022 S.n11797 VSUBS 0.14fF $ **FLOATING
C13023 S.n11799 VSUBS 1.88fF $ **FLOATING
C13024 S.n11800 VSUBS 2.67fF $ **FLOATING
C13025 S.t411 VSUBS 0.02fF
C13026 S.n11801 VSUBS 0.24fF $ **FLOATING
C13027 S.n11802 VSUBS 0.36fF $ **FLOATING
C13028 S.n11803 VSUBS 0.61fF $ **FLOATING
C13029 S.n11804 VSUBS 0.12fF $ **FLOATING
C13030 S.t2117 VSUBS 0.02fF
C13031 S.n11805 VSUBS 0.14fF $ **FLOATING
C13032 S.n11807 VSUBS 5.17fF $ **FLOATING
C13033 S.t686 VSUBS 0.02fF
C13034 S.n11808 VSUBS 0.24fF $ **FLOATING
C13035 S.n11809 VSUBS 0.91fF $ **FLOATING
C13036 S.n11810 VSUBS 0.05fF $ **FLOATING
C13037 S.t463 VSUBS 0.02fF
C13038 S.n11811 VSUBS 0.12fF $ **FLOATING
C13039 S.n11812 VSUBS 0.14fF $ **FLOATING
C13040 S.n11814 VSUBS 1.88fF $ **FLOATING
C13041 S.n11815 VSUBS 0.12fF $ **FLOATING
C13042 S.t1330 VSUBS 0.02fF
C13043 S.n11816 VSUBS 0.14fF $ **FLOATING
C13044 S.t2144 VSUBS 0.02fF
C13045 S.n11818 VSUBS 0.24fF $ **FLOATING
C13046 S.n11819 VSUBS 0.36fF $ **FLOATING
C13047 S.n11820 VSUBS 0.61fF $ **FLOATING
C13048 S.n11821 VSUBS 2.67fF $ **FLOATING
C13049 S.n11822 VSUBS 5.17fF $ **FLOATING
C13050 S.t2421 VSUBS 0.02fF
C13051 S.n11823 VSUBS 0.24fF $ **FLOATING
C13052 S.n11824 VSUBS 0.91fF $ **FLOATING
C13053 S.n11825 VSUBS 0.05fF $ **FLOATING
C13054 S.t2197 VSUBS 0.02fF
C13055 S.n11826 VSUBS 0.12fF $ **FLOATING
C13056 S.n11827 VSUBS 0.14fF $ **FLOATING
C13057 S.n11829 VSUBS 1.88fF $ **FLOATING
C13058 S.n11830 VSUBS 2.67fF $ **FLOATING
C13059 S.t1360 VSUBS 0.02fF
C13060 S.n11831 VSUBS 0.24fF $ **FLOATING
C13061 S.n11832 VSUBS 0.36fF $ **FLOATING
C13062 S.n11833 VSUBS 0.61fF $ **FLOATING
C13063 S.n11834 VSUBS 0.12fF $ **FLOATING
C13064 S.t544 VSUBS 0.02fF
C13065 S.n11835 VSUBS 0.14fF $ **FLOATING
C13066 S.n11837 VSUBS 5.17fF $ **FLOATING
C13067 S.t1637 VSUBS 0.02fF
C13068 S.n11838 VSUBS 0.24fF $ **FLOATING
C13069 S.n11839 VSUBS 0.91fF $ **FLOATING
C13070 S.n11840 VSUBS 0.05fF $ **FLOATING
C13071 S.t2578 VSUBS 0.02fF
C13072 S.n11841 VSUBS 0.12fF $ **FLOATING
C13073 S.n11842 VSUBS 0.14fF $ **FLOATING
C13074 S.n11844 VSUBS 1.88fF $ **FLOATING
C13075 S.n11845 VSUBS 2.67fF $ **FLOATING
C13076 S.t1742 VSUBS 0.02fF
C13077 S.n11846 VSUBS 0.24fF $ **FLOATING
C13078 S.n11847 VSUBS 0.36fF $ **FLOATING
C13079 S.n11848 VSUBS 0.61fF $ **FLOATING
C13080 S.n11849 VSUBS 0.12fF $ **FLOATING
C13081 S.t932 VSUBS 0.02fF
C13082 S.n11850 VSUBS 0.14fF $ **FLOATING
C13083 S.n11852 VSUBS 5.16fF $ **FLOATING
C13084 S.t2035 VSUBS 0.02fF
C13085 S.n11853 VSUBS 0.24fF $ **FLOATING
C13086 S.n11854 VSUBS 0.91fF $ **FLOATING
C13087 S.n11855 VSUBS 0.05fF $ **FLOATING
C13088 S.t1796 VSUBS 0.02fF
C13089 S.n11856 VSUBS 0.12fF $ **FLOATING
C13090 S.n11857 VSUBS 0.14fF $ **FLOATING
C13091 S.n11859 VSUBS 1.88fF $ **FLOATING
C13092 S.n11860 VSUBS 0.12fF $ **FLOATING
C13093 S.t2534 VSUBS 0.02fF
C13094 S.n11861 VSUBS 0.14fF $ **FLOATING
C13095 S.t829 VSUBS 0.02fF
C13096 S.n11863 VSUBS 0.24fF $ **FLOATING
C13097 S.n11864 VSUBS 0.36fF $ **FLOATING
C13098 S.n11865 VSUBS 0.61fF $ **FLOATING
C13099 S.n11866 VSUBS 0.32fF $ **FLOATING
C13100 S.n11867 VSUBS 0.92fF $ **FLOATING
C13101 S.n11868 VSUBS 1.09fF $ **FLOATING
C13102 S.n11869 VSUBS 0.15fF $ **FLOATING
C13103 S.n11870 VSUBS 4.96fF $ **FLOATING
C13104 S.t1134 VSUBS 0.02fF
C13105 S.n11871 VSUBS 0.24fF $ **FLOATING
C13106 S.n11872 VSUBS 0.91fF $ **FLOATING
C13107 S.n11873 VSUBS 0.05fF $ **FLOATING
C13108 S.t883 VSUBS 0.02fF
C13109 S.n11874 VSUBS 0.12fF $ **FLOATING
C13110 S.n11875 VSUBS 0.14fF $ **FLOATING
C13111 S.t1225 VSUBS 0.02fF
C13112 S.n11877 VSUBS 0.95fF $ **FLOATING
C13113 S.n11878 VSUBS 0.71fF $ **FLOATING
C13114 S.n11879 VSUBS 1.78fF $ **FLOATING
C13115 S.n11880 VSUBS 3.05fF $ **FLOATING
C13116 S.t2563 VSUBS 0.02fF
C13117 S.n11881 VSUBS 0.24fF $ **FLOATING
C13118 S.n11882 VSUBS 0.36fF $ **FLOATING
C13119 S.n11883 VSUBS 0.61fF $ **FLOATING
C13120 S.n11884 VSUBS 0.12fF $ **FLOATING
C13121 S.t1750 VSUBS 0.02fF
C13122 S.n11885 VSUBS 0.14fF $ **FLOATING
C13123 S.n11887 VSUBS 0.23fF $ **FLOATING
C13124 S.n11888 VSUBS 0.66fF $ **FLOATING
C13125 S.n11889 VSUBS 0.91fF $ **FLOATING
C13126 S.n11890 VSUBS 0.23fF $ **FLOATING
C13127 S.n11891 VSUBS 1.99fF $ **FLOATING
C13128 S.t345 VSUBS 0.02fF
C13129 S.n11892 VSUBS 0.24fF $ **FLOATING
C13130 S.n11893 VSUBS 0.91fF $ **FLOATING
C13131 S.n11894 VSUBS 0.05fF $ **FLOATING
C13132 S.t66 VSUBS 0.02fF
C13133 S.n11895 VSUBS 0.12fF $ **FLOATING
C13134 S.n11896 VSUBS 0.14fF $ **FLOATING
C13135 S.n11898 VSUBS 0.25fF $ **FLOATING
C13136 S.n11899 VSUBS 0.09fF $ **FLOATING
C13137 S.n11900 VSUBS 0.20fF $ **FLOATING
C13138 S.n11901 VSUBS 0.78fF $ **FLOATING
C13139 S.n11902 VSUBS 1.93fF $ **FLOATING
C13140 S.n11903 VSUBS 1.88fF $ **FLOATING
C13141 S.n11904 VSUBS 0.12fF $ **FLOATING
C13142 S.t1806 VSUBS 0.02fF
C13143 S.n11905 VSUBS 0.14fF $ **FLOATING
C13144 S.t1596 VSUBS 0.02fF
C13145 S.n11907 VSUBS 0.24fF $ **FLOATING
C13146 S.n11908 VSUBS 0.36fF $ **FLOATING
C13147 S.n11909 VSUBS 0.61fF $ **FLOATING
C13148 S.n11910 VSUBS 2.67fF $ **FLOATING
C13149 S.n11911 VSUBS 2.99fF $ **FLOATING
C13150 S.t143 VSUBS 0.02fF
C13151 S.n11912 VSUBS 0.12fF $ **FLOATING
C13152 S.n11913 VSUBS 0.14fF $ **FLOATING
C13153 S.t2438 VSUBS 0.02fF
C13154 S.n11915 VSUBS 0.24fF $ **FLOATING
C13155 S.n11916 VSUBS 0.91fF $ **FLOATING
C13156 S.n11917 VSUBS 0.05fF $ **FLOATING
C13157 S.t1598 VSUBS 0.02fF
C13158 S.n11918 VSUBS 0.01fF $ **FLOATING
C13159 S.n11919 VSUBS 0.26fF $ **FLOATING
C13160 S.t65 VSUBS 48.27fF
C13161 S.n11920 VSUBS 0.25fF $ **FLOATING
C13162 S.n11921 VSUBS 2.92fF $ **FLOATING
C13163 S.n11922 VSUBS 2.33fF $ **FLOATING
C13164 S.n11923 VSUBS 4.57fF $ **FLOATING
C13165 S.t379 VSUBS 0.02fF
C13166 S.n11924 VSUBS 1.28fF $ **FLOATING
C13167 S.t266 VSUBS 0.02fF
C13168 S.n11925 VSUBS 0.44fF $ **FLOATING
C13169 S.t1973 VSUBS 0.02fF
C13170 S.n11926 VSUBS 0.89fF $ **FLOATING
C13171 S.t2295 VSUBS 0.02fF
C13172 S.n11927 VSUBS 0.02fF $ **FLOATING
C13173 S.n11928 VSUBS 0.37fF $ **FLOATING
C13174 S.t1110 VSUBS 0.02fF
C13175 S.n11929 VSUBS 0.89fF $ **FLOATING
C13176 S.t2540 VSUBS 0.02fF
C13177 S.n11930 VSUBS 0.89fF $ **FLOATING
C13178 S.t890 VSUBS 0.02fF
C13179 S.n11931 VSUBS 0.89fF $ **FLOATING
C13180 S.t2017 VSUBS 0.02fF
C13181 S.n11932 VSUBS 0.02fF $ **FLOATING
C13182 S.n11933 VSUBS 0.37fF $ **FLOATING
C13183 S.t1673 VSUBS 0.02fF
C13184 S.n11934 VSUBS 0.89fF $ **FLOATING
C13185 S.t807 VSUBS 0.02fF
C13186 S.n11935 VSUBS 0.89fF $ **FLOATING
C13187 S.t289 VSUBS 0.02fF
C13188 S.n11936 VSUBS 0.02fF $ **FLOATING
C13189 S.n11937 VSUBS 0.37fF $ **FLOATING
C13190 S.t6 VSUBS 0.02fF
C13191 S.n11938 VSUBS 0.89fF $ **FLOATING
C13192 S.t1715 VSUBS 0.02fF
C13193 S.n11939 VSUBS 0.89fF $ **FLOATING
C13194 S.t1204 VSUBS 0.02fF
C13195 S.n11940 VSUBS 0.02fF $ **FLOATING
C13196 S.n11941 VSUBS 0.37fF $ **FLOATING
C13197 S.t852 VSUBS 0.02fF
C13198 S.n11942 VSUBS 0.89fF $ **FLOATING
C13199 S.t1336 VSUBS 0.02fF
C13200 S.n11943 VSUBS 0.89fF $ **FLOATING
C13201 S.t794 VSUBS 0.02fF
C13202 S.n11944 VSUBS 0.02fF $ **FLOATING
C13203 S.n11945 VSUBS 0.37fF $ **FLOATING
C13204 S.t469 VSUBS 0.02fF
C13205 S.n11946 VSUBS 0.89fF $ **FLOATING
C13206 S.t2122 VSUBS 0.02fF
C13207 S.n11947 VSUBS 0.89fF $ **FLOATING
C13208 S.t1576 VSUBS 0.02fF
C13209 S.n11948 VSUBS 0.02fF $ **FLOATING
C13210 S.n11949 VSUBS 0.37fF $ **FLOATING
C13211 S.t1258 VSUBS 0.02fF
C13212 S.n11950 VSUBS 0.89fF $ **FLOATING
C13213 S.t389 VSUBS 0.02fF
C13214 S.n11951 VSUBS 0.89fF $ **FLOATING
C13215 S.t2365 VSUBS 0.02fF
C13216 S.n11952 VSUBS 0.02fF $ **FLOATING
C13217 S.n11953 VSUBS 0.37fF $ **FLOATING
C13218 S.t2042 VSUBS 0.02fF
C13219 S.n11954 VSUBS 0.89fF $ **FLOATING
C13220 S.t1181 VSUBS 0.02fF
C13221 S.n11955 VSUBS 0.89fF $ **FLOATING
C13222 S.t633 VSUBS 0.02fF
C13223 S.n11956 VSUBS 0.02fF $ **FLOATING
C13224 S.n11957 VSUBS 0.37fF $ **FLOATING
C13225 S.t432 VSUBS 0.02fF
C13226 S.n11958 VSUBS 0.89fF $ **FLOATING
C13227 S.t2085 VSUBS 0.02fF
C13228 S.n11959 VSUBS 0.89fF $ **FLOATING
C13229 S.t1543 VSUBS 0.02fF
C13230 S.n11960 VSUBS 0.02fF $ **FLOATING
C13231 S.n11961 VSUBS 0.37fF $ **FLOATING
C13232 S.t2554 VSUBS 0.02fF
C13233 S.n11962 VSUBS 0.89fF $ **FLOATING
C13234 S.t1686 VSUBS 0.02fF
C13235 S.n11963 VSUBS 0.89fF $ **FLOATING
C13236 S.t1173 VSUBS 0.02fF
C13237 S.n11964 VSUBS 0.02fF $ **FLOATING
C13238 S.n11965 VSUBS 0.37fF $ **FLOATING
C13239 S.t819 VSUBS 0.02fF
C13240 S.n11966 VSUBS 0.89fF $ **FLOATING
C13241 S.t2472 VSUBS 0.02fF
C13242 S.n11967 VSUBS 0.89fF $ **FLOATING
C13243 S.t1955 VSUBS 0.02fF
C13244 S.n11968 VSUBS 0.02fF $ **FLOATING
C13245 S.n11969 VSUBS 0.37fF $ **FLOATING
C13246 S.t1601 VSUBS 0.02fF
C13247 S.n11970 VSUBS 0.89fF $ **FLOATING
C13248 S.t730 VSUBS 0.02fF
C13249 S.n11971 VSUBS 0.89fF $ **FLOATING
C13250 S.t215 VSUBS 0.02fF
C13251 S.n11972 VSUBS 0.02fF $ **FLOATING
C13252 S.n11973 VSUBS 0.37fF $ **FLOATING
C13253 S.t2389 VSUBS 0.02fF
C13254 S.n11974 VSUBS 0.89fF $ **FLOATING
C13255 S.t1523 VSUBS 0.02fF
C13256 S.n11975 VSUBS 0.89fF $ **FLOATING
C13257 S.t1003 VSUBS 0.02fF
C13258 S.n11976 VSUBS 0.02fF $ **FLOATING
C13259 S.n11977 VSUBS 0.37fF $ **FLOATING
C13260 S.t778 VSUBS 0.02fF
C13261 S.n11978 VSUBS 0.89fF $ **FLOATING
C13262 S.t478 VSUBS 0.02fF
C13263 S.n11979 VSUBS 0.89fF $ **FLOATING
C13264 S.t1668 VSUBS 0.02fF
C13265 S.n11980 VSUBS 0.02fF $ **FLOATING
C13266 S.n11981 VSUBS 0.37fF $ **FLOATING
C13267 S.t2134 VSUBS 0.02fF
C13268 S.n11982 VSUBS 0.89fF $ **FLOATING
C13269 S.t1265 VSUBS 0.02fF
C13270 S.n11983 VSUBS 0.89fF $ **FLOATING
C13271 S.t2459 VSUBS 0.02fF
C13272 S.n11984 VSUBS 0.02fF $ **FLOATING
C13273 S.n11985 VSUBS 0.37fF $ **FLOATING
C13274 S.t2055 VSUBS 0.02fF
C13275 S.n11986 VSUBS 0.89fF $ **FLOATING
C13276 S.t400 VSUBS 0.02fF
C13277 S.n11987 VSUBS 0.89fF $ **FLOATING
C13278 S.t717 VSUBS 0.02fF
C13279 S.n11988 VSUBS 0.02fF $ **FLOATING
C13280 S.n11989 VSUBS 0.37fF $ **FLOATING
C13281 S.t322 VSUBS 0.02fF
C13282 S.n11990 VSUBS 0.89fF $ **FLOATING
C13283 S.t1191 VSUBS 0.02fF
C13284 S.n11991 VSUBS 0.89fF $ **FLOATING
C13285 S.t1509 VSUBS 0.02fF
C13286 S.n11992 VSUBS 0.02fF $ **FLOATING
C13287 S.n11993 VSUBS 0.37fF $ **FLOATING
C13288 S.t0 VSUBS 1373.26fF
C13289 S.n11994 VSUBS 0.47fF $ **FLOATING
C13290 S.n11995 VSUBS 6.92fF $ **FLOATING
C13291 S.n11996 VSUBS 16.14fF $ **FLOATING
C13292 S.n11997 VSUBS 2.81fF $ **FLOATING
C13293 S.n11998 VSUBS 1.89fF $ **FLOATING
C13294 S.n11999 VSUBS 0.06fF $ **FLOATING
C13295 S.n12000 VSUBS 0.03fF $ **FLOATING
C13296 S.n12001 VSUBS 0.04fF $ **FLOATING
C13297 S.n12002 VSUBS 0.99fF $ **FLOATING
C13298 S.n12003 VSUBS 0.02fF $ **FLOATING
C13299 S.n12004 VSUBS 0.01fF $ **FLOATING
C13300 S.n12005 VSUBS 0.02fF $ **FLOATING
C13301 S.n12006 VSUBS 0.08fF $ **FLOATING
C13302 S.n12007 VSUBS 0.36fF $ **FLOATING
C13303 S.n12008 VSUBS 1.85fF $ **FLOATING
C13304 S.t1406 VSUBS 0.02fF
C13305 S.n12009 VSUBS 0.24fF $ **FLOATING
C13306 S.n12010 VSUBS 0.36fF $ **FLOATING
C13307 S.n12011 VSUBS 0.61fF $ **FLOATING
C13308 S.n12012 VSUBS 0.12fF $ **FLOATING
C13309 S.t584 VSUBS 0.02fF
C13310 S.n12013 VSUBS 0.14fF $ **FLOATING
C13311 S.n12015 VSUBS 0.70fF $ **FLOATING
C13312 S.n12016 VSUBS 0.23fF $ **FLOATING
C13313 S.n12017 VSUBS 0.23fF $ **FLOATING
C13314 S.n12018 VSUBS 0.70fF $ **FLOATING
C13315 S.n12019 VSUBS 1.16fF $ **FLOATING
C13316 S.n12020 VSUBS 0.22fF $ **FLOATING
C13317 S.n12021 VSUBS 0.25fF $ **FLOATING
C13318 S.n12022 VSUBS 0.09fF $ **FLOATING
C13319 S.n12023 VSUBS 1.88fF $ **FLOATING
C13320 S.t1683 VSUBS 0.02fF
C13321 S.n12024 VSUBS 0.24fF $ **FLOATING
C13322 S.n12025 VSUBS 0.91fF $ **FLOATING
C13323 S.n12026 VSUBS 0.05fF $ **FLOATING
C13324 S.t1453 VSUBS 0.02fF
C13325 S.n12027 VSUBS 0.12fF $ **FLOATING
C13326 S.n12028 VSUBS 0.14fF $ **FLOATING
C13327 S.n12030 VSUBS 0.09fF $ **FLOATING
C13328 S.n12031 VSUBS 0.21fF $ **FLOATING
C13329 S.n12032 VSUBS 0.07fF $ **FLOATING
C13330 S.n12033 VSUBS 0.06fF $ **FLOATING
C13331 S.n12034 VSUBS 0.07fF $ **FLOATING
C13332 S.n12035 VSUBS 0.18fF $ **FLOATING
C13333 S.n12036 VSUBS 0.20fF $ **FLOATING
C13334 S.n12037 VSUBS 1.04fF $ **FLOATING
C13335 S.n12038 VSUBS 0.54fF $ **FLOATING
C13336 S.n12039 VSUBS 2.33fF $ **FLOATING
C13337 S.n12040 VSUBS 0.12fF $ **FLOATING
C13338 S.t2321 VSUBS 0.02fF
C13339 S.n12041 VSUBS 0.14fF $ **FLOATING
C13340 S.t615 VSUBS 0.02fF
C13341 S.n12043 VSUBS 0.24fF $ **FLOATING
C13342 S.n12044 VSUBS 0.36fF $ **FLOATING
C13343 S.n12045 VSUBS 0.61fF $ **FLOATING
C13344 S.n12046 VSUBS 1.73fF $ **FLOATING
C13345 S.n12047 VSUBS 2.44fF $ **FLOATING
C13346 S.t663 VSUBS 0.02fF
C13347 S.n12048 VSUBS 0.12fF $ **FLOATING
C13348 S.n12049 VSUBS 0.14fF $ **FLOATING
C13349 S.t904 VSUBS 0.02fF
C13350 S.n12051 VSUBS 0.24fF $ **FLOATING
C13351 S.n12052 VSUBS 0.91fF $ **FLOATING
C13352 S.n12053 VSUBS 0.05fF $ **FLOATING
C13353 S.n12054 VSUBS 2.94fF $ **FLOATING
C13354 S.n12055 VSUBS 1.88fF $ **FLOATING
C13355 S.n12056 VSUBS 0.12fF $ **FLOATING
C13356 S.t1497 VSUBS 0.02fF
C13357 S.n12057 VSUBS 0.14fF $ **FLOATING
C13358 S.t2314 VSUBS 0.02fF
C13359 S.n12059 VSUBS 0.24fF $ **FLOATING
C13360 S.n12060 VSUBS 0.36fF $ **FLOATING
C13361 S.n12061 VSUBS 0.61fF $ **FLOATING
C13362 S.n12062 VSUBS 0.92fF $ **FLOATING
C13363 S.n12063 VSUBS 0.32fF $ **FLOATING
C13364 S.n12064 VSUBS 0.92fF $ **FLOATING
C13365 S.n12065 VSUBS 1.09fF $ **FLOATING
C13366 S.n12066 VSUBS 0.15fF $ **FLOATING
C13367 S.n12067 VSUBS 4.96fF $ **FLOATING
C13368 S.t2360 VSUBS 0.02fF
C13369 S.n12068 VSUBS 0.12fF $ **FLOATING
C13370 S.n12069 VSUBS 0.14fF $ **FLOATING
C13371 S.t37 VSUBS 0.02fF
C13372 S.n12071 VSUBS 0.24fF $ **FLOATING
C13373 S.n12072 VSUBS 0.91fF $ **FLOATING
C13374 S.n12073 VSUBS 0.05fF $ **FLOATING
C13375 S.n12074 VSUBS 1.88fF $ **FLOATING
C13376 S.n12075 VSUBS 2.67fF $ **FLOATING
C13377 S.t1938 VSUBS 0.02fF
C13378 S.n12076 VSUBS 0.24fF $ **FLOATING
C13379 S.n12077 VSUBS 0.36fF $ **FLOATING
C13380 S.n12078 VSUBS 0.61fF $ **FLOATING
C13381 S.n12079 VSUBS 0.12fF $ **FLOATING
C13382 S.t1124 VSUBS 0.02fF
C13383 S.n12080 VSUBS 0.14fF $ **FLOATING
C13384 S.n12082 VSUBS 2.94fF $ **FLOATING
C13385 S.n12083 VSUBS 5.16fF $ **FLOATING
C13386 S.t630 VSUBS 0.02fF
C13387 S.n12084 VSUBS 0.12fF $ **FLOATING
C13388 S.n12085 VSUBS 0.14fF $ **FLOATING
C13389 S.t2214 VSUBS 0.02fF
C13390 S.n12087 VSUBS 0.24fF $ **FLOATING
C13391 S.n12088 VSUBS 0.91fF $ **FLOATING
C13392 S.n12089 VSUBS 0.05fF $ **FLOATING
C13393 S.n12090 VSUBS 1.88fF $ **FLOATING
C13394 S.n12091 VSUBS 2.67fF $ **FLOATING
C13395 S.t197 VSUBS 0.02fF
C13396 S.n12092 VSUBS 0.24fF $ **FLOATING
C13397 S.n12093 VSUBS 0.36fF $ **FLOATING
C13398 S.n12094 VSUBS 0.61fF $ **FLOATING
C13399 S.n12095 VSUBS 0.12fF $ **FLOATING
C13400 S.t1907 VSUBS 0.02fF
C13401 S.n12096 VSUBS 0.14fF $ **FLOATING
C13402 S.n12098 VSUBS 5.17fF $ **FLOATING
C13403 S.t254 VSUBS 0.02fF
C13404 S.n12099 VSUBS 0.12fF $ **FLOATING
C13405 S.n12100 VSUBS 0.14fF $ **FLOATING
C13406 S.t482 VSUBS 0.02fF
C13407 S.n12102 VSUBS 0.24fF $ **FLOATING
C13408 S.n12103 VSUBS 0.91fF $ **FLOATING
C13409 S.n12104 VSUBS 0.05fF $ **FLOATING
C13410 S.n12105 VSUBS 1.88fF $ **FLOATING
C13411 S.n12106 VSUBS 0.12fF $ **FLOATING
C13412 S.t158 VSUBS 0.02fF
C13413 S.n12107 VSUBS 0.14fF $ **FLOATING
C13414 S.t984 VSUBS 0.02fF
C13415 S.n12109 VSUBS 0.24fF $ **FLOATING
C13416 S.n12110 VSUBS 0.36fF $ **FLOATING
C13417 S.n12111 VSUBS 0.61fF $ **FLOATING
C13418 S.n12112 VSUBS 2.67fF $ **FLOATING
C13419 S.n12113 VSUBS 5.17fF $ **FLOATING
C13420 S.t1039 VSUBS 0.02fF
C13421 S.n12114 VSUBS 0.12fF $ **FLOATING
C13422 S.n12115 VSUBS 0.14fF $ **FLOATING
C13423 S.t1268 VSUBS 0.02fF
C13424 S.n12117 VSUBS 0.24fF $ **FLOATING
C13425 S.n12118 VSUBS 0.91fF $ **FLOATING
C13426 S.n12119 VSUBS 0.05fF $ **FLOATING
C13427 S.n12120 VSUBS 1.88fF $ **FLOATING
C13428 S.n12121 VSUBS 2.67fF $ **FLOATING
C13429 S.t1766 VSUBS 0.02fF
C13430 S.n12122 VSUBS 0.24fF $ **FLOATING
C13431 S.n12123 VSUBS 0.36fF $ **FLOATING
C13432 S.n12124 VSUBS 0.61fF $ **FLOATING
C13433 S.n12125 VSUBS 0.12fF $ **FLOATING
C13434 S.t949 VSUBS 0.02fF
C13435 S.n12126 VSUBS 0.14fF $ **FLOATING
C13436 S.n12128 VSUBS 5.17fF $ **FLOATING
C13437 S.t1819 VSUBS 0.02fF
C13438 S.n12129 VSUBS 0.12fF $ **FLOATING
C13439 S.n12130 VSUBS 0.14fF $ **FLOATING
C13440 S.t2058 VSUBS 0.02fF
C13441 S.n12132 VSUBS 0.24fF $ **FLOATING
C13442 S.n12133 VSUBS 0.91fF $ **FLOATING
C13443 S.n12134 VSUBS 0.05fF $ **FLOATING
C13444 S.n12135 VSUBS 1.88fF $ **FLOATING
C13445 S.n12136 VSUBS 2.67fF $ **FLOATING
C13446 S.t146 VSUBS 0.02fF
C13447 S.n12137 VSUBS 0.24fF $ **FLOATING
C13448 S.n12138 VSUBS 0.36fF $ **FLOATING
C13449 S.n12139 VSUBS 0.61fF $ **FLOATING
C13450 S.n12140 VSUBS 0.12fF $ **FLOATING
C13451 S.t1862 VSUBS 0.02fF
C13452 S.n12141 VSUBS 0.14fF $ **FLOATING
C13453 S.n12143 VSUBS 5.17fF $ **FLOATING
C13454 S.t208 VSUBS 0.02fF
C13455 S.n12144 VSUBS 0.12fF $ **FLOATING
C13456 S.n12145 VSUBS 0.14fF $ **FLOATING
C13457 S.t442 VSUBS 0.02fF
C13458 S.n12147 VSUBS 0.24fF $ **FLOATING
C13459 S.n12148 VSUBS 0.91fF $ **FLOATING
C13460 S.n12149 VSUBS 0.05fF $ **FLOATING
C13461 S.n12150 VSUBS 1.88fF $ **FLOATING
C13462 S.n12151 VSUBS 2.67fF $ **FLOATING
C13463 S.t2282 VSUBS 0.02fF
C13464 S.n12152 VSUBS 0.24fF $ **FLOATING
C13465 S.n12153 VSUBS 0.36fF $ **FLOATING
C13466 S.n12154 VSUBS 0.61fF $ **FLOATING
C13467 S.n12155 VSUBS 0.12fF $ **FLOATING
C13468 S.t1467 VSUBS 0.02fF
C13469 S.n12156 VSUBS 0.14fF $ **FLOATING
C13470 S.n12158 VSUBS 5.17fF $ **FLOATING
C13471 S.t2334 VSUBS 0.02fF
C13472 S.n12159 VSUBS 0.12fF $ **FLOATING
C13473 S.n12160 VSUBS 0.14fF $ **FLOATING
C13474 S.t2570 VSUBS 0.02fF
C13475 S.n12162 VSUBS 0.24fF $ **FLOATING
C13476 S.n12163 VSUBS 0.91fF $ **FLOATING
C13477 S.n12164 VSUBS 0.05fF $ **FLOATING
C13478 S.n12165 VSUBS 1.88fF $ **FLOATING
C13479 S.n12166 VSUBS 2.67fF $ **FLOATING
C13480 S.t554 VSUBS 0.02fF
C13481 S.n12167 VSUBS 0.24fF $ **FLOATING
C13482 S.n12168 VSUBS 0.36fF $ **FLOATING
C13483 S.n12169 VSUBS 0.61fF $ **FLOATING
C13484 S.n12170 VSUBS 0.12fF $ **FLOATING
C13485 S.t2255 VSUBS 0.02fF
C13486 S.n12171 VSUBS 0.14fF $ **FLOATING
C13487 S.n12173 VSUBS 5.17fF $ **FLOATING
C13488 S.t598 VSUBS 0.02fF
C13489 S.n12174 VSUBS 0.12fF $ **FLOATING
C13490 S.n12175 VSUBS 0.14fF $ **FLOATING
C13491 S.t835 VSUBS 0.02fF
C13492 S.n12177 VSUBS 0.24fF $ **FLOATING
C13493 S.n12178 VSUBS 0.91fF $ **FLOATING
C13494 S.n12179 VSUBS 0.05fF $ **FLOATING
C13495 S.n12180 VSUBS 1.88fF $ **FLOATING
C13496 S.n12181 VSUBS 2.67fF $ **FLOATING
C13497 S.t1342 VSUBS 0.02fF
C13498 S.n12182 VSUBS 0.24fF $ **FLOATING
C13499 S.n12183 VSUBS 0.36fF $ **FLOATING
C13500 S.n12184 VSUBS 0.61fF $ **FLOATING
C13501 S.n12185 VSUBS 0.12fF $ **FLOATING
C13502 S.t523 VSUBS 0.02fF
C13503 S.n12186 VSUBS 0.14fF $ **FLOATING
C13504 S.n12188 VSUBS 5.17fF $ **FLOATING
C13505 S.t1391 VSUBS 0.02fF
C13506 S.n12189 VSUBS 0.12fF $ **FLOATING
C13507 S.n12190 VSUBS 0.14fF $ **FLOATING
C13508 S.t1618 VSUBS 0.02fF
C13509 S.n12192 VSUBS 0.24fF $ **FLOATING
C13510 S.n12193 VSUBS 0.91fF $ **FLOATING
C13511 S.n12194 VSUBS 0.05fF $ **FLOATING
C13512 S.n12195 VSUBS 1.88fF $ **FLOATING
C13513 S.n12196 VSUBS 2.67fF $ **FLOATING
C13514 S.t2129 VSUBS 0.02fF
C13515 S.n12197 VSUBS 0.24fF $ **FLOATING
C13516 S.n12198 VSUBS 0.36fF $ **FLOATING
C13517 S.n12199 VSUBS 0.61fF $ **FLOATING
C13518 S.n12200 VSUBS 0.12fF $ **FLOATING
C13519 S.t1311 VSUBS 0.02fF
C13520 S.n12201 VSUBS 0.14fF $ **FLOATING
C13521 S.n12203 VSUBS 5.17fF $ **FLOATING
C13522 S.t2181 VSUBS 0.02fF
C13523 S.n12204 VSUBS 0.12fF $ **FLOATING
C13524 S.n12205 VSUBS 0.14fF $ **FLOATING
C13525 S.t2404 VSUBS 0.02fF
C13526 S.n12207 VSUBS 0.24fF $ **FLOATING
C13527 S.n12208 VSUBS 0.91fF $ **FLOATING
C13528 S.n12209 VSUBS 0.05fF $ **FLOATING
C13529 S.n12210 VSUBS 1.88fF $ **FLOATING
C13530 S.n12211 VSUBS 2.67fF $ **FLOATING
C13531 S.t137 VSUBS 0.02fF
C13532 S.n12212 VSUBS 0.24fF $ **FLOATING
C13533 S.n12213 VSUBS 0.36fF $ **FLOATING
C13534 S.n12214 VSUBS 0.61fF $ **FLOATING
C13535 S.n12215 VSUBS 0.12fF $ **FLOATING
C13536 S.t358 VSUBS 0.02fF
C13537 S.n12216 VSUBS 0.14fF $ **FLOATING
C13538 S.n12218 VSUBS 5.17fF $ **FLOATING
C13539 S.t566 VSUBS 0.02fF
C13540 S.n12219 VSUBS 0.12fF $ **FLOATING
C13541 S.n12220 VSUBS 0.14fF $ **FLOATING
C13542 S.t993 VSUBS 0.02fF
C13543 S.n12222 VSUBS 0.24fF $ **FLOATING
C13544 S.n12223 VSUBS 0.91fF $ **FLOATING
C13545 S.n12224 VSUBS 0.05fF $ **FLOATING
C13546 S.n12225 VSUBS 1.88fF $ **FLOATING
C13547 S.n12226 VSUBS 2.67fF $ **FLOATING
C13548 S.t934 VSUBS 0.02fF
C13549 S.n12227 VSUBS 0.24fF $ **FLOATING
C13550 S.n12228 VSUBS 0.36fF $ **FLOATING
C13551 S.n12229 VSUBS 0.61fF $ **FLOATING
C13552 S.n12230 VSUBS 0.12fF $ **FLOATING
C13553 S.t1144 VSUBS 0.02fF
C13554 S.n12231 VSUBS 0.14fF $ **FLOATING
C13555 S.n12233 VSUBS 5.17fF $ **FLOATING
C13556 S.t2007 VSUBS 0.02fF
C13557 S.n12234 VSUBS 0.12fF $ **FLOATING
C13558 S.n12235 VSUBS 0.14fF $ **FLOATING
C13559 S.t1776 VSUBS 0.02fF
C13560 S.n12237 VSUBS 0.24fF $ **FLOATING
C13561 S.n12238 VSUBS 0.91fF $ **FLOATING
C13562 S.n12239 VSUBS 0.05fF $ **FLOATING
C13563 S.n12240 VSUBS 1.88fF $ **FLOATING
C13564 S.n12241 VSUBS 2.67fF $ **FLOATING
C13565 S.t1713 VSUBS 0.02fF
C13566 S.n12242 VSUBS 0.24fF $ **FLOATING
C13567 S.n12243 VSUBS 0.36fF $ **FLOATING
C13568 S.n12244 VSUBS 0.61fF $ **FLOATING
C13569 S.n12245 VSUBS 0.12fF $ **FLOATING
C13570 S.t1926 VSUBS 0.02fF
C13571 S.n12246 VSUBS 0.14fF $ **FLOATING
C13572 S.n12248 VSUBS 5.17fF $ **FLOATING
C13573 S.t277 VSUBS 0.02fF
C13574 S.n12249 VSUBS 0.12fF $ **FLOATING
C13575 S.n12250 VSUBS 0.14fF $ **FLOATING
C13576 S.t2556 VSUBS 0.02fF
C13577 S.n12252 VSUBS 0.24fF $ **FLOATING
C13578 S.n12253 VSUBS 0.91fF $ **FLOATING
C13579 S.n12254 VSUBS 0.05fF $ **FLOATING
C13580 S.n12255 VSUBS 1.88fF $ **FLOATING
C13581 S.n12256 VSUBS 2.67fF $ **FLOATING
C13582 S.t2501 VSUBS 0.02fF
C13583 S.n12257 VSUBS 0.24fF $ **FLOATING
C13584 S.n12258 VSUBS 0.36fF $ **FLOATING
C13585 S.n12259 VSUBS 0.61fF $ **FLOATING
C13586 S.n12260 VSUBS 0.12fF $ **FLOATING
C13587 S.t182 VSUBS 0.02fF
C13588 S.n12261 VSUBS 0.14fF $ **FLOATING
C13589 S.n12263 VSUBS 4.89fF $ **FLOATING
C13590 S.t1057 VSUBS 0.02fF
C13591 S.n12264 VSUBS 0.12fF $ **FLOATING
C13592 S.n12265 VSUBS 0.14fF $ **FLOATING
C13593 S.t821 VSUBS 0.02fF
C13594 S.n12267 VSUBS 0.24fF $ **FLOATING
C13595 S.n12268 VSUBS 0.91fF $ **FLOATING
C13596 S.n12269 VSUBS 0.05fF $ **FLOATING
C13597 S.n12270 VSUBS 0.11fF $ **FLOATING
C13598 S.n12271 VSUBS 0.12fF $ **FLOATING
C13599 S.n12272 VSUBS 0.09fF $ **FLOATING
C13600 S.n12273 VSUBS 0.12fF $ **FLOATING
C13601 S.n12274 VSUBS 0.18fF $ **FLOATING
C13602 S.n12275 VSUBS 1.88fF $ **FLOATING
C13603 S.n12276 VSUBS 0.12fF $ **FLOATING
C13604 S.t999 VSUBS 0.02fF
C13605 S.n12277 VSUBS 0.14fF $ **FLOATING
C13606 S.t1215 VSUBS 0.02fF
C13607 S.n12279 VSUBS 1.22fF $ **FLOATING
C13608 S.n12280 VSUBS 0.06fF $ **FLOATING
C13609 S.n12281 VSUBS 0.10fF $ **FLOATING
C13610 S.n12282 VSUBS 0.61fF $ **FLOATING
C13611 S.n12283 VSUBS 2.42fF $ **FLOATING
C13612 S.n12284 VSUBS 2.47fF $ **FLOATING
C13613 S.n12285 VSUBS 4.29fF $ **FLOATING
C13614 S.n12286 VSUBS 0.25fF $ **FLOATING
C13615 S.n12287 VSUBS 0.01fF $ **FLOATING
C13616 S.t392 VSUBS 0.02fF
C13617 S.n12288 VSUBS 0.26fF $ **FLOATING
C13618 S.t1484 VSUBS 0.02fF
C13619 S.n12289 VSUBS 0.95fF $ **FLOATING
C13620 S.n12290 VSUBS 0.71fF $ **FLOATING
C13621 S.n12291 VSUBS 1.89fF $ **FLOATING
C13622 S.n12292 VSUBS 1.88fF $ **FLOATING
C13623 S.t1993 VSUBS 0.02fF
C13624 S.n12293 VSUBS 0.24fF $ **FLOATING
C13625 S.n12294 VSUBS 0.36fF $ **FLOATING
C13626 S.n12295 VSUBS 0.61fF $ **FLOATING
C13627 S.n12296 VSUBS 0.12fF $ **FLOATING
C13628 S.t1185 VSUBS 0.02fF
C13629 S.n12297 VSUBS 0.14fF $ **FLOATING
C13630 S.n12299 VSUBS 1.16fF $ **FLOATING
C13631 S.n12300 VSUBS 0.22fF $ **FLOATING
C13632 S.n12301 VSUBS 0.25fF $ **FLOATING
C13633 S.n12302 VSUBS 0.09fF $ **FLOATING
C13634 S.n12303 VSUBS 1.88fF $ **FLOATING
C13635 S.t2268 VSUBS 0.02fF
C13636 S.n12304 VSUBS 0.24fF $ **FLOATING
C13637 S.n12305 VSUBS 0.91fF $ **FLOATING
C13638 S.n12306 VSUBS 0.05fF $ **FLOATING
C13639 S.t2046 VSUBS 0.02fF
C13640 S.n12307 VSUBS 0.12fF $ **FLOATING
C13641 S.n12308 VSUBS 0.14fF $ **FLOATING
C13642 S.n12310 VSUBS 0.77fF $ **FLOATING
C13643 S.n12311 VSUBS 0.44fF $ **FLOATING
C13644 S.n12312 VSUBS 1.58fF $ **FLOATING
C13645 S.n12313 VSUBS 0.12fF $ **FLOATING
C13646 S.t459 VSUBS 0.02fF
C13647 S.n12314 VSUBS 0.14fF $ **FLOATING
C13648 S.t265 VSUBS 0.02fF
C13649 S.n12316 VSUBS 0.24fF $ **FLOATING
C13650 S.n12317 VSUBS 0.36fF $ **FLOATING
C13651 S.n12318 VSUBS 0.61fF $ **FLOATING
C13652 S.n12319 VSUBS 0.01fF $ **FLOATING
C13653 S.n12320 VSUBS 0.07fF $ **FLOATING
C13654 S.n12321 VSUBS 0.01fF $ **FLOATING
C13655 S.n12322 VSUBS 0.02fF $ **FLOATING
C13656 S.n12323 VSUBS 0.01fF $ **FLOATING
C13657 S.n12324 VSUBS 0.24fF $ **FLOATING
C13658 S.n12325 VSUBS 1.16fF $ **FLOATING
C13659 S.n12326 VSUBS 1.34fF $ **FLOATING
C13660 S.n12327 VSUBS 1.99fF $ **FLOATING
C13661 S.t1646 VSUBS 0.02fF
C13662 S.n12328 VSUBS 0.24fF $ **FLOATING
C13663 S.n12329 VSUBS 0.91fF $ **FLOATING
C13664 S.n12330 VSUBS 0.05fF $ **FLOATING
C13665 S.t107 VSUBS 0.02fF
C13666 S.n12331 VSUBS 0.12fF $ **FLOATING
C13667 S.n12332 VSUBS 0.14fF $ **FLOATING
C13668 S.n12334 VSUBS 1.88fF $ **FLOATING
C13669 S.n12335 VSUBS 0.12fF $ **FLOATING
C13670 S.t2087 VSUBS 0.02fF
C13671 S.n12336 VSUBS 0.14fF $ **FLOATING
C13672 S.t264 VSUBS 0.02fF
C13673 S.n12338 VSUBS 0.24fF $ **FLOATING
C13674 S.n12339 VSUBS 0.36fF $ **FLOATING
C13675 S.n12340 VSUBS 0.61fF $ **FLOATING
C13676 S.n12341 VSUBS 0.32fF $ **FLOATING
C13677 S.n12342 VSUBS 1.09fF $ **FLOATING
C13678 S.n12343 VSUBS 0.15fF $ **FLOATING
C13679 S.n12344 VSUBS 2.10fF $ **FLOATING
C13680 S.t314 VSUBS 0.02fF
C13681 S.n12345 VSUBS 0.12fF $ **FLOATING
C13682 S.n12346 VSUBS 0.14fF $ **FLOATING
C13683 S.t539 VSUBS 0.02fF
C13684 S.n12348 VSUBS 0.24fF $ **FLOATING
C13685 S.n12349 VSUBS 0.91fF $ **FLOATING
C13686 S.n12350 VSUBS 0.05fF $ **FLOATING
C13687 S.n12351 VSUBS 1.88fF $ **FLOATING
C13688 S.n12352 VSUBS 2.67fF $ **FLOATING
C13689 S.t1171 VSUBS 0.02fF
C13690 S.n12353 VSUBS 0.24fF $ **FLOATING
C13691 S.n12354 VSUBS 0.36fF $ **FLOATING
C13692 S.n12355 VSUBS 0.61fF $ **FLOATING
C13693 S.n12356 VSUBS 0.12fF $ **FLOATING
C13694 S.t361 VSUBS 0.02fF
C13695 S.n12357 VSUBS 0.14fF $ **FLOATING
C13696 S.n12359 VSUBS 2.30fF $ **FLOATING
C13697 S.t1229 VSUBS 0.02fF
C13698 S.n12360 VSUBS 0.12fF $ **FLOATING
C13699 S.n12361 VSUBS 0.14fF $ **FLOATING
C13700 S.t1448 VSUBS 0.02fF
C13701 S.n12363 VSUBS 0.24fF $ **FLOATING
C13702 S.n12364 VSUBS 0.91fF $ **FLOATING
C13703 S.n12365 VSUBS 0.05fF $ **FLOATING
C13704 S.n12366 VSUBS 1.88fF $ **FLOATING
C13705 S.n12367 VSUBS 2.67fF $ **FLOATING
C13706 S.t766 VSUBS 0.02fF
C13707 S.n12368 VSUBS 0.24fF $ **FLOATING
C13708 S.n12369 VSUBS 0.36fF $ **FLOATING
C13709 S.n12370 VSUBS 0.61fF $ **FLOATING
C13710 S.n12371 VSUBS 0.12fF $ **FLOATING
C13711 S.t2475 VSUBS 0.02fF
C13712 S.n12372 VSUBS 0.14fF $ **FLOATING
C13713 S.n12374 VSUBS 2.80fF $ **FLOATING
C13714 S.n12375 VSUBS 2.30fF $ **FLOATING
C13715 S.t822 VSUBS 0.02fF
C13716 S.n12376 VSUBS 0.12fF $ **FLOATING
C13717 S.n12377 VSUBS 0.14fF $ **FLOATING
C13718 S.t1069 VSUBS 0.02fF
C13719 S.n12379 VSUBS 0.24fF $ **FLOATING
C13720 S.n12380 VSUBS 0.91fF $ **FLOATING
C13721 S.n12381 VSUBS 0.05fF $ **FLOATING
C13722 S.n12382 VSUBS 2.80fF $ **FLOATING
C13723 S.n12383 VSUBS 1.88fF $ **FLOATING
C13724 S.n12384 VSUBS 0.12fF $ **FLOATING
C13725 S.t734 VSUBS 0.02fF
C13726 S.n12385 VSUBS 0.14fF $ **FLOATING
C13727 S.t1555 VSUBS 0.02fF
C13728 S.n12387 VSUBS 0.24fF $ **FLOATING
C13729 S.n12388 VSUBS 0.36fF $ **FLOATING
C13730 S.n12389 VSUBS 0.61fF $ **FLOATING
C13731 S.n12390 VSUBS 2.67fF $ **FLOATING
C13732 S.n12391 VSUBS 2.30fF $ **FLOATING
C13733 S.t1604 VSUBS 0.02fF
C13734 S.n12392 VSUBS 0.12fF $ **FLOATING
C13735 S.n12393 VSUBS 0.14fF $ **FLOATING
C13736 S.t1855 VSUBS 0.02fF
C13737 S.n12395 VSUBS 0.24fF $ **FLOATING
C13738 S.n12396 VSUBS 0.91fF $ **FLOATING
C13739 S.n12397 VSUBS 0.05fF $ **FLOATING
C13740 S.n12398 VSUBS 1.88fF $ **FLOATING
C13741 S.n12399 VSUBS 2.67fF $ **FLOATING
C13742 S.t2343 VSUBS 0.02fF
C13743 S.n12400 VSUBS 0.24fF $ **FLOATING
C13744 S.n12401 VSUBS 0.36fF $ **FLOATING
C13745 S.n12402 VSUBS 0.61fF $ **FLOATING
C13746 S.n12403 VSUBS 0.12fF $ **FLOATING
C13747 S.t1525 VSUBS 0.02fF
C13748 S.n12404 VSUBS 0.14fF $ **FLOATING
C13749 S.n12406 VSUBS 2.80fF $ **FLOATING
C13750 S.n12407 VSUBS 2.30fF $ **FLOATING
C13751 S.t2393 VSUBS 0.02fF
C13752 S.n12408 VSUBS 0.12fF $ **FLOATING
C13753 S.n12409 VSUBS 0.14fF $ **FLOATING
C13754 S.t86 VSUBS 0.02fF
C13755 S.n12411 VSUBS 0.24fF $ **FLOATING
C13756 S.n12412 VSUBS 0.91fF $ **FLOATING
C13757 S.n12413 VSUBS 0.05fF $ **FLOATING
C13758 S.n12414 VSUBS 1.88fF $ **FLOATING
C13759 S.n12415 VSUBS 2.67fF $ **FLOATING
C13760 S.t605 VSUBS 0.02fF
C13761 S.n12416 VSUBS 0.24fF $ **FLOATING
C13762 S.n12417 VSUBS 0.36fF $ **FLOATING
C13763 S.n12418 VSUBS 0.61fF $ **FLOATING
C13764 S.n12419 VSUBS 0.12fF $ **FLOATING
C13765 S.t2433 VSUBS 0.02fF
C13766 S.n12420 VSUBS 0.14fF $ **FLOATING
C13767 S.n12422 VSUBS 2.80fF $ **FLOATING
C13768 S.n12423 VSUBS 2.30fF $ **FLOATING
C13769 S.t656 VSUBS 0.02fF
C13770 S.n12424 VSUBS 0.12fF $ **FLOATING
C13771 S.n12425 VSUBS 0.14fF $ **FLOATING
C13772 S.t895 VSUBS 0.02fF
C13773 S.n12427 VSUBS 0.24fF $ **FLOATING
C13774 S.n12428 VSUBS 0.91fF $ **FLOATING
C13775 S.n12429 VSUBS 0.05fF $ **FLOATING
C13776 S.n12430 VSUBS 1.88fF $ **FLOATING
C13777 S.n12431 VSUBS 2.67fF $ **FLOATING
C13778 S.t359 VSUBS 0.02fF
C13779 S.n12432 VSUBS 0.24fF $ **FLOATING
C13780 S.n12433 VSUBS 0.36fF $ **FLOATING
C13781 S.n12434 VSUBS 0.61fF $ **FLOATING
C13782 S.n12435 VSUBS 0.12fF $ **FLOATING
C13783 S.t2061 VSUBS 0.02fF
C13784 S.n12436 VSUBS 0.14fF $ **FLOATING
C13785 S.n12438 VSUBS 2.80fF $ **FLOATING
C13786 S.n12439 VSUBS 2.30fF $ **FLOATING
C13787 S.t1564 VSUBS 0.02fF
C13788 S.n12440 VSUBS 0.12fF $ **FLOATING
C13789 S.n12441 VSUBS 0.14fF $ **FLOATING
C13790 S.t628 VSUBS 0.02fF
C13791 S.n12443 VSUBS 0.24fF $ **FLOATING
C13792 S.n12444 VSUBS 0.91fF $ **FLOATING
C13793 S.n12445 VSUBS 0.05fF $ **FLOATING
C13794 S.n12446 VSUBS 1.88fF $ **FLOATING
C13795 S.n12447 VSUBS 2.67fF $ **FLOATING
C13796 S.t1145 VSUBS 0.02fF
C13797 S.n12448 VSUBS 0.24fF $ **FLOATING
C13798 S.n12449 VSUBS 0.36fF $ **FLOATING
C13799 S.n12450 VSUBS 0.61fF $ **FLOATING
C13800 S.n12451 VSUBS 0.12fF $ **FLOATING
C13801 S.t326 VSUBS 0.02fF
C13802 S.n12452 VSUBS 0.14fF $ **FLOATING
C13803 S.n12454 VSUBS 2.80fF $ **FLOATING
C13804 S.n12455 VSUBS 2.30fF $ **FLOATING
C13805 S.t1199 VSUBS 0.02fF
C13806 S.n12456 VSUBS 0.12fF $ **FLOATING
C13807 S.n12457 VSUBS 0.14fF $ **FLOATING
C13808 S.t1418 VSUBS 0.02fF
C13809 S.n12459 VSUBS 0.24fF $ **FLOATING
C13810 S.n12460 VSUBS 0.91fF $ **FLOATING
C13811 S.n12461 VSUBS 0.05fF $ **FLOATING
C13812 S.n12462 VSUBS 1.88fF $ **FLOATING
C13813 S.n12463 VSUBS 2.67fF $ **FLOATING
C13814 S.t1927 VSUBS 0.02fF
C13815 S.n12464 VSUBS 0.24fF $ **FLOATING
C13816 S.n12465 VSUBS 0.36fF $ **FLOATING
C13817 S.n12466 VSUBS 0.61fF $ **FLOATING
C13818 S.n12467 VSUBS 0.12fF $ **FLOATING
C13819 S.t1115 VSUBS 0.02fF
C13820 S.n12468 VSUBS 0.14fF $ **FLOATING
C13821 S.n12470 VSUBS 2.80fF $ **FLOATING
C13822 S.n12471 VSUBS 2.30fF $ **FLOATING
C13823 S.t1979 VSUBS 0.02fF
C13824 S.n12472 VSUBS 0.12fF $ **FLOATING
C13825 S.n12473 VSUBS 0.14fF $ **FLOATING
C13826 S.t2207 VSUBS 0.02fF
C13827 S.n12475 VSUBS 0.24fF $ **FLOATING
C13828 S.n12476 VSUBS 0.91fF $ **FLOATING
C13829 S.n12477 VSUBS 0.05fF $ **FLOATING
C13830 S.n12478 VSUBS 1.88fF $ **FLOATING
C13831 S.n12479 VSUBS 2.67fF $ **FLOATING
C13832 S.t183 VSUBS 0.02fF
C13833 S.n12480 VSUBS 0.24fF $ **FLOATING
C13834 S.n12481 VSUBS 0.36fF $ **FLOATING
C13835 S.n12482 VSUBS 0.61fF $ **FLOATING
C13836 S.n12483 VSUBS 0.12fF $ **FLOATING
C13837 S.t1897 VSUBS 0.02fF
C13838 S.n12484 VSUBS 0.14fF $ **FLOATING
C13839 S.n12486 VSUBS 2.80fF $ **FLOATING
C13840 S.n12487 VSUBS 2.30fF $ **FLOATING
C13841 S.t243 VSUBS 0.02fF
C13842 S.n12488 VSUBS 0.12fF $ **FLOATING
C13843 S.n12489 VSUBS 0.14fF $ **FLOATING
C13844 S.t474 VSUBS 0.02fF
C13845 S.n12491 VSUBS 0.24fF $ **FLOATING
C13846 S.n12492 VSUBS 0.91fF $ **FLOATING
C13847 S.n12493 VSUBS 0.05fF $ **FLOATING
C13848 S.n12494 VSUBS 1.88fF $ **FLOATING
C13849 S.n12495 VSUBS 2.67fF $ **FLOATING
C13850 S.t974 VSUBS 0.02fF
C13851 S.n12496 VSUBS 0.24fF $ **FLOATING
C13852 S.n12497 VSUBS 0.36fF $ **FLOATING
C13853 S.n12498 VSUBS 0.61fF $ **FLOATING
C13854 S.n12499 VSUBS 0.12fF $ **FLOATING
C13855 S.t292 VSUBS 0.02fF
C13856 S.n12500 VSUBS 0.14fF $ **FLOATING
C13857 S.n12502 VSUBS 2.80fF $ **FLOATING
C13858 S.n12503 VSUBS 2.30fF $ **FLOATING
C13859 S.t1030 VSUBS 0.02fF
C13860 S.n12504 VSUBS 0.12fF $ **FLOATING
C13861 S.n12505 VSUBS 0.14fF $ **FLOATING
C13862 S.t1263 VSUBS 0.02fF
C13863 S.n12507 VSUBS 0.24fF $ **FLOATING
C13864 S.n12508 VSUBS 0.91fF $ **FLOATING
C13865 S.n12509 VSUBS 0.05fF $ **FLOATING
C13866 S.n12510 VSUBS 1.88fF $ **FLOATING
C13867 S.n12511 VSUBS 2.67fF $ **FLOATING
C13868 S.t958 VSUBS 0.02fF
C13869 S.n12512 VSUBS 0.24fF $ **FLOATING
C13870 S.n12513 VSUBS 0.36fF $ **FLOATING
C13871 S.n12514 VSUBS 0.61fF $ **FLOATING
C13872 S.n12515 VSUBS 0.12fF $ **FLOATING
C13873 S.t1165 VSUBS 0.02fF
C13874 S.n12516 VSUBS 0.14fF $ **FLOATING
C13875 S.n12518 VSUBS 2.80fF $ **FLOATING
C13876 S.n12519 VSUBS 2.30fF $ **FLOATING
C13877 S.t2028 VSUBS 0.02fF
C13878 S.n12520 VSUBS 0.12fF $ **FLOATING
C13879 S.n12521 VSUBS 0.14fF $ **FLOATING
C13880 S.t1799 VSUBS 0.02fF
C13881 S.n12523 VSUBS 0.24fF $ **FLOATING
C13882 S.n12524 VSUBS 0.91fF $ **FLOATING
C13883 S.n12525 VSUBS 0.05fF $ **FLOATING
C13884 S.n12526 VSUBS 1.88fF $ **FLOATING
C13885 S.n12527 VSUBS 2.67fF $ **FLOATING
C13886 S.t1740 VSUBS 0.02fF
C13887 S.n12528 VSUBS 0.24fF $ **FLOATING
C13888 S.n12529 VSUBS 0.36fF $ **FLOATING
C13889 S.n12530 VSUBS 0.61fF $ **FLOATING
C13890 S.n12531 VSUBS 0.12fF $ **FLOATING
C13891 S.t1952 VSUBS 0.02fF
C13892 S.n12532 VSUBS 0.14fF $ **FLOATING
C13893 S.n12534 VSUBS 2.80fF $ **FLOATING
C13894 S.n12535 VSUBS 2.30fF $ **FLOATING
C13895 S.t299 VSUBS 0.02fF
C13896 S.n12536 VSUBS 0.12fF $ **FLOATING
C13897 S.n12537 VSUBS 0.14fF $ **FLOATING
C13898 S.t1 VSUBS 0.02fF
C13899 S.n12539 VSUBS 0.24fF $ **FLOATING
C13900 S.n12540 VSUBS 0.91fF $ **FLOATING
C13901 S.n12541 VSUBS 0.05fF $ **FLOATING
C13902 S.n12542 VSUBS 1.88fF $ **FLOATING
C13903 S.n12543 VSUBS 2.67fF $ **FLOATING
C13904 S.t2524 VSUBS 0.02fF
C13905 S.n12544 VSUBS 0.24fF $ **FLOATING
C13906 S.n12545 VSUBS 0.36fF $ **FLOATING
C13907 S.n12546 VSUBS 0.61fF $ **FLOATING
C13908 S.n12547 VSUBS 0.12fF $ **FLOATING
C13909 S.t210 VSUBS 0.02fF
C13910 S.n12548 VSUBS 0.14fF $ **FLOATING
C13911 S.n12550 VSUBS 2.80fF $ **FLOATING
C13912 S.n12551 VSUBS 2.30fF $ **FLOATING
C13913 S.t1084 VSUBS 0.02fF
C13914 S.n12552 VSUBS 0.12fF $ **FLOATING
C13915 S.n12553 VSUBS 0.14fF $ **FLOATING
C13916 S.t845 VSUBS 0.02fF
C13917 S.n12555 VSUBS 0.24fF $ **FLOATING
C13918 S.n12556 VSUBS 0.91fF $ **FLOATING
C13919 S.n12557 VSUBS 0.05fF $ **FLOATING
C13920 S.t106 VSUBS 48.27fF
C13921 S.t1866 VSUBS 0.02fF
C13922 S.n12558 VSUBS 0.12fF $ **FLOATING
C13923 S.n12559 VSUBS 0.14fF $ **FLOATING
C13924 S.t1630 VSUBS 0.02fF
C13925 S.n12561 VSUBS 0.24fF $ **FLOATING
C13926 S.n12562 VSUBS 0.91fF $ **FLOATING
C13927 S.n12563 VSUBS 0.05fF $ **FLOATING
C13928 S.t785 VSUBS 0.02fF
C13929 S.n12564 VSUBS 0.24fF $ **FLOATING
C13930 S.n12565 VSUBS 0.36fF $ **FLOATING
C13931 S.n12566 VSUBS 0.61fF $ **FLOATING
C13932 S.n12567 VSUBS 2.66fF $ **FLOATING
C13933 S.n12568 VSUBS 3.27fF $ **FLOATING
C13934 S.n12569 VSUBS 0.11fF $ **FLOATING
C13935 S.n12570 VSUBS 0.36fF $ **FLOATING
C13936 S.n12571 VSUBS 0.47fF $ **FLOATING
C13937 S.n12572 VSUBS 1.14fF $ **FLOATING
C13938 S.n12573 VSUBS 1.87fF $ **FLOATING
C13939 S.n12574 VSUBS 0.12fF $ **FLOATING
C13940 S.t973 VSUBS 0.02fF
C13941 S.n12575 VSUBS 0.14fF $ **FLOATING
C13942 S.t759 VSUBS 0.02fF
C13943 S.n12577 VSUBS 0.24fF $ **FLOATING
C13944 S.n12578 VSUBS 0.36fF $ **FLOATING
C13945 S.n12579 VSUBS 0.61fF $ **FLOATING
C13946 S.n12580 VSUBS 1.27fF $ **FLOATING
C13947 S.n12581 VSUBS 2.38fF $ **FLOATING
C13948 S.n12582 VSUBS 4.20fF $ **FLOATING
C13949 S.t1842 VSUBS 0.02fF
C13950 S.n12583 VSUBS 0.12fF $ **FLOATING
C13951 S.n12584 VSUBS 0.14fF $ **FLOATING
C13952 S.t1603 VSUBS 0.02fF
C13953 S.n12586 VSUBS 0.24fF $ **FLOATING
C13954 S.n12587 VSUBS 0.91fF $ **FLOATING
C13955 S.n12588 VSUBS 0.05fF $ **FLOATING
C13956 S.t157 VSUBS 47.89fF
C13957 S.t1825 VSUBS 0.02fF
C13958 S.n12589 VSUBS 0.01fF $ **FLOATING
C13959 S.n12590 VSUBS 0.26fF $ **FLOATING
C13960 S.t1782 VSUBS 0.02fF
C13961 S.n12592 VSUBS 1.19fF $ **FLOATING
C13962 S.n12593 VSUBS 0.05fF $ **FLOATING
C13963 S.t1492 VSUBS 0.02fF
C13964 S.n12594 VSUBS 0.64fF $ **FLOATING
C13965 S.n12595 VSUBS 0.61fF $ **FLOATING
C13966 S.n12596 VSUBS 1.50fF $ **FLOATING
C13967 S.n12597 VSUBS 0.02fF $ **FLOATING
C13968 S.n12598 VSUBS 0.01fF $ **FLOATING
C13969 S.n12599 VSUBS 0.01fF $ **FLOATING
C13970 S.n12600 VSUBS 0.01fF $ **FLOATING
C13971 S.n12601 VSUBS 0.01fF $ **FLOATING
C13972 S.n12602 VSUBS 0.02fF $ **FLOATING
C13973 S.n12603 VSUBS 0.03fF $ **FLOATING
C13974 S.n12604 VSUBS 0.04fF $ **FLOATING
C13975 S.n12605 VSUBS 0.16fF $ **FLOATING
C13976 S.n12606 VSUBS 0.10fF $ **FLOATING
C13977 S.n12607 VSUBS 0.17fF $ **FLOATING
C13978 S.n12608 VSUBS 0.15fF $ **FLOATING
C13979 S.n12609 VSUBS 0.28fF $ **FLOATING
C13980 S.n12610 VSUBS 0.24fF $ **FLOATING
C13981 S.n12611 VSUBS 4.69fF $ **FLOATING
C13982 S.n12612 VSUBS 9.29fF $ **FLOATING
C13983 S.n12613 VSUBS 9.29fF $ **FLOATING
C13984 S.n12614 VSUBS 9.29fF $ **FLOATING
C13985 S.n12615 VSUBS 9.29fF $ **FLOATING
C13986 S.n12616 VSUBS 9.29fF $ **FLOATING
C13987 S.n12617 VSUBS 9.29fF $ **FLOATING
C13988 S.n12618 VSUBS 9.29fF $ **FLOATING
C13989 S.n12619 VSUBS 9.29fF $ **FLOATING
C13990 S.n12620 VSUBS 9.29fF $ **FLOATING
C13991 S.n12621 VSUBS 9.29fF $ **FLOATING
C13992 S.n12622 VSUBS 9.29fF $ **FLOATING
C13993 S.n12623 VSUBS 9.29fF $ **FLOATING
C13994 S.n12624 VSUBS 9.28fF $ **FLOATING
C13995 S.n12625 VSUBS 9.29fF $ **FLOATING
C13996 S.n12626 VSUBS 9.35fF $ **FLOATING
C13997 S.n12627 VSUBS 12.13fF $ **FLOATING
.ends

