* NGSPICE file created from mag_files/POSTLAYOUT/power_stage_flat.ext - technology: sky130A

.subckt power_stage_flat s1 s2 s3 s4 fc1 fc2 out VP VN
X0 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7 VN.t2590 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11 VN.t2589 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X15 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X16 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X17 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X18 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X19 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X20 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X21 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X22 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X23 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X24 fc2 s4 VN.t2588 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X25 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X26 VN.t2587 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X27 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X28 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X29 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X30 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X31 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X32 fc2 s4 VN.t2586 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X33 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X34 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X35 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X36 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X37 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X38 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X39 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X40 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X41 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X42 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X43 VN.t2585 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X44 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X45 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X46 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X47 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X48 VN.t2584 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X49 VN.t2583 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X50 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X51 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X52 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X53 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X54 VN.t2582 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X55 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X56 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X57 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X58 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X59 VN.t2581 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X60 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X61 VN.t2580 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X62 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X63 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X64 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X65 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X66 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X67 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X68 fc2 s4 VN.t2579 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X69 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X70 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X71 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X72 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X73 VN.t2578 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X74 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X75 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X76 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X77 VN.t2577 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X78 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X79 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X80 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X81 fc2 s4 VN.t2576 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X82 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X83 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X84 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X85 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X86 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X87 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X88 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X89 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X90 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X91 fc2 s4 VN.t2575 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X92 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X93 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X94 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X95 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X96 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X97 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X98 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X99 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X100 VN.t2574 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X101 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X102 VN.t2573 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X103 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X104 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X105 fc2 s4 VN.t2572 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X106 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X107 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X108 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X109 fc2 s4 VN.t2571 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X110 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X111 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X112 VN.t2570 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X113 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X114 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X115 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X116 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X117 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X119 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X120 fc2 s4 VN.t2569 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X121 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X122 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X123 VN.t2568 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X124 fc2 s4 VN.t2567 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X125 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X126 VN.t2566 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X127 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X128 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X129 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X130 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X131 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X132 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X133 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X134 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X136 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X137 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X138 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X139 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X140 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X141 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X142 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X143 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X144 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X145 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X146 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X147 fc2 s4 VN.t2565 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X148 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X149 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X150 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X151 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X152 VN.t2564 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X153 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X154 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X155 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X156 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X157 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X158 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X159 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X160 VN.t2563 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X161 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X162 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X163 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X164 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X165 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X166 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X167 VN.t2562 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X168 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X169 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X170 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X171 fc2 s4 VN.t2561 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X172 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X173 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X174 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X175 fc2 s4 VN.t2560 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X176 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X177 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X178 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X180 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X181 VN.t2559 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X182 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X183 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X184 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X185 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X186 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X187 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X188 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X189 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X190 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X191 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X192 fc2 s4 VN.t2558 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X193 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X194 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X195 VN.t2557 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X196 VN.t2556 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X197 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X198 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X199 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X200 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X201 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X202 VN.t2555 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X203 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X204 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X205 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X206 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X208 VN.t2554 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X209 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X210 VN.t2553 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X211 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X212 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X213 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X214 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X215 fc2 s4 VN.t2552 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X216 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X217 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X218 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X219 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X220 VN.t2551 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X221 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X222 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X223 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X224 VN.t2550 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X225 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X226 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X227 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X228 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X229 fc2 s4 VN.t2549 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X230 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X231 fc2 s4 VN.t2548 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X232 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X234 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X235 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X236 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X237 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X238 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X239 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X240 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X241 VN.t2547 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X242 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X243 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X244 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X245 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X246 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X247 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X248 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X249 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X250 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X251 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X252 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X253 VN.t2546 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X254 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X255 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X256 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X257 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X258 fc2 s4 VN.t2545 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X259 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X260 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X261 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X262 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X263 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X264 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X265 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X266 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X267 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X268 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X269 VN.t2544 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X270 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X271 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X272 VN.t2543 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X273 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X274 fc2 s4 VN.t2542 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X275 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X276 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X278 VN.t2541 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X279 VN.t2540 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X280 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X281 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X282 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X283 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X284 VN.t2539 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X285 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X286 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X287 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X288 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X289 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X290 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X291 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X292 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X293 fc2 s4 VN.t2538 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X295 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X296 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X297 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X298 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X299 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X300 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X301 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X302 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X303 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X304 fc2 s4 VN.t2537 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X305 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X306 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X307 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X308 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X309 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X310 VN.t2536 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X311 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X312 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X313 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X314 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X315 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X316 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X317 VN.t2535 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X318 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X319 fc2 s4 VN.t2534 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X320 VN.t2533 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X321 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X322 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X323 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X324 fc2 s4 VN.t2532 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X325 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X326 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X327 fc2 s4 VN.t2531 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X328 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X329 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X330 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X331 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X332 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X333 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X334 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X335 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X336 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X337 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X338 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X339 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X340 VN.t2530 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X341 fc2 s4 VN.t2529 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X342 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X343 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X344 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X345 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X346 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X347 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X348 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X349 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X350 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X351 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X352 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X353 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X354 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X355 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X356 fc2 s4 VN.t2528 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X357 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X358 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X359 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X360 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X361 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X362 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X363 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X364 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X365 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X366 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X367 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X368 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X369 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X370 fc2 s4 VN.t2527 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X372 fc2 s4 VN.t2526 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X373 VN.t2525 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X374 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X375 VN.t2524 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X376 VN.t2523 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X377 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X378 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X379 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X380 fc2 s4 VN.t2522 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X381 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X382 fc2 s4 VN.t2521 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X383 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X384 fc2 s4 VN.t2520 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X385 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X386 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X387 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X388 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X389 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X390 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X391 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X392 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X393 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X394 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X395 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X396 fc2 s4 VN.t2519 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X397 fc2 s4 VN.t2518 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X398 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X399 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X400 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X401 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X402 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X403 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X404 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X405 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X406 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X407 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X408 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X409 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X410 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X411 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X412 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X413 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X414 fc2 s4 VN.t2517 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X415 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X416 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X417 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X418 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X419 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X420 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X421 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X422 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X423 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X424 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X425 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X426 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X427 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X428 VN.t2516 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X429 fc2 s4 VN.t2515 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X430 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X431 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X432 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X433 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X434 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X435 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X436 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X437 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X438 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X439 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X440 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X441 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X442 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X443 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X444 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X445 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X446 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X447 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X448 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X449 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X450 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X451 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X452 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X453 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X454 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X455 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X456 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X457 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X458 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X459 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X460 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X461 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X462 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X463 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X464 VN.t2514 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X465 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X466 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X467 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X468 fc2 s4 VN.t2513 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X469 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X470 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X471 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X472 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X473 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X474 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X475 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X476 VN.t2512 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X477 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X478 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X479 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X480 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X481 fc2 s4 VN.t2511 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X482 fc2 s4 VN.t2510 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X483 fc2 s4 VN.t2509 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X484 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X485 VN.t2508 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X486 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X487 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X488 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X489 fc2 s4 VN.t2507 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X490 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X491 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X492 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X493 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X494 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X495 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X496 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X497 fc2 s4 VN.t2506 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X498 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X499 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X500 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X502 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X503 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X504 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X505 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X506 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X507 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X508 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X509 fc2 s4 VN.t2505 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X510 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X511 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X512 VN.t2504 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X513 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X514 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X515 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X516 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X517 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X518 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X519 fc2 s4 VN.t2503 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X520 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X521 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X522 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X523 VN.t2502 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X524 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X525 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X526 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X527 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X528 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X529 VN.t2501 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X530 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X531 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X532 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X533 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X534 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X535 fc2 s4 VN.t2500 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X536 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X537 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X538 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X539 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X540 fc2 s4 VN.t2499 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X541 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X542 fc2 s4 VN.t2498 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X543 fc2 s4 VN.t2497 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X544 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X545 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X546 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X547 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X548 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X549 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X550 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X551 VN.t2496 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X552 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X553 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X554 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X555 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X556 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X557 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X558 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X559 VN.t2495 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X560 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X561 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X562 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X563 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X564 VN.t2494 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X565 fc2 s4 VN.t2493 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X566 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X567 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X568 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X569 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X570 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X571 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X572 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X573 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X574 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X575 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X576 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X577 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X578 VN.t2492 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X579 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X580 fc2 s4 VN.t2491 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X581 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X582 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X583 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X584 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X585 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X586 VN.t2490 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X587 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X588 VN.t2489 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X590 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X591 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X592 fc2 s4 VN.t2488 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X593 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X594 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X595 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X596 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X597 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X598 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X599 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X600 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X601 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X602 VN.t2487 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X603 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X604 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X605 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X606 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X607 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X608 fc2 s4 VN.t2486 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X609 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X610 VN.t2485 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X611 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X612 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X613 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X614 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X615 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X616 fc2 s4 VN.t2484 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X617 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X618 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X619 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X620 fc2 s4 VN.t2483 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X622 fc2 s4 VN.t2482 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X623 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X624 fc2 s4 VN.t2481 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X625 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X626 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X627 VN.t2480 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X628 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X629 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X630 VN.t2479 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X631 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X632 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X633 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X634 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X635 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X636 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X637 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X638 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X639 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X640 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X641 fc2 s4 VN.t2478 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X643 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X644 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X645 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X646 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X647 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X648 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X649 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X650 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X651 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X652 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X653 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X654 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X655 fc2 s4 VN.t2477 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X656 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X657 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X658 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X659 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X660 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X661 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X663 VN.t2476 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X664 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X665 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X666 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X667 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X668 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X669 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X670 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X671 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X672 fc2 s4 VN.t2475 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X673 fc2 s4 VN.t2474 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X674 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X675 VN.t2473 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X676 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X677 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X678 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X679 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X680 VN.t2472 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X681 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X682 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X683 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X684 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X685 fc2 s4 VN.t2471 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X686 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X687 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X688 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X689 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X690 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X691 VN.t2470 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X692 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X693 VN.t2469 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X694 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X695 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X696 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X697 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X698 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X699 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X700 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X701 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X702 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X703 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X704 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X705 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X706 fc2 s4 VN.t2468 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X707 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X708 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X709 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X710 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X711 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X712 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X713 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X714 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X715 VN.t2467 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X716 VN.t2466 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X717 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X718 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X719 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X720 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X721 VN.t2465 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X722 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X723 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X724 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X725 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X726 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X727 VN.t2464 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X728 fc2 s4 VN.t2463 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X729 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X730 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X731 VN.t2462 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X732 fc2 s4 VN.t2461 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X733 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X734 fc2 s4 VN.t2460 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X735 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X736 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X737 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X739 fc2 s4 VN.t2459 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X740 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X741 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X742 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X743 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X744 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X745 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X746 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X747 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X748 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X749 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X750 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X751 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X752 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X753 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X754 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X755 VN.t2458 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X756 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X757 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X758 fc2 s4 VN.t2457 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X760 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X761 fc2 s4 VN.t2456 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X762 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X763 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X764 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X765 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X766 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X767 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X768 fc2 s4 VN.t2455 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X769 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X770 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X771 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X772 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X773 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X774 fc2 s4 VN.t2454 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X775 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X776 VN.t2453 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X777 fc2 s4 VN.t2452 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X778 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X779 fc2 s4 VN.t2451 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X780 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X781 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X782 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X783 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X784 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X785 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X786 fc2 s4 VN.t2450 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X787 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X788 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X789 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X790 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X791 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X792 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X793 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X794 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X795 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X796 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X797 fc2 s4 VN.t2449 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X798 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X799 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X800 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X801 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X802 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X803 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X804 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X805 VN.t2448 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X806 fc2 s4 VN.t2447 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X807 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X808 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X809 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X810 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X811 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X812 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X813 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X814 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X815 fc2 s4 VN.t2446 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X816 fc2 s4 VN.t2445 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X817 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X818 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X819 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X820 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X821 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X822 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X823 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X824 fc2 s4 VN.t2444 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X825 fc2 s4 VN.t2443 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X826 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X827 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X828 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X829 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X830 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X831 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X832 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X833 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X834 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X835 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X836 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X837 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X838 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X839 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X840 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X841 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X842 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X843 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X844 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X845 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X846 fc2 s4 VN.t2442 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X847 fc2 s4 VN.t2441 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X848 VN.t2440 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X849 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X850 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X851 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X852 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X853 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X854 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X855 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X856 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X857 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X858 VN.t2439 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X859 fc2 s4 VN.t2438 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X860 fc2 s4 VN.t2437 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X861 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X862 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X863 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X864 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X865 VN.t2436 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X866 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X867 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X868 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X869 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X870 VN.t2435 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X871 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X872 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X873 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X874 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X875 fc2 s4 VN.t2434 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X876 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X877 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X878 fc2 s4 VN.t2433 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X879 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X880 VN.t2432 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X881 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X882 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X883 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X884 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X885 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X886 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X887 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X888 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X889 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X890 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X891 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X892 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X893 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X894 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X895 VN.t2431 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X896 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X897 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X898 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X899 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X900 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X901 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X902 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X904 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X905 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X906 VN.t2430 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X907 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X908 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X909 fc2 s4 VN.t2429 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X910 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X911 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X912 VN.t2428 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X913 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X914 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X915 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X916 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X917 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X918 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X919 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X920 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X921 fc2 s4 VN.t2427 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X922 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X923 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X924 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X925 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X926 VN.t2426 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X927 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X928 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X929 VN.t2425 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X930 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X931 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X932 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X933 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X934 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X935 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X936 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X937 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X938 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X939 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X940 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X941 fc2 s4 VN.t2424 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X942 VN.t2423 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X943 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X944 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X945 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X946 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X947 fc2 s4 VN.t2422 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X948 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X949 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X950 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X951 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X952 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X953 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X954 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X955 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X956 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X957 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X958 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X959 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X960 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X961 VN.t2421 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X962 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X963 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X964 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X965 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X966 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X967 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X968 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X969 fc2 s4 VN.t2420 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X970 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X971 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X972 fc2 s4 VN.t2419 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X973 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X974 VN.t2418 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X975 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X976 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X977 VN.t2417 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X978 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X979 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X980 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X981 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X982 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X983 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X984 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X985 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X986 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X987 VN.t2416 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X988 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X989 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X990 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X991 VN.t2415 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X992 fc2 s4 VN.t2414 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X993 VN.t2413 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X994 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X995 fc2 s4 VN.t2412 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X996 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X998 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X999 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1000 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1001 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1002 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1003 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1004 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1005 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1007 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1009 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1010 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1011 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1012 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1013 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1014 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1015 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1016 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1017 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1018 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1019 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1020 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1021 fc2 s4 VN.t2411 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1022 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1023 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1024 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1025 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1026 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1027 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1028 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1029 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1030 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1031 VN.t2410 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1032 VN.t2409 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1033 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1034 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1035 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1036 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1037 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1038 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1039 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1040 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1041 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1042 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1043 fc2 s4 VN.t2408 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1044 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1045 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1046 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1047 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1048 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1049 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1050 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1051 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1052 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1053 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1054 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1055 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1056 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1057 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1058 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1059 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1060 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1061 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1062 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1063 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1064 VN.t2407 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1065 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1066 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1067 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1068 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1069 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1070 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1071 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1072 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1073 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1074 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1075 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1076 fc2 s4 VN.t2406 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1077 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1078 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1079 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1080 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1081 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1082 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1083 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1084 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1085 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1086 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1088 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1089 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1090 fc2 s4 VN.t2405 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1091 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1092 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1093 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1094 VN.t2404 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1095 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1096 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1097 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1098 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1099 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1100 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1101 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1102 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1103 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1104 fc2 s4 VN.t2403 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1105 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1106 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1107 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1108 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1109 VN.t2402 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1110 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1111 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1112 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1113 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1114 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1115 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1116 VN.t2401 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1117 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1118 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1119 fc2 s4 VN.t2400 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1120 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1121 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1122 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1123 fc2 s4 VN.t2399 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1124 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1125 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1126 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1127 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1128 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1129 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1130 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1131 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1132 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1133 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1134 VN.t2398 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1135 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1136 VN.t2397 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1137 fc2 s4 VN.t2396 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1138 fc2 s4 VN.t2395 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1139 VN.t2394 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1140 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1141 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1142 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1143 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1144 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1145 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1146 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1147 fc2 s4 VN.t2393 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1148 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1149 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1150 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1151 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1152 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1153 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1154 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1156 fc2 s4 VN.t2392 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1157 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1158 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1159 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1160 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1161 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1162 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1163 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1164 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1165 fc2 s4 VN.t2391 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1166 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1167 VN.t2390 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1168 fc2 s4 VN.t2389 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1169 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1170 VN.t2388 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1171 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1172 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1173 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1174 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1175 VN.t2387 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1176 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1177 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1178 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1180 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1181 VN.t2386 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1182 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1183 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1184 VN.t2385 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1185 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1186 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1187 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1188 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1189 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1190 fc2 s4 VN.t2384 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1191 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1192 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1193 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1194 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1195 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1196 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1198 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1199 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1200 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1201 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1202 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1203 VN.t2383 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1204 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1205 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1206 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1207 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1208 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1209 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1210 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1211 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1212 VN.t2382 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1213 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1214 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1215 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1216 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1217 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1218 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1219 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1220 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1221 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1222 VN.t2381 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1223 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1224 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1225 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1226 VN.t2380 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1227 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1228 fc2 s4 VN.t2379 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1229 fc2 s4 VN.t2378 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1230 VN.t2377 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1231 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1232 fc2 s4 VN.t2376 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1233 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1234 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1235 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1236 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1237 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1238 VN.t2375 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1239 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1240 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1241 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1242 fc2 s4 VN.t2374 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1243 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1244 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1245 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1246 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1247 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1248 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1249 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1250 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1251 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1252 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1253 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1254 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1255 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1256 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1257 VN.t2373 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1258 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1259 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1260 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1261 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1262 VN.t2372 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1263 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1264 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1265 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1266 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X1267 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1268 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1269 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1270 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1271 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1272 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1273 VN.t2371 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1274 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1275 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1276 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1278 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1279 VN.t2370 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1280 VN.t2369 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1281 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1282 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1283 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1284 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1285 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1286 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1287 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1288 fc2 s4 VN.t2368 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1290 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1291 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1292 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1293 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1294 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1295 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1296 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1297 fc2 s4 VN.t2367 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1298 VN.t2366 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1299 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1300 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1301 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1302 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1303 fc2 s4 VN.t2365 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1304 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1305 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1306 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1307 VN.t2364 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1308 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1309 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1310 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1311 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1312 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1313 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1314 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1315 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1316 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1317 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1318 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1319 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1320 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1321 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1322 VN.t2363 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1323 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1324 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1325 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1326 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1327 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1328 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1329 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1330 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1331 fc2 s4 VN.t2362 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1332 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1333 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1334 VN.t2361 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1335 VN.t2360 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1336 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1337 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1339 fc2 s4 VN.t2359 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1340 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1341 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1342 fc2 s4 VN.t2358 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1343 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1344 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1345 VN.t2357 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1346 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1347 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1348 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1349 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1350 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1351 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1352 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1353 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1354 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1355 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1356 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1357 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1358 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1359 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1360 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1361 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1362 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1363 VN.t2356 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1364 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1365 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1366 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1367 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1368 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1369 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1370 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1371 fc2 s4 VN.t2355 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1372 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1373 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1374 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1375 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1377 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1378 fc2 s4 VN.t2354 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1379 VN.t2353 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1380 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1381 fc2 s4 VN.t2352 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1382 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1383 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1384 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1385 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1386 VN.t2351 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1387 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1388 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1389 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1390 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1391 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1392 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1393 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1394 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1395 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1396 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1397 fc2 s4 VN.t2350 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1398 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1399 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1400 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1401 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1402 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1403 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1404 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1405 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1406 fc2 s4 VN.t2349 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1407 VN.t2348 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1408 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1409 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1410 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1411 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1412 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1413 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1414 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1415 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1416 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1417 VN.t2347 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1418 VN.t2346 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1419 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1420 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1421 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1422 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1423 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1424 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1425 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1426 fc2 s4 VN.t2345 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1427 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1428 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1429 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1430 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1431 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1432 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1433 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1434 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1435 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1436 VN.t2344 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1437 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1438 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1439 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1440 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1441 fc2 s4 VN.t2343 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1442 fc2 s4 VN.t2342 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1443 fc2 s4 VN.t2341 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1444 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1445 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1446 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1447 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1448 VN.t2340 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1449 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1450 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1451 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1452 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1453 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1454 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1455 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1456 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X1457 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1458 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1459 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1460 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1461 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1462 VN.t2339 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1463 fc2 s4 VN.t2338 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1464 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1465 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1466 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1467 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1468 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1469 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1470 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1471 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1472 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1473 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1474 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1475 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1476 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1477 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1478 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1479 fc2 s4 VN.t2337 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1480 fc2 s4 VN.t2336 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1481 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1482 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1483 VN.t2335 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1484 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1485 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1486 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1487 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1488 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1489 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1490 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1491 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1492 VN.t2334 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1493 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1494 fc2 s4 VN.t2333 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1495 VN.t2332 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1496 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1497 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1498 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1499 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1500 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1501 fc2 s4 VN.t2331 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1502 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1503 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1504 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1505 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1506 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1507 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1508 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1509 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1510 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1511 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1512 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1513 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1514 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1515 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1516 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1517 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1518 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1519 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1520 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1521 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1522 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1523 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1524 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1525 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1526 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1527 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1528 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1529 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1530 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1531 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1532 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1533 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1534 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1535 VN.t2330 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1536 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1537 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1538 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1539 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1540 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1541 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1542 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1543 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1544 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1545 fc2 s4 VN.t2329 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1546 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1547 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1548 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1549 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1550 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1551 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1552 VN.t2328 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1553 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1554 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1555 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1556 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1557 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1558 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1559 fc2 s4 VN.t2327 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1560 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1561 VN.t2326 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1562 fc2 s4 VN.t2325 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1563 VN.t2324 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1564 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1565 fc2 s4 VN.t2323 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1566 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1567 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1568 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1569 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1570 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1571 VN.t2322 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1572 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1573 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1574 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1575 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1576 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1577 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1578 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1579 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1580 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1582 VN.t2321 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1583 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1584 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1585 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1586 fc2 s4 VN.t2320 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1587 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1588 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1590 VN.t2319 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1591 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1592 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1593 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1594 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1595 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1596 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1597 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1598 VN.t2318 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1599 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1600 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1601 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1602 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1603 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1604 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1605 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1606 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1607 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1608 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1609 VN.t2317 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1610 VN.t2316 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1611 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1612 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1613 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1614 fc2 s4 VN.t2315 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1615 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1616 VN.t2314 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1617 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1618 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1619 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1620 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1622 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1623 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1624 fc2 s4 VN.t2313 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1625 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1626 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1627 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1628 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1629 VN.t2312 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1630 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1631 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1632 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1633 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1634 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1635 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1636 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1637 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1638 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1639 VN.t2311 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1640 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1641 VN.t2310 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1642 fc2 s4 VN.t2309 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1643 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1644 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1645 VN.t2308 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1646 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1647 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1648 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1649 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1650 VN.t2307 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1651 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1652 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1653 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1654 fc2 s4 VN.t2306 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1655 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1656 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1657 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1658 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1659 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1660 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1661 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1663 VN.t2305 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1664 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1665 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1666 fc2 s4 VN.t2304 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1667 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1668 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1669 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1670 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1671 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1672 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1673 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1674 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1675 fc2 s4 VN.t2303 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1676 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1677 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1678 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1679 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1680 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1681 VN.t2302 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1682 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1683 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1684 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1685 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1686 fc2 s4 VN.t2301 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1687 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1688 VN.t2300 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1689 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1690 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1691 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1692 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1693 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1694 VN.t2299 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1695 fc2 s4 VN.t2298 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1696 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1697 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1698 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1699 fc2 s4 VN.t2297 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1700 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1701 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1702 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1703 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1704 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1705 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1706 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1707 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1708 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1709 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1710 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1711 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1712 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1713 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1714 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1715 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1716 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1717 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1718 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1719 fc2 s4 VN.t2296 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1720 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1721 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1722 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1723 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1724 VN.t2295 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1725 VN.t2294 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1726 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1727 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1728 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1729 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1730 fc2 s4 VN.t2293 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1731 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1732 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1733 fc2 s4 VN.t2292 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1734 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1735 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1736 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1737 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1738 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1739 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1740 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1741 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1742 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1743 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1744 VN.t2291 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1745 VN.t2290 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1746 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1747 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1748 VN.t2289 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1749 fc2 s4 VN.t2288 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1750 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1751 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1752 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1753 fc2 s4 VN.t2287 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1754 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1755 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1756 VN.t2286 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1757 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1758 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1759 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1760 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1761 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1762 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1763 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1764 VN.t2285 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1765 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1766 fc2 s4 VN.t2284 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1767 VN.t2283 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1768 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1769 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1770 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1771 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1772 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1773 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1774 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1775 fc2 s4 VN.t2282 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1776 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1777 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1778 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1779 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1780 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1781 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1782 VN.t2281 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1783 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1784 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1785 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1786 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1787 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1788 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1789 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1790 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1791 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1792 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1793 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1794 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1795 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1796 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1797 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1798 fc2 s4 VN.t2280 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1799 VN.t2279 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1800 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1801 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1802 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1803 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1804 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1805 fc2 s4 VN.t2278 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1806 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1807 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1808 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1809 fc2 s4 VN.t2277 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1810 VN.t2276 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1811 fc2 s4 VN.t2275 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1812 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1813 VN.t2274 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1814 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1815 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1816 fc2 s4 VN.t2273 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1817 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1818 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1819 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1820 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1821 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1822 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1823 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1824 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1825 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1826 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1827 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1828 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1829 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1830 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1831 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1832 VN.t2272 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1833 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1834 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1835 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1836 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1837 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1838 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1839 fc2 s4 VN.t2271 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1840 VN.t2270 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1841 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1842 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1844 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1845 fc2 s4 VN.t2269 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1846 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1847 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1848 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1849 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1850 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1851 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1852 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1853 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1854 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1855 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1856 VN.t2268 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1857 fc2 s4 VN.t2267 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1858 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1859 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1860 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1861 VN.t2266 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1862 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1863 VN.t2265 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1864 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1865 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1866 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1867 VN.t2264 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1868 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1869 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1870 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1871 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1872 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1873 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1874 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1875 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1876 fc2 s4 VN.t2263 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1877 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1878 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1879 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1880 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1881 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1882 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1883 fc2 s4 VN.t2262 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1884 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1885 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1886 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1887 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1888 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1889 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1890 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1891 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1892 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1894 VN.t2261 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1895 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1896 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1897 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1898 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1899 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1900 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1901 fc2 s4 VN.t2260 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1902 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1903 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1904 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1905 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1906 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1907 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1908 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1909 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1910 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1911 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1912 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1913 fc2 s4 VN.t2259 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1914 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1915 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1916 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1917 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1918 fc2 s4 VN.t2258 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1919 VN.t2257 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1920 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1921 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1922 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1923 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1924 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1925 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1926 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1927 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1928 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1929 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1930 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1931 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1932 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1933 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1934 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1935 fc2 s4 VN.t2256 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1936 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1937 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1938 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1939 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1940 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1941 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1942 fc2 s4 VN.t2255 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1943 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1944 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1945 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1946 VN.t2254 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1947 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1948 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1949 VN.t2253 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1950 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1951 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1952 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1953 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1954 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1955 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1956 fc2 s4 VN.t2252 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1957 fc2 s4 VN.t2251 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1958 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1959 fc2 s4 VN.t2250 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1960 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1961 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1962 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1963 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1964 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1965 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1966 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1967 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1968 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1969 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1970 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1971 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1972 fc2 s4 VN.t2249 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1973 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1974 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1975 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1976 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1977 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1978 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1980 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1981 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1982 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1983 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1984 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1985 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1986 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1987 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1988 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1989 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1990 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1991 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1992 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1993 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1994 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1995 fc2 s4 VN.t2248 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1996 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1997 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1998 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1999 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2000 fc2 s4 VN.t2247 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2001 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2002 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2003 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2004 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2005 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2006 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2007 VN.t2246 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2009 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2010 VN.t2245 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2011 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2012 VN.t2244 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2013 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2014 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2015 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2017 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2018 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2019 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2020 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2021 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2022 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2023 fc2 s4 VN.t2243 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2024 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2025 fc2 s4 VN.t2242 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2026 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2027 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2028 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2029 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2030 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2031 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2032 fc2 s4 VN.t2241 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2033 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2034 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2035 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2036 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2037 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2038 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2039 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2040 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2041 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2042 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2043 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2044 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2045 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2047 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2048 fc2 s4 VN.t2240 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2049 VN.t2239 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2050 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2051 fc2 s4 VN.t2238 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2052 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2053 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2054 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2055 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2056 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2057 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2058 VN.t2237 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2059 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2060 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2061 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2062 fc2 s4 VN.t2236 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2063 VN.t2235 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2064 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2065 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2066 fc2 s4 VN.t2234 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2067 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2068 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2069 VN.t2233 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2070 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2071 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2072 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2073 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2074 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2075 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2076 VN.t2232 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2077 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2078 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2079 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2080 fc2 s4 VN.t2231 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2081 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2082 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2083 fc2 s4 VN.t2230 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2084 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2085 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2086 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2088 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2089 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2090 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2091 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2092 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2093 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2094 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2095 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2096 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2097 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2098 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2099 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2100 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2101 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2102 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2103 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2104 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2105 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2106 VN.t2229 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2107 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2108 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2109 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2111 VN.t2228 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2112 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2113 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2114 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2116 fc2 s4 VN.t2227 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2117 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2119 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2120 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2121 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2122 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2123 fc2 s4 VN.t2226 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2124 fc2 s4 VN.t2225 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2125 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2126 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2127 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2128 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2129 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2130 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2131 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2132 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2133 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2134 VN.t2224 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2135 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2136 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2137 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2138 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2139 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2140 VN.t2223 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2141 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2142 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2143 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2144 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2145 fc2 s4 VN.t2222 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2146 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2147 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2148 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2149 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2150 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2151 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2152 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2153 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2154 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2155 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2156 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2157 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2158 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2159 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2160 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2161 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2162 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2163 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2164 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2165 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2166 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2167 fc2 s4 VN.t2221 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2168 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2169 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2170 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2171 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2172 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2173 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2174 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2175 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2176 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2177 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2178 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2179 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2180 fc2 s4 VN.t2220 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2181 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2182 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2183 VN.t2219 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2184 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2185 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2186 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2187 fc2 s4 VN.t2218 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2188 fc2 s4 VN.t2217 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2189 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2190 VN.t2216 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2191 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2192 fc2 s4 VN.t2215 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2193 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2194 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2195 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2196 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2197 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2198 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2199 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2200 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2201 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2202 fc2 s4 VN.t2214 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2203 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2205 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2206 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2207 fc2 s4 VN.t2213 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2208 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2209 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2210 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2211 VN.t2212 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2212 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2213 VN.t2211 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2214 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2215 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2216 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2217 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2218 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2219 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2220 VN.t2210 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2221 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2222 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2223 fc2 s4 VN.t2209 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2224 VN.t2208 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2225 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2226 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2227 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2228 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2229 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2230 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2231 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2232 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2234 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2235 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2236 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2237 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2238 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2239 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2240 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2241 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2242 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2243 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2244 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2245 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2246 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2247 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2248 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2249 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2250 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2251 fc2 s4 VN.t2207 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2252 VN.t2206 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2253 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2254 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2255 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2256 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2257 fc2 s4 VN.t2205 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2258 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2259 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2260 fc2 s4 VN.t2204 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2261 fc2 s4 VN.t2203 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2262 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2263 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2264 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2265 fc2 s4 VN.t2202 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2266 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2267 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2268 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2269 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2270 VN.t2201 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2271 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2272 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2273 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2274 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2275 VN.t2200 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2276 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2277 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2278 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2279 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2280 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2281 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2282 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2283 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2284 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2285 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2286 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2287 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2288 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2289 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2290 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2291 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2292 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2293 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2294 fc2 s4 VN.t2199 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2295 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2296 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2297 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2298 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2299 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2300 VN.t2198 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2301 fc2 s4 VN.t2197 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2302 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2303 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2304 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2305 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2306 VN.t2196 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2307 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2308 VN.t2195 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2309 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2310 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2311 VN.t2194 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2312 fc2 s4 VN.t2193 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2313 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2314 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2315 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2316 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2317 fc2 s4 VN.t2192 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2318 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2319 VN.t2191 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2320 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2321 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2322 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2323 fc2 s4 VN.t2190 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2324 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2325 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2326 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2327 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2328 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2329 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2330 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2331 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2332 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2333 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2334 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2335 VN.t2189 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2336 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2337 fc2 s4 VN.t2188 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2338 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2339 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2340 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2341 fc2 s4 VN.t2187 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2342 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2343 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2344 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2345 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2346 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X2347 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2348 fc2 s4 VN.t2186 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2349 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2350 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2351 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2352 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2353 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2354 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X2355 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2356 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2357 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2358 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2359 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2360 fc2 s4 VN.t2185 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2361 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2362 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2363 VN.t2184 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2364 fc2 s4 VN.t2183 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2365 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2366 fc2 s4 VN.t2182 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2367 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2368 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2369 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2370 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2371 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2372 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2373 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2374 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2375 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2377 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2378 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2379 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2380 fc2 s4 VN.t2181 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2381 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2382 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2383 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2384 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2385 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2386 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2387 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2388 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2389 VN.t2180 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2390 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2391 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2392 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2393 VN.t2179 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2394 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2395 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2396 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2397 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2398 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2399 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2400 VN.t2178 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2401 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2402 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2403 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2404 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2405 fc2 s4 VN.t2177 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2406 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2407 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2408 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2409 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2410 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2411 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2412 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2413 fc2 s4 VN.t2176 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2414 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2415 fc2 s4 VN.t2175 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2416 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2417 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2418 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2419 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2420 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2421 VN.t2174 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2422 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2423 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2424 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2425 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2426 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2427 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2428 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2429 fc2 s4 VN.t2173 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2430 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2431 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2432 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2433 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2434 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2435 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2436 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2437 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2438 fc2 s4 VN.t2172 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2439 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2440 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2441 fc2 s4 VN.t2171 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2442 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2443 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2444 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2445 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2446 fc2 s4 VN.t2170 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2447 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2448 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2449 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2450 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2451 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2452 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2453 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2454 VN.t2169 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2455 fc2 s4 VN.t2168 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2456 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2457 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2458 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2459 VN.t2167 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2460 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2461 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2462 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2463 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2464 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2465 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2466 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2467 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2468 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2469 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2470 fc2 s4 VN.t2166 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2471 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2472 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2473 VN.t2165 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2474 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2475 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2476 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2477 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2478 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2479 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2480 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2481 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2482 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2483 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2484 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2485 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2486 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2487 VN.t2164 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2488 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2489 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2490 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2491 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2492 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2493 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2494 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2495 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2496 fc2 s4 VN.t2163 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2497 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2498 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2499 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2500 fc2 s4 VN.t2162 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2501 VN.t2161 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2502 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2503 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2504 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2505 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2506 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2507 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2508 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2509 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2510 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2511 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2512 fc2 s4 VN.t2160 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2513 VN.t2159 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2514 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2515 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2516 VN.t2158 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2517 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2518 VN.t2157 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2519 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2520 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2521 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2522 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2523 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2524 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2525 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2526 fc2 s4 VN.t2156 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2527 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2528 VN.t2155 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2529 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2530 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2531 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2532 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2533 VN.t2154 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2534 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2535 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2536 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2537 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2538 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2539 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2540 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2541 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2542 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2543 VN.t2153 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2544 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2545 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2546 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2547 VN.t2152 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2548 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2549 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2550 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2551 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2552 fc2 s4 VN.t2151 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2553 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2554 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2555 VN.t2150 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2556 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2557 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2558 VN.t2149 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2559 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2560 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2561 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2562 VN.t2148 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2563 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2564 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2565 VN.t2147 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2566 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2567 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2568 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2569 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2570 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2571 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2572 VN.t2146 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2573 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2574 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2575 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2576 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2577 fc2 s4 VN.t2145 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2578 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2579 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2580 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2581 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2582 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2583 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2584 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2585 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2586 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2587 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2588 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2589 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2590 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2591 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2592 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2593 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2594 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2595 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2596 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2597 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2598 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2599 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2600 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2601 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2602 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2603 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2604 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2605 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2606 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2607 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2608 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2609 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2610 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2611 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2612 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2613 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2614 VN.t2144 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2615 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2616 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2618 VN.t2143 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2619 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2620 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2621 fc2 s4 VN.t2142 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2622 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2623 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2624 VN.t2141 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2625 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2626 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2627 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2628 VN.t2140 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2629 fc2 s4 VN.t2139 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2630 VN.t2138 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2631 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2632 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2633 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2634 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2635 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2636 fc2 s4 VN.t2137 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2637 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2638 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2639 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2640 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2641 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2643 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2644 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2645 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2646 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2647 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2648 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2649 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2650 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2651 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2652 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2653 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2654 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2655 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2656 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2657 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2658 fc2 s4 VN.t2136 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2659 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2660 VN.t2135 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2661 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2662 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2663 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2664 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2665 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2666 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2667 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2668 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2669 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2670 VN.t2134 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2671 fc2 s4 VN.t2133 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2672 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2673 fc2 s4 VN.t2132 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2674 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2675 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2676 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2677 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2678 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2679 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2680 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2681 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2682 fc2 s4 VN.t2131 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2683 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2684 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2685 VN.t2130 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2686 VN.t2129 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2687 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2688 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2689 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2690 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2691 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2692 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2693 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2694 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2695 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2696 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2697 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2698 fc2 s4 VN.t2128 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2699 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2700 fc2 s4 VN.t2127 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2701 VN.t2126 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2702 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2703 fc2 s4 VN.t2125 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2704 VN.t2124 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2705 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2706 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2707 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2708 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2709 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2710 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2711 fc2 s4 VN.t2123 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2712 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2713 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2714 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2715 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2716 fc2 s4 VN.t2122 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2717 VN.t2121 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2718 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2719 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2720 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2721 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2722 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2723 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2724 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2725 VN.t2120 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2726 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2727 fc2 s4 VN.t2119 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2728 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2729 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2730 VN.t2118 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2731 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2732 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2733 fc2 s4 VN.t2117 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2734 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2735 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2736 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2737 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2738 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2739 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2740 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2741 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2742 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2743 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2744 fc2 s4 VN.t2116 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2745 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2746 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2747 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2748 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X2749 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2750 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2751 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2752 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2753 fc2 s4 VN.t2115 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2754 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2755 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2756 fc2 s4 VN.t2114 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2757 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2758 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2759 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2760 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2761 VN.t2113 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2762 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2763 VN.t2112 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2764 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2765 VN.t2111 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2766 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2767 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2768 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2769 fc2 s4 VN.t2110 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2770 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2771 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2772 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2773 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2774 VN.t2109 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2775 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2776 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2777 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2778 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2779 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2780 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2781 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2782 VN.t2108 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2783 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2784 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2785 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2786 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2787 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2788 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2789 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2790 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2791 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2792 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2793 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2794 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2795 VN.t2107 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2796 VN.t2106 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2797 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2798 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2799 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2800 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2801 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2802 fc2 s4 VN.t2105 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2803 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2804 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2805 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2806 VN.t2104 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2807 VN.t2103 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2808 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2809 fc2 s4 VN.t2102 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2810 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2811 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2812 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2813 VN.t2101 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2814 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2815 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2816 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2817 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2818 VN.t2100 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2819 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2820 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2821 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2822 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2823 fc2 s4 VN.t2099 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2824 fc2 s4 VN.t2098 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2825 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2826 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2827 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2828 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2829 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2830 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2831 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2832 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2833 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2834 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2835 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2836 VN.t2097 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2837 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2838 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2839 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2840 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2841 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2842 VN.t2096 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2844 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2845 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2846 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2847 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2848 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2849 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2850 VN.t2095 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2851 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2852 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2853 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2854 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2855 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2856 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2857 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2858 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2859 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2860 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2861 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2862 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2863 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2864 fc2 s4 VN.t2094 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2865 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2866 VN.t2093 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2867 VN.t2092 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2868 VN.t2091 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2869 VN.t2090 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2870 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2871 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2872 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2873 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2874 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2875 fc2 s4 VN.t2089 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2876 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2877 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2878 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2879 VN.t2088 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2880 fc2 s4 VN.t2087 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2881 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2882 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2883 fc2 s4 VN.t2086 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2884 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2886 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2887 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2888 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2889 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2890 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2891 fc2 s4 VN.t2085 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2892 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2893 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2894 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2895 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2896 fc2 s4 VN.t2084 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2897 VN.t2083 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2898 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2899 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2900 VN.t2082 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2901 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2902 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2903 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2904 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2905 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2906 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2907 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2908 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2909 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2910 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2911 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2912 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2913 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2914 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2915 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2916 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2917 fc2 s4 VN.t2081 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2918 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2919 VN.t2080 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2920 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2921 VN.t2079 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2922 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2923 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2924 fc2 s4 VN.t2078 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2925 fc2 s4 VN.t2077 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2926 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2927 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2928 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2929 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2930 VN.t2076 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2931 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2932 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2933 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2934 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2935 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2936 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2937 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2938 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2939 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2940 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2941 fc2 s4 VN.t2075 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2942 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2943 VN.t2074 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2944 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2945 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2946 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2947 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2948 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2949 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2950 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2951 VN.t2073 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2952 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2953 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2954 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2955 fc2 s4 VN.t2072 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2956 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2957 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2958 fc2 s4 VN.t2071 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2959 VN.t2070 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2960 VN.t2069 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2961 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2962 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2963 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2964 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2965 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2966 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2967 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2968 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2969 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2970 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2971 fc2 s4 VN.t2068 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2972 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2973 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2974 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2975 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2976 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2977 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2978 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2980 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2981 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2982 fc2 s4 VN.t2067 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2983 VN.t2066 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2984 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2985 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2986 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2987 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2988 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2989 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2990 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2991 VN.t2065 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2992 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2993 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2994 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2995 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2996 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2998 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2999 fc2 s4 VN.t2064 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3000 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3001 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3002 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3003 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3004 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3005 VN.t2063 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3006 VN.t2062 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3007 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3008 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3009 VN.t2061 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3010 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3011 fc2 s4 VN.t2060 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3012 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3013 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3014 fc2 s4 VN.t2059 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3015 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3017 fc2 s4 VN.t2058 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3019 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3020 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3021 VN.t2057 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3022 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3023 VN.t2056 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3024 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3025 fc2 s4 VN.t2055 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3026 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3027 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3028 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3029 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3030 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3031 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3032 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3033 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3034 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3035 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3036 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3037 VN.t2054 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3038 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3039 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3040 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3041 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3042 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3043 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3044 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3045 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3046 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3047 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3048 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3049 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3050 fc2 s4 VN.t2053 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3051 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3052 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3053 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3054 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3055 fc2 s4 VN.t2052 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3056 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3057 VN.t2051 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3058 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3059 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3060 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3061 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3062 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3063 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3064 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3065 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3066 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3067 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3068 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3069 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3070 VN.t2050 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3071 fc2 s4 VN.t2049 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3072 VN.t2048 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3073 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3074 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3075 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3076 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3077 VN.t2047 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3078 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3079 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3080 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3081 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3082 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3083 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3084 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3085 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3086 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3087 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3088 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3089 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3090 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3091 VN.t2046 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3092 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3093 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3094 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3095 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3096 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3097 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3098 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3099 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3101 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3102 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3103 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3104 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3105 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3106 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3107 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3108 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3109 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3110 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3111 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3112 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3113 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3114 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3116 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3117 VN.t2045 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3118 VN.t2044 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3119 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3120 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3121 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3122 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3123 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3124 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3125 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3126 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3127 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3128 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3129 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3130 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3131 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3132 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3133 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3134 VN.t2043 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3135 fc2 s4 VN.t2042 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3136 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3137 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3138 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3139 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3140 VN.t2041 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3141 VN.t2040 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3142 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3143 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3144 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3145 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3146 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3147 fc2 s4 VN.t2039 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3148 VN.t2038 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3149 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3150 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3151 fc2 s4 VN.t2037 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3152 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3153 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3154 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3155 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3156 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3157 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3158 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3159 VN.t2036 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3160 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3161 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3162 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3163 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3164 VN.t2035 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3165 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3166 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3167 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3168 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3169 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3170 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3171 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3172 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3173 fc2 s4 VN.t2034 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3174 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3175 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3176 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3177 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3178 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3180 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3181 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3182 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3183 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3184 fc2 s4 VN.t2033 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3185 VN.t2032 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3186 VN.t2031 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3187 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3188 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3189 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3190 VN.t2030 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3191 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3192 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3193 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3194 VN.t2029 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3195 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3196 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3198 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3199 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3200 VN.t2028 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3201 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3202 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3203 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3204 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3205 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3206 fc2 s4 VN.t2027 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3207 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3208 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3209 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3210 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3211 VN.t2026 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3212 VN.t2025 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3213 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3214 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3215 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3216 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3217 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3218 VN.t2024 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3219 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3220 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3221 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3222 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3223 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3224 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3225 VN.t2023 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3226 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3227 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3228 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3229 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3230 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3231 VN.t2022 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3232 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3233 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3234 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3235 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3236 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3237 fc2 s4 VN.t2021 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3238 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3239 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3240 VN.t2020 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3241 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3242 fc2 s4 VN.t2019 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3243 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3244 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3246 VN.t2018 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3247 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3248 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3249 fc2 s4 VN.t2017 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3250 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3251 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3252 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3253 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3254 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3255 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3256 VN.t2016 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3257 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3258 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3259 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3260 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3261 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3262 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3263 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3264 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3265 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3266 VN.t2015 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3267 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3268 fc2 s4 VN.t2014 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3269 VN.t2013 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3270 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3271 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3272 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3273 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3274 fc2 s4 VN.t2012 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3275 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3276 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3277 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3278 VN.t2011 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3279 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3280 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3281 VN.t2010 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3282 VN.t2009 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3283 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3284 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3285 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3286 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3287 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3288 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3290 VN.t2008 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3291 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3292 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3293 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3294 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3295 fc2 s4 VN.t2007 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3296 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3297 fc2 s4 VN.t2006 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3298 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3299 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3300 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3301 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3302 fc2 s4 VN.t2005 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3303 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3304 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3305 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3306 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3307 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3308 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3309 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3310 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3311 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3312 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3313 fc2 s4 VN.t2004 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3314 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3315 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3316 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3317 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3318 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3319 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3320 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3321 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3322 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3323 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3324 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3325 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3326 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3327 fc2 s4 VN.t2003 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3328 fc2 s4 VN.t2002 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3329 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3330 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3331 fc2 s4 VN.t2001 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3332 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3333 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3334 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3335 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3336 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3337 fc2 s4 VN.t2000 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3338 VN.t1999 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3339 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3340 VN.t1998 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3341 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3342 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3343 fc2 s4 VN.t1997 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3344 VN.t1996 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3345 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3346 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3347 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3348 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3349 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3350 fc2 s4 VN.t1995 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3351 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3352 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3353 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3354 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3355 fc2 s4 VN.t1994 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3356 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3357 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3358 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3359 VN.t1993 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3360 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3361 VN.t1992 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3362 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3363 VN.t1991 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3364 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3365 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3366 fc2 s4 VN.t1990 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3367 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3368 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3369 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3370 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3372 VN.t1989 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3373 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3374 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3375 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3376 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3377 VN.t1988 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3378 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3379 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3380 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3381 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3382 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3383 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3384 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3385 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3386 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3387 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3388 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3389 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3390 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3391 VN.t1987 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3392 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3393 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3394 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3395 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3396 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3397 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3398 fc2 s4 VN.t1986 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3399 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3400 fc2 s4 VN.t1985 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3401 VN.t1984 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3402 fc2 s4 VN.t1983 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3403 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3404 VN.t1982 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3405 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3406 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3407 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3408 fc2 s4 VN.t1981 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3409 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3410 fc2 s4 VN.t1980 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3411 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3412 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3413 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3414 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3415 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3416 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3417 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3418 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3419 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3420 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3421 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3422 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3423 VN.t1979 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3424 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3425 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3426 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3427 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3428 fc2 s4 VN.t1978 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3429 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3430 VN.t1977 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3431 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3432 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3433 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3434 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3435 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3436 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3437 fc2 s4 VN.t1976 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3438 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3439 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3440 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3441 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3442 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3443 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3444 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3445 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3446 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3447 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3448 fc2 s4 VN.t1975 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3449 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3450 fc2 s4 VN.t1974 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3451 VN.t1973 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3452 VN.t1972 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3453 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3454 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3455 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3456 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3457 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3458 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3459 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3460 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3461 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3462 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3463 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3464 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3465 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3466 fc2 s4 VN.t1971 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3467 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3468 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3469 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3470 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3471 fc2 s4 VN.t1970 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3472 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3473 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3474 fc2 s4 VN.t1969 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3475 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3476 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3477 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3478 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3479 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3480 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3481 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3482 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3483 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3484 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3485 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3486 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3487 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3488 fc2 s4 VN.t1968 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3489 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3490 fc2 s4 VN.t1967 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3491 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3492 fc2 s4 VN.t1966 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3493 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3494 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3495 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3496 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3497 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3498 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3499 fc2 s4 VN.t1965 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3500 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3501 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3502 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3503 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3504 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3505 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3506 VN.t1964 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3507 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3508 fc2 s4 VN.t1963 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3509 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3510 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3511 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3512 VN.t1962 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3513 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3514 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3515 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3516 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3517 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3518 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3519 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3520 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3521 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3522 fc2 s4 VN.t1961 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3523 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3524 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3525 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3526 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3527 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3528 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3529 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3530 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3531 VN.t1960 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3532 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3533 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3534 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3535 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3536 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3537 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3538 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3539 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3540 VN.t1959 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3541 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3542 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3543 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3544 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3545 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3546 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3547 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3548 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3549 fc2 s4 VN.t1958 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3550 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3551 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3552 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3553 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3554 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3555 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3556 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3557 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3558 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3559 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3560 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3561 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3562 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3563 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3564 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3565 fc2 s4 VN.t1957 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3566 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3567 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3568 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3569 VN.t1956 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3570 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3571 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3572 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3573 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3574 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3575 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3576 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3577 fc2 s4 VN.t1955 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3578 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3579 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3580 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3582 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3583 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3584 fc2 s4 VN.t1954 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3585 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3586 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3587 fc2 s4 VN.t1953 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3588 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3589 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3590 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3591 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3592 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3593 fc2 s4 VN.t1952 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3594 fc2 s4 VN.t1951 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3595 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3596 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3597 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3598 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3599 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3600 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3601 VN.t1950 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3602 VN.t1949 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3603 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3604 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3605 VN.t1948 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3606 fc2 s4 VN.t1947 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3607 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3608 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3609 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3610 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3611 fc2 s4 VN.t1946 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3612 fc2 s4 VN.t1945 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3613 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3614 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3615 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3616 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3618 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3619 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3620 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3621 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3622 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3623 fc2 s4 VN.t1944 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3624 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3625 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3626 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3627 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3628 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3629 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3630 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3631 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3632 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3633 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3634 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3635 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3636 fc2 s4 VN.t1943 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3637 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3638 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3639 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3640 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3641 fc2 s4 VN.t1942 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3643 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3644 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3645 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3646 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3647 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3648 VN.t1941 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3649 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3650 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3651 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3652 fc2 s4 VN.t1940 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3653 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3654 VN.t1939 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3655 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3656 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3657 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3658 VN.t1938 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3659 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3660 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3661 fc2 s4 VN.t1937 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3663 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3664 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3665 fc2 s4 VN.t1936 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3666 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3667 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3668 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3669 VN.t1935 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3670 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3671 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3672 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3673 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3674 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3675 fc2 s4 VN.t1934 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3676 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3677 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3678 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3679 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3680 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3681 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3682 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3683 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3684 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3685 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3686 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3687 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3688 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3689 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3690 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3691 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3692 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3693 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3694 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3695 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3696 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3697 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3698 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3699 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3700 VN.t1933 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3701 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3702 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3703 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3704 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3705 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3706 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3707 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3708 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3709 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3710 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3711 fc2 s4 VN.t1932 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3712 fc2 s4 VN.t1931 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3713 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3714 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3715 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3716 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3717 VN.t1930 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3718 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3719 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3720 VN.t1929 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3721 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3722 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3723 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3724 fc2 s4 VN.t1928 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3725 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3726 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3727 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3728 VN.t1927 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3729 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3730 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3731 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3732 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3733 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3734 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3735 fc2 s4 VN.t1926 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3736 fc2 s4 VN.t1925 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3737 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3739 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3740 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3741 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3742 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3743 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3744 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3745 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3746 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3747 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X3748 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3749 VN.t1924 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3750 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3751 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3752 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3753 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3754 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3755 fc2 s4 VN.t1923 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3756 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3757 VN.t1922 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3758 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3759 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3760 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3761 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3762 VN.t1921 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3763 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3764 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3765 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3766 fc2 s4 VN.t1920 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3767 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3768 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3769 fc2 s4 VN.t1919 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3770 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3771 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3772 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3773 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3774 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3775 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3776 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3777 VN.t1918 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3778 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3779 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3780 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3781 VN.t1917 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3782 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3783 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3784 VN.t1916 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3785 fc2 s4 VN.t1915 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3786 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3787 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3788 fc2 s4 VN.t1914 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3789 fc2 s4 VN.t1913 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3790 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3791 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3792 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3793 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3794 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3795 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3796 fc2 s4 VN.t1912 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3797 VN.t1911 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3798 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3799 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3800 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3801 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3802 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3803 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3804 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3805 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3806 fc2 s4 VN.t1910 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3807 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3808 fc2 s4 VN.t1909 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3809 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3810 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3811 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3812 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3813 fc2 s4 VN.t1908 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3814 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3815 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3816 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3817 fc2 s4 VN.t1907 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3818 VN.t1906 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3819 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3820 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3821 VN.t1905 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3822 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3823 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3824 VN.t1904 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3825 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3826 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3827 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3828 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3829 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3830 fc2 s4 VN.t1903 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3831 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3832 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3833 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3834 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3835 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3836 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3837 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3838 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3839 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3840 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3841 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3842 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3843 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3844 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3845 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3846 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3847 VN.t1902 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3848 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3849 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3850 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3851 fc2 s4 VN.t1901 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3852 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3853 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3854 VN.t1900 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3855 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3856 VN.t1899 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3857 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3858 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3859 fc2 s4 VN.t1898 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3860 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3861 fc2 s4 VN.t1897 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3862 fc2 s4 VN.t1896 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3863 VN.t1895 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3864 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3865 fc2 s4 VN.t1894 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3866 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3867 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3868 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3869 VN.t1893 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3870 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3871 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3872 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3873 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3874 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3875 VN.t1892 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3876 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3877 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3878 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3879 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3880 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3881 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3882 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3883 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3884 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3885 VN.t1891 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3886 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3887 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3888 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3889 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3890 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3891 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3892 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3894 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3895 fc2 s4 VN.t1890 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3896 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3897 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3898 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3899 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3900 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3901 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3902 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3904 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3905 fc2 s4 VN.t1889 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3906 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3907 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3908 VN.t1888 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3909 fc2 s4 VN.t1887 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3910 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3911 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3912 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3913 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3914 VN.t1886 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3915 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3916 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3917 fc2 s4 VN.t1885 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3918 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3919 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3920 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3921 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3922 fc2 s4 VN.t1884 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3923 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3924 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3925 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3926 fc2 s4 VN.t1883 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3927 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3929 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3930 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3931 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3932 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3933 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3934 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3935 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3936 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3937 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3938 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3939 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3940 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3941 fc2 s4 VN.t1882 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3942 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3943 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3944 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3945 fc2 s4 VN.t1881 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3946 fc2 s4 VN.t1880 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3947 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3948 fc2 s4 VN.t1879 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3949 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3950 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3951 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3952 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3953 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3954 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3955 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3956 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3957 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3958 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3959 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3960 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3961 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3962 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3963 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3964 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3965 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3966 fc2 s4 VN.t1878 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3967 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3968 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3969 VN.t1877 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3970 fc2 s4 VN.t1876 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3971 fc2 s4 VN.t1875 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3972 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3973 fc2 s4 VN.t1874 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3974 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3975 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3976 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3977 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3978 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3979 fc2 s4 VN.t1873 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3980 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3981 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3982 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3983 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3984 fc2 s4 VN.t1872 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3985 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3986 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3987 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3988 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3989 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3990 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3991 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3992 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3993 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3994 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3995 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3996 fc2 s4 VN.t1871 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3997 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3998 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3999 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4000 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4001 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4002 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4003 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4004 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4005 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4007 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4008 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4009 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4010 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4011 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4012 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4013 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4014 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4015 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4017 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4018 fc2 s4 VN.t1870 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4019 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4020 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X4021 VN.t1869 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4022 fc2 s4 VN.t1868 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4023 fc2 s4 VN.t1867 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4024 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4025 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4026 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4027 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4028 VN.t1866 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4029 fc2 s4 VN.t1865 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4030 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4031 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4032 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4033 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4034 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4035 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4036 fc2 s4 VN.t1864 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4037 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4038 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4039 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4040 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4041 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4042 fc2 s4 VN.t1863 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4043 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4044 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4045 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4047 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4048 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4049 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4050 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4051 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4052 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4053 fc2 s4 VN.t1862 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4054 fc2 s4 VN.t1861 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4055 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4056 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4057 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4058 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4059 fc2 s4 VN.t1860 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4060 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4061 VN.t1859 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4062 VN.t1858 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4063 fc2 s4 VN.t1857 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4064 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4065 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4066 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4067 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4068 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4069 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4070 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4071 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4072 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4073 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4074 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4075 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4076 VN.t1856 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4077 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4078 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4079 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4080 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4081 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4082 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4083 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4084 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4085 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4086 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4087 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4088 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4089 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4090 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4091 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4092 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4093 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4094 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4095 fc2 s4 VN.t1855 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4096 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4097 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4098 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4099 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4101 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4102 fc2 s4 VN.t1854 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4103 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4104 VN.t1853 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4105 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4106 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4107 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4108 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4109 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4111 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4112 fc2 s4 VN.t1852 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4113 fc2 s4 VN.t1851 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4114 VN.t1850 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4115 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4116 VN.t1849 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4117 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4119 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4120 VN.t1848 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4121 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4122 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4123 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4124 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4125 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4126 VN.t1847 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4127 fc2 s4 VN.t1846 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4128 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4129 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4130 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4131 fc2 s4 VN.t1845 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4132 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4133 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4134 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4136 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4137 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4138 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4139 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4140 VN.t1844 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4141 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4142 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4143 fc2 s4 VN.t1843 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4144 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4145 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4146 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4147 VN.t1842 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4148 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4149 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4150 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4151 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4152 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4153 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4154 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4155 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4156 VN.t1841 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4157 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4158 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4159 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4160 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4161 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4162 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4163 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4164 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4165 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4166 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4167 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4168 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4169 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4170 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4171 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4172 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4173 VN.t1840 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4174 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4175 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4176 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4177 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4178 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4179 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4180 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4181 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4182 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4183 VN.t1839 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4184 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4185 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4186 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4187 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4188 fc2 s4 VN.t1838 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4189 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4190 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4191 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4192 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4193 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4194 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4195 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4196 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4198 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4199 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4200 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4201 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4202 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4203 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4204 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4205 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4206 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4207 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4208 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4209 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4210 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4211 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4212 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4213 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4214 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4215 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4216 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4217 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4218 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4219 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4220 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4221 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4222 fc2 s4 VN.t1837 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4223 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4224 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4225 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4226 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4227 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4228 VN.t1836 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4229 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4230 VN.t1835 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4231 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4232 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4234 VN.t1834 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4235 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4236 fc2 s4 VN.t1833 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4237 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4238 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4239 fc2 s4 VN.t1832 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4240 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4241 VN.t1831 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4242 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4243 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4244 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4246 VN.t1830 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4247 fc2 s4 VN.t1829 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4248 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4249 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4250 fc2 s4 VN.t1828 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4251 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4252 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4253 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4254 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4255 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4256 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4257 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4258 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4259 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4260 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4261 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4262 fc2 s4 VN.t1827 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4263 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4264 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4265 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4266 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4267 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4268 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4269 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4270 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4271 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4272 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4273 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4274 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4275 fc2 s4 VN.t1826 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4276 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4277 fc2 s4 VN.t1825 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4278 VN.t1824 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4279 fc2 s4 VN.t1823 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4280 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4281 VN.t1822 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4282 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4283 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4284 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4285 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4286 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4287 fc2 s4 VN.t1821 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4288 VN.t1820 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4289 VN.t1819 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4290 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4291 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4292 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4293 fc2 s4 VN.t1818 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4294 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4295 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4296 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4297 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4298 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4299 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4300 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4301 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4302 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4303 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4304 fc2 s4 VN.t1817 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4305 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4306 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4307 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4308 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4309 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4310 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4311 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4312 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4313 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4314 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4315 VN.t1816 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4316 fc2 s4 VN.t1815 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4317 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4318 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4319 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4320 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4321 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4322 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4323 fc2 s4 VN.t1814 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4324 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4325 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4326 fc2 s4 VN.t1813 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4327 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4328 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4329 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4330 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4331 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4332 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4333 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4334 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4335 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4336 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4337 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4339 VN.t1812 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4340 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4341 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4342 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4343 fc2 s4 VN.t1811 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4344 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4345 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4346 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4347 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4348 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4349 fc2 s4 VN.t1810 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4350 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4351 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4352 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4353 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4354 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4355 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4356 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4357 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4358 fc2 s4 VN.t1809 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4359 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4360 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4361 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4362 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4363 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4364 fc2 s4 VN.t1808 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4365 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4366 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4367 VN.t1807 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4368 fc2 s4 VN.t1806 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4369 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4370 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4371 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4372 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4373 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4374 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4375 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4376 VN.t1805 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4377 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4378 VN.t1804 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4379 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4380 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4381 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4382 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4383 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4384 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4385 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X4386 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4387 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4388 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4389 VN.t1803 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4390 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4391 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4392 VN.t1802 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4393 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4394 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4395 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4396 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4397 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4398 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4399 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4400 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4401 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4402 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4403 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4404 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4405 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4406 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4407 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4408 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4409 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4410 fc2 s4 VN.t1801 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4411 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4412 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4413 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4414 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4415 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4416 VN.t1800 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4417 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4418 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4419 VN.t1799 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4420 fc2 s4 VN.t1798 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4421 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4422 VN.t1797 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4423 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4424 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4425 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4426 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4427 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4428 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4429 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4430 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4431 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4432 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4433 VN.t1796 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4434 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4435 fc2 s4 VN.t1795 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4436 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4437 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4438 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4439 VN.t1794 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4440 VN.t1793 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4441 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4442 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4443 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4444 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4445 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4446 VN.t1792 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4447 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4448 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4449 fc2 s4 VN.t1791 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4450 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4451 fc2 s4 VN.t1790 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4452 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4453 VN.t1789 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4454 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4455 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4456 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4457 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4458 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4459 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4460 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4461 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4462 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4463 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4464 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4465 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4466 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4467 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4468 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4469 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4470 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4471 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4472 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4473 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4474 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4475 fc2 s4 VN.t1788 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4476 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4477 VN.t1787 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4478 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4479 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4480 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4481 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4482 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4483 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4484 fc2 s4 VN.t1786 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4485 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4486 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4487 VN.t1785 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4488 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4489 VN.t1784 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4490 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4491 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4492 fc2 s4 VN.t1783 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4493 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4494 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4495 fc2 s4 VN.t1782 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4496 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4497 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4498 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4499 VN.t1781 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4500 fc2 s4 VN.t1780 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4501 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4502 VN.t1779 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4503 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4504 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4505 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4506 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4507 fc2 s4 VN.t1778 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4508 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4509 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4510 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4511 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4512 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4513 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4514 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4515 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4516 fc2 s4 VN.t1777 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4517 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4518 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4519 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4520 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4521 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4522 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4523 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4524 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4525 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4526 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4527 VN.t1776 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4528 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4529 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4530 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4531 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4532 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4533 VN.t1775 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4534 VN.t1774 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4535 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4536 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4537 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4538 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4539 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4540 VN.t1773 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4541 VN.t1772 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4542 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4543 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4544 fc2 s4 VN.t1771 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4545 fc2 s4 VN.t1770 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4546 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4547 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4548 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4549 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4550 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4551 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4552 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4553 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4554 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4555 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4556 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4557 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4558 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4559 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4560 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4561 VN.t1769 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4562 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4563 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4564 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4565 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4566 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4567 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4568 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4569 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4570 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4571 VN.t1768 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4572 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4573 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4574 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4575 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4576 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4577 fc2 s4 VN.t1767 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4578 VN.t1766 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4579 VN.t1765 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4580 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4582 VN.t1764 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4583 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4584 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4585 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4586 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4587 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4588 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4590 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4591 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4592 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4593 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4594 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4595 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4596 VN.t1763 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4597 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4598 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4599 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4600 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4601 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4602 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4603 fc2 s4 VN.t1762 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4604 VN.t1761 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4605 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4606 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4607 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4608 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4609 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4610 VN.t1760 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4611 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4612 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4613 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4614 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4615 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4616 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4618 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4619 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4620 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4622 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4623 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4624 VN.t1759 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4625 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4626 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4627 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4628 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4629 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4630 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4631 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4632 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4633 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4634 VN.t1758 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4635 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4636 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4637 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4638 fc2 s4 VN.t1757 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4639 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4640 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4641 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4642 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4643 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4644 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4645 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4646 VN.t1756 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4647 VN.t1755 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4648 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4649 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4650 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4651 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X4652 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4653 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4654 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4655 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4656 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4657 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4658 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4659 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4660 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4661 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4663 VN.t1754 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4664 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4665 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4666 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4667 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4668 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4669 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4670 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4671 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4672 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4673 fc2 s4 VN.t1753 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4674 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4675 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4676 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4677 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4678 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4679 fc2 s4 VN.t1752 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4680 VN.t1751 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4681 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4682 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4683 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4684 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4685 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4686 fc2 s4 VN.t1750 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4687 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4688 VN.t1749 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4689 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4690 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4691 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4692 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4693 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4694 VN.t1748 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4695 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4696 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4697 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4698 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4699 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4700 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4701 VN.t1747 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4702 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4703 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4704 fc2 s4 VN.t1746 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4705 fc2 s4 VN.t1745 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4706 fc2 s4 VN.t1744 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4707 VN.t1743 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4708 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4709 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4710 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4711 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4712 VN.t1742 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4713 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4714 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4715 VN.t1741 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4716 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4717 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4718 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4719 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4720 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4721 VN.t1740 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4722 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4723 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4724 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X4725 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4726 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4727 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4728 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4729 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4730 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4731 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4732 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4733 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4734 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4735 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4736 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4737 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4739 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4740 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4741 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4742 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4743 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4744 fc2 s4 VN.t1739 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4745 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4746 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4747 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4748 VN.t1738 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4749 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4750 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4751 VN.t1737 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4752 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4753 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4754 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4755 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4756 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4757 VN.t1736 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4758 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4760 VN.t1735 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4761 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4762 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4763 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4764 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4765 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4766 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4767 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4768 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4769 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4770 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4771 fc2 s4 VN.t1734 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4772 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4773 fc2 s4 VN.t1733 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4774 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4775 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4776 VN.t1732 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4777 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4778 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4779 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4780 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4781 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4782 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4783 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4784 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4785 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4786 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4787 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4788 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4789 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4790 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4791 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4792 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4793 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4794 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4795 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4796 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4797 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4798 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4799 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4800 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4801 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4802 VN.t1731 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4803 VN.t1730 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4804 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4805 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4806 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4807 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4808 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4809 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4810 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4811 VN.t1729 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4812 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4813 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4814 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4815 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4816 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4817 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4818 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4819 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4820 fc2 s4 VN.t1728 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4821 VN.t1727 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4822 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4823 VN.t1726 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4824 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4825 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4826 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4827 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4828 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4829 VN.t1725 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4830 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4831 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4832 VN.t1724 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4833 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4834 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4835 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4836 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4837 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4838 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4839 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4840 VN.t1723 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4841 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4842 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4843 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4844 VN.t1722 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4845 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4846 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4847 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4848 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4849 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4850 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4851 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4852 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4853 VN.t1721 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4854 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4855 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4856 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4857 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4858 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4859 VN.t1720 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4860 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4861 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4862 fc2 s4 VN.t1719 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4863 fc2 s4 VN.t1718 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4864 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4865 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4866 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4867 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4868 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4869 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4870 VN.t1717 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4871 fc2 s4 VN.t1716 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4872 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4873 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4874 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4875 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4876 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4877 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4878 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4879 VN.t1715 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4880 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4881 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4882 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4883 VN.t1714 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4884 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X4885 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4886 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4887 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4888 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4889 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4890 VN.t1713 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4891 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4892 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4894 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4895 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4896 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4897 VN.t1712 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4898 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4899 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4900 VN.t1711 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4901 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4902 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4903 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4904 fc2 s4 VN.t1710 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4905 fc2 s4 VN.t1709 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4906 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4907 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4908 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4909 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4910 VN.t1708 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4911 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4912 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4913 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4914 fc2 s4 VN.t1707 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4915 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4916 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4917 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4918 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4919 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4920 VN.t1706 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4921 fc2 s4 VN.t1705 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4922 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4923 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4924 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4925 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4926 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4927 fc2 s4 VN.t1704 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4928 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4929 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4930 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4931 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4932 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4933 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4934 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4935 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4936 fc2 s4 VN.t1703 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4937 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4938 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4939 VN.t1702 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4940 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4941 fc2 s4 VN.t1701 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4942 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4943 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4944 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4945 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4946 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4947 fc2 s4 VN.t1700 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4948 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4949 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4950 VN.t1699 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4951 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4952 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4953 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4954 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4955 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4956 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4957 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4958 fc2 s4 VN.t1698 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4959 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4960 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4961 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4962 VN.t1697 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4963 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4964 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4965 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4966 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4967 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4968 VN.t1696 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4969 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4970 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4971 VN.t1695 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4972 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4973 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4974 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4975 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4976 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4977 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4978 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4979 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4980 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4981 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4982 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4983 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4984 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4985 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4986 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4987 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4988 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4989 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4990 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4991 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4992 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4993 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4994 VN.t1694 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4995 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4996 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4997 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4998 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4999 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5000 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5001 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5002 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5003 fc2 s4 VN.t1693 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5004 VN.t1692 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5005 fc2 s4 VN.t1691 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5007 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5009 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5010 fc2 s4 VN.t1690 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5011 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5012 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5013 fc2 s4 VN.t1689 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5014 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5015 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5016 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5017 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5018 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5019 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5020 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5021 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5022 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5023 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5024 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5025 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5026 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5027 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5028 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5029 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5030 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5031 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5032 fc2 s4 VN.t1688 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5033 VN.t1687 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5034 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5035 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5036 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5037 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5038 fc2 s4 VN.t1686 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5039 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5040 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5041 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5042 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5043 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5044 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5045 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5047 VN.t1685 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5048 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5049 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5050 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5051 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5052 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5053 fc2 s4 VN.t1684 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5054 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5055 fc2 s4 VN.t1683 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5056 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5057 VN.t1682 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5058 VN.t1681 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5059 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5060 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5061 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5062 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5063 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5064 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5065 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5066 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5067 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5068 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5069 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5070 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5071 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5072 fc2 s4 VN.t1680 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5073 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5074 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5075 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5076 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5077 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5078 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5079 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5080 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5081 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5082 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5083 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5084 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5085 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5086 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5087 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5088 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5089 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5090 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5091 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5092 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5093 fc2 s4 VN.t1679 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5094 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5095 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5096 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5097 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5098 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5099 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5101 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5102 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5103 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5104 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5105 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5106 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5107 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5108 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5109 fc2 s4 VN.t1678 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5111 VN.t1677 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5112 VN.t1676 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5113 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5114 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5115 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5116 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5117 VN.t1675 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5118 VN.t1674 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5119 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5120 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5121 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5122 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5123 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5124 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5125 fc2 s4 VN.t1673 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5126 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5127 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5128 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5129 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5130 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5131 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5132 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5133 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5134 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5135 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5136 fc2 s4 VN.t1672 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5137 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5138 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5139 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5140 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5141 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5142 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5143 VN.t1671 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5144 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5145 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5146 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5147 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5148 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5149 fc2 s4 VN.t1670 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5150 VN.t1669 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5151 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5152 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5153 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5154 fc2 s4 VN.t1668 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5156 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5157 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5158 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5159 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5160 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5161 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5162 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5163 fc2 s4 VN.t1667 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5164 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5165 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5166 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5167 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5168 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5169 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5170 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5171 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5172 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5173 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5174 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5175 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5176 VN.t1666 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5177 fc2 s4 VN.t1665 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5178 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5180 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5181 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5182 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5183 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5184 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5185 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5186 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5187 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5188 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5189 fc2 s4 VN.t1664 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5190 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5191 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5192 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5193 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5194 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5195 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5196 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5198 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5199 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5200 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5201 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5202 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5203 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5205 fc2 s4 VN.t1663 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5206 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5208 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5209 VN.t1662 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5210 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5211 VN.t1661 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5212 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5213 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5214 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5215 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5216 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5217 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5218 fc2 s4 VN.t1660 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5219 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5220 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5221 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5222 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5223 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5224 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5225 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5226 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5227 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5228 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5229 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5230 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5231 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5232 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5233 fc2 s4 VN.t1659 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5234 fc2 s4 VN.t1658 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5235 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5236 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5237 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5238 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5239 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5240 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5241 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5242 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5243 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5244 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5246 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5247 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5248 fc2 s4 VN.t1657 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5249 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5250 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5251 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5252 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5253 VN.t1656 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5254 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5255 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5256 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5257 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5258 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5259 fc2 s4 VN.t1655 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5260 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5261 VN.t1654 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5262 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5263 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5264 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5265 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5266 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5267 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5268 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5269 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5270 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5271 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5272 fc2 s4 VN.t1653 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5273 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5274 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5275 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5276 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5278 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5279 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5280 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5281 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5282 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5283 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5284 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5285 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5286 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5287 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5288 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5290 fc2 s4 VN.t1652 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5291 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5292 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5293 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5295 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5296 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5297 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5298 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5299 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5300 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5301 VN.t1651 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5302 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5303 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5304 fc2 s4 VN.t1650 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5305 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5306 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5307 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5308 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5309 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5310 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5311 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5312 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5313 fc2 s4 VN.t1649 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5314 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5315 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5316 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5317 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5318 fc2 s4 VN.t1648 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5319 fc2 s4 VN.t1647 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5320 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5321 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5322 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5323 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5324 VN.t1646 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5325 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5326 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5327 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5328 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5329 VN.t1645 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5330 fc2 s4 VN.t1644 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5331 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5332 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5333 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5334 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5335 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5336 fc2 s4 VN.t1643 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5337 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5339 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5340 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5341 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5342 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5343 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5344 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5345 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5346 fc2 s4 VN.t1642 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5347 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5348 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5349 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5350 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5351 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5352 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5353 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5354 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5355 fc2 s4 VN.t1641 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5356 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5357 VN.t1640 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5358 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5359 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5360 fc2 s4 VN.t1639 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5361 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5362 VN.t1638 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5363 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5364 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5365 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5366 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5367 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5368 fc2 s4 VN.t1637 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5369 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5370 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5371 fc2 s4 VN.t1636 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5372 fc2 s4 VN.t1635 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5373 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5374 VN.t1634 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5375 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5377 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5378 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5379 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5380 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5381 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5382 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5383 VN.t1633 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5384 fc2 s4 VN.t1632 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5385 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5386 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5387 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5388 VN.t1631 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5389 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5390 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5391 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5392 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5393 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5394 VN.t1630 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5395 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5396 fc2 s4 VN.t1629 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5397 VN.t1628 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5398 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5399 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5400 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5401 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5402 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5403 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5404 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5405 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5406 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5407 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5408 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5409 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5410 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5411 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5412 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5413 VN.t1627 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5414 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5415 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5416 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5417 VN.t1626 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5418 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5419 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5420 VN.t1625 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5421 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5422 VN.t1624 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5423 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5424 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5425 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5426 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5427 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5428 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5429 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5430 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5431 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5432 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5433 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5435 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5436 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5437 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5438 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5439 VN.t1623 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5440 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5441 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5442 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5443 fc2 s4 VN.t1622 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5444 VN.t1621 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5445 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5446 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5447 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5448 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5449 fc2 s4 VN.t1620 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5450 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5451 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5452 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5453 fc2 s4 VN.t1619 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5454 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5455 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5456 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5457 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5458 fc2 s4 VN.t1618 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5459 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5460 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5461 VN.t1617 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5462 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5463 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5464 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5465 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5466 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5467 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5468 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5469 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5470 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5471 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5472 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5473 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5474 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5475 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5476 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5477 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5478 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5479 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5480 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5481 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5482 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5483 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5484 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5485 fc2 s4 VN.t1616 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5486 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5487 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5488 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5489 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5490 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5491 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5492 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5493 VN.t1615 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5494 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5495 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5496 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5497 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5498 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5499 fc2 s4 VN.t1614 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5500 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5502 fc2 s4 VN.t1613 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5503 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5504 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5505 VN.t1612 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5506 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5507 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5508 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5509 VN.t1611 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5510 VN.t1610 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5511 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5512 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5513 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5514 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5515 fc2 s4 VN.t1609 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5516 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5517 fc2 s4 VN.t1608 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5518 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5519 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5520 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5521 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5522 VN.t1607 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5523 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5524 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5525 fc2 s4 VN.t1606 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5526 VN.t1605 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5527 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5528 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5529 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5530 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X5531 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5532 fc2 s4 VN.t1604 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5533 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5534 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5535 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5536 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5537 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5538 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5539 fc2 s4 VN.t1603 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5540 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5541 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5542 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5543 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5544 fc2 s4 VN.t1602 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5545 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5546 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5547 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5548 fc2 s4 VN.t1601 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5549 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5550 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5551 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5552 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5553 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5554 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5555 fc2 s4 VN.t1600 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5556 VN.t1599 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5557 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5558 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5559 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5560 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5561 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5562 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5563 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5564 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5565 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5566 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5567 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5568 VN.t1598 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5569 fc2 s4 VN.t1597 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5570 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5571 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5572 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5573 VN.t1596 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5574 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5575 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5576 fc2 s4 VN.t1595 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5577 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5578 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5579 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5580 fc2 s4 VN.t1594 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5581 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5582 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5583 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5584 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5585 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5586 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5587 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5588 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5589 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5590 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5591 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5592 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5593 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5594 VN.t1593 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5595 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5596 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5597 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5598 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5599 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5600 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5601 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5602 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5603 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5604 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5605 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5606 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5607 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5608 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5609 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5610 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5611 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5612 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5613 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5614 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5615 fc2 s4 VN.t1592 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5616 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5617 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5618 VN.t1591 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5619 fc2 s4 VN.t1590 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5620 fc2 s4 VN.t1589 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5622 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5623 VN.t1588 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5624 fc2 s4 VN.t1587 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5625 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5626 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5627 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5628 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5629 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5630 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5631 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5632 fc2 s4 VN.t1586 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5633 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5634 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5635 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5636 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5637 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5638 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5639 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5640 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5641 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5642 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5643 fc2 s4 VN.t1585 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5644 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5645 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5646 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5647 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5648 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5649 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5650 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5651 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5652 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5653 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5654 fc2 s4 VN.t1584 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5655 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5656 VN.t1583 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5657 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5658 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5659 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5660 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5661 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5662 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5663 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5664 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5665 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5666 fc2 s4 VN.t1582 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5667 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5668 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5669 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5670 VN.t1581 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5671 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5672 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5673 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5674 VN.t1580 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5675 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5676 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5677 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5678 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5679 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5680 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5681 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5682 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5683 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5684 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5685 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5686 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5687 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5688 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5689 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5690 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5691 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5692 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5693 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5694 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5695 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5696 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5697 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5698 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5699 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5700 fc2 s4 VN.t1579 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5701 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5702 VN.t1578 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5703 fc2 s4 VN.t1577 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5704 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5705 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5706 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5707 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5708 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5709 VN.t1576 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5710 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5711 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5712 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5713 VN.t1575 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5714 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5715 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5716 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5717 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5718 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5719 fc2 s4 VN.t1574 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5720 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5721 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5722 fc2 s4 VN.t1573 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5723 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5724 VN.t1572 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5725 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5726 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5727 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5728 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5729 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5730 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5731 VN.t1571 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5732 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5733 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5734 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5735 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5736 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5737 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5738 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5739 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5740 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5741 VN.t1570 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5742 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5743 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5744 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5745 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5746 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5747 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5748 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5749 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5750 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5751 VN.t1569 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5752 fc2 s4 VN.t1568 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5753 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5754 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5755 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5756 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5757 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5758 VN.t1567 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5760 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5761 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5762 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5763 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5764 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5765 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5766 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5767 VN.t1566 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5768 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5769 fc2 s4 VN.t1565 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5770 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5771 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5772 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5773 VN.t1564 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5774 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5775 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5776 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5777 VN.t1563 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5778 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5779 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5780 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5781 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5782 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5783 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5784 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5785 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5786 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5787 fc2 s4 VN.t1562 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5788 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5789 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5790 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5791 VN.t1561 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5792 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5793 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5794 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5795 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5796 fc2 s4 VN.t1560 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5797 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5798 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5799 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5800 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5801 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5802 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5803 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5804 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5805 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5806 VN.t1559 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5807 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5808 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5809 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5810 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5811 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5812 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5813 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5814 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5815 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5816 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5817 fc2 s4 VN.t1558 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5818 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5819 fc2 s4 VN.t1557 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5820 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5821 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5822 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5823 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5824 VN.t1556 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5825 VN.t1555 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5826 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5827 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5828 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5829 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5830 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5831 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5832 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5833 VN.t1554 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5834 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5835 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5836 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5837 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5838 VN.t1553 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5839 fc2 s4 VN.t1552 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5840 fc2 s4 VN.t1551 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5841 VN.t1550 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5842 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5844 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5845 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5846 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5847 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5848 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5849 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5850 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5851 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5852 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5853 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5854 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5855 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5856 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5857 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5858 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5859 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5860 fc2 s4 VN.t1549 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5861 fc2 s4 VN.t1548 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5862 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5863 VN.t1547 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5864 fc2 s4 VN.t1546 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5865 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5866 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5867 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5868 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5869 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5870 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5871 VN.t1545 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5872 VN.t1544 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5873 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5874 fc2 s4 VN.t1543 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5875 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5876 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5877 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5878 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5879 VN.t1542 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X5880 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5881 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5882 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5883 fc2 s4 VN.t1541 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5884 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5886 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5887 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5888 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5889 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5890 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5891 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5892 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5893 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5894 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5895 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5896 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5897 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5898 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5899 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5900 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5901 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5902 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5904 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5905 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5906 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5907 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5908 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5909 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5910 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5911 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5912 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5913 VN.t1540 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5914 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5915 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5916 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5917 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5918 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5919 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5920 fc2 s4 VN.t1539 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5921 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5922 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5923 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5924 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5925 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5926 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5927 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5929 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5930 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5931 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5932 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5933 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5934 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5935 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5936 fc2 s4 VN.t1538 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5937 fc2 s4 VN.t1537 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5938 VN.t1536 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5939 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X5940 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5941 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5942 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5943 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5944 fc2 s4 VN.t1535 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5945 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5946 fc2 s4 VN.t1534 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5947 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5948 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5949 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5950 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5951 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5952 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5953 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5954 VN.t1533 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5955 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5956 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5957 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5958 VN.t1532 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5959 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5960 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5961 fc2 s4 VN.t1531 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5962 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5963 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5964 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5965 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5966 fc2 s4 VN.t1530 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5967 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5968 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X5969 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5970 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5971 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5972 VN.t1529 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X5973 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5974 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5975 VN.t1528 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X5976 fc2 s4 VN.t1527 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5977 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5978 VN.t1526 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5979 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5980 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5981 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5982 fc2 s4 VN.t1525 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5983 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5984 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5985 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5986 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5987 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5988 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5989 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5990 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5991 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5992 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5993 fc2 s4 VN.t1524 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5994 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5995 VN.t1523 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5996 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5997 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5998 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X5999 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6000 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6001 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6002 fc2 s4 VN.t1522 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6003 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6004 VN.t1521 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6005 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6007 VN.t1520 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6009 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6010 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6011 fc2 s4 VN.t1519 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6012 VN.t1518 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6013 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6014 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6015 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6017 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6018 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6019 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6020 VN.t1517 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6021 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6022 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6023 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6024 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6025 VN.t1516 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6026 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6027 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6028 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6029 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6030 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6031 fc2 s4 VN.t1515 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6032 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6033 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6034 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6035 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6036 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6037 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6038 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6039 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6040 VN.t1514 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6041 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6042 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6043 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6044 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6045 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6046 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6047 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6048 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6049 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6050 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6051 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6052 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6053 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6054 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6055 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6056 fc2 s4 VN.t1513 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6057 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6058 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6059 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6060 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6061 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6062 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6063 VN.t1512 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6064 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6065 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6066 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6067 fc2 s4 VN.t1511 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6068 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6069 VN.t1510 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6070 fc2 s4 VN.t1509 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6071 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6072 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6073 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6074 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6075 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6076 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6077 VN.t1508 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6078 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6079 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6080 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6081 VN.t1507 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6082 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6083 fc2 s4 VN.t1506 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6084 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6085 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6086 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6087 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6088 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6089 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6090 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6091 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6092 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6093 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6094 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6095 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6096 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6097 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6098 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6099 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6100 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6101 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6102 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6103 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6104 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6105 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6106 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6107 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6108 VN.t1505 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6109 VN.t1504 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6110 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6111 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6112 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6113 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6114 VN.t1503 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6115 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6116 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6117 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6118 VN.t1502 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6119 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6120 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6121 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6122 VN.t1501 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6123 VN.t1500 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6124 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6125 VN.t1499 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6126 fc2 s4 VN.t1498 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6127 fc2 s4 VN.t1497 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6128 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6129 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6130 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6131 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6132 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6133 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6134 fc2 s4 VN.t1496 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6136 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6137 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6138 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6139 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6140 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6141 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6142 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6143 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6144 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6145 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6146 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6147 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6148 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6149 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6150 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6151 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6152 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6153 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6154 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6155 fc2 s4 VN.t1495 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6156 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6157 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6158 VN.t1494 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6159 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6160 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6161 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6162 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6163 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6164 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6165 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6166 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6167 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6168 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6169 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6170 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6171 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6172 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6173 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6174 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6175 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6176 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6177 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6178 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6180 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6181 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6182 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6183 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6184 VN.t1493 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6185 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6186 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6187 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6188 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6189 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6190 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6191 fc2 s4 VN.t1492 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6192 VN.t1491 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6193 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6194 fc2 s4 VN.t1490 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6195 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6196 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6198 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6199 VN.t1489 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6200 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6201 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6202 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6203 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6205 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6206 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6207 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6208 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6209 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6210 VN.t1488 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6211 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6212 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6213 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6214 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6215 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6216 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6217 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6218 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6219 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6220 fc2 s4 VN.t1487 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6221 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6222 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6223 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6224 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6225 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6226 fc2 s4 VN.t1486 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6227 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6228 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6229 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6230 VN.t1485 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6231 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6232 fc2 s4 VN.t1484 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6233 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6234 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6235 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6236 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6237 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6238 fc2 s4 VN.t1483 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6239 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6240 VN.t1482 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6241 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6242 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6243 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6244 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6245 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6246 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6247 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6248 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6249 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6250 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6251 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6252 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6253 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6254 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6255 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6256 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6257 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6258 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6259 VN.t1481 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6260 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6261 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6262 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6263 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6264 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6265 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6266 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6267 fc2 s4 VN.t1480 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6268 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6269 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6270 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6271 fc2 s4 VN.t1479 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6272 VN.t1478 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6273 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6274 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6275 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6276 VN.t1477 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6277 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6278 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6279 fc2 s4 VN.t1476 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6280 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6281 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6282 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6283 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6284 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6285 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6286 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6287 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6288 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6290 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6291 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6292 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6293 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6294 fc2 s4 VN.t1475 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6295 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6296 fc2 s4 VN.t1474 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6297 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6298 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6299 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6300 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6301 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6302 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6303 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6304 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6305 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6306 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6307 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6308 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6309 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6310 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6311 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6312 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6313 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6314 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6315 fc2 s4 VN.t1473 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6316 VN.t1472 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6317 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6318 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6319 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6320 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6321 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6322 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6323 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6324 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6325 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6326 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X6327 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6328 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6329 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6330 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6331 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6332 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6333 fc2 s4 VN.t1471 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6334 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6335 VN.t1470 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6336 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6337 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6338 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6339 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6340 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6341 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6342 VN.t1469 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6343 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6344 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6345 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6346 VN.t1468 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6347 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6348 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6349 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6350 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6351 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6352 fc2 s4 VN.t1467 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6353 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6354 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6355 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6356 fc2 s4 VN.t1466 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6357 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6358 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6359 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6360 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6361 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6362 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6363 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6364 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6365 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6366 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6367 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6368 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6369 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6370 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6372 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6373 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6374 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6375 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6377 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6378 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6379 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6380 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6381 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6382 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6383 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6384 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6385 VN.t1465 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6386 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6387 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6388 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6389 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6390 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6391 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6392 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6393 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6394 VN.t1464 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6395 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6396 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6397 VN.t1463 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6398 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6399 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6400 fc2 s4 VN.t1462 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6401 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6402 fc2 s4 VN.t1461 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6403 VN.t1460 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6404 fc2 s4 VN.t1459 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6405 VN.t1458 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6406 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6407 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6408 fc2 s4 VN.t1457 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6409 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6410 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6411 fc2 s4 VN.t1456 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6412 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6413 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6414 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6415 VN.t1455 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6416 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6417 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6418 fc2 s4 VN.t1454 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6419 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6420 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6421 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6422 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6423 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6424 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6425 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6426 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6427 VN.t1453 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6428 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6429 fc2 s4 VN.t1452 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6430 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6431 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6432 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6433 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6435 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6436 VN.t1451 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6437 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6438 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6439 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6440 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6441 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6442 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6443 fc2 s4 VN.t1450 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6444 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6445 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6446 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6447 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6448 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6449 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6450 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6451 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6452 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6453 VN.t1449 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6454 VN.t1448 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6455 VN.t1447 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6456 fc2 s4 VN.t1446 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6457 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6458 fc2 s4 VN.t1445 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6459 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6460 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6461 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6462 VN.t1444 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6463 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6464 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6465 fc2 s4 VN.t1443 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6466 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6467 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6468 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6469 VN.t1442 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6470 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6471 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6472 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6473 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6474 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6475 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6476 fc2 s4 VN.t1441 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6477 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6478 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6479 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6480 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6481 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6482 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6483 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6484 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6485 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6486 VN.t1440 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6487 fc2 s4 VN.t1439 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6488 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6489 VN.t1438 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6490 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6491 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6492 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6493 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6494 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6495 VN.t1437 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6496 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6497 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6498 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6499 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6500 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6501 fc2 s4 VN.t1436 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6502 fc2 s4 VN.t1435 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6503 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6504 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6505 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6506 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6507 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6508 fc2 s4 VN.t1434 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6509 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6510 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6511 VN.t1433 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6512 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6513 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6514 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6515 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6516 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6517 fc2 s4 VN.t1432 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6518 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6519 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6520 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6521 fc2 s4 VN.t1431 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6522 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6523 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6524 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6525 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6526 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6527 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6528 fc2 s4 VN.t1430 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6529 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6530 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6531 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6532 fc2 s4 VN.t1429 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6533 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6534 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6535 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6536 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6537 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6538 fc2 s4 VN.t1428 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6539 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6540 VN.t1427 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6541 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6542 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6543 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6544 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6545 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6546 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6547 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6548 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6549 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6550 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6551 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6552 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6553 fc2 s4 VN.t1426 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6554 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6555 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6556 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6557 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6558 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6559 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6560 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6561 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6562 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6563 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6564 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6565 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6566 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6567 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6568 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6569 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6570 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6571 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6572 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6573 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6574 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6575 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6576 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6577 fc2 s4 VN.t1425 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6578 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6579 VN.t1424 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6580 fc2 s4 VN.t1423 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6581 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6582 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6583 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6584 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6585 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6586 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6587 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6588 VN.t1422 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6589 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6590 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6591 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6592 fc2 s4 VN.t1421 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6593 VN.t1420 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6594 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6595 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6596 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6597 fc2 s4 VN.t1419 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6598 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6599 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6600 fc2 s4 VN.t1418 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6601 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6602 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6603 VN.t1417 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6604 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6605 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6606 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6607 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6608 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6609 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6610 VN.t1416 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6611 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6612 fc2 s4 VN.t1415 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6613 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6614 VN.t1414 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6615 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6616 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6617 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6618 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6619 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6620 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6622 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6623 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6624 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6625 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6626 fc2 s4 VN.t1413 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6627 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6628 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6629 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6630 VN.t1412 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6631 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6632 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6633 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6634 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6635 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6636 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6637 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6638 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6639 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6640 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6641 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6643 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6644 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6645 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6646 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6647 VN.t1411 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6648 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6649 fc2 s4 VN.t1410 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6650 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6651 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6652 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6653 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6654 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6655 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6656 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6657 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6658 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6659 fc2 s4 VN.t1409 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6660 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6661 VN.t1408 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6662 fc2 s4 VN.t1407 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6663 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6664 fc2 s4 VN.t1406 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6665 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6666 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6667 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6668 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6669 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6670 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6671 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6672 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6673 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6674 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6675 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6676 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6677 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6678 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6679 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6680 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6681 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6682 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6683 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6684 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6685 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6686 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6687 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6688 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6689 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6690 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6691 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6692 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6693 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6694 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6695 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6696 fc2 s4 VN.t1405 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6697 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6698 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6699 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6700 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6701 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6702 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6703 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6704 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6705 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6706 fc2 s4 VN.t1404 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6707 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6708 fc2 s4 VN.t1403 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6709 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6710 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6711 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6712 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6713 VN.t1402 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6714 VN.t1401 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6715 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6716 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6717 VN.t1400 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6718 VN.t1399 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6719 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6720 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6721 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6722 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6723 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6724 fc2 s4 VN.t1398 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6725 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6726 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6727 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6728 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6729 fc2 s4 VN.t1397 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6730 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6731 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6732 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6733 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6734 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6735 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6736 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6737 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6739 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6740 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6741 VN.t1396 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6742 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6743 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6744 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6745 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6746 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6747 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6748 fc2 s4 VN.t1395 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6749 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6750 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6751 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6752 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6753 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6754 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6755 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6756 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6757 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X6758 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6759 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6760 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6761 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6762 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6763 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6764 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6765 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6766 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6767 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6768 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6769 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6770 VN.t1394 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6771 fc2 s4 VN.t1393 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6772 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6773 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6774 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6775 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6776 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6777 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6778 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6779 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6780 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6781 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6782 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6783 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6784 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6785 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6786 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6787 fc2 s4 VN.t1392 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6788 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6789 fc2 s4 VN.t1391 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6790 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6791 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6792 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6793 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6794 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6795 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6796 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6797 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6798 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6799 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6800 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6801 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6802 VN.t1390 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6803 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6804 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6805 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6806 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6807 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6808 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6809 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6810 fc2 s4 VN.t1389 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6811 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6812 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6813 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6814 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6815 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6816 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6817 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6818 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6819 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6820 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6821 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6822 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6823 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6824 fc2 s4 VN.t1388 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6825 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6826 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6827 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6828 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6829 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6830 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6831 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6832 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6833 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6834 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6835 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6836 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6837 fc2 s4 VN.t1387 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6838 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6839 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6840 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6841 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6842 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6843 VN.t1386 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6844 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6845 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6846 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X6847 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6848 fc2 s4 VN.t1385 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6849 VN.t1384 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6850 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6851 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6852 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6853 VN.t1383 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6854 VN.t1382 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6855 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6856 fc2 s4 VN.t1381 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6857 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6858 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6859 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6860 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6861 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6862 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6863 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6864 fc2 s4 VN.t1380 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6865 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X6866 fc2 s4 VN.t1379 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6867 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6868 fc2 s4 VN.t1378 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6869 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6870 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6871 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6872 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6873 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6874 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6875 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6876 fc2 s4 VN.t1377 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6877 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6878 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6879 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6880 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6881 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X6882 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6883 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6884 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6886 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6887 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6888 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6889 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6890 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6891 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6892 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6893 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6894 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6895 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6896 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6897 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6898 fc2 s4 VN.t1376 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6899 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6900 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6901 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6902 fc2 s4 VN.t1375 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6903 VN.t1374 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6904 fc2 s4 VN.t1373 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6905 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6906 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6907 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6908 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6909 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6910 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6911 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6912 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6913 VN.t1372 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6914 fc2 s4 VN.t1371 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6915 fc2 s4 VN.t1370 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6916 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6917 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6918 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6919 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6920 VN.t1369 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6921 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6922 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6923 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6924 VN.t1368 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6925 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6926 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6927 VN.t1367 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6928 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6929 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6930 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6931 fc2 s4 VN.t1366 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6932 fc2 s4 VN.t1365 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6933 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6934 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6935 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6936 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6937 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6938 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6939 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X6940 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6941 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6942 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6943 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6944 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6945 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6946 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6947 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6948 VN.t1364 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6949 fc2 s4 VN.t1363 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6950 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6951 VN.t1362 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6952 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X6953 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6954 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6955 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6956 fc2 s4 VN.t1361 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6957 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6958 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6959 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6960 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6961 fc2 s4 VN.t1360 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6962 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6963 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6964 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6965 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6966 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6967 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6968 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6969 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6970 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6971 VN.t1359 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6972 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6973 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6974 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6975 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6976 VN.t1358 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6977 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6978 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6979 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6980 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6981 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6982 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6983 fc2 s4 VN.t1357 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6984 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6985 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6986 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6987 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6988 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X6989 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6990 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6991 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6992 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6993 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6994 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6995 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6996 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6998 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6999 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7000 VN.t1356 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7001 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7002 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7003 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7004 fc2 s4 VN.t1355 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X7005 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7006 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7007 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7008 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7009 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7010 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7011 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7012 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7013 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7014 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7015 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7016 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7017 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7018 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7019 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7020 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7021 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7022 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7023 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7024 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7025 VN.t1354 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7026 VN.t1353 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7027 fc2 s4 VN.t1352 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7028 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7029 fc2 s4 VN.t1351 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7030 fc2 s4 VN.t1350 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7031 VN.t1349 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7032 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7033 fc2 s4 VN.t1348 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7034 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7035 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7036 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7037 fc2 s4 VN.t1347 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7038 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7039 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7040 fc2 s4 VN.t1346 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7041 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7042 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7043 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7044 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7045 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7046 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7047 VN.t1345 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7048 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7049 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7050 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7051 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7052 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7053 VN.t1344 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7054 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7055 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7056 VN.t1343 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7057 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7058 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7059 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7060 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7061 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7062 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7063 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7064 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7065 VN.t1342 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7066 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7068 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7069 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7070 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7071 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7072 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7073 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7074 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7075 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7076 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7077 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7078 VN.t1341 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7079 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7080 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7081 fc2 s4 VN.t1340 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7082 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7083 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7084 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7085 VN.t1339 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7086 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7088 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7089 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7090 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7091 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7092 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7093 VN.t1338 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7094 fc2 s4 VN.t1337 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7095 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7096 fc2 s4 VN.t1336 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7097 fc2 s4 VN.t1335 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7098 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7099 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7100 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7101 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7102 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7103 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7104 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7105 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7106 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7107 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7108 VN.t1334 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7109 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7111 VN.t1333 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7112 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7113 fc2 s4 VN.t1332 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7114 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7116 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7117 VN.t1331 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7118 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7119 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7120 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7121 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7122 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7123 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7124 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7125 fc2 s4 VN.t1330 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7126 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7127 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7128 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7129 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7130 fc2 s4 VN.t1329 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7131 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7132 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7133 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7134 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7135 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7136 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7137 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7138 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7139 fc2 s4 VN.t1328 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7140 fc2 s4 VN.t1327 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7141 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7142 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7143 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7144 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7145 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7146 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7147 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7148 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7149 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7150 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7151 fc2 s4 VN.t1326 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7152 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7153 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7154 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7156 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7157 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7158 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7159 VN.t1325 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7160 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7161 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7162 VN.t1324 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7163 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7164 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7165 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7166 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7167 fc2 s4 VN.t1323 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7168 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7169 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7170 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7171 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7172 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7173 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7174 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7175 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7176 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7177 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7178 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7179 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7180 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7181 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7182 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7183 VN.t1322 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7184 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7185 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7186 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7187 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7188 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7189 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7190 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7191 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7192 fc2 s4 VN.t1321 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7193 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7194 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7195 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7196 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7197 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7198 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7199 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7200 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7201 fc2 s4 VN.t1320 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7202 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7203 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7204 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7205 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7206 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7207 VN.t1319 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7208 fc2 s4 VN.t1318 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7209 fc2 s4 VN.t1317 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7210 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7211 fc2 s4 VN.t1316 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7212 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7213 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7214 VN.t1315 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7215 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7216 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7217 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7218 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7219 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7220 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7221 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7222 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7223 fc2 s4 VN.t1314 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7224 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7225 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7226 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7227 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7228 fc2 s4 VN.t1313 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7229 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7230 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7231 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7232 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7234 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7235 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7236 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7237 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7238 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7239 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7240 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7241 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7242 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7243 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7244 VN.t1312 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7246 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7247 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7248 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7249 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7250 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7251 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7252 VN.t1311 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7253 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7254 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7255 VN.t1310 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7256 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7257 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7258 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7259 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7260 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7261 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7262 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7263 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7264 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7265 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7266 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7267 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7268 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7269 fc2 s4 VN.t1309 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7270 VN.t1308 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7271 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7272 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7273 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7274 VN.t1307 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7275 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7276 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7278 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7279 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7280 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7281 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7282 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7283 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7284 fc2 s4 VN.t1306 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7285 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7286 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7287 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7288 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7289 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7290 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7291 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7292 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7293 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7295 fc2 s4 VN.t1305 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7296 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7297 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7298 fc2 s4 VN.t1304 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7299 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7300 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7301 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7302 fc2 s4 VN.t1303 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7303 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7304 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7305 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7306 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7307 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7308 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7309 VN.t1302 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7310 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7311 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7312 VN.t1301 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7313 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7314 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7315 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7316 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7317 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7318 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7319 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7320 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7321 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7322 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7323 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7324 fc2 s4 VN.t1300 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7325 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7326 VN.t1299 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7327 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7328 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7329 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7330 VN.t1298 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7331 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7332 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7333 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7334 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7335 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7336 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7337 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7339 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7340 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7341 VN.t1297 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7342 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7343 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7344 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7345 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7346 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7347 fc2 s4 VN.t1296 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7348 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7349 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7350 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7351 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7352 VN.t1295 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7353 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7354 fc2 s4 VN.t1294 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7355 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7356 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7357 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7358 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7359 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7360 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7361 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7362 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7363 VN.t1293 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7364 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7365 fc2 s4 VN.t1292 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7366 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7367 VN.t1291 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7368 VN.t1290 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7369 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7370 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7372 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7373 VN.t1289 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7374 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7375 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7376 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7377 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7378 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7379 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7380 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7381 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7382 fc2 s4 VN.t1288 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7383 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7384 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7385 VN.t1287 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7386 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7387 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7388 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7389 VN.t1286 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7390 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7391 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7392 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7393 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7394 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7395 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7396 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7397 VN.t1285 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7398 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7399 VN.t1284 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7400 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7401 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7402 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7403 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7404 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7405 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7406 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7407 fc2 s4 VN.t1283 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7408 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7409 VN.t1282 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7410 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7411 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7412 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7413 VN.t1281 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7414 VN.t1280 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7415 VN.t1279 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7416 VN.t1278 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7417 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7418 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7419 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7420 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7421 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7422 VN.t1277 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7423 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7424 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7425 VN.t1276 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7426 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7427 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7428 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7429 fc2 s4 VN.t1275 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7430 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7431 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7432 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7433 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7435 VN.t1274 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7436 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7437 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7438 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7439 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7440 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7441 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7442 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7443 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7444 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7445 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7446 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7447 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7448 fc2 s4 VN.t1273 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7449 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7450 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7451 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7452 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7453 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7454 fc2 s4 VN.t1272 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7455 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7456 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7457 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7458 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7459 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7460 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7461 VN.t1271 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7462 VN.t1270 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7463 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7464 fc2 s4 VN.t1269 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7465 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7466 fc2 s4 VN.t1268 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7467 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7468 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7469 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7470 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7471 VN.t1267 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7472 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7473 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7474 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7475 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7476 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7477 VN.t1266 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7478 VN.t1265 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7479 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7480 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7481 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7482 VN.t1264 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7483 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7484 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7485 fc2 s4 VN.t1263 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7486 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7487 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7488 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7489 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7490 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7491 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7492 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7493 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7494 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7495 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7496 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7497 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7498 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7499 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7500 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7502 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7503 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7504 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7505 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7506 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7507 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7508 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7509 fc2 s4 VN.t1262 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7510 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7511 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7512 VN.t1261 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7513 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7514 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7515 VN.t1260 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7516 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7517 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7518 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7519 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7520 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7521 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7522 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7523 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7524 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7525 fc2 s4 VN.t1259 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7526 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7527 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7528 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7529 VN.t1258 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7530 fc2 s4 VN.t1257 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7531 VN.t1256 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X7532 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7533 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7534 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7535 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7536 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7537 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7538 fc2 s4 VN.t1255 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7539 VN.t1254 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7540 VN.t1253 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7541 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7542 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7543 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7544 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7545 fc2 s4 VN.t1252 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7546 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7547 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7548 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7549 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7550 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7551 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7552 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7553 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7554 fc2 s4 VN.t1251 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7555 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7556 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7557 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7558 VN.t1250 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7559 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7560 VN.t1249 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7561 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7562 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7563 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7564 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7565 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7566 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7567 fc2 s4 VN.t1248 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7568 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7569 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7570 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7571 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7572 fc2 s4 VN.t1247 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7573 VN.t1246 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7574 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7575 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7576 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7577 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7578 VN.t1245 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7579 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7580 VN.t1244 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7581 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7582 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7583 fc2 s4 VN.t1243 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7584 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7585 VN.t1242 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7586 VN.t1241 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7587 fc2 s4 VN.t1240 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7588 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7589 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7590 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7591 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7592 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7593 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7594 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7595 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7596 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7597 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7598 fc2 s4 VN.t1239 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7599 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7600 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7601 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7602 VN.t1238 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7603 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7604 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7605 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7606 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7607 fc2 s4 VN.t1237 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7608 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7609 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7610 VN.t1236 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7611 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7612 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7613 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7614 VN.t1235 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7615 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7616 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7618 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7619 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7620 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7621 VN.t1234 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7622 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7623 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7624 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7625 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7626 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7627 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7628 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7629 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7630 fc2 s4 VN.t1233 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7631 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7632 VN.t1232 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7633 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7634 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7635 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7636 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7637 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7638 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7639 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7640 VN.t1231 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7641 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7643 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7644 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7645 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7646 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7647 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7648 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7649 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7650 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7651 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7652 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7653 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7654 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7655 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7656 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7657 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7658 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7659 VN.t1230 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7660 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7661 VN.t1229 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7662 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7663 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7664 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7665 fc2 s4 VN.t1228 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7666 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7667 VN.t1227 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7668 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7669 VN.t1226 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7670 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7671 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7672 fc2 s4 VN.t1225 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7673 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7674 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7675 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7676 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7677 VN.t1224 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7678 VN.t1223 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7679 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7680 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7681 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7682 fc2 s4 VN.t1222 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7683 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7684 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7685 fc2 s4 VN.t1221 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7686 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7687 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7688 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7689 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7690 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7691 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7692 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7693 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7694 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7695 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7696 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7697 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7698 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7699 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7700 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7701 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7702 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7703 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7704 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7705 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7706 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7707 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7708 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7709 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7710 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7711 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7712 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7713 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7714 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7715 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7716 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7717 fc2 s4 VN.t1220 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7718 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7719 VN.t1219 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7720 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7721 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7722 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7723 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7724 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7725 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7726 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7727 fc2 s4 VN.t1218 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7728 VN.t1217 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7729 VN.t1216 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7730 VN.t1215 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7731 VN.t1214 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7732 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7733 fc2 s4 VN.t1213 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7734 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7735 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7736 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7737 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7738 fc2 s4 VN.t1212 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7739 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7740 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7741 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7742 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7743 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7744 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7745 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7746 fc2 s4 VN.t1211 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7747 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7748 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7749 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7750 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7751 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7752 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7753 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7754 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7755 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7756 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7757 fc2 s4 VN.t1210 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7758 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7759 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7760 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7761 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7762 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7763 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7764 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7765 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7766 VN.t1209 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7767 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7768 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7769 VN.t1208 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7770 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7771 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7772 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7773 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7774 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7775 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7776 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7777 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7778 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7779 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7780 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7781 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7782 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7783 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7784 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7785 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7786 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7787 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7788 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7789 VN.t1207 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7790 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7791 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7792 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7793 fc2 s4 VN.t1206 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7794 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7795 fc2 s4 VN.t1205 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7796 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7797 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7798 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7799 VN.t1204 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7800 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7801 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7802 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7803 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7804 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7805 fc2 s4 VN.t1203 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7806 VN.t1202 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7807 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7808 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7809 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7810 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7811 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7812 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7813 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7814 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7815 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7816 fc2 s4 VN.t1201 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7817 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7818 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7819 fc2 s4 VN.t1200 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7820 VN.t1199 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7821 VN.t1198 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7822 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X7823 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7824 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7825 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7826 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7827 fc2 s4 VN.t1197 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7828 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7829 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7830 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7831 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7832 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7833 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7834 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7835 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7836 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7837 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7838 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7839 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7840 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7841 VN.t1196 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7842 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7843 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7844 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7845 fc2 s4 VN.t1195 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7846 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7847 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7848 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7849 fc2 s4 VN.t1194 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7850 VN.t1193 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7851 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7852 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7853 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7854 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7855 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7856 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7857 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7858 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7859 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7860 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7861 fc2 s4 VN.t1192 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7862 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7863 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7864 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7865 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7866 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7867 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7868 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7869 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7870 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7871 VN.t1191 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7872 VN.t1190 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7873 fc2 s4 VN.t1189 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7874 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7875 fc2 s4 VN.t1188 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7876 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7877 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7878 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7879 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7880 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7881 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7882 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7883 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7884 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7885 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7886 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X7887 fc2 s4 VN.t1187 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7888 VN.t1186 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7889 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7890 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7891 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7892 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7893 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7894 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7895 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7896 VN.t1185 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7897 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7898 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7899 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7900 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7901 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7902 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7903 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7904 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7905 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7906 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7907 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7908 fc2 s4 VN.t1184 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7909 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7910 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7911 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7912 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7913 VN.t1183 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7914 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7915 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7916 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7917 fc2 s4 VN.t1182 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7918 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7919 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7920 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7921 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7922 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7923 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X7924 VN.t1181 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7925 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7926 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7927 VN.t1180 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7929 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7930 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7931 VN.t1179 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7932 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7933 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7934 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7935 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7936 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X7937 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7938 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X7939 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7940 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7941 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7942 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7943 VN.t1178 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7944 fc2 s4 VN.t1177 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7945 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7946 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7947 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7948 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7949 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7950 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7951 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7952 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7953 VN.t1176 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7954 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7955 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X7956 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7957 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7958 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7959 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7960 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7961 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7962 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7963 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7964 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7965 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7966 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7967 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7968 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7969 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7970 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X7971 VN.t1175 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7972 VN.t1174 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7973 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7974 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7975 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7976 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7977 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7978 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7979 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7980 fc2 s4 VN.t1173 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7981 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7982 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7983 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7984 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7985 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7986 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7987 fc2 s4 VN.t1172 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7988 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7989 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7990 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7991 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7992 VN.t1171 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7993 VN.t1170 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7994 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7995 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X7996 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X7997 VN.t1169 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X7998 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7999 VN.t1168 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8000 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8001 fc2 s4 VN.t1167 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8002 fc2 s4 VN.t1166 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8003 VN.t1165 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8004 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8005 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8006 fc2 s4 VN.t1164 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8007 fc2 s4 VN.t1163 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8009 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8010 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8011 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8012 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8013 VN.t1162 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8014 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8015 fc2 s4 VN.t1161 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8016 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8017 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8018 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8019 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8020 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8021 VN.t1160 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8022 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8023 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8024 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8025 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8026 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8027 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8028 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8029 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8030 fc2 s4 VN.t1159 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8031 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8032 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8033 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8034 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8035 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8036 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8037 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8038 VN.t1158 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8039 fc2 s4 VN.t1157 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8040 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8041 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8042 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8043 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8044 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8045 VN.t1156 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8046 VN.t1155 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8047 fc2 s4 VN.t1154 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8048 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8049 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8050 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8051 VN.t1153 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8052 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8053 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8054 fc2 s4 VN.t1152 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8055 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8056 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8057 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8058 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8059 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8060 VN.t1151 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8061 VN.t1150 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8062 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8063 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8064 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8065 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8066 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8068 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8069 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8070 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8071 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8072 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8073 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8074 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8075 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8076 VN.t1149 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8077 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8078 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8079 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8080 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8081 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8082 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8083 VN.t1148 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8084 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8085 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8086 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8088 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8089 fc2 s4 VN.t1147 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8090 fc2 s4 VN.t1146 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8091 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8092 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8093 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8094 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8095 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8096 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8097 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8098 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8099 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8100 VN.t1145 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8101 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8102 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8103 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8104 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8105 fc2 s4 VN.t1144 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8106 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8107 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8108 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8109 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8110 VN.t1143 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8111 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8112 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8113 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8114 fc2 s4 VN.t1142 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8115 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8116 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8117 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8119 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8120 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8121 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8122 fc2 s4 VN.t1141 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8123 fc2 s4 VN.t1140 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8124 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8125 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8126 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8127 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8128 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8129 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8130 fc2 s4 VN.t1139 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8131 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8132 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8133 VN.t1138 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8134 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8136 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8137 VN.t1137 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8138 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8139 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8140 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8141 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8142 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8143 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8144 fc2 s4 VN.t1136 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8145 VN.t1135 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8146 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8147 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8148 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8149 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8150 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8151 VN.t1134 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8152 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8153 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8154 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8155 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8156 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8157 fc2 s4 VN.t1133 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8158 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8159 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8160 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8161 fc2 s4 VN.t1132 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8162 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8163 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8164 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8165 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8166 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8167 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8168 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8169 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8170 fc2 s4 VN.t1131 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8171 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8172 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8173 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8174 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8175 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8176 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8177 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8178 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8179 fc2 s4 VN.t1130 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8180 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8181 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8182 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8183 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8184 fc2 s4 VN.t1129 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8185 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8186 fc2 s4 VN.t1128 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8187 VN.t1127 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8188 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8189 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8190 fc2 s4 VN.t1126 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8191 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8192 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8193 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8194 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8195 VN.t1125 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8196 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8198 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8199 VN.t1124 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8200 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8201 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8202 fc2 s4 VN.t1123 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8203 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8205 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8206 fc2 s4 VN.t1122 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8208 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8209 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8210 fc2 s4 VN.t1121 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8211 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8212 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8213 VN.t1120 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8214 fc2 s4 VN.t1119 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8215 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8216 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8217 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8218 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8219 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8220 VN.t1118 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8221 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8222 VN.t1117 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8223 fc2 s4 VN.t1116 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8224 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8225 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8226 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8227 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8228 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8229 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8230 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8231 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8232 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8234 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8235 VN.t1115 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8236 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8237 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8238 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8239 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8240 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8241 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8242 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8243 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8244 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8245 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8246 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8247 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8248 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8249 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8250 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8251 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8252 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8253 VN.t1114 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8254 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8255 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8256 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8257 VN.t1113 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8258 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8259 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8260 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8261 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8262 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8263 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8264 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8265 fc2 s4 VN.t1112 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8266 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8267 fc2 s4 VN.t1111 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8268 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8269 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8270 fc2 s4 VN.t1110 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8271 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8272 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8273 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8274 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8275 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8276 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8277 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8278 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8279 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8280 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8281 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8282 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8283 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8284 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8285 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8286 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8287 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8288 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8289 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8290 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8291 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8292 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8293 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8295 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8296 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8297 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8298 fc2 s4 VN.t1109 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8299 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8300 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8301 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8302 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8303 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8304 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8305 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8306 fc2 s4 VN.t1108 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8307 fc2 s4 VN.t1107 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8308 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8309 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8310 VN.t1106 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8311 VN.t1105 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8312 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8313 VN.t1104 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8314 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8315 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8316 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8317 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8318 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8319 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8320 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8321 fc2 s4 VN.t1103 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8322 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8323 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8324 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8325 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8326 fc2 s4 VN.t1102 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8327 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8328 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8329 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8330 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8331 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8332 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8333 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8334 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8335 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8336 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8337 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8339 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8340 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8341 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8342 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8343 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8344 fc2 s4 VN.t1101 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8345 fc2 s4 VN.t1100 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8346 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8347 fc2 s4 VN.t1099 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8348 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8349 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8350 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8351 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8352 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8353 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8354 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8355 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8356 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8357 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8358 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8359 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8360 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8361 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8362 VN.t1098 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8363 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8364 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8365 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8366 VN.t1097 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8367 fc2 s4 VN.t1096 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8368 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8369 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8370 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8372 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8373 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8374 fc2 s4 VN.t1095 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8375 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8376 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8377 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8378 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8379 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8380 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8381 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8382 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8383 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8384 fc2 s4 VN.t1094 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8385 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8386 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8387 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8388 fc2 s4 VN.t1093 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8389 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8390 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8391 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8392 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8393 VN.t1092 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8394 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8395 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8396 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8397 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8398 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8399 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8400 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8401 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8402 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8403 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8404 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8405 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8406 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8407 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8408 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8409 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8410 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8411 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8412 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8413 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8414 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8415 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8416 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8417 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8418 fc2 s4 VN.t1091 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8419 fc2 s4 VN.t1090 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8420 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8421 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8422 VN.t1089 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8423 fc2 s4 VN.t1088 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8424 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8425 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8426 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8427 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8428 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8429 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8430 fc2 s4 VN.t1087 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8431 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8432 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8433 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8434 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8435 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8436 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8437 fc2 s4 VN.t1086 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8438 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8439 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8440 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8441 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8442 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8443 fc2 s4 VN.t1085 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8444 VN.t1084 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8445 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8446 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8447 fc2 s4 VN.t1083 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8448 fc2 s4 VN.t1082 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8449 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8450 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8451 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8452 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8453 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8454 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8455 VN.t1081 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8456 VN.t1080 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8457 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8458 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8459 VN.t1079 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8460 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8461 fc2 s4 VN.t1078 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8462 fc2 s4 VN.t1077 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8463 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8464 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8465 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8466 fc2 s4 VN.t1076 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8467 fc2 s4 VN.t1075 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8468 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8469 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8470 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8471 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8472 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8473 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8474 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8475 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8476 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8477 fc2 s4 VN.t1074 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8478 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8479 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8480 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8481 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8482 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8483 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8484 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8485 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8486 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8487 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8488 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8489 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8490 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8491 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8492 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8493 fc2 s4 VN.t1073 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8494 fc2 s4 VN.t1072 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8495 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8496 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8497 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8498 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8499 fc2 s4 VN.t1071 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8500 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8502 VN.t1070 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8503 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8504 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8505 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8506 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8507 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8508 fc2 s4 VN.t1069 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8509 VN.t1068 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8510 fc2 s4 VN.t1067 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8511 fc2 s4 VN.t1066 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8512 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8513 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8514 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8515 VN.t1065 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8516 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8517 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8518 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8519 fc2 s4 VN.t1064 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8520 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8521 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8522 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8523 VN.t1063 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8524 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8525 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8526 VN.t1062 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8527 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8528 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8529 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8530 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8531 fc2 s4 VN.t1061 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8532 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8533 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8534 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8535 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8536 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8537 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8538 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8539 fc2 s4 VN.t1060 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8540 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8541 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8542 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8543 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8544 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8545 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8546 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8547 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8548 fc2 s4 VN.t1059 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8549 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8550 VN.t1058 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8551 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8552 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8553 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8554 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8555 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8556 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8557 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8558 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8559 VN.t1057 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8560 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8561 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8562 fc2 s4 VN.t1056 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8563 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8564 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8565 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8566 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8567 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8568 VN.t1055 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8569 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8570 VN.t1054 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8571 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8572 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8573 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8574 fc2 s4 VN.t1053 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8575 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8576 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8577 VN.t1052 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8578 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8579 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8580 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8581 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8582 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8583 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8584 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8585 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8586 fc2 s4 VN.t1051 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8587 fc2 s4 VN.t1050 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8588 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8589 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8590 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8591 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8592 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8593 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8594 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8595 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8596 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8597 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8598 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8599 VN.t1049 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8600 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8601 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8602 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8603 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8604 fc2 s4 VN.t1048 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8605 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8606 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8607 VN.t1047 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8608 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8609 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8610 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8611 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8612 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8613 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8614 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8615 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X8616 VN.t1046 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8617 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8618 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8619 fc2 s4 VN.t1045 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8620 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8621 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8622 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8623 fc2 s4 VN.t1044 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8624 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8625 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8626 VN.t1043 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8627 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8628 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8629 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8630 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8631 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8632 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8633 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8634 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8635 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8636 VN.t1042 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8637 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8638 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8639 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8640 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8641 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8642 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8643 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8644 VN.t1041 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8645 fc2 s4 VN.t1040 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8646 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8647 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8648 fc2 s4 VN.t1039 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8649 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8650 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8651 VN.t1038 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8652 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8653 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8654 fc2 s4 VN.t1037 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8655 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8656 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8657 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8658 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8659 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8660 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8661 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8662 fc2 s4 VN.t1036 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8663 fc2 s4 VN.t1035 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8664 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8665 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8666 fc2 s4 VN.t1034 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8667 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8668 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8669 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8670 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8671 fc2 s4 VN.t1033 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8672 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8673 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8674 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8675 VN.t1032 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8676 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8677 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8678 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8679 fc2 s4 VN.t1031 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8680 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8681 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8682 VN.t1030 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8683 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8684 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8685 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8686 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8687 fc2 s4 VN.t1029 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8688 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8689 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8690 VN.t1028 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8691 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8692 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8693 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8694 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8695 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8696 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8697 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8698 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8699 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8700 VN.t1027 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8701 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8702 fc2 s4 VN.t1026 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8703 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8704 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8705 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8706 VN.t1025 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8707 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8708 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8709 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8710 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8711 VN.t1024 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8712 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8713 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8714 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8715 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8716 fc2 s4 VN.t1023 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8717 fc2 s4 VN.t1022 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8718 fc2 s4 VN.t1021 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8719 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8720 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8721 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8722 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8723 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8724 VN.t1020 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8725 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8726 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8727 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8728 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8729 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8730 VN.t1019 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8731 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8732 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8733 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8734 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8735 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8736 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8737 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8738 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8739 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8740 fc2 s4 VN.t1018 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8741 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8742 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8743 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8744 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8745 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8746 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8747 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8748 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8749 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8750 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8751 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8752 fc2 s4 VN.t1017 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8753 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8754 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8755 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8756 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8757 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8758 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8760 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8761 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8762 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8763 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8764 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8765 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X8766 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8767 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8768 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8769 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8770 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8771 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8772 VN.t1016 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8773 fc2 s4 VN.t1015 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8774 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8775 VN.t1014 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8776 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8777 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8778 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8779 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8780 fc2 s4 VN.t1013 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8781 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8782 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8783 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8784 fc2 s4 VN.t1012 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8785 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8786 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8787 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8788 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8789 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8790 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8791 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8792 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8793 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8794 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8795 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8796 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8797 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8798 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8799 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8800 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8801 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8802 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8803 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8804 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8805 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8806 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8807 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8808 fc2 s4 VN.t1011 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8809 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8810 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8811 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8812 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8813 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8814 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8815 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8816 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8817 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8818 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8819 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8820 VN.t1010 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8821 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8822 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8823 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8824 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8825 fc2 s4 VN.t1009 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8826 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8827 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8828 VN.t1008 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8829 fc2 s4 VN.t1007 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8830 fc2 s4 VN.t1006 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8831 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8832 VN.t1005 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8833 fc2 s4 VN.t1004 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8834 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8835 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8836 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8837 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8838 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8839 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8840 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8841 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8842 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8844 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8845 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8846 fc2 s4 VN.t1003 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8847 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8848 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8849 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8850 fc2 s4 VN.t1002 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8851 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8852 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8853 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8854 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8855 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8856 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8857 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8858 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8859 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8860 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8861 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8862 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8863 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8864 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8865 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8866 fc2 s4 VN.t1001 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8867 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8868 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8869 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8870 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8871 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8872 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8873 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8874 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8875 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8876 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8877 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8878 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8879 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8880 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8881 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8882 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8883 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8884 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8886 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8887 fc2 s4 VN.t1000 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8888 fc2 s4 VN.t999 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8889 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8890 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X8891 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8892 VN.t998 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8893 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8894 VN.t997 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8895 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8896 VN.t996 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8897 fc2 s4 VN.t995 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8898 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8899 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8900 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8901 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8902 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8904 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8905 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8906 fc2 s4 VN.t994 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8907 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8908 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8909 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8910 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8911 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8912 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8913 fc2 s4 VN.t993 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8914 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8915 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8916 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8917 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8918 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8919 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8920 fc2 s4 VN.t992 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8921 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8922 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8923 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8924 fc2 s4 VN.t991 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8925 VN.t990 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8926 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8927 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8929 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8930 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8931 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8932 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8933 VN.t989 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8934 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8935 VN.t988 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8936 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8937 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8938 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8939 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8940 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8941 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8942 VN.t987 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8943 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8944 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8945 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8946 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8947 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8948 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8949 fc2 s4 VN.t986 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8950 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8951 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8952 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8953 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8954 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8955 fc2 s4 VN.t985 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8956 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8957 VN.t984 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8958 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8959 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8960 VN.t983 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X8961 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X8962 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8963 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8964 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8965 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8966 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8967 VN.t982 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8968 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8969 fc2 s4 VN.t981 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8970 fc2 s4 VN.t980 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8971 VN.t979 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8972 VN.t978 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8973 VN.t977 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8974 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8975 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8976 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8977 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8978 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8980 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8981 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8982 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8983 fc2 s4 VN.t976 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8984 VN.t975 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8985 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8986 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8987 VN.t974 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X8988 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8989 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8990 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8991 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8992 fc2 s4 VN.t973 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8993 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8994 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X8995 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8996 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X8998 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8999 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9000 VN.t972 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9001 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9002 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9003 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9004 fc2 s4 VN.t971 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9005 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9007 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9008 VN.t970 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9009 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9010 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9011 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9012 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9013 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9014 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9015 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9017 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9019 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9020 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9021 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9022 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9023 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9024 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9025 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9026 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9027 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9028 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9029 VN.t969 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9030 VN.t968 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9031 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9032 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9033 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9034 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9035 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9036 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9037 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9038 VN.t967 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9039 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9040 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9041 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9042 fc2 s4 VN.t966 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9043 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9044 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9045 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9046 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9047 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9048 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9049 fc2 s4 VN.t965 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9050 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9051 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9052 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9053 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9054 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9055 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9056 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9057 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9058 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9059 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9060 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9061 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9062 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9063 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9064 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9065 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9066 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9067 fc2 s4 VN.t964 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9068 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9069 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9070 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9071 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9072 VN.t963 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9073 fc2 s4 VN.t962 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9074 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9075 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9076 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9077 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9078 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9079 VN.t961 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9080 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9081 VN.t960 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9082 VN.t959 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9083 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9084 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9085 fc2 s4 VN.t958 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9086 fc2 s4 VN.t957 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9087 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9088 fc2 s4 VN.t956 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9089 fc2 s4 VN.t955 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9090 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9091 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9092 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9093 VN.t954 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9094 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9095 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9096 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9097 VN.t953 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9098 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9099 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9100 VN.t952 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9101 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9102 fc2 s4 VN.t951 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9103 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9104 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9105 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9106 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9107 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9108 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9109 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9111 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9112 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9113 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9114 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9115 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9116 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9117 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9119 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9120 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9121 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9122 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9123 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9124 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9125 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9126 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9127 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9128 fc2 s4 VN.t950 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9129 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9130 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9131 VN.t949 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9132 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9133 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9134 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9135 VN.t948 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9136 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9137 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9138 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9139 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9140 VN.t947 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9141 fc2 s4 VN.t946 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9142 VN.t945 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9143 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9144 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9145 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9146 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9147 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9148 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9149 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9150 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9151 fc2 s4 VN.t944 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9152 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9153 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9154 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9155 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9156 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9157 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9158 VN.t943 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9159 fc2 s4 VN.t942 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9160 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9161 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9162 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9163 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9164 VN.t941 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9165 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9166 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9167 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9168 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9169 fc2 s4 VN.t940 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9170 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9171 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9172 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9173 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9174 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9175 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9176 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9177 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9178 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9179 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9180 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9181 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9182 fc2 s4 VN.t939 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9183 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9184 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9185 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9186 VN.t938 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9187 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9188 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9189 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9190 VN.t937 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9191 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9192 fc2 s4 VN.t936 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9193 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9194 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9195 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9196 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9197 fc2 s4 VN.t935 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9198 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9199 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9200 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9201 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9202 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9203 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9204 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9205 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9206 fc2 s4 VN.t934 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9207 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9208 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9209 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9210 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9211 VN.t933 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9212 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9213 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9214 fc2 s4 VN.t932 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9215 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9216 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9217 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9218 VN.t931 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9219 VN.t930 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9220 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9221 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9222 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9223 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9224 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9225 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9226 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9227 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9228 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9229 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9230 VN.t929 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9231 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9232 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9234 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9235 VN.t928 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9236 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9237 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9238 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9239 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9240 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9241 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9242 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9243 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9244 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9245 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9246 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9247 VN.t927 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9248 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9249 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9250 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9251 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9252 VN.t926 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9253 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9254 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9255 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9256 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9257 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9258 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9260 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9261 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9262 fc2 s4 VN.t925 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9263 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9264 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9265 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9266 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9267 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9268 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9269 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9270 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9271 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9272 fc2 s4 VN.t924 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9273 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9274 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9275 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9276 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9277 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9278 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9279 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9280 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9281 VN.t923 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9282 VN.t922 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9283 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9284 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9285 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9286 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9287 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9288 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9289 VN.t921 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9290 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9291 fc2 s4 VN.t920 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9292 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9293 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9295 VN.t919 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9296 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9297 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9298 VN.t918 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9299 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9300 VN.t917 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9301 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9302 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9303 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9304 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9305 fc2 s4 VN.t916 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9306 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9307 fc2 s4 VN.t915 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9308 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9309 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9310 VN.t914 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9311 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9312 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9313 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9314 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9315 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9316 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9317 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9318 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9319 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9320 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9321 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9322 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9323 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9324 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9325 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9326 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9327 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9328 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9329 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9330 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9331 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9332 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9333 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9334 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9335 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9336 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9337 fc2 s4 VN.t913 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9338 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9339 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9340 VN.t912 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9341 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9342 VN.t911 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9343 fc2 s4 VN.t910 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9344 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9345 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9346 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9347 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9348 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9349 fc2 s4 VN.t909 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9350 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9351 VN.t908 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9352 VN.t907 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9353 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9354 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9355 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9356 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9357 fc2 s4 VN.t906 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9358 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9359 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9360 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9361 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9362 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9363 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9364 fc2 s4 VN.t905 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9365 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9366 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9367 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9368 VN.t904 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9369 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9370 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9371 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9372 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9373 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9374 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9375 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9376 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9377 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9378 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9379 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9380 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9381 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9382 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9383 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9384 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9385 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9386 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9387 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9388 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9389 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9390 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9391 VN.t903 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9392 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9393 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9394 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9395 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9396 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9397 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9398 VN.t902 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9399 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9400 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9401 VN.t901 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9402 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9403 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9404 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9405 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9406 VN.t900 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9407 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9408 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9409 fc2 s4 VN.t899 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9410 fc2 s4 VN.t898 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9411 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9412 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9413 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9414 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9415 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9416 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9417 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9418 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9419 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9420 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9421 VN.t897 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9422 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9423 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9424 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9425 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9426 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9427 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9428 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9429 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9430 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9431 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9432 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9433 fc2 s4 VN.t896 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9434 VN.t895 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9435 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9436 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9437 VN.t894 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9438 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9439 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9440 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9441 VN.t893 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9442 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9443 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9444 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9445 fc2 s4 VN.t892 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9446 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9447 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9448 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9449 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9450 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9451 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9452 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9453 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9454 VN.t891 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9455 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9456 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9457 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9458 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9459 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9460 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9461 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9462 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9463 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9464 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9465 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9466 VN.t890 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9467 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9468 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9469 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9470 VN.t889 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9471 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9472 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9473 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9474 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9475 fc2 s4 VN.t888 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9476 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9477 fc2 s4 VN.t887 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9478 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9479 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9480 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9481 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9482 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9483 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9484 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9485 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9486 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9487 VN.t886 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9488 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9489 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9490 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9491 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9492 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9493 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9494 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9495 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9496 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9497 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9498 VN.t885 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9499 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9500 fc2 s4 VN.t884 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9501 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9502 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9503 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9504 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9505 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9506 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9507 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9508 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9509 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9510 VN.t883 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9511 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9512 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9513 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9514 fc2 s4 VN.t882 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9515 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9516 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9517 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9518 VN.t881 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9519 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9520 VN.t880 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9521 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9522 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9523 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9524 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9525 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9526 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9527 fc2 s4 VN.t879 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9528 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9529 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9530 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9531 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9532 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9533 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9534 fc2 s4 VN.t878 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9535 VN.t877 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9536 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9537 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9538 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9539 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9540 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9541 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9542 VN.t876 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9543 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9544 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9545 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9546 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9547 VN.t875 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9548 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9549 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9550 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9551 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9552 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9553 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9554 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9555 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9556 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9557 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9558 VN.t874 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9559 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9560 fc2 s4 VN.t873 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9561 fc2 s4 VN.t872 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9562 VN.t871 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9563 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9564 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9565 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9566 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9567 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9568 VN.t870 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9569 VN.t869 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9570 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9571 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9572 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9573 VN.t868 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9574 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9575 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9576 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9577 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9578 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9579 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9580 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9581 VN.t867 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9582 VN.t866 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9583 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9584 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9585 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9586 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9587 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9588 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9589 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9590 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9591 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9592 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9593 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9594 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9595 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9596 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9597 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9598 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9599 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9600 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9601 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9602 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9603 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9604 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9605 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9606 VN.t865 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9607 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9608 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9609 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9610 fc2 s4 VN.t864 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9611 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9612 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9613 VN.t863 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9614 VN.t862 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9615 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9616 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9617 VN.t861 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9618 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9619 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9620 fc2 s4 VN.t860 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9622 fc2 s4 VN.t859 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9623 fc2 s4 VN.t858 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9624 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9625 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9626 VN.t857 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9627 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9628 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9629 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9630 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9631 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9632 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9633 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9634 fc2 s4 VN.t856 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9635 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9636 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9637 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9638 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9639 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9640 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9641 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9643 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9644 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9645 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9646 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9647 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9648 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9649 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9650 VN.t855 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9651 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9652 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9653 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9654 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9655 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9656 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9657 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9658 VN.t854 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9659 fc2 s4 VN.t853 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9660 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9661 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9662 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9663 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9664 fc2 s4 VN.t852 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9665 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9666 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9667 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9668 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9669 VN.t851 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9670 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9671 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9672 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9673 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9674 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9675 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9676 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9677 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9678 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9679 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9680 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9681 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9682 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9683 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9684 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9685 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9686 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9687 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9688 VN.t850 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9689 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9690 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9691 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9692 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9693 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9694 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9695 fc2 s4 VN.t849 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9696 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9697 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9698 fc2 s4 VN.t848 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9699 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9700 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9701 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9702 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9703 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9704 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9705 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9706 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9707 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9708 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9709 VN.t847 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9710 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9711 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9712 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9713 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9714 fc2 s4 VN.t846 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9715 fc2 s4 VN.t845 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9716 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9717 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9718 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9719 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9720 VN.t844 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9721 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9722 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9723 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9724 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9725 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9726 fc2 s4 VN.t843 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9727 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9728 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9729 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9730 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9731 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9732 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9733 fc2 s4 VN.t842 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9734 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9735 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9736 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9737 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9738 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9739 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9740 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9741 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9742 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9743 VN.t841 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9744 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9745 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9746 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9747 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9748 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9749 fc2 s4 VN.t840 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9750 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9751 VN.t839 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9752 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9753 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9754 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9755 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9756 VN.t838 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9757 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9758 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9759 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9760 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9761 fc2 s4 VN.t837 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9762 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9763 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9764 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9765 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9766 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9767 fc2 s4 VN.t836 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9768 VN.t835 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9769 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9770 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9771 fc2 s4 VN.t834 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9772 fc2 s4 VN.t833 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9773 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9774 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9775 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9776 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9777 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9778 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9779 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9780 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9781 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9782 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9783 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9784 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9785 fc2 s4 VN.t832 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9786 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9787 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9788 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9789 VN.t831 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9790 fc2 s4 VN.t830 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9791 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9792 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9793 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9794 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9795 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9796 VN.t829 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9797 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9798 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9799 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9800 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9801 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9802 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9803 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9804 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9805 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9806 fc2 s4 VN.t828 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9807 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9808 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9809 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9810 VN.t827 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9811 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9812 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9813 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9814 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9815 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9816 VN.t826 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9817 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9818 VN.t825 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9819 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9820 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9821 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9822 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9823 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9824 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9825 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9826 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9827 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9828 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9829 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9830 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9831 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9832 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9833 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9834 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9835 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9836 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9837 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9838 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9839 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9840 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9841 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9842 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9843 VN.t824 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9844 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9845 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9846 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9847 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9848 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9849 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9850 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9851 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9852 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9853 fc2 s4 VN.t823 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9854 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9855 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9856 fc2 s4 VN.t822 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9857 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9858 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9859 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9860 fc2 s4 VN.t821 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9861 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9862 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9863 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9864 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9865 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9866 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9867 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9868 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9869 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9870 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9871 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9872 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9873 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9874 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9875 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9876 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9877 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9878 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9879 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9880 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9881 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9882 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9883 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9884 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9885 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9886 fc2 s4 VN.t820 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9887 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9888 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9889 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9890 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9891 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9892 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9893 VN.t819 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9894 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9895 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9896 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9897 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9898 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9899 fc2 s4 VN.t818 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9900 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9901 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9902 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9903 fc2 s4 VN.t817 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9904 VN.t816 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9905 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9906 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9907 VN.t815 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9908 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9909 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9910 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9911 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9912 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9913 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9914 fc2 s4 VN.t814 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9915 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9916 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9917 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9918 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9919 VN.t813 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9920 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9921 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9922 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9923 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9924 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9925 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9926 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9927 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9928 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9929 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9930 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9931 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9932 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9933 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9934 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X9935 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9936 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9937 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9938 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9939 fc2 s4 VN.t812 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9940 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9941 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9942 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9943 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9944 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9945 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9946 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9947 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9948 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9949 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9950 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X9951 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9952 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9953 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9954 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9955 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9956 VN.t811 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9957 VN.t810 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9958 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9959 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9960 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9961 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X9962 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9963 VN.t809 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9964 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9965 fc2 s4 VN.t808 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9966 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9967 fc2 s4 VN.t807 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9968 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9969 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9970 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9971 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9972 fc2 s4 VN.t806 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9973 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9974 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9975 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9976 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9977 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9978 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9979 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9980 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9981 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9982 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9983 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9984 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9985 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9986 VN.t805 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9987 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9988 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9989 fc2 s4 VN.t804 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X9990 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9991 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9992 fc2 s4 VN.t803 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X9993 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9994 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9995 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9996 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X9998 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9999 fc2 s4 VN.t802 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10000 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10001 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10002 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10003 VN.t801 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10004 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10005 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10006 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10007 fc2 s4 VN.t800 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10008 fc2 s4 VN.t799 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10009 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10010 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10011 VN.t798 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10012 fc2 s4 VN.t797 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10013 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10014 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10015 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10016 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10017 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10019 fc2 s4 VN.t796 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10020 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10021 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10022 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10023 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10024 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10025 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10026 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10027 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10028 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10029 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10030 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10031 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10032 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10033 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10034 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10035 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10036 fc2 s4 VN.t795 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10037 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10038 VN.t794 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10039 VN.t793 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10040 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10041 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10042 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10043 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10044 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10045 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10046 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10047 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10048 fc2 s4 VN.t792 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10049 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10050 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10051 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10052 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10053 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10054 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10055 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10056 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10057 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10058 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10059 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10060 fc2 s4 VN.t791 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10061 fc2 s4 VN.t790 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10062 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10063 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10064 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10065 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10066 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10068 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10069 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10070 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10071 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10072 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10073 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10074 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10075 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10076 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10077 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10078 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10079 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X10080 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10081 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10082 fc2 s4 VN.t789 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10083 VN.t788 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10084 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10085 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10086 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10087 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10088 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10089 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10090 VN.t787 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10091 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10092 fc2 s4 VN.t786 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10093 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10094 VN.t785 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10095 fc2 s4 VN.t784 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10096 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10097 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10098 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10099 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10100 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10101 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10102 VN.t783 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10103 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10104 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10105 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10106 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10107 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10108 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10109 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10110 fc2 s4 VN.t782 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10111 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10112 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10113 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10114 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10115 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10116 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10117 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10119 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10120 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10121 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10122 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10123 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10124 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10125 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10126 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10127 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10128 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10129 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10130 fc2 s4 VN.t781 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10131 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10132 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10133 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10134 fc2 s4 VN.t780 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10135 VN.t779 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10136 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10137 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10138 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10139 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10140 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10141 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10142 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10143 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10144 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10145 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10146 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10147 fc2 s4 VN.t778 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10148 fc2 s4 VN.t777 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10149 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10150 VN.t776 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10151 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10152 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10153 VN.t775 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10154 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10156 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10157 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10158 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10159 VN.t774 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10160 fc2 s4 VN.t773 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10161 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10162 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10163 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10164 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10165 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10166 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10167 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10168 fc2 s4 VN.t772 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10169 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10170 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10171 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10172 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10173 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10174 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10175 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10176 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10177 fc2 s4 VN.t771 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10178 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10179 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10180 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10181 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10182 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10183 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10184 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10185 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10186 VN.t770 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10187 fc2 s4 VN.t769 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10188 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10189 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10190 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10191 VN.t768 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10192 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10193 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10194 VN.t767 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10195 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10196 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10198 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10199 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10200 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10201 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10202 fc2 s4 VN.t766 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10203 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10204 fc2 s4 VN.t765 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10205 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10206 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10207 fc2 s4 VN.t764 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10208 VN.t763 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10209 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10210 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10211 VN.t762 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10212 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10213 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10214 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10215 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10216 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10217 fc2 s4 VN.t761 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10218 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10219 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10220 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10221 VN.t760 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10222 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10223 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10224 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10225 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10226 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10227 fc2 s4 VN.t759 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10228 fc2 s4 VN.t758 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10229 VN.t757 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10230 VN.t756 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10231 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10232 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10233 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10234 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10235 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10236 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10237 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10238 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10239 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10240 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10241 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10242 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10243 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10244 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10245 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10246 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10247 VN.t755 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10248 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10249 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10250 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10251 fc2 s4 VN.t754 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10252 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10253 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10254 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10255 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10256 VN.t753 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10257 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10258 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10260 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10261 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10262 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10263 VN.t752 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10264 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10265 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10266 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10267 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10268 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10269 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10270 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10271 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10272 VN.t751 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10273 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10274 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10275 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10276 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10277 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10278 VN.t750 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10279 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10280 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10281 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10282 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10283 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10284 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10285 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10286 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10287 fc2 s4 VN.t749 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10288 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10290 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10291 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10292 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10293 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10295 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10296 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10297 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10298 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10299 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10300 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10301 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10302 VN.t748 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10303 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10304 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10305 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10306 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10307 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10308 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10309 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10310 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10311 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10312 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10313 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10314 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10315 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10316 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10317 fc2 s4 VN.t747 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10318 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10319 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10320 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10321 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10322 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10323 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10324 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10325 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10326 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10327 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10328 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10329 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10330 fc2 s4 VN.t746 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10331 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10332 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10333 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10334 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10335 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10336 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10337 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10339 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10340 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10341 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10342 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10343 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10344 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10345 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10346 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10347 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10348 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10349 VN.t745 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10350 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10351 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10352 VN.t744 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10353 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10354 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10355 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10356 fc2 s4 VN.t743 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10357 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10358 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10359 fc2 s4 VN.t742 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10360 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10361 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10362 VN.t741 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10363 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10364 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10365 VN.t740 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10366 fc2 s4 VN.t739 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10367 fc2 s4 VN.t738 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10368 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10369 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10370 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10371 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10372 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10373 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10374 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10375 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10376 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10377 fc2 s4 VN.t737 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10378 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10379 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10380 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10381 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10382 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10383 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10384 fc2 s4 VN.t736 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10385 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10386 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10387 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10388 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10389 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10390 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10391 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10392 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10393 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10394 VN.t735 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10395 fc2 s4 VN.t734 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10396 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10397 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10398 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10399 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10400 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10401 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10402 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10403 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10404 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10405 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10406 VN.t733 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10407 fc2 s4 VN.t732 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10408 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10409 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10410 VN.t731 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10411 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10412 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10413 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10414 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10415 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10416 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10417 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10418 fc2 s4 VN.t730 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10419 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10420 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10421 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10422 fc2 s4 VN.t729 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10423 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10424 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10425 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10426 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10427 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10428 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10429 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10430 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10431 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10432 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10433 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10434 VN.t728 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10435 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10436 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10437 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10438 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10439 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10440 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10441 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10442 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10443 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10444 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10445 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10446 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10447 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10448 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10449 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10450 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10451 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10452 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10453 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10454 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10455 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10456 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10457 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10458 fc2 s4 VN.t727 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10459 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10460 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10461 fc2 s4 VN.t726 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10462 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10463 VN.t725 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10464 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10465 VN.t724 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10466 VN.t723 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10467 fc2 s4 VN.t722 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10468 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10469 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10470 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10471 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10472 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10473 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10474 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10475 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10476 fc2 s4 VN.t721 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10477 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10478 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10479 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10480 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10481 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10482 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10483 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10484 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10485 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10486 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10487 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10488 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10489 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10490 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10491 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10492 fc2 s4 VN.t720 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10493 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10494 VN.t719 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10495 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10496 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10497 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10498 VN.t718 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10499 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10500 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10501 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10502 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10503 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10504 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10505 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10506 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10507 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10508 fc2 s4 VN.t717 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10509 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10510 VN.t716 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10511 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10512 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10513 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10514 VN.t715 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10515 VN.t714 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10516 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10517 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10518 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10519 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10520 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10521 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10522 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10523 VN.t713 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10524 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10525 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10526 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10527 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10528 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10529 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10530 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10531 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10532 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10533 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10534 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10535 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10536 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10537 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10538 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10539 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10540 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10541 fc2 s4 VN.t712 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10542 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10543 VN.t711 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10544 fc2 s4 VN.t710 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10545 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10546 VN.t709 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10547 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10548 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10549 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10550 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10551 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10552 VN.t708 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10553 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10554 VN.t707 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10555 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10556 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10557 VN.t706 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10558 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10559 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10560 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10561 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10562 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10563 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10564 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10565 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10566 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10567 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10568 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10569 fc2 s4 VN.t705 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10570 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10571 VN.t704 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10572 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10573 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10574 fc2 s4 VN.t703 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10575 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10576 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10577 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10578 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10579 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10580 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10582 VN.t702 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10583 VN.t701 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10584 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10585 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10586 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10587 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10588 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10589 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10590 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10591 VN.t700 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10592 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10593 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10594 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10595 VN.t699 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10596 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10597 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10598 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10599 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10600 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10601 fc2 s4 VN.t698 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10602 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10603 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10604 VN.t697 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10605 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10606 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10607 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10608 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10609 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10610 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10611 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10612 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10613 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10614 VN.t696 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10615 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10616 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10617 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10618 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10619 fc2 s4 VN.t695 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10620 VN.t694 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10621 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10622 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10623 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10624 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10625 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10626 VN.t693 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10627 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10628 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10629 fc2 s4 VN.t692 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10630 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10631 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10632 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10633 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10634 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10635 VN.t691 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10636 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10637 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10638 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10639 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10640 fc2 s4 VN.t690 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10641 fc2 s4 VN.t689 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10642 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10643 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10644 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10645 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10646 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10647 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10648 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10649 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10650 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10651 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10652 VN.t688 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10653 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10654 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10655 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10656 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10657 fc2 s4 VN.t687 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10658 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10659 fc2 s4 VN.t686 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10660 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10661 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10662 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10663 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10664 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10665 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10666 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10667 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10668 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10669 VN.t685 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10670 VN.t684 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10671 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10672 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10673 fc2 s4 VN.t683 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10674 fc2 s4 VN.t682 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10675 fc2 s4 VN.t681 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10676 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10677 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10678 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10679 VN.t680 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10680 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10681 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10682 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10683 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10684 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10685 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10686 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10687 VN.t679 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10688 fc2 s4 VN.t678 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10689 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10690 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10691 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10692 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10693 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10694 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10695 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10696 fc2 s4 VN.t677 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10697 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10698 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10699 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10700 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10701 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10702 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10703 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10704 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10705 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10706 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10707 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10708 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10709 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10710 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10711 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10712 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10713 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10714 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10715 fc2 s4 VN.t676 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10716 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10717 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10718 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10719 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10720 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10721 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10722 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10723 VN.t675 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10724 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10725 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10726 fc2 s4 VN.t674 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10727 VN.t673 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10728 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10729 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10730 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10731 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10732 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10733 fc2 s4 VN.t672 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10734 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10735 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10736 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10737 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10738 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10739 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10740 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10741 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10742 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10743 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10744 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10745 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10746 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10747 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10748 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10749 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10750 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10751 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10752 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10753 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10754 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10755 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10756 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10757 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10758 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10760 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10761 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10762 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10763 VN.t671 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10764 VN.t670 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10765 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10766 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10767 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10768 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10769 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10770 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10771 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10772 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10773 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10774 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10775 fc2 s4 VN.t669 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10776 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10777 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10778 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10779 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10780 VN.t668 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10781 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10782 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10783 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10784 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10785 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10786 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10787 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10788 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10789 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10790 fc2 s4 VN.t667 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10791 VN.t666 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10792 fc2 s4 VN.t665 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10793 VN.t664 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10794 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10795 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10796 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10797 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10798 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10799 fc2 s4 VN.t663 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10800 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10801 VN.t662 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10802 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10803 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10804 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10805 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10806 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10807 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10808 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10809 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10810 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10811 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10812 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10813 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10814 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10815 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10816 VN.t661 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10817 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10818 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10819 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10820 fc2 s4 VN.t660 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10821 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10822 VN.t659 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10823 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10824 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10825 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10826 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10827 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10828 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10829 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10830 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10831 VN.t658 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10832 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10833 VN.t657 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10834 fc2 s4 VN.t656 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10835 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10836 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10837 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10838 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10839 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10840 fc2 s4 VN.t655 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X10841 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10842 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10844 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10845 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10846 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10847 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10848 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10849 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10850 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10851 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10852 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10853 fc2 s4 VN.t654 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10854 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10855 VN.t653 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10856 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10857 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10858 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10859 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10860 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10861 VN.t652 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10862 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10863 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10864 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10865 VN.t651 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10866 fc2 s4 VN.t650 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10867 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10868 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10869 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10870 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10871 VN.t649 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10872 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10873 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10874 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10875 VN.t648 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10876 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10877 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10878 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10879 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10880 fc2 s4 VN.t647 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10881 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10882 VN.t646 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10883 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10884 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10886 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10887 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10888 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10889 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10890 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10891 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10892 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10893 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10894 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10895 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10896 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10897 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10898 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10899 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10900 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10901 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10902 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10903 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10904 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10905 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10906 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10907 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10908 fc2 s4 VN.t645 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10909 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X10910 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10911 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10912 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10913 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10914 VN.t644 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10915 VN.t643 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10916 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10917 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10918 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10919 fc2 s4 VN.t642 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10920 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10921 VN.t641 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10922 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10923 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10924 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10925 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10926 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10927 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10928 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10929 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10930 VN.t640 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10931 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10932 fc2 s4 VN.t639 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10933 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10934 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10935 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10936 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10937 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10938 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10939 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10940 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10941 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10942 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10943 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10944 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10945 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10946 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10947 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10948 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10949 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10950 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10951 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10952 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10953 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10954 VN.t638 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10955 VN.t637 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10956 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10957 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10958 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10959 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X10960 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10961 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10962 VN.t636 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10963 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10964 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10965 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10966 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10967 VN.t635 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10968 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10969 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10970 VN.t634 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10971 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10972 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10973 VN.t633 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10974 fc2 s4 VN.t632 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10975 fc2 s4 VN.t631 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10976 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10977 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10978 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10980 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10981 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10982 fc2 s4 VN.t630 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10983 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10984 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10985 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10986 VN.t629 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10987 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10988 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X10989 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10990 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10991 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10992 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10993 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X10994 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10995 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10996 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10997 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10998 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X10999 fc2 s4 VN.t628 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11000 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11001 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11002 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11003 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11004 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11005 VN.t627 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11006 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11007 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11008 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11009 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11010 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11011 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11012 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11013 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11014 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11015 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11017 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11019 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11020 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11021 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11022 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11023 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11024 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11025 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11026 fc2 s4 VN.t626 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11027 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11028 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11029 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11030 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11031 fc2 s4 VN.t625 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11032 VN.t624 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11033 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11034 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11035 VN.t623 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11036 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11037 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11038 fc2 s4 VN.t622 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11039 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11040 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11041 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11042 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11043 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11044 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11045 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11046 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11047 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11048 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11049 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11050 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11051 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11052 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11053 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11054 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11055 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11056 VN.t621 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11057 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11058 fc2 s4 VN.t620 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11059 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11060 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11061 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11062 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11063 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11064 fc2 s4 VN.t619 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11065 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11066 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11068 VN.t618 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11069 fc2 s4 VN.t617 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11070 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11071 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11072 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11073 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11074 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11075 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11076 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11077 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11078 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11079 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11080 VN.t616 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11081 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11082 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11083 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11084 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11085 fc2 s4 VN.t615 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11086 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11088 VN.t614 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11089 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11090 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11091 VN.t613 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11092 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11093 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11094 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11095 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11096 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11097 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11098 fc2 s4 VN.t612 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11099 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11101 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11102 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11103 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11104 fc2 s4 VN.t611 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11105 VN.t610 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11106 VN.t609 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11107 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11108 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11109 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11111 fc2 s4 VN.t608 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11112 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11113 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11114 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11115 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11116 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11117 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11119 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11120 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11121 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11122 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11123 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11124 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11125 fc2 s4 VN.t607 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11126 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11127 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11128 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11129 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11130 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11131 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11132 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11133 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11134 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11135 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11136 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11137 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11138 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11139 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11140 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11141 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11142 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11143 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11144 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11145 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11146 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11147 fc2 s4 VN.t606 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11148 VN.t605 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11149 VN.t604 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11150 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11151 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11152 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11153 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11154 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11155 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11156 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11157 VN.t603 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11158 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11159 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11160 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11161 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11162 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11163 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11164 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11165 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11166 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11167 fc2 s4 VN.t602 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11168 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11169 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11170 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11171 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11172 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11173 fc2 s4 VN.t601 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11174 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11175 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11176 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11177 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11178 VN.t600 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11179 VN.t599 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11180 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11181 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11182 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11183 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11184 VN.t598 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11185 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11186 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11187 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11188 fc2 s4 VN.t597 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11189 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11190 fc2 s4 VN.t596 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11191 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11192 fc2 s4 VN.t595 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11193 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11194 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11195 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11196 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11197 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11198 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11199 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11200 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11201 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11202 fc2 s4 VN.t594 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11203 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11204 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11205 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11206 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11208 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11209 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11210 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11211 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11212 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11213 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11214 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11215 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11216 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11217 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11218 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11219 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11220 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11221 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11222 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11223 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11224 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11225 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11226 VN.t593 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11227 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11228 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11229 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11230 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11231 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11232 VN.t592 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11233 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11234 VN.t591 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11235 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11236 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11237 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11238 fc2 s4 VN.t590 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11239 fc2 s4 VN.t589 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11240 fc2 s4 VN.t588 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X11241 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11242 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11243 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11244 fc2 s4 VN.t587 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11245 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11246 fc2 s4 VN.t586 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11247 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11248 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11249 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11250 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11251 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11252 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11253 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11254 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11255 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11256 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11257 fc2 s4 VN.t585 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11258 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11260 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11261 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11262 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11263 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11264 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11265 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11266 VN.t584 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11267 fc2 s4 VN.t583 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11268 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11269 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11270 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11271 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11272 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11273 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11274 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11275 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11276 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11277 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11278 fc2 s4 VN.t582 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11279 fc2 s4 VN.t581 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11280 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11281 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11282 fc2 s4 VN.t580 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11283 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11284 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11285 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11286 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11287 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11288 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11290 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11291 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11292 VN.t579 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11293 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11294 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11295 fc2 s4 VN.t578 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11296 VN.t577 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11297 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11298 fc2 s4 VN.t576 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11299 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11300 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11301 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11302 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11303 VN.t575 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11304 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11305 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11306 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11307 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11308 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11309 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11310 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11311 VN.t574 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11312 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11313 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11314 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11315 fc2 s4 VN.t573 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11316 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11317 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11318 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11319 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11320 fc2 s4 VN.t572 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11321 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11322 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11323 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11324 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11325 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11326 fc2 s4 VN.t571 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11327 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11328 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11329 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11330 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11331 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11332 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11333 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11334 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11335 VN.t570 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11336 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11337 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11338 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11339 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11340 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11341 VN.t569 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11342 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11343 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11344 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11345 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11346 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11347 fc2 s4 VN.t568 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11348 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11349 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11350 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11351 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11352 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11353 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11354 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11355 VN.t567 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11356 fc2 s4 VN.t566 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11357 fc2 s4 VN.t565 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11358 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11359 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11360 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11361 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11362 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11363 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11364 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11365 fc2 s4 VN.t564 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11366 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11367 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11368 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11369 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11370 fc2 s4 VN.t563 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11371 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11372 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11373 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11374 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11375 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11377 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11378 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11379 VN.t562 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11380 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11381 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11382 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11383 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11384 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11385 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11386 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11387 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11388 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11389 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11390 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11391 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11392 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11393 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11394 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11395 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11396 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11397 fc2 s4 VN.t561 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11398 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11399 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11400 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11401 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11402 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11403 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11404 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11405 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11406 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11407 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11408 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11409 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11410 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11411 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11412 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11413 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11414 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11415 VN.t560 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11416 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11417 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11418 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11419 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11420 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11421 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11422 fc2 s4 VN.t559 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11423 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11424 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11425 fc2 s4 VN.t558 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11426 VN.t557 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11427 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11428 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11429 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11430 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11431 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11432 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11433 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11435 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11436 fc2 s4 VN.t556 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11437 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11438 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11439 fc2 s4 VN.t555 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11440 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11441 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11442 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11443 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11444 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11445 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11446 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11447 VN.t554 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11448 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11449 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11450 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11451 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11452 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11453 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11454 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11455 fc2 s4 VN.t553 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11456 VN.t552 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11457 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11458 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X11459 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11460 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11461 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11462 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11463 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11464 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11465 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11466 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11467 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11468 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11469 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11470 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11471 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11472 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11473 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11474 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11475 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11476 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11477 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11478 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11479 VN.t551 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11480 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11481 fc2 s4 VN.t550 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11482 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11483 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11484 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11485 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11486 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11487 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11488 fc2 s4 VN.t549 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11489 VN.t548 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11490 fc2 s4 VN.t547 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11491 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11492 fc2 s4 VN.t546 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11493 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11494 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11495 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11496 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11497 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11498 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11499 VN.t545 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11500 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11501 VN.t544 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11502 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11503 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11504 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11505 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11506 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11507 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11508 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11509 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11510 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11511 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11512 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11513 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11514 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11515 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11516 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11517 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11518 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11519 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11520 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11521 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11522 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11523 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11524 fc2 s4 VN.t543 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11525 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11526 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11527 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11528 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11529 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11530 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11531 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11532 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11533 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11534 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11535 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11536 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11537 fc2 s4 VN.t542 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11538 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11539 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11540 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11541 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11542 VN.t541 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11543 VN.t540 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11544 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11545 VN.t539 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11546 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11547 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11548 fc2 s4 VN.t538 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11549 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11550 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11551 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11552 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11553 fc2 s4 VN.t537 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11554 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11555 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11556 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11557 VN.t536 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11558 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11559 fc2 s4 VN.t535 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11560 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11561 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11562 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11563 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11564 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11565 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11566 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11567 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11568 VN.t534 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11569 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11570 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11571 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11572 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11573 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11574 fc2 s4 VN.t533 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11575 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11576 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11577 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11578 fc2 s4 VN.t532 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11579 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11580 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11582 VN.t531 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11583 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11584 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11585 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11586 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11587 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11588 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11589 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11590 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11591 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11592 fc2 s4 VN.t530 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11593 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11594 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11595 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11596 VN.t529 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11597 fc2 s4 VN.t528 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11598 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11599 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11600 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11601 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11602 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11603 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11604 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11605 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11606 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11607 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11608 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11609 fc2 s4 VN.t527 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11610 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11611 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11612 fc2 s4 VN.t526 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11613 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11614 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11615 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11616 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11618 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11619 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11620 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11621 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11622 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11623 fc2 s4 VN.t525 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11624 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11625 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11626 VN.t524 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11627 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11628 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11629 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11630 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11631 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11632 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11633 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11634 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11635 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11636 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11637 fc2 s4 VN.t523 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11638 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11639 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11640 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11641 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11642 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11643 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11644 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11645 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11646 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11647 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11648 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11649 fc2 s4 VN.t522 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11650 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11651 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11652 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11653 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11654 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11655 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11656 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11657 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11658 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11659 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11660 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11661 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11662 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11663 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11664 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11665 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11666 fc2 s4 VN.t521 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11667 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11668 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11669 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11670 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11671 VN.t520 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11672 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11673 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11674 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11675 fc2 s4 VN.t519 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11676 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11677 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11678 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11679 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11680 VN.t518 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11681 fc2 s4 VN.t517 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11682 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11683 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11684 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11685 VN.t516 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11686 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11687 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11688 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11689 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11690 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X11691 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11692 fc2 s4 VN.t515 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11693 fc2 s4 VN.t514 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11694 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11695 fc2 s4 VN.t513 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11696 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11697 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11698 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11699 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11700 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11701 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11702 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11703 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11704 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11705 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11706 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11707 fc2 s4 VN.t512 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11708 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11709 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11710 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11711 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11712 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11713 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11714 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11715 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11716 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11717 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11718 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11719 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11720 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11721 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11722 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11723 fc2 s4 VN.t511 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11724 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11725 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11726 fc2 s4 VN.t510 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11727 fc2 s4 VN.t509 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11728 VN.t508 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11729 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11730 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11731 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11732 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11733 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11734 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11735 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11736 fc2 s4 VN.t507 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11737 fc2 s4 VN.t506 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11738 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11739 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11740 VN.t505 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11741 fc2 s4 VN.t504 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11742 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11743 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11744 VN.t503 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11745 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11746 VN.t502 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11747 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11748 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11749 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11750 VN.t501 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11751 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11752 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11753 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11754 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11755 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11756 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11757 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11758 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11759 fc2 s4 VN.t500 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11760 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11761 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11762 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11763 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11764 VN.t499 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11765 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11766 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11767 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11768 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11769 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11770 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11771 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11772 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11773 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11774 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11775 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11776 VN.t498 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11777 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11778 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11779 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11780 VN.t497 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11781 VN.t496 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11782 VN.t495 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11783 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11784 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11785 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11786 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11787 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11788 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11789 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11790 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11791 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11792 fc2 s4 VN.t494 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11793 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11794 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11795 VN.t493 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11796 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11797 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11798 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11799 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11800 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11801 VN.t492 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11802 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11803 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11804 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11805 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11806 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11807 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11808 VN.t491 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11809 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11810 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11811 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11812 fc2 s4 VN.t490 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11813 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11814 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11815 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11816 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11817 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11818 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11819 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11820 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11821 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11822 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11823 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11824 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11825 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11826 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11827 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11828 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11829 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11830 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11831 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11832 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11833 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11834 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11835 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11836 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11837 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11838 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11839 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11840 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11841 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11842 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11843 VN.t489 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11844 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11845 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11846 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11847 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11848 fc2 s4 VN.t488 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11849 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11850 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11851 VN.t487 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11852 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11853 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11854 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11855 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11856 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11857 VN.t486 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11858 VN.t485 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X11859 fc2 s4 VN.t484 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11860 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11861 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11862 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11863 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11864 fc2 s4 VN.t483 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11865 VN.t482 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11866 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11867 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11868 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11869 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11870 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11871 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11872 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11873 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11874 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11875 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11876 fc2 s4 VN.t481 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11877 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11878 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11879 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11880 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11881 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11882 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11883 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11884 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11885 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11886 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11887 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11888 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11889 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11890 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11891 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11892 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11893 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11894 VN.t480 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11895 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11896 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11897 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11898 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11899 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11900 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11901 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11902 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11903 VN.t479 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11904 fc2 s4 VN.t478 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X11905 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11906 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11907 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11908 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11909 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11910 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11911 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X11912 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11913 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11914 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11915 fc2 s4 VN.t477 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11916 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11917 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11918 VN.t476 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11919 fc2 s4 VN.t475 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11920 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11921 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11922 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11923 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11924 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11925 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11926 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11927 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11929 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11930 VN.t474 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11931 fc2 s4 VN.t473 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11932 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11933 fc2 s4 VN.t472 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11934 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11935 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11936 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11937 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11938 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11939 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11940 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11941 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11942 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11943 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11944 VN.t471 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11945 fc2 s4 VN.t470 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11946 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11947 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11948 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11949 VN.t469 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11950 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11951 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11952 fc2 s4 VN.t468 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11953 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11954 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11955 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11956 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11957 fc2 s4 VN.t467 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11958 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11959 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11960 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11961 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11962 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11963 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11964 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11965 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11966 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11967 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11968 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11969 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11970 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11971 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11972 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11973 fc2 s4 VN.t466 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11974 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11975 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11976 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11977 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11978 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11979 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11980 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11981 fc2 s4 VN.t465 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11982 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11983 fc2 s4 VN.t464 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X11984 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11985 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X11986 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11987 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X11988 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11989 VN.t463 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11990 VN.t462 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11991 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11992 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11993 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11994 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11995 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11996 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X11997 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11998 fc2 s4 VN.t461 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11999 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12000 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12001 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12002 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12003 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12004 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12005 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12006 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12007 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12009 VN.t460 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12010 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12011 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12012 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12013 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12014 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12015 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12016 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12017 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12018 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12019 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12020 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12021 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12022 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12023 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12024 fc2 s4 VN.t459 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12025 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12026 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12027 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12028 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12029 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12030 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12031 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12032 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12033 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12034 VN.t458 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12035 fc2 s4 VN.t457 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12036 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12037 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12038 VN.t456 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12039 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12040 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12041 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12042 VN.t455 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12043 fc2 s4 VN.t454 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12044 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12045 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12046 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12047 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12048 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12049 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12050 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12051 fc2 s4 VN.t453 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12052 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12053 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12054 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12055 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12056 fc2 s4 VN.t452 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12057 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12058 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12059 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12060 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12061 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12062 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12063 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12064 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12065 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12066 VN.t451 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12067 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12068 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12069 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12070 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12071 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12072 VN.t450 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12073 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12074 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12075 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12076 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12077 VN.t449 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12078 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12079 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12080 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12081 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12082 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12083 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12084 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12085 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12086 fc2 s4 VN.t448 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12087 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12088 VN.t447 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12089 VN.t446 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12090 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12091 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12092 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12093 VN.t445 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12094 VN.t444 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12095 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12096 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12097 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12098 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12099 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12100 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12101 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12102 VN.t443 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12103 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12104 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12105 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12106 fc2 s4 VN.t442 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12107 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12108 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12109 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12110 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12111 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12112 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12113 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12114 fc2 s4 VN.t441 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12115 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12116 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12117 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12118 fc2 s4 VN.t440 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12119 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12120 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12121 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12122 fc2 s4 VN.t439 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12123 VN.t438 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12124 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12125 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12126 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12127 VN.t437 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12128 VN.t436 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12129 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12130 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12131 VN.t435 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12132 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12133 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12134 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12135 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12136 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12137 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12138 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12139 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12140 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12141 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12142 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12143 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12144 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12145 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12146 fc2 s4 VN.t434 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12147 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12148 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12149 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12150 VN.t433 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12151 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12152 VN.t432 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12153 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12154 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12155 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12156 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12157 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12158 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12159 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12160 VN.t431 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12161 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12162 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12163 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12164 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12165 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12166 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12167 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12168 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12169 fc2 s4 VN.t430 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12170 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12171 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12172 fc2 s4 VN.t429 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12173 VN.t428 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12174 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12175 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12176 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12177 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12178 VN.t427 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12180 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12181 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12182 VN.t426 s4 fc2 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12183 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12184 fc2 s4 VN.t425 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12185 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12186 VN.t424 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12187 VN.t423 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12188 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12189 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12190 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12191 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12192 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12193 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12194 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12195 VN.t422 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12196 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12197 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12198 fc2 s4 VN.t421 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12199 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12200 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12201 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12202 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12203 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12204 VN.t420 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12205 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12206 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12208 VN.t419 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12209 fc2 s4 VN.t418 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12210 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12211 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12212 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12213 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12214 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12215 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12216 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12217 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12218 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12219 VN.t417 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12220 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12221 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12222 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12223 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12224 VN.t416 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12225 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12226 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12227 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12228 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12229 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12230 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12231 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12232 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12233 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12234 VN.t415 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12235 VN.t414 s4 fc2 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12236 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12237 VN.t413 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12238 VN.t412 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12239 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12240 fc2 s4 VN.t411 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12241 fc2 s4 VN.t410 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12242 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12243 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12244 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12245 fc2 s4 VN.t409 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12246 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12247 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12248 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12249 VN.t408 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12250 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12251 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12252 VN.t407 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12253 VN.t406 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12254 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12255 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12256 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12257 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12258 fc2 s4 VN.t405 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12260 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12261 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12262 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12263 VN.t404 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12264 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12265 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12266 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12267 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12268 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12269 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12270 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12271 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12272 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12273 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12274 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12275 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12276 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12277 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12278 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12279 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12280 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12281 fc2 s4 VN.t403 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12282 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12283 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12284 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12285 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12286 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12287 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12288 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12289 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12290 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12291 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12292 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12293 VN.t402 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12294 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12295 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12296 fc2 s4 VN.t401 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12297 VN.t400 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12298 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12299 fc2 s4 VN.t399 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12300 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12301 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12302 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12303 VN.t398 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12304 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12305 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12306 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12307 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12308 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12309 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12310 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12311 VN.t397 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12312 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12313 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12314 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12315 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12316 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12317 VN.t396 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12318 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12319 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12320 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12321 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12322 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12323 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12324 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12325 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12326 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12327 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12328 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12329 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12330 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12331 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12332 fc2 s4 VN.t395 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12333 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12334 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12335 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12336 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12337 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12338 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12339 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12340 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12341 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12342 fc2 s4 VN.t394 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12343 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12344 VN.t393 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12345 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12346 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12347 VN.t392 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12348 VN.t391 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12349 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12350 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12351 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12352 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12353 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12354 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12355 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12356 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12357 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12358 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12359 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12360 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12361 VN.t390 s4 fc2 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12362 fc2 s4 VN.t389 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12363 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12364 fc2 s4 VN.t388 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12365 VN.t387 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12366 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12367 VN.t386 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12368 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12369 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12370 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12371 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12372 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12373 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12374 fc2 s4 VN.t385 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12375 VN.t384 s4 fc2 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12376 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12377 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12378 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12379 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12380 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12381 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12382 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12383 fc2 s4 VN.t383 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12384 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12385 VN.t382 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12386 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12387 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12388 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12389 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12390 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12391 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12392 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12393 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12394 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12395 VN.t381 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12396 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12397 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12398 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12399 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12400 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12401 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12402 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12403 fc2 s4 VN.t380 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12404 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12405 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12406 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12407 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12408 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12409 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12410 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12411 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12412 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12413 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12414 fc2 s4 VN.t379 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12415 VN.t378 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12416 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12417 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12418 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12419 VN.t377 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12420 VN.t376 s4 fc2 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12421 fc2 s4 VN.t375 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12422 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12423 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12424 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12425 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12426 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12427 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12428 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12429 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12430 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12431 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12432 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12433 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12435 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12436 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12437 fc2 s4 VN.t374 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12438 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12439 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12440 VN.t373 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12441 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12442 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12443 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12444 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12445 VN.t372 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12446 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12447 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12448 VN.t371 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12449 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12450 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12451 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12452 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12453 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12454 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12455 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12456 VN.t370 s4 fc2 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12457 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12458 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12459 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12460 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12461 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12462 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12463 fc2 s4 VN.t369 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12464 VN.t368 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12465 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12466 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12467 VN.t367 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12468 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12469 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12470 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12471 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12472 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12473 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12474 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12475 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12476 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12477 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12478 VN.t366 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12479 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12480 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12481 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12482 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12483 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12484 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12485 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12486 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12487 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12488 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12489 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12490 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12491 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12492 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12493 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12494 VN.t365 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12495 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12496 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12497 VN.t364 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12498 VN.t363 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12499 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12500 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12501 fc2 s4 VN.t362 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12502 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12503 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12504 VN.t361 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12505 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12506 VN.t360 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12507 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12508 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12509 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12510 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12511 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12512 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12513 VN.t359 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12514 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12515 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12516 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12517 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12518 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12519 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12520 fc2 s4 VN.t358 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12521 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12522 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12523 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12524 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12525 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12526 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12527 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12528 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12529 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12530 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12531 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12532 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12533 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12534 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12535 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12536 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12537 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12538 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12539 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12540 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12541 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12542 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12543 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12544 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12545 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12546 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12547 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12548 fc2 s4 VN.t357 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12549 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12550 VN.t356 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12551 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12552 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12553 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12554 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12555 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12556 fc2 s4 VN.t355 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12557 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12558 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12559 VN.t354 s4 fc2 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12560 VN.t353 s4 fc2 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12561 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12562 fc2 s4 VN.t352 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12563 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12564 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12565 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12566 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12567 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12568 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12569 fc2 s4 VN.t351 VN.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12570 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12571 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12572 VN.t349 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12573 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12574 fc2 s4 VN.t348 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12575 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12576 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12577 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12578 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12579 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12580 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12581 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12582 fc2 s4 VN.t347 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12583 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12584 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12585 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12586 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12587 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12588 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12589 VN.t346 s4 fc2 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12590 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12591 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12592 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12593 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12594 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12595 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12596 VN.t345 s4 fc2 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12597 fc2 s4 VN.t344 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12598 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12599 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12600 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12601 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12602 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12603 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12604 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12605 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12606 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12607 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12608 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12609 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12610 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12611 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12612 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12613 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12614 fc2 s4 VN.t343 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12615 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12616 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12617 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12618 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12619 fc2 s4 VN.t342 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12620 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12621 fc2 s4 VN.t341 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12622 VN.t340 s4 fc2 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12623 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12624 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12625 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12626 VN.t339 s4 fc2 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12627 fc2 s4 VN.t338 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12628 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12629 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12630 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12631 fc2 s4 VN.t337 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12632 VN.t336 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12633 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12634 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12635 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12636 fc2 s4 VN.t335 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X12637 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12638 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12639 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12640 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12641 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12642 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12643 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12644 VN.t334 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12645 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12646 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12647 fc2 s4 VN.t333 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12648 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12649 fc2 s4 VN.t332 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12650 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12651 VN.t331 s4 fc2 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12652 VN.t330 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12653 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12654 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12655 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12656 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12657 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12658 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12659 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12660 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12661 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12662 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12663 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12664 fc2 s4 VN.t329 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12665 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12666 fc2 s4 VN.t328 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12667 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12668 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12669 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12670 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12671 VN.t327 s4 fc2 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12672 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12673 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12674 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12675 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12676 fc2 s4 VN.t326 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12677 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12678 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12679 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12680 fc2 s4 VN.t325 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12681 VN.t324 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12682 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12683 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12684 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12685 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12686 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12687 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12688 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12689 fc2 s4 VN.t323 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12690 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12691 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12692 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12693 fc2 s4 VN.t322 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12694 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12695 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12696 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12697 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12698 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12699 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12700 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12701 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12702 VN.t321 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12703 VN.t320 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12704 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12705 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12706 fc2 s4 VN.t319 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12707 fc2 s4 VN.t318 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12708 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12709 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12710 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12711 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12712 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12713 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12714 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12715 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12716 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12717 VN.t317 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12718 fc2 s4 VN.t316 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12719 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12720 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12721 VN.t315 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12722 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12723 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12724 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12725 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12726 VN.t314 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12727 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12728 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12729 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12730 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12731 VN.t313 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12732 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12733 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12734 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12735 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12736 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12737 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12738 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12739 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12740 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12741 fc2 s4 VN.t312 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12742 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12743 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12744 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12745 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12746 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12747 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12748 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12749 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12750 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12751 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12752 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12753 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12754 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12755 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12756 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12757 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12758 VN.t311 s4 fc2 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12759 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12760 VN.t310 s4 fc2 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12761 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12762 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12763 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12764 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12765 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12766 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12767 fc2 s4 VN.t309 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12768 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12769 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12770 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12771 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12772 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12773 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12774 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12775 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12776 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12777 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12778 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12779 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12780 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12781 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12782 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12783 VN.t308 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12784 fc2 s4 VN.t307 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12785 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12786 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12787 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12788 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12789 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12790 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12791 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12792 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12793 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12794 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12795 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12796 fc2 s4 VN.t306 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12797 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12798 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12799 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12800 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12801 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12802 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12803 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12804 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12805 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X12806 fc2 s4 VN.t305 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12807 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12808 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12809 fc2 s4 VN.t304 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12810 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12811 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12812 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12813 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12814 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12815 fc2 s4 VN.t303 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12816 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12817 VN.t302 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12818 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12819 VN.t301 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12820 VN.t300 s4 fc2 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12821 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12822 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12823 VN.t299 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12824 fc2 s4 VN.t298 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12825 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12826 fc2 s4 VN.t297 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12827 fc2 s4 VN.t296 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12828 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12829 fc2 s4 VN.t295 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12830 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12831 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12832 fc2 s4 VN.t294 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12833 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12834 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12835 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12836 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12837 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12838 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12839 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12840 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12841 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12842 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12844 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12845 fc2 s4 VN.t293 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12846 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12847 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12848 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12849 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12850 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12851 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12852 fc2 s4 VN.t292 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12853 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12854 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12855 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12856 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12857 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12858 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12859 fc2 s4 VN.t291 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12860 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12861 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12862 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12863 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12864 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12865 fc2 s4 VN.t290 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12866 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12867 fc2 s4 VN.t289 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12868 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12869 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12870 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12871 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12872 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12873 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12874 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12875 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12876 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12877 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12878 fc2 s4 VN.t288 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12879 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12880 VN.t287 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12881 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12882 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12883 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12884 VN.t286 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12886 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12887 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12888 fc2 s4 VN.t285 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12889 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12890 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12891 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12892 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12893 VN.t284 s4 fc2 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12894 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12895 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12896 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12897 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12898 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12899 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12900 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12901 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12902 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12904 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12905 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12906 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12907 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12908 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12909 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12910 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12911 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12912 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12913 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12914 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12915 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12916 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12917 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12918 VN.t283 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X12919 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12920 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12921 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12922 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12923 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12924 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12925 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12926 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12927 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12928 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12929 VN.t282 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12930 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12931 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12932 fc2 s4 VN.t281 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12933 fc2 s4 VN.t280 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12934 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12935 VN.t279 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12936 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12937 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12938 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12939 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12940 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12941 fc2 s4 VN.t278 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X12942 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12943 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12944 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12945 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12946 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12947 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12948 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12949 fc2 s4 VN.t277 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12950 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12951 fc2 s4 VN.t276 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12952 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12953 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12954 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12955 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12956 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12957 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12958 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12959 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12960 VN.t275 s4 fc2 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12961 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12962 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X12963 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12964 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12965 VN.t274 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12966 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12967 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12968 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12969 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12970 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12971 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12972 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12973 fc2 s4 VN.t273 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12974 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X12975 VN.t272 s4 fc2 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12976 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12977 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12978 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12979 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12980 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12981 VN.t271 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12982 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12983 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12984 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12985 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12986 fc2 s4 VN.t270 VN.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12987 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12988 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12989 fc2 s4 VN.t268 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12990 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12991 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12992 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12993 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12994 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12995 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12996 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12997 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12998 fc2 s4 VN.t267 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X12999 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13000 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13001 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13002 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13003 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13004 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13005 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13006 VN.t266 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13007 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13008 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13009 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13010 VN.t265 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13011 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13012 fc2 s4 VN.t264 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13013 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13014 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13015 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13016 fc2 s4 VN.t263 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13017 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13019 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13020 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13021 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13022 fc2 s4 VN.t262 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13023 VN.t261 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13024 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13025 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13026 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13027 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13028 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13029 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13030 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13031 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13032 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13033 fc2 s4 VN.t260 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13034 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13035 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13036 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13037 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13038 fc2 s4 VN.t259 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13039 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13040 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13041 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13042 VN.t258 s4 fc2 VN.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13043 fc2 s4 VN.t256 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13044 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13045 fc2 s4 VN.t255 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13046 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13047 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13048 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13049 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13050 VN.t254 s4 fc2 VN.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13051 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13052 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13053 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13054 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13055 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13056 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13057 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13058 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13059 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13060 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13061 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13062 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13063 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13064 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13065 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13066 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13067 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13068 VN.t252 s4 fc2 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13069 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13070 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13071 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13072 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13073 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13074 fc2 s4 VN.t251 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13075 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13076 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13077 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13078 VN.t250 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13079 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13080 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13081 VN.t249 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13082 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13083 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13084 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13085 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13086 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13087 fc2 s4 VN.t248 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13088 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13089 fc2 s4 VN.t247 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13090 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13091 fc2 s4 VN.t246 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13092 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13093 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13094 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13095 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13096 VN.t245 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13097 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13098 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13099 VN.t244 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13100 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13101 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13102 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13103 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13104 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13105 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13106 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13107 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13108 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13109 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13110 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13111 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13112 fc2 s4 VN.t243 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13113 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13114 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13115 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13116 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13117 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13118 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13119 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13120 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13121 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13122 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13123 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13124 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13125 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13126 fc2 s4 VN.t242 VN.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13127 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13128 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13129 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13130 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13131 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13132 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13133 fc2 s4 VN.t240 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13134 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13135 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13136 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13137 VN.t239 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13138 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13139 VN.t238 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13140 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13141 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13142 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13143 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13144 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13145 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13146 fc2 s4 VN.t237 VN.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13147 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13148 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13149 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13150 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13151 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13152 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13153 fc2 s4 VN.t235 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13154 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13155 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13156 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13157 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13158 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13159 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13160 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13161 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13162 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13163 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13164 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13165 fc2 s4 VN.t234 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13166 fc2 s4 VN.t233 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13167 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13168 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13169 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13170 fc2 s4 VN.t232 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13171 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13172 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13173 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13174 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13175 VN.t231 s4 fc2 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13176 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13177 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13178 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13179 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13180 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13181 VN.t230 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13182 fc2 s4 VN.t229 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13183 fc2 s4 VN.t228 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13184 fc2 s4 VN.t227 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13185 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13186 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13187 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13188 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13189 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13190 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13191 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13192 fc2 s4 VN.t226 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13193 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13194 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13195 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13196 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13197 fc2 s4 VN.t225 VN.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13198 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13199 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13200 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13201 fc2 s4 VN.t223 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13202 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13203 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13204 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13205 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13206 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13207 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13208 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13209 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13210 VN.t222 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13211 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13212 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13213 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13214 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13215 fc2 s4 VN.t221 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13216 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13217 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13218 fc2 s4 VN.t220 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13219 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13220 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13221 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13222 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13223 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13224 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13225 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13226 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13227 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13228 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13229 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13230 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13231 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13232 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13233 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13234 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13235 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13236 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13237 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13238 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13239 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13240 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13241 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13242 VN.t219 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13243 VN.t218 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13244 fc2 s4 VN.t217 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13245 fc2 s4 VN.t216 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13246 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13247 fc2 s4 VN.t215 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13248 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13249 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13250 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13251 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13252 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13253 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13254 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13255 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13256 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13257 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13258 fc2 s4 VN.t214 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13259 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13260 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13261 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13262 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13263 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13264 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13265 fc2 s4 VN.t213 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13266 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13267 fc2 s4 VN.t212 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13268 VN.t211 s4 fc2 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13269 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13270 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13271 fc2 s4 VN.t210 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13272 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13273 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13274 fc2 s4 VN.t209 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13275 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13276 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13277 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13278 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13279 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13280 VN.t208 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13281 fc2 s4 VN.t207 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13282 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13283 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13284 VN.t206 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13285 fc2 s4 VN.t205 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13286 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13287 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13288 VN.t204 s4 fc2 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13289 fc2 s4 VN.t203 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13290 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13291 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13292 fc2 s4 VN.t202 VN.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13293 fc2 s4 VN.t200 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13294 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13295 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13296 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13297 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13298 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13299 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13300 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13301 fc2 s4 VN.t199 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13302 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13303 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13304 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13305 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13306 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13307 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13308 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13309 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13310 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13311 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13312 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13313 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13314 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13315 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13316 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13317 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13318 fc2 s4 VN.t198 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13319 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13320 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13321 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13322 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13323 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13324 fc2 s4 VN.t197 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13325 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13326 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13327 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13328 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13329 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13330 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13331 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13332 fc2 s4 VN.t196 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13333 fc2 s4 VN.t195 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13334 VN.t194 s4 fc2 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13335 fc2 s4 VN.t193 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13336 fc2 s4 VN.t192 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13337 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13338 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13339 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13340 VN.t191 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13341 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13342 VN.t190 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13343 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13344 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13345 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13346 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13347 VN.t189 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13348 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13349 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13350 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13351 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13352 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13353 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13354 fc2 s4 VN.t188 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13355 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13356 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13357 fc2 s4 VN.t187 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13358 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13359 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13360 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13361 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13362 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13363 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13364 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13365 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13366 fc2 s4 VN.t186 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13367 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13368 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13369 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13370 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13371 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13372 VN.t185 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13373 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13374 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13375 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13376 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13377 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13378 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13379 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13380 VN.t184 s4 fc2 VN.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13381 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13382 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13383 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13384 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13385 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13386 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13387 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13388 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13389 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13390 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13391 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13392 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13393 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13394 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13395 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13396 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13397 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13398 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13399 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13400 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13401 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13402 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13403 VN.t182 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13404 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13405 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13406 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13407 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13408 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13409 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13410 VN.t181 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13411 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13412 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13413 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13414 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13415 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13416 fc2 s4 VN.t180 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13417 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13418 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13419 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13420 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13421 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13422 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13423 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13424 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13425 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13426 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13427 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13428 VN.t179 s4 fc2 VN.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13429 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13430 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13431 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13432 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13433 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13434 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13435 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13436 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13437 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13438 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13439 VN.t177 s4 fc2 VN.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13440 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13441 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13442 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13443 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13444 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13445 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13446 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13447 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13448 fc2 s4 VN.t175 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13449 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13450 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13451 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13452 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13453 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13454 VN.t174 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13455 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13456 VN.t173 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13457 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13458 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13459 VN.t172 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13460 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13461 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13462 fc2 s4 VN.t171 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13463 VN.t170 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13464 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13465 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13466 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13467 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13468 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13469 VN.t169 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13470 fc2 s4 VN.t168 VN.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13471 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13472 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13473 VN.t166 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13474 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13475 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13476 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13477 fc2 s4 VN.t165 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13478 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13479 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13480 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13481 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13482 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13483 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13484 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13485 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13486 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13487 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13488 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13489 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13490 fc2 s4 VN.t164 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13491 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13492 fc2 s4 VN.t163 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13493 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13494 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13495 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13496 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13497 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13498 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13499 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13500 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13501 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13502 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13503 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13504 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13505 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13506 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13507 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13508 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13509 VN.t162 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13510 fc2 s4 VN.t161 VN.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13511 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13512 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13513 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13514 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13515 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13516 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13517 fc2 s4 VN.t159 VN.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13518 VN.t157 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13519 VN.t156 s4 fc2 VN.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13520 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13521 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13522 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13523 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13524 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13525 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13526 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13527 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13528 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13529 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13530 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13531 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13532 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13533 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13534 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13535 fc2 s4 VN.t154 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13536 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13537 fc2 s4 VN.t153 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13538 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13539 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13540 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13541 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13542 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13543 VN.t152 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13544 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13545 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13546 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13547 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13548 fc2 s4 VN.t151 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13549 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13550 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13551 fc2 s4 VN.t150 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13552 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13553 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13554 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13555 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13556 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13557 VN.t149 s4 fc2 VN.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13558 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13559 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13560 fc2 s4 VN.t147 VN.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13561 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13562 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13563 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13564 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13565 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13566 fc2 s4 VN.t145 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13567 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13568 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13569 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13570 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13571 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13572 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13573 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13574 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13575 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13576 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13577 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13578 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13579 fc2 s4 VN.t144 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13580 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13581 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13582 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13583 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13584 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13585 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13586 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13587 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13588 fc2 s4 VN.t143 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13589 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13590 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13591 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13592 VN.t142 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13593 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13594 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13595 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13596 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13597 fc2 s4 VN.t141 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13598 VN.t140 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13599 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13600 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13601 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13602 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13603 fc2 s4 VN.t139 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13604 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13605 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13606 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13607 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13608 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13609 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13610 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13611 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13612 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13613 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13614 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13615 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13616 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13617 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13618 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13619 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13620 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13621 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13622 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13623 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13624 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13625 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13626 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13627 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13628 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13629 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13630 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13631 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13632 fc2 s4 VN.t138 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13633 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13634 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13635 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13636 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13637 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13638 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13639 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13640 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13641 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13642 fc2 s4 VN.t137 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13643 VN.t136 s4 fc2 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13644 VN.t135 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13645 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13646 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13647 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13648 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13649 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13650 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13651 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13652 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13653 VN.t134 s4 fc2 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13654 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13655 VN.t133 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13656 fc2 s4 VN.t132 VN.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13657 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13658 fc2 s4 VN.t130 VN.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13659 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13660 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13661 VN.t128 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13662 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13663 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13664 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13665 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13666 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13667 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13668 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13669 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13670 fc2 s4 VN.t127 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13671 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13672 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13673 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13674 fc2 s4 VN.t126 VN.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13675 VN.t124 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13676 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13677 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13678 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13679 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13680 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13681 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13682 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13683 fc2 s4 VN.t123 VN.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13684 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13685 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13686 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13687 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13688 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13689 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13690 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13691 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13692 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13693 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13694 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13695 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13696 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13697 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13698 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13699 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13700 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13701 VN.t121 s4 fc2 VN.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13702 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13703 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13704 fc2 s4 VN.t119 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13705 fc2 s4 VN.t118 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13706 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13707 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13708 VN.t117 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13709 VN.t116 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13710 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13711 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13712 fc2 s4 VN.t115 VN.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13713 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13714 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13715 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13716 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13717 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13718 VN.t113 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13719 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13720 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13721 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13722 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13723 fc2 s4 VN.t112 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13724 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13725 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13726 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13727 VN.t111 s4 fc2 VN.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13728 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13729 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13730 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13731 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13732 fc2 s4 VN.t109 VN.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13733 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13734 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13735 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13736 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13737 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13738 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13739 fc2 s4 VN.t107 VN.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13740 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13741 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13742 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13743 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13744 VN.t105 s4 fc2 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13745 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13746 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13747 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13748 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13749 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13750 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13751 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13752 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13753 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13754 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13755 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13756 VN.t104 s4 fc2 VN.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13757 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13758 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13759 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13760 VN.t102 s4 fc2 VN.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13761 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13762 VN.t100 s4 fc2 VN.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13763 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13764 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13765 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13766 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13767 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13768 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13769 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13770 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13771 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13772 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13773 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13774 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13775 VN.t98 s4 fc2 VN.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13776 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13777 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13778 fc2 s4 VN.t96 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13779 VN.t95 s4 fc2 VN.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13780 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13781 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13782 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13783 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13784 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13785 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13786 VN.t93 s4 fc2 VN.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13787 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13788 VN.t91 s4 fc2 VN.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13789 fc2 s4 VN.t89 VN.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13790 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13791 VN.t87 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13792 VN.t86 s4 fc2 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13793 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13794 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13795 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13796 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13797 VN.t85 s4 fc2 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13798 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13799 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13800 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13801 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13802 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13803 VN.t84 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13804 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13805 VN.t83 s4 fc2 VN.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13806 VN.t81 s4 fc2 VN.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13807 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13808 fc2 s4 VN.t79 VN.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13809 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13810 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13811 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13812 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13813 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13814 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13815 VN.t77 s4 fc2 VN.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13816 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13817 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13818 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13819 fc2 s4 VN.t75 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13820 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13821 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13822 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13823 VN.t74 s4 fc2 VN.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13824 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13825 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13826 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13827 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13828 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13829 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13830 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13831 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13832 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13833 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13834 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13835 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13836 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13837 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13838 VN.t72 s4 fc2 VN.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13839 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13840 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13841 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13842 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13843 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13844 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13845 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13846 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13847 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13848 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13849 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13850 VN.t70 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13851 VN.t69 s4 fc2 VN.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13852 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13853 fc2 s4 VN.t67 VN.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13854 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13855 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13856 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13857 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13858 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13859 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13860 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13861 VN.t65 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13862 VN.t64 s4 fc2 VN.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13863 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13864 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13865 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13866 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13867 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13868 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13869 fc2 s4 VN.t62 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13870 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13871 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13872 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13873 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13874 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13875 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13876 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13877 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13878 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13879 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13880 fc2 s4 VN.t61 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13881 VN.t60 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X13882 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13883 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13884 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13885 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13886 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13887 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13888 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13889 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X13890 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13891 VN.t59 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13892 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13893 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13894 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13895 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13896 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13897 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13898 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13899 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13900 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13901 fc2 s4 VN.t58 VN.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13902 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13903 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13904 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13905 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13906 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13907 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13908 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13909 VN.t56 s4 fc2 VN.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13910 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13911 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13912 VN.t54 s4 fc2 VN.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13913 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13914 VN.t52 s4 fc2 VN.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13915 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13916 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13917 fc2 s4 VN.t50 VN.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13918 fc2 s4 VN.t48 VN.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13919 VN.t46 s4 fc2 VN.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13920 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13921 fc2 s4 VN.t44 VN.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13922 fc2 s4 VN.t42 VN.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13923 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13924 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13925 VN.t40 s4 fc2 VN.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13926 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13927 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13928 VN.t38 s4 fc2 VN.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13929 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13930 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13931 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13932 VN.t36 s4 fc2 VN.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13933 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13934 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13935 VN.t34 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13936 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13937 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X13938 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13939 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13940 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13941 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13942 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13943 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X13944 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13945 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13946 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13947 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13948 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13949 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13950 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13951 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13952 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13953 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13954 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13955 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13956 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13957 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13958 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13959 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13960 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13961 fc2 s4 VN.t33 VN.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13962 fc2 s4 VN.t31 VN.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13963 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X13964 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13965 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13966 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13967 VN.t29 s4 fc2 VN.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13968 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13969 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13970 VN.t27 s4 fc2 VN.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13971 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13972 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13973 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13974 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13975 VN.t25 s4 fc2 VN.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13976 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13977 fc2 s4 VN.t23 VN.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13978 VN.t21 s4 fc2 VN.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13979 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13980 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13981 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13982 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13983 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13984 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13985 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13986 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13987 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13988 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13989 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13990 fc2 s4 VN.t19 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13991 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13992 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13993 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13994 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X13995 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13996 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13997 VN.t18 s4 fc2 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13998 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X13999 fc2 s4 VN.t17 VN.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14000 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14001 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14002 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14003 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14004 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14005 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14006 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14007 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14008 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14009 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14010 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X14011 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14012 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14013 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X14014 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14015 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14016 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14017 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14018 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14019 VN.t15 s4 fc2 VN.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14020 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14021 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14022 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14023 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14024 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14025 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14026 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14027 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14028 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14029 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14030 fc2 s4 VN.t13 VN.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14031 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14032 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14033 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14034 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14035 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14036 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14037 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14038 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14039 fc2 s4 VN.t11 VN.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14040 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14041 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14042 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14043 VN.t9 s4 fc2 VN.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X14044 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14045 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X14046 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14047 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14048 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14049 VN.t7 s4 fc2 VN.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14050 VN.t5 s4 fc2 VN.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14051 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14052 VP s1 fc1 VP sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14053 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14054 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14055 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X14056 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14057 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14058 VN.t3 s4 fc2 VN.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14059 fc2 s3 out fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14060 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X14061 fc1 s2 out fc1 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14062 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X14063 VN.t1 s4 fc2 VN.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
R0 VN.n11534 VN.n11533 169.353
R1 VN.n11536 VN.n11535 137.98
R2 VN.n10716 VN.n10715 137.98
R3 VN.n9856 VN.n9855 137.98
R4 VN.n9008 VN.n9007 137.98
R5 VN.n8175 VN.n8174 137.98
R6 VN.n7364 VN.n7363 137.98
R7 VN.n6571 VN.n6570 137.98
R8 VN.n5795 VN.n5794 137.98
R9 VN.n5032 VN.n5031 137.98
R10 VN.n4291 VN.n4290 137.98
R11 VN.n3563 VN.n3562 137.98
R12 VN.n2857 VN.n2856 137.98
R13 VN.n2164 VN.n2163 137.98
R14 VN.n1490 VN.n1489 137.98
R15 VN.n840 VN.n839 137.98
R16 VN.n813 VN.n812 137.98
R17 VN.n13129 VN.n13128 137.98
R18 VN.n10710 VN.n10709 137.754
R19 VN.n9850 VN.n9849 137.754
R20 VN.n9002 VN.n9001 137.754
R21 VN.n8169 VN.n8168 137.754
R22 VN.n7358 VN.n7357 137.754
R23 VN.n6565 VN.n6564 137.754
R24 VN.n5789 VN.n5788 137.754
R25 VN.n5026 VN.n5025 137.754
R26 VN.n4285 VN.n4284 137.754
R27 VN.n3557 VN.n3556 137.754
R28 VN.n2851 VN.n2850 137.754
R29 VN.n2158 VN.n2157 137.754
R30 VN.n1484 VN.n1483 137.754
R31 VN.n834 VN.n833 137.754
R32 VN.n807 VN.n806 137.754
R33 VN.n13123 VN.n13122 137.754
R34 VN.n12358 VN.n12357 135.611
R35 VN.n11532 VN.n11531 129.387
R36 VN.n10713 VN.n10712 129.387
R37 VN.n9853 VN.n9852 129.387
R38 VN.n9005 VN.n9004 129.387
R39 VN.n8172 VN.n8171 129.387
R40 VN.n7361 VN.n7360 129.387
R41 VN.n6568 VN.n6567 129.387
R42 VN.n5792 VN.n5791 129.387
R43 VN.n5029 VN.n5028 129.387
R44 VN.n4288 VN.n4287 129.387
R45 VN.n3560 VN.n3559 129.387
R46 VN.n2854 VN.n2853 129.387
R47 VN.n2161 VN.n2160 129.387
R48 VN.n1487 VN.n1486 129.387
R49 VN.n837 VN.n836 129.387
R50 VN.n810 VN.n809 129.387
R51 VN.n13126 VN.n13125 129.387
R52 VN.n11382 VN.n11381 91.65
R53 VN.n12369 VN.n12368 91.65
R54 VN.n2510 VN.n2509 91.65
R55 VN.n1818 VN.n1817 91.65
R56 VN.n1145 VN.n1144 91.65
R57 VN.n492 VN.n491 91.65
R58 VN.n12700 VN.n12699 91.65
R59 VN.n3942 VN.n3941 91.65
R60 VN.n3215 VN.n3214 91.65
R61 VN.n5444 VN.n5443 91.65
R62 VN.n4682 VN.n4681 91.65
R63 VN.n6219 VN.n6218 91.65
R64 VN.n6647 VN.n6646 91.65
R65 VN.n8653 VN.n8652 91.65
R66 VN.n7821 VN.n7820 91.65
R67 VN.n10354 VN.n10353 91.65
R68 VN.n9498 VN.n9497 91.65
R69 VN.n13112 VN.n13111 91.389
R70 VN.n12176 VN.n12175 91.389
R71 VN.n11514 VN.n11513 91.389
R72 VN.n10701 VN.n10700 91.389
R73 VN.n9821 VN.n9820 91.389
R74 VN.n8975 VN.n8974 91.389
R75 VN.n8142 VN.n8141 91.389
R76 VN.n7331 VN.n7330 91.389
R77 VN.n6538 VN.n6537 91.389
R78 VN.n5762 VN.n5761 91.389
R79 VN.n4999 VN.n4998 91.389
R80 VN.n4258 VN.n4257 91.389
R81 VN.n3530 VN.n3529 91.389
R82 VN.n2824 VN.n2823 91.389
R83 VN.n2131 VN.n2130 91.389
R84 VN.n1457 VN.n1456 91.389
R85 VN.n804 VN.n803 91.389
R86 VN.n11666 VN.n11665 87.222
R87 VN.n11676 VN.n11675 87.222
R88 VN.n11722 VN.n11721 87.222
R89 VN.n11858 VN.n11857 87.222
R90 VN.n11711 VN.n11710 87.222
R91 VN.n11698 VN.n11697 87.222
R92 VN.n11685 VN.n11684 87.222
R93 VN.n11733 VN.n11732 87.222
R94 VN.n11834 VN.n11833 87.222
R95 VN.n11744 VN.n11743 87.222
R96 VN.n11823 VN.n11822 87.222
R97 VN.n11861 VN.n11860 87.222
R98 VN.n11755 VN.n11754 87.222
R99 VN.n11766 VN.n11765 87.222
R100 VN.n11812 VN.n11811 87.222
R101 VN.n11775 VN.n11774 87.222
R102 VN.n11801 VN.n11800 87.222
R103 VN.n102 VN.n101 86.961
R104 VN.n106 VN.n105 86.961
R105 VN.n110 VN.n109 86.961
R106 VN.n114 VN.n113 86.961
R107 VN.n118 VN.n117 86.961
R108 VN.n122 VN.n121 86.961
R109 VN.n126 VN.n125 86.961
R110 VN.n130 VN.n129 86.961
R111 VN.n134 VN.n133 86.961
R112 VN.n138 VN.n137 86.961
R113 VN.n142 VN.n141 86.961
R114 VN.n146 VN.n145 86.961
R115 VN.n150 VN.n149 86.961
R116 VN.n154 VN.n153 86.961
R117 VN.n158 VN.n157 86.961
R118 VN.n162 VN.n161 86.961
R119 VN.n166 VN.n165 86.961
R120 VN.n11539 VN.t110 50.285
R121 VN.n11371 VN.t20 50.285
R122 VN.n10719 VN.t78 50.285
R123 VN.n10344 VN.t148 50.285
R124 VN.n9859 VN.t350 50.285
R125 VN.n9489 VN.t66 50.285
R126 VN.n9011 VN.t90 50.285
R127 VN.n8643 VN.t45 50.285
R128 VN.n8178 VN.t155 50.285
R129 VN.n7812 VN.t30 50.285
R130 VN.n7367 VN.t22 50.285
R131 VN.n6637 VN.t37 50.285
R132 VN.n6574 VN.t131 50.285
R133 VN.n6208 VN.t6 50.285
R134 VN.n5798 VN.t158 50.285
R135 VN.n5434 VN.t55 50.285
R136 VN.n5035 VN.t47 50.285
R137 VN.n4673 VN.t103 50.285
R138 VN.n4294 VN.t122 50.285
R139 VN.n3932 VN.t269 50.285
R140 VN.n3566 VN.t68 50.285
R141 VN.n3206 VN.t4 50.285
R142 VN.n2860 VN.t167 50.285
R143 VN.n2500 VN.t97 50.285
R144 VN.n2167 VN.t92 50.285
R145 VN.n1809 VN.t16 50.285
R146 VN.n1493 VN.t114 50.285
R147 VN.n1135 VN.t53 50.285
R148 VN.n843 VN.t201 50.285
R149 VN.n483 VN.t257 50.285
R150 VN.n816 VN.t2 50.285
R151 VN.n12690 VN.t88 50.285
R152 VN.n13132 VN.t129 50.285
R153 VN.n12360 VN.t178 50.285
R154 VN.t160 VN.n12172 48.609
R155 VN.t35 VN.n11107 48.609
R156 VN.t106 VN.n11472 48.609
R157 VN.t241 VN.n10634 48.609
R158 VN.t120 VN.n10304 48.609
R159 VN.t0 VN.n9746 48.609
R160 VN.t125 VN.n9421 48.609
R161 VN.t39 VN.n8884 48.609
R162 VN.t26 VN.n8559 48.609
R163 VN.t73 VN.n8035 48.609
R164 VN.t80 VN.n7714 48.609
R165 VN.t253 VN.n6844 48.609
R166 VN.t76 VN.n7325 48.609
R167 VN.t146 VN.n6399 48.609
R168 VN.t10 VN.n6082 48.609
R169 VN.t176 VN.n5607 48.609
R170 VN.t71 VN.n5290 48.609
R171 VN.t32 VN.n4828 48.609
R172 VN.t99 VN.n4515 48.609
R173 VN.t28 VN.n4071 48.609
R174 VN.t14 VN.n3758 48.609
R175 VN.t183 VN.n3327 48.609
R176 VN.t63 VN.n3018 48.609
R177 VN.t57 VN.n2605 48.609
R178 VN.t49 VN.n2296 48.609
R179 VN.t108 VN.n1896 48.609
R180 VN.t224 VN.n1588 48.609
R181 VN.t94 VN.n1206 48.609
R182 VN.t24 VN.n905 48.609
R183 VN.t41 VN.n531 48.609
R184 VN.t12 VN.n234 48.609
R185 VN.t101 VN.n12744 48.609
R186 VN.t236 VN.n12237 48.609
R187 VN.t82 VN.n12412 48.609
R188 VN.t51 VN.n103 48.609
R189 VN.n12172 VN.t43 9.009
R190 VN.n6603 VN.t856 3.904
R191 VN.n7327 VN.n7326 3.904
R192 VN.n11364 VN.t430 3.904
R193 VN.n11664 VN.t1823 3.904
R194 VN.n11574 VN.n11573 3.904
R195 VN.n11577 VN.t1788 3.904
R196 VN.n11569 VN.n11568 3.904
R197 VN.n11547 VN.t464 3.904
R198 VN.n12407 VN.n12406 3.904
R199 VN.n12410 VN.t1965 3.904
R200 VN.n168 VN.t335 3.904
R201 VN.n169 VN.t588 3.904
R202 VN.n13112 VN.t1177 3.904
R203 VN.n13114 VN.t571 3.904
R204 VN.n102 VN.t1459 3.904
R205 VN.n85 VN.t1064 3.904
R206 VN.n11674 VN.t1053 3.904
R207 VN.n12157 VN.n12156 3.904
R208 VN.n12170 VN.t1825 3.904
R209 VN.n12167 VN.t2221 3.904
R210 VN.n12154 VN.n12153 3.904
R211 VN.n12370 VN.t1874 3.904
R212 VN.n12244 VN.n12243 3.904
R213 VN.n12261 VN.t747 3.904
R214 VN.n12264 VN.t2217 3.904
R215 VN.n12241 VN.n12240 3.904
R216 VN.n12709 VN.n12708 3.904
R217 VN.n12718 VN.t1059 3.904
R218 VN.n12715 VN.t1316 3.904
R219 VN.n12706 VN.n12705 3.904
R220 VN.n215 VN.n214 3.904
R221 VN.n232 VN.t145 3.904
R222 VN.n229 VN.t1622 3.904
R223 VN.n212 VN.n211 3.904
R224 VN.n520 VN.n519 3.904
R225 VN.n529 VN.t615 3.904
R226 VN.n526 VN.t722 3.904
R227 VN.n517 VN.n516 3.904
R228 VN.n886 VN.n885 3.904
R229 VN.n903 VN.t2117 3.904
R230 VN.n900 VN.t1172 3.904
R231 VN.n883 VN.n882 3.904
R232 VN.n1195 VN.n1194 3.904
R233 VN.n1204 VN.t2542 3.904
R234 VN.n1201 VN.t115 3.904
R235 VN.n1192 VN.n1191 3.904
R236 VN.n1569 VN.n1568 3.904
R237 VN.n1586 VN.t1525 3.904
R238 VN.n1583 VN.t17 3.904
R239 VN.n1566 VN.n1565 3.904
R240 VN.n1885 VN.n1884 3.904
R241 VN.n1894 VN.t1476 3.904
R242 VN.n1891 VN.t1585 3.904
R243 VN.n1882 VN.n1881 3.904
R244 VN.n2277 VN.n2276 3.904
R245 VN.n2294 VN.t465 3.904
R246 VN.n2291 VN.t842 3.904
R247 VN.n2274 VN.n2273 3.904
R248 VN.n2594 VN.n2593 3.904
R249 VN.n2603 VN.t2248 3.904
R250 VN.n2600 VN.t2355 3.904
R251 VN.n2591 VN.n2590 3.904
R252 VN.n2999 VN.n2998 3.904
R253 VN.n3016 VN.t1498 3.904
R254 VN.n3013 VN.t277 3.904
R255 VN.n2996 VN.n2995 3.904
R256 VN.n3316 VN.n3315 3.904
R257 VN.n3325 VN.t1657 3.904
R258 VN.n3322 VN.t2060 3.904
R259 VN.n3313 VN.n3312 3.904
R260 VN.n3739 VN.n3738 3.904
R261 VN.n3756 VN.t899 3.904
R262 VN.n3753 VN.t2222 3.904
R263 VN.n3736 VN.n3735 3.904
R264 VN.n4060 VN.n4059 3.904
R265 VN.n4069 VN.t1071 3.904
R266 VN.n4066 VN.t1475 3.904
R267 VN.n4057 VN.n4056 3.904
R268 VN.n4496 VN.n4495 3.904
R269 VN.n4513 VN.t477 3.904
R270 VN.n4510 VN.t1629 3.904
R271 VN.n4493 VN.n4492 3.904
R272 VN.n4817 VN.n4816 3.904
R273 VN.n4826 VN.t510 3.904
R274 VN.n4823 VN.t1003 3.904
R275 VN.n4814 VN.n4813 3.904
R276 VN.n5271 VN.n5270 3.904
R277 VN.n5288 VN.t2405 3.904
R278 VN.n5285 VN.t1037 3.904
R279 VN.n5268 VN.n5267 3.904
R280 VN.n5596 VN.n5595 3.904
R281 VN.n5605 VN.t2429 3.904
R282 VN.n5602 VN.t453 3.904
R283 VN.n5593 VN.n5592 3.904
R284 VN.n6063 VN.n6062 3.904
R285 VN.n6080 VN.t1809 3.904
R286 VN.n6077 VN.t483 3.904
R287 VN.n6060 VN.n6059 3.904
R288 VN.n6388 VN.n6387 3.904
R289 VN.n6397 VN.t2151 3.904
R290 VN.n6394 VN.t2374 3.904
R291 VN.n6385 VN.n6384 3.904
R292 VN.n7306 VN.n7305 3.904
R293 VN.n7323 VN.t1239 3.904
R294 VN.n7320 VN.t150 3.904
R295 VN.n7303 VN.n7302 3.904
R296 VN.n6833 VN.n6832 3.904
R297 VN.n6842 VN.t1557 3.904
R298 VN.n6839 VN.t1780 3.904
R299 VN.n6830 VN.n6829 3.904
R300 VN.n7695 VN.n7694 3.904
R301 VN.n7712 VN.t654 3.904
R302 VN.n7709 VN.t2125 3.904
R303 VN.n7692 VN.n7691 3.904
R304 VN.n8024 VN.n8023 3.904
R305 VN.n8033 VN.t1095 3.904
R306 VN.n8030 VN.t1211 3.904
R307 VN.n8021 VN.n8020 3.904
R308 VN.n8540 VN.n8539 3.904
R309 VN.n8557 VN.t2586 3.904
R310 VN.n8554 VN.t580 3.904
R311 VN.n8537 VN.n8536 3.904
R312 VN.n8873 VN.n8872 3.904
R313 VN.n8882 VN.t1958 3.904
R314 VN.n8879 VN.t2081 3.904
R315 VN.n8870 VN.n8869 3.904
R316 VN.n9402 VN.n9401 3.904
R317 VN.n9419 VN.t915 3.904
R318 VN.n9416 VN.t2293 3.904
R319 VN.n9399 VN.n9398 3.904
R320 VN.n9735 VN.n9734 3.904
R321 VN.n9744 VN.t1136 3.904
R322 VN.n9741 VN.t1376 3.904
R323 VN.n9732 VN.n9731 3.904
R324 VN.n10285 VN.n10284 3.904
R325 VN.n10302 VN.t207 3.904
R326 VN.n10299 VN.t2262 3.904
R327 VN.n10282 VN.n10281 3.904
R328 VN.n10622 VN.n10621 3.904
R329 VN.n10632 VN.t1109 3.904
R330 VN.n10629 VN.t1352 3.904
R331 VN.n10619 VN.n10618 3.904
R332 VN.n11454 VN.n11453 3.904
R333 VN.n11470 VN.t1846 3.904
R334 VN.n11467 VN.t2242 3.904
R335 VN.n11451 VN.n11450 3.904
R336 VN.n11114 VN.n11113 3.904
R337 VN.n11120 VN.t1087 3.904
R338 VN.n11123 VN.t473 3.904
R339 VN.n11111 VN.n11110 3.904
R340 VN.n11720 VN.t1461 3.904
R341 VN.n12030 VN.n12029 3.904
R342 VN.n12041 VN.t1303 3.904
R343 VN.n12038 VN.t2456 3.904
R344 VN.n12033 VN.n12032 3.904
R345 VN.n2511 VN.t304 3.904
R346 VN.n3025 VN.n3024 3.904
R347 VN.n3041 VN.t1963 3.904
R348 VN.n3044 VN.t622 3.904
R349 VN.n3022 VN.n3021 3.904
R350 VN.n3224 VN.n3223 3.904
R351 VN.n3233 VN.t2004 3.904
R352 VN.n3230 VN.t2515 3.904
R353 VN.n3221 VN.n3220 3.904
R354 VN.n3588 VN.n3587 3.904
R355 VN.n3605 VN.t1393 3.904
R356 VN.n3602 VN.t2549 3.904
R357 VN.n3585 VN.n3584 3.904
R358 VN.n3968 VN.n3967 3.904
R359 VN.n3977 VN.t1549 3.904
R360 VN.n3974 VN.t1940 3.904
R361 VN.n3965 VN.n3964 3.904
R362 VN.n4345 VN.n4344 3.904
R363 VN.n4362 VN.t799 3.904
R364 VN.n4359 VN.t2115 3.904
R365 VN.n4342 VN.n4341 3.904
R366 VN.n4725 VN.n4724 3.904
R367 VN.n4734 VN.t950 3.904
R368 VN.n4731 VN.t1371 3.904
R369 VN.n4722 VN.n4721 3.904
R370 VN.n5120 VN.n5119 3.904
R371 VN.n5137 VN.t217 3.904
R372 VN.n5134 VN.t1522 3.904
R373 VN.n5117 VN.n5116 3.904
R374 VN.n5504 VN.n5503 3.904
R375 VN.n5513 VN.t394 3.904
R376 VN.n5510 VN.t777 3.904
R377 VN.n5501 VN.n5500 3.904
R378 VN.n5912 VN.n5911 3.904
R379 VN.n5929 VN.t2175 3.904
R380 VN.n5926 VN.t2292 3.904
R381 VN.n5909 VN.n5908 3.904
R382 VN.n6296 VN.n6295 3.904
R383 VN.n6305 VN.t1434 3.904
R384 VN.n6302 VN.t1543 3.904
R385 VN.n6293 VN.n6292 3.904
R386 VN.n7155 VN.n7154 3.904
R387 VN.n7172 VN.t418 3.904
R388 VN.n7169 VN.t1986 3.904
R389 VN.n7152 VN.n7151 3.904
R390 VN.n6741 VN.n6740 3.904
R391 VN.n6750 VN.t837 3.904
R392 VN.n6747 VN.t946 3.904
R393 VN.n6738 VN.n6737 3.904
R394 VN.n7544 VN.n7543 3.904
R395 VN.n7561 VN.t2349 3.904
R396 VN.n7558 VN.t1409 3.904
R397 VN.n7541 VN.n7540 3.904
R398 VN.n7932 VN.n7931 3.904
R399 VN.n7941 VN.t268 3.904
R400 VN.n7938 VN.t388 3.904
R401 VN.n7929 VN.n7928 3.904
R402 VN.n8389 VN.n8388 3.904
R403 VN.n8406 VN.t1879 3.904
R404 VN.n8403 VN.t2269 3.904
R405 VN.n8386 VN.n8385 3.904
R406 VN.n8781 VN.n8780 3.904
R407 VN.n8790 VN.t1123 3.904
R408 VN.n8787 VN.t1378 3.904
R409 VN.n8778 VN.n8777 3.904
R410 VN.n9251 VN.n9250 3.904
R411 VN.n9268 VN.t223 3.904
R412 VN.n9265 VN.t1679 3.904
R413 VN.n9248 VN.n9247 3.904
R414 VN.n9643 VN.n9642 3.904
R415 VN.n9652 VN.t556 3.904
R416 VN.n9649 VN.t782 3.904
R417 VN.n9640 VN.n9639 3.904
R418 VN.n10133 VN.n10132 3.904
R419 VN.n10150 VN.t2181 3.904
R420 VN.n10147 VN.t1101 3.904
R421 VN.n10130 VN.n10129 3.904
R422 VN.n10520 VN.n10519 3.904
R423 VN.n10530 VN.t2483 3.904
R424 VN.n10527 VN.t187 3.904
R425 VN.n10517 VN.n10516 3.904
R426 VN.n11002 VN.n11001 3.904
R427 VN.n11014 VN.t1862 3.904
R428 VN.n11011 VN.t533 3.904
R429 VN.n10999 VN.n10998 3.904
R430 VN.n11184 VN.n11183 3.904
R431 VN.n11190 VN.t1894 3.904
R432 VN.n11193 VN.t2422 3.904
R433 VN.n11181 VN.n11180 3.904
R434 VN.n11856 VN.t590 3.904
R435 VN.n12053 VN.n12052 3.904
R436 VN.n12064 VN.t439 3.904
R437 VN.n12061 VN.t1710 3.904
R438 VN.n12056 VN.n12055 3.904
R439 VN.n1819 VN.t2527 3.904
R440 VN.n2307 VN.n2306 3.904
R441 VN.n2322 VN.t1404 3.904
R442 VN.n2325 VN.t338 3.904
R443 VN.n2310 VN.n2309 3.904
R444 VN.n2517 VN.n2516 3.904
R445 VN.n2528 VN.t1704 3.904
R446 VN.n2525 VN.t1951 3.904
R447 VN.n2520 VN.n2519 3.904
R448 VN.n2874 VN.n2873 3.904
R449 VN.n2894 VN.t1096 3.904
R450 VN.n2891 VN.t2273 3.904
R451 VN.n2877 VN.n2876 3.904
R452 VN.n3239 VN.n3238 3.904
R453 VN.n3250 VN.t1273 3.904
R454 VN.n3247 VN.t1655 3.904
R455 VN.n3242 VN.n3241 3.904
R456 VN.n3614 VN.n3613 3.904
R457 VN.n3634 VN.t530 3.904
R458 VN.n3631 VN.t1808 3.904
R459 VN.n3617 VN.n3616 3.904
R460 VN.n3983 VN.n3982 3.904
R461 VN.n3994 VN.t676 3.904
R462 VN.n3991 VN.t1067 3.904
R463 VN.n3986 VN.n3985 3.904
R464 VN.n4371 VN.n4370 3.904
R465 VN.n4391 VN.t2454 3.904
R466 VN.n4388 VN.t1237 3.904
R467 VN.n4374 VN.n4373 3.904
R468 VN.n4740 VN.n4739 3.904
R469 VN.n4751 VN.t33 3.904
R470 VN.n4748 VN.t506 3.904
R471 VN.n4743 VN.n4742 3.904
R472 VN.n5146 VN.n5145 3.904
R473 VN.n5166 VN.t1868 3.904
R474 VN.n5163 VN.t2001 3.904
R475 VN.n5149 VN.n5148 3.904
R476 VN.n5519 VN.n5518 3.904
R477 VN.n5530 VN.t849 3.904
R478 VN.n5527 VN.t1269 3.904
R479 VN.n5522 VN.n5521 3.904
R480 VN.n5938 VN.n5937 3.904
R481 VN.n5958 VN.t75 3.904
R482 VN.n5955 VN.t1423 3.904
R483 VN.n5941 VN.n5940 3.904
R484 VN.n6311 VN.n6310 3.904
R485 VN.n6322 VN.t568 3.904
R486 VN.n6319 VN.t674 3.904
R487 VN.n6314 VN.n6313 3.904
R488 VN.n7181 VN.n7180 3.904
R489 VN.n7201 VN.t2067 3.904
R490 VN.n7198 VN.t1112 3.904
R491 VN.n7184 VN.n7183 3.904
R492 VN.n6756 VN.n6755 3.904
R493 VN.n6767 VN.t2500 3.904
R494 VN.n6764 VN.t23 3.904
R495 VN.n6759 VN.n6758 3.904
R496 VN.n7570 VN.n7569 3.904
R497 VN.n7590 VN.t1601 3.904
R498 VN.n7587 VN.t549 3.904
R499 VN.n7573 VN.n7572 3.904
R500 VN.n7947 VN.n7946 3.904
R501 VN.n7958 VN.t1919 3.904
R502 VN.n7955 VN.t2173 3.904
R503 VN.n7950 VN.n7949 3.904
R504 VN.n8415 VN.n8414 3.904
R505 VN.n8435 VN.t1011 3.904
R506 VN.n8432 VN.t1405 3.904
R507 VN.n8418 VN.n8417 3.904
R508 VN.n8796 VN.n8795 3.904
R509 VN.n8807 VN.t260 3.904
R510 VN.n8804 VN.t513 3.904
R511 VN.n8799 VN.n8798 3.904
R512 VN.n9277 VN.n9276 3.904
R513 VN.n9297 VN.t1872 3.904
R514 VN.n9294 VN.t812 3.904
R515 VN.n9280 VN.n9279 3.904
R516 VN.n9658 VN.n9657 3.904
R517 VN.n9669 VN.t2214 3.904
R518 VN.n9666 VN.t2433 3.904
R519 VN.n9661 VN.n9660 3.904
R520 VN.n10159 VN.n10158 3.904
R521 VN.n10179 VN.t1313 3.904
R522 VN.n10176 VN.t234 3.904
R523 VN.n10162 VN.n10161 3.904
R524 VN.n10536 VN.n10535 3.904
R525 VN.n10550 VN.t1619 3.904
R526 VN.n10547 VN.t1845 3.904
R527 VN.n10539 VN.n10538 3.904
R528 VN.n10557 VN.n10556 3.904
R529 VN.n10571 VN.t859 3.904
R530 VN.n10568 VN.t973 3.904
R531 VN.n10560 VN.n10559 3.904
R532 VN.n11050 VN.n11049 3.904
R533 VN.n11074 VN.t107 3.904
R534 VN.n11071 VN.t1436 3.904
R535 VN.n11053 VN.n11052 3.904
R536 VN.n11148 VN.n11147 3.904
R537 VN.n11156 VN.t297 3.904
R538 VN.n11159 VN.t690 3.904
R539 VN.n11151 VN.n11150 3.904
R540 VN.n12070 VN.n12069 3.904
R541 VN.n12086 VN.t2084 3.904
R542 VN.n12083 VN.t2297 3.904
R543 VN.n12073 VN.n12072 3.904
R544 VN.n11709 VN.t1142 3.904
R545 VN.n10197 VN.n10196 3.904
R546 VN.n10214 VN.t452 3.904
R547 VN.n10211 VN.t1881 3.904
R548 VN.n10194 VN.n10193 3.904
R549 VN.n9314 VN.n9313 3.904
R550 VN.n9331 VN.t1002 3.904
R551 VN.n9328 VN.t2468 3.904
R552 VN.n9311 VN.n9310 3.904
R553 VN.n8452 VN.n8451 3.904
R554 VN.n8469 VN.t138 3.904
R555 VN.n8466 VN.t543 3.904
R556 VN.n8449 VN.n8448 3.904
R557 VN.n7607 VN.n7606 3.904
R558 VN.n7624 VN.t736 3.904
R559 VN.n7621 VN.t2204 3.904
R560 VN.n7604 VN.n7603 3.904
R561 VN.n7218 VN.n7217 3.904
R562 VN.n7235 VN.t1328 3.904
R563 VN.n7232 VN.t248 3.904
R564 VN.n7215 VN.n7214 3.904
R565 VN.n5975 VN.n5974 3.904
R566 VN.n5992 VN.t1762 3.904
R567 VN.n5989 VN.t558 3.904
R568 VN.n5972 VN.n5971 3.904
R569 VN.n5183 VN.n5182 3.904
R570 VN.n5200 VN.t2359 3.904
R571 VN.n5197 VN.t1126 3.904
R572 VN.n5180 VN.n5179 3.904
R573 VN.n4408 VN.n4407 3.904
R574 VN.n4425 VN.t1590 3.904
R575 VN.n4422 VN.t1701 3.904
R576 VN.n4405 VN.n4404 3.904
R577 VN.n3651 VN.n3650 3.904
R578 VN.n3668 VN.t2185 3.904
R579 VN.n3665 VN.t932 3.904
R580 VN.n3648 VN.n3647 3.904
R581 VN.n2911 VN.n2910 3.904
R582 VN.n2928 VN.t228 3.904
R583 VN.n2925 VN.t1535 3.904
R584 VN.n2908 VN.n2907 3.904
R585 VN.n2189 VN.n2188 3.904
R586 VN.n2206 VN.t542 3.904
R587 VN.n2203 VN.t1981 3.904
R588 VN.n2186 VN.n2185 3.904
R589 VN.n1598 VN.n1597 3.904
R590 VN.n1614 VN.t1604 3.904
R591 VN.n1617 VN.t2560 3.904
R592 VN.n1595 VN.n1594 3.904
R593 VN.n1146 VN.t215 3.904
R594 VN.n1827 VN.n1826 3.904
R595 VN.n1836 VN.t1431 3.904
R596 VN.n1833 VN.t1663 3.904
R597 VN.n1824 VN.n1823 3.904
R598 VN.n2536 VN.n2535 3.904
R599 VN.n2545 VN.t964 3.904
R600 VN.n2542 VN.t1082 3.904
R601 VN.n2533 VN.n2532 3.904
R602 VN.n3258 VN.n3257 3.904
R603 VN.n3267 VN.t403 3.904
R604 VN.n3264 VN.t786 3.904
R605 VN.n3255 VN.n3254 3.904
R606 VN.n4002 VN.n4001 3.904
R607 VN.n4011 VN.t2337 3.904
R608 VN.n4008 VN.t193 3.904
R609 VN.n3999 VN.n3998 3.904
R610 VN.n4759 VN.n4758 3.904
R611 VN.n4768 VN.t581 3.904
R612 VN.n4765 VN.t957 3.904
R613 VN.n4756 VN.n4755 3.904
R614 VN.n5538 VN.n5537 3.904
R615 VN.n5547 VN.t2513 3.904
R616 VN.n5544 VN.t401 3.904
R617 VN.n5535 VN.n5534 3.904
R618 VN.n6330 VN.n6329 3.904
R619 VN.n6339 VN.t2227 3.904
R620 VN.n6336 VN.t2333 3.904
R621 VN.n6327 VN.n6326 3.904
R622 VN.n6775 VN.n6774 3.904
R623 VN.n6784 VN.t1637 3.904
R624 VN.n6781 VN.t1864 3.904
R625 VN.n6772 VN.n6771 3.904
R626 VN.n7966 VN.n7965 3.904
R627 VN.n7975 VN.t1044 3.904
R628 VN.n7972 VN.t1306 3.904
R629 VN.n7963 VN.n7962 3.904
R630 VN.n8815 VN.n8814 3.904
R631 VN.n8824 VN.t1909 3.904
R632 VN.n8821 VN.t2166 3.904
R633 VN.n8812 VN.n8811 3.904
R634 VN.n9677 VN.n9676 3.904
R635 VN.n9686 VN.t1346 3.904
R636 VN.n9683 VN.t1573 3.904
R637 VN.n9674 VN.n9673 3.904
R638 VN.n11401 VN.n11400 3.904
R639 VN.n11419 VN.t1777 3.904
R640 VN.n11416 VN.t1456 3.904
R641 VN.n11404 VN.n11403 3.904
R642 VN.n11089 VN.n11088 3.904
R643 VN.n11384 VN.t306 3.904
R644 VN.n11387 VN.t2205 3.904
R645 VN.n11390 VN.n11389 3.904
R646 VN.n12104 VN.n12103 3.904
R647 VN.n12120 VN.t1031 3.904
R648 VN.n12117 VN.t1426 3.904
R649 VN.n12107 VN.n12106 3.904
R650 VN.n11696 VN.t278 3.904
R651 VN.n493 VN.t2451 3.904
R652 VN.n919 VN.n918 3.904
R653 VN.n927 VN.t1330 3.904
R654 VN.n930 VN.t251 3.904
R655 VN.n916 VN.n915 3.904
R656 VN.n1160 VN.n1159 3.904
R657 VN.n1168 VN.t1639 3.904
R658 VN.n1165 VN.t1865 3.904
R659 VN.n1157 VN.n1156 3.904
R660 VN.n1513 VN.n1512 3.904
R661 VN.n1531 VN.t737 3.904
R662 VN.n1528 VN.t1690 3.904
R663 VN.n1510 VN.n1509 3.904
R664 VN.n1850 VN.n1849 3.904
R665 VN.n1858 VN.t687 3.904
R666 VN.n1855 VN.t795 3.904
R667 VN.n1847 VN.n1846 3.904
R668 VN.n2221 VN.n2220 3.904
R669 VN.n2239 VN.t2197 3.904
R670 VN.n2236 VN.t1252 3.904
R671 VN.n2218 VN.n2217 3.904
R672 VN.n2559 VN.n2558 3.904
R673 VN.n2567 VN.t58 3.904
R674 VN.n2564 VN.t210 3.904
R675 VN.n2556 VN.n2555 3.904
R676 VN.n2943 VN.n2942 3.904
R677 VN.n2961 VN.t1878 3.904
R678 VN.n2958 VN.t663 3.904
R679 VN.n2940 VN.n2939 3.904
R680 VN.n3281 VN.n3280 3.904
R681 VN.n3289 VN.t2052 3.904
R682 VN.n3286 VN.t2438 3.904
R683 VN.n3278 VN.n3277 3.904
R684 VN.n3683 VN.n3682 3.904
R685 VN.n3701 VN.t1318 3.904
R686 VN.n3698 VN.t1429 3.904
R687 VN.n3680 VN.n3679 3.904
R688 VN.n4025 VN.n4024 3.904
R689 VN.n4033 VN.t290 3.904
R690 VN.n4030 VN.t683 3.904
R691 VN.n4022 VN.n4021 3.904
R692 VN.n4440 VN.n4439 3.904
R693 VN.n4458 VN.t2078 3.904
R694 VN.n4455 VN.t830 3.904
R695 VN.n4437 VN.n4436 3.904
R696 VN.n4782 VN.n4781 3.904
R697 VN.n4790 VN.t2238 3.904
R698 VN.n4787 VN.t48 3.904
R699 VN.n4779 VN.n4778 3.904
R700 VN.n5215 VN.n5214 3.904
R701 VN.n5233 VN.t1492 3.904
R702 VN.n5230 VN.t262 3.904
R703 VN.n5212 VN.n5211 3.904
R704 VN.n5561 VN.n5560 3.904
R705 VN.n5569 VN.t1650 3.904
R706 VN.n5566 VN.t2049 3.904
R707 VN.n5558 VN.n5557 3.904
R708 VN.n6007 VN.n6006 3.904
R709 VN.n6025 VN.t1017 3.904
R710 VN.n6022 VN.t2215 3.904
R711 VN.n6004 VN.n6003 3.904
R712 VN.n6353 VN.n6352 3.904
R713 VN.n6361 VN.t1361 3.904
R714 VN.n6358 VN.t1586 3.904
R715 VN.n6350 VN.n6349 3.904
R716 VN.n7250 VN.n7249 3.904
R717 VN.n7268 VN.t466 3.904
R718 VN.n7265 VN.t1897 3.904
R719 VN.n7247 VN.n7246 3.904
R720 VN.n6798 VN.n6797 3.904
R721 VN.n6806 VN.t765 3.904
R722 VN.n6803 VN.t994 3.904
R723 VN.n6795 VN.n6794 3.904
R724 VN.n7639 VN.n7638 3.904
R725 VN.n7657 VN.t2392 3.904
R726 VN.n7654 VN.t1336 3.904
R727 VN.n7636 VN.n7635 3.904
R728 VN.n7989 VN.n7988 3.904
R729 VN.n7997 VN.t175 3.904
R730 VN.n7994 VN.t442 3.904
R731 VN.n7986 VN.n7985 3.904
R732 VN.n8484 VN.n8483 3.904
R733 VN.n8502 VN.t1801 3.904
R734 VN.n8499 VN.t2199 3.904
R735 VN.n8481 VN.n8480 3.904
R736 VN.n8838 VN.n8837 3.904
R737 VN.n8846 VN.t1034 3.904
R738 VN.n8843 VN.t1300 3.904
R739 VN.n8835 VN.n8834 3.904
R740 VN.n9346 VN.n9345 3.904
R741 VN.n9364 VN.t126 3.904
R742 VN.n9361 VN.t1602 3.904
R743 VN.n9343 VN.n9342 3.904
R744 VN.n9700 VN.n9699 3.904
R745 VN.n9708 VN.t596 3.904
R746 VN.n9705 VN.t703 3.904
R747 VN.n9697 VN.n9696 3.904
R748 VN.n10229 VN.n10228 3.904
R749 VN.n10247 VN.t2098 3.904
R750 VN.n10244 VN.t1147 3.904
R751 VN.n10226 VN.n10225 3.904
R752 VN.n10585 VN.n10584 3.904
R753 VN.n10593 VN.t2521 3.904
R754 VN.n10590 VN.t79 3.904
R755 VN.n10582 VN.n10581 3.904
R756 VN.n11428 VN.n11427 3.904
R757 VN.n11446 VN.t188 3.904
R758 VN.n11443 VN.t586 3.904
R759 VN.n11431 VN.n11430 3.904
R760 VN.n11129 VN.n11128 3.904
R761 VN.n11140 VN.t1955 3.904
R762 VN.n11143 VN.t1337 3.904
R763 VN.n11132 VN.n11131 3.904
R764 VN.n10605 VN.n10604 3.904
R765 VN.n10614 VN.t1976 3.904
R766 VN.n10611 VN.t2220 3.904
R767 VN.n10602 VN.n10601 3.904
R768 VN.n10256 VN.n10255 3.904
R769 VN.n10268 VN.t1221 3.904
R770 VN.n10265 VN.t608 3.904
R771 VN.n10259 VN.n10258 3.904
R772 VN.n9714 VN.n9713 3.904
R773 VN.n9727 VN.t2251 3.904
R774 VN.n9724 VN.t2362 3.904
R775 VN.n9717 VN.n9716 3.904
R776 VN.n9373 VN.n9372 3.904
R777 VN.n9385 VN.t1790 3.904
R778 VN.n9382 VN.t848 3.904
R779 VN.n9376 VN.n9375 3.904
R780 VN.n8852 VN.n8851 3.904
R781 VN.n8865 VN.t309 3.904
R782 VN.n8862 VN.t434 3.904
R783 VN.n8855 VN.n8854 3.904
R784 VN.n8511 VN.n8510 3.904
R785 VN.n8523 VN.t924 3.904
R786 VN.n8520 VN.t1327 3.904
R787 VN.n8514 VN.n8513 3.904
R788 VN.n8003 VN.n8002 3.904
R789 VN.n8016 VN.t1837 3.904
R790 VN.n8013 VN.t2087 3.904
R791 VN.n8006 VN.n8005 3.904
R792 VN.n7666 VN.n7665 3.904
R793 VN.n7678 VN.t1524 3.904
R794 VN.n7675 VN.t472 3.904
R795 VN.n7669 VN.n7668 3.904
R796 VN.n6812 VN.n6811 3.904
R797 VN.n6825 VN.t2419 3.904
R798 VN.n6822 VN.t112 3.904
R799 VN.n6815 VN.n6814 3.904
R800 VN.n7277 VN.n7276 3.904
R801 VN.n7289 VN.t2116 3.904
R802 VN.n7286 VN.t1022 3.904
R803 VN.n7280 VN.n7279 3.904
R804 VN.n6367 VN.n6366 3.904
R805 VN.n6380 VN.t494 3.904
R806 VN.n6377 VN.t721 3.904
R807 VN.n6370 VN.n6369 3.904
R808 VN.n6034 VN.n6033 3.904
R809 VN.n6046 VN.t144 3.904
R810 VN.n6043 VN.t1348 3.904
R811 VN.n6037 VN.n6036 3.904
R812 VN.n5575 VN.n5574 3.904
R813 VN.n5588 VN.t780 3.904
R814 VN.n5585 VN.t1314 3.904
R815 VN.n5578 VN.n5577 3.904
R816 VN.n5242 VN.n5241 3.904
R817 VN.n5254 VN.t746 3.904
R818 VN.n5251 VN.t1912 3.904
R819 VN.n5245 VN.n5244 3.904
R820 VN.n4796 VN.n4795 3.904
R821 VN.n4809 VN.t1373 3.904
R822 VN.n4806 VN.t1745 3.904
R823 VN.n4799 VN.n4798 3.904
R824 VN.n4467 VN.n4466 3.904
R825 VN.n4479 VN.t1206 3.904
R826 VN.n4476 VN.t2493 3.904
R827 VN.n4470 VN.n4469 3.904
R828 VN.n4039 VN.n4038 3.904
R829 VN.n4052 VN.t1942 3.904
R830 VN.n4049 VN.t2343 3.904
R831 VN.n4042 VN.n4041 3.904
R832 VN.n3710 VN.n3709 3.904
R833 VN.n3722 VN.t1771 3.904
R834 VN.n3719 VN.t563 3.904
R835 VN.n3713 VN.n3712 3.904
R836 VN.n3295 VN.n3294 3.904
R837 VN.n3308 VN.t2517 3.904
R838 VN.n3305 VN.t411 3.904
R839 VN.n3298 VN.n3297 3.904
R840 VN.n2970 VN.n2969 3.904
R841 VN.n2982 VN.t1009 3.904
R842 VN.n2979 VN.t1140 3.904
R843 VN.n2973 VN.n2972 3.904
R844 VN.n2573 VN.n2572 3.904
R845 VN.n2586 VN.t1750 3.904
R846 VN.n2583 VN.t1861 3.904
R847 VN.n2576 VN.n2575 3.904
R848 VN.n2248 VN.n2247 3.904
R849 VN.n2260 VN.t1326 3.904
R850 VN.n2257 VN.t383 3.904
R851 VN.n2251 VN.n2250 3.904
R852 VN.n1864 VN.n1863 3.904
R853 VN.n1877 VN.t2345 3.904
R854 VN.n1874 VN.t2449 3.904
R855 VN.n1867 VN.n1866 3.904
R856 VN.n1543 VN.n1542 3.904
R857 VN.n1552 VN.t2393 3.904
R858 VN.n1534 VN.t942 3.904
R859 VN.n1546 VN.n1545 3.904
R860 VN.n1174 VN.n1173 3.904
R861 VN.n1187 VN.t882 3.904
R862 VN.n1184 VN.t995 3.904
R863 VN.n1177 VN.n1176 3.904
R864 VN.n857 VN.n856 3.904
R865 VN.n869 VN.t467 3.904
R866 VN.n866 VN.t1901 3.904
R867 VN.n860 VN.n859 3.904
R868 VN.n499 VN.n498 3.904
R869 VN.n512 VN.t1363 3.904
R870 VN.n509 VN.t1587 3.904
R871 VN.n502 VN.n501 3.904
R872 VN.n246 VN.n245 3.904
R873 VN.n255 VN.t1018 3.904
R874 VN.n258 VN.t2486 3.904
R875 VN.n249 VN.n248 3.904
R876 VN.n12701 VN.t2182 3.904
R877 VN.n11683 VN.t1928 3.904
R878 VN.n12130 VN.n12129 3.904
R879 VN.n12149 VN.t161 3.904
R880 VN.n12146 VN.t561 3.904
R881 VN.n12133 VN.n12132 3.904
R882 VN.n11023 VN.n11022 3.904
R883 VN.n11041 VN.t992 3.904
R884 VN.n11038 VN.t2187 3.904
R885 VN.n11026 VN.n11025 3.904
R886 VN.n11166 VN.n11165 3.904
R887 VN.n11174 VN.t1166 3.904
R888 VN.n11177 VN.t1560 3.904
R889 VN.n11169 VN.n11168 3.904
R890 VN.n11731 VN.t547 3.904
R891 VN.n11985 VN.n11984 3.904
R892 VN.n11996 VN.t519 3.904
R893 VN.n11993 VN.t1668 3.904
R894 VN.n11988 VN.n11987 3.904
R895 VN.n3943 VN.t1154 3.904
R896 VN.n4522 VN.n4521 3.904
R897 VN.n4538 VN.t2529 3.904
R898 VN.n4541 VN.t1195 3.904
R899 VN.n4519 VN.n4518 3.904
R900 VN.n4691 VN.n4690 3.904
R901 VN.n4700 VN.t2565 3.904
R902 VN.n4697 VN.t578 3.904
R903 VN.n4688 VN.n4687 3.904
R904 VN.n5057 VN.n5056 3.904
R905 VN.n5074 VN.t1957 3.904
R906 VN.n5071 VN.t612 3.904
R907 VN.n5054 VN.n5053 3.904
R908 VN.n5470 VN.n5469 3.904
R909 VN.n5479 VN.t2136 3.904
R910 VN.n5476 VN.t2510 3.904
R911 VN.n5467 VN.n5466 3.904
R912 VN.n5849 VN.n5848 3.904
R913 VN.n5866 VN.t1388 3.904
R914 VN.n5863 VN.t137 3.904
R915 VN.n5846 VN.n5845 3.904
R916 VN.n6262 VN.n6261 3.904
R917 VN.n6271 VN.t1811 3.904
R918 VN.n6268 VN.t1931 3.904
R919 VN.n6259 VN.n6258 3.904
R920 VN.n7092 VN.n7091 3.904
R921 VN.n7109 VN.t790 3.904
R922 VN.n7106 VN.t2378 3.904
R923 VN.n7089 VN.n7088 3.904
R924 VN.n6707 VN.n6706 3.904
R925 VN.n6716 VN.t1243 3.904
R926 VN.n6713 VN.t1360 3.904
R927 VN.n6704 VN.n6703 3.904
R928 VN.n7481 VN.n7480 3.904
R929 VN.n7498 VN.t199 3.904
R930 VN.n7495 VN.t626 3.904
R931 VN.n7478 VN.n7477 3.904
R932 VN.n7898 VN.n7897 3.904
R933 VN.n7907 VN.t2005 3.904
R934 VN.n7904 VN.t2132 3.904
R935 VN.n7895 VN.n7894 3.904
R936 VN.n8326 VN.n8325 3.904
R937 VN.n8343 VN.t965 3.904
R938 VN.n8340 VN.t1484 3.904
R939 VN.n8323 VN.n8322 3.904
R940 VN.n8747 VN.n8746 3.904
R941 VN.n8756 VN.t352 3.904
R942 VN.n8753 VN.t470 3.904
R943 VN.n8744 VN.n8743 3.904
R944 VN.n9188 VN.n9187 3.904
R945 VN.n9205 VN.t1832 3.904
R946 VN.n9202 VN.t884 3.904
R947 VN.n9185 VN.n9184 3.904
R948 VN.n9609 VN.n9608 3.904
R949 VN.n9618 VN.t2288 3.904
R950 VN.n9615 VN.t2399 3.904
R951 VN.n9606 VN.n9605 3.904
R952 VN.n10070 VN.n10069 3.904
R953 VN.n10087 VN.t1392 3.904
R954 VN.n10084 VN.t319 3.904
R955 VN.n10067 VN.n10066 3.904
R956 VN.n10485 VN.n10484 3.904
R957 VN.n10495 VN.t1693 3.904
R958 VN.n10492 VN.t1934 3.904
R959 VN.n10482 VN.n10481 3.904
R960 VN.n10944 VN.n10943 3.904
R961 VN.n10956 VN.t1083 3.904
R962 VN.n10953 VN.t2260 3.904
R963 VN.n10941 VN.n10940 3.904
R964 VN.n11218 VN.n11217 3.904
R965 VN.n11224 VN.t1111 3.904
R966 VN.n11227 VN.t1642 3.904
R967 VN.n11215 VN.n11214 3.904
R968 VN.n11832 VN.t2202 3.904
R969 VN.n12008 VN.n12007 3.904
R970 VN.n12019 VN.t2170 3.904
R971 VN.n12016 VN.t803 3.904
R972 VN.n12011 VN.n12010 3.904
R973 VN.n3216 VN.t853 3.904
R974 VN.n3769 VN.n3768 3.904
R975 VN.n3784 VN.t2259 3.904
R976 VN.n3787 VN.t888 3.904
R977 VN.n3772 VN.n3771 3.904
R978 VN.n3949 VN.n3948 3.904
R979 VN.n3960 VN.t2296 3.904
R980 VN.n3957 VN.t288 3.904
R981 VN.n3952 VN.n3951 3.904
R982 VN.n4308 VN.n4307 3.904
R983 VN.n4328 VN.t1665 3.904
R984 VN.n4325 VN.t326 3.904
R985 VN.n4311 VN.n4310 3.904
R986 VN.n4706 VN.n4705 3.904
R987 VN.n4717 VN.t1826 3.904
R988 VN.n4714 VN.t2236 3.904
R989 VN.n4709 VN.n4708 3.904
R990 VN.n5083 VN.n5082 3.904
R991 VN.n5103 VN.t1090 3.904
R992 VN.n5100 VN.t2391 3.904
R993 VN.n5086 VN.n5085 3.904
R994 VN.n5485 VN.n5484 3.904
R995 VN.n5496 VN.t1262 3.904
R996 VN.n5493 VN.t1647 3.904
R997 VN.n5488 VN.n5487 3.904
R998 VN.n5875 VN.n5874 3.904
R999 VN.n5895 VN.t522 3.904
R1000 VN.n5892 VN.t1798 3.904
R1001 VN.n5878 VN.n5877 3.904
R1002 VN.n6277 VN.n6276 3.904
R1003 VN.n6288 VN.t936 3.904
R1004 VN.n6285 VN.t1056 3.904
R1005 VN.n6280 VN.n6279 3.904
R1006 VN.n7118 VN.n7117 3.904
R1007 VN.n7138 VN.t2443 3.904
R1008 VN.n7135 VN.t342 3.904
R1009 VN.n7121 VN.n7120 3.904
R1010 VN.n6722 VN.n6721 3.904
R1011 VN.n6733 VN.t1707 3.904
R1012 VN.n6730 VN.t1818 3.904
R1013 VN.n6725 VN.n6724 3.904
R1014 VN.n7507 VN.n7506 3.904
R1015 VN.n7527 VN.t689 3.904
R1016 VN.n7524 VN.t2278 3.904
R1017 VN.n7510 VN.n7509 3.904
R1018 VN.n7913 VN.n7912 3.904
R1019 VN.n7924 VN.t1132 3.904
R1020 VN.n7921 VN.t1257 3.904
R1021 VN.n7916 VN.n7915 3.904
R1022 VN.n8352 VN.n8351 3.904
R1023 VN.n8372 VN.t61 3.904
R1024 VN.n8369 VN.t617 3.904
R1025 VN.n8355 VN.n8354 3.904
R1026 VN.n8762 VN.n8761 3.904
R1027 VN.n8773 VN.t1997 3.904
R1028 VN.n8770 VN.t2122 3.904
R1029 VN.n8765 VN.n8764 3.904
R1030 VN.n9214 VN.n9213 3.904
R1031 VN.n9234 VN.t1093 3.904
R1032 VN.n9231 VN.t2545 3.904
R1033 VN.n9217 VN.n9216 3.904
R1034 VN.n9624 VN.n9623 3.904
R1035 VN.n9635 VN.t1421 3.904
R1036 VN.n9632 VN.t1653 3.904
R1037 VN.n9627 VN.n9626 3.904
R1038 VN.n10096 VN.n10095 3.904
R1039 VN.n10116 VN.t527 3.904
R1040 VN.n10113 VN.t1968 3.904
R1041 VN.n10099 VN.n10098 3.904
R1042 VN.n10501 VN.n10500 3.904
R1043 VN.n10512 VN.t823 3.904
R1044 VN.n10509 VN.t1061 3.904
R1045 VN.n10504 VN.n10503 3.904
R1046 VN.n10965 VN.n10964 3.904
R1047 VN.n10985 VN.t209 3.904
R1048 VN.n10982 VN.t1395 3.904
R1049 VN.n10968 VN.n10967 3.904
R1050 VN.n11200 VN.n11199 3.904
R1051 VN.n11208 VN.t247 3.904
R1052 VN.n11211 VN.t771 3.904
R1053 VN.n11203 VN.n11202 3.904
R1054 VN.n11742 VN.t2277 3.904
R1055 VN.n11940 VN.n11939 3.904
R1056 VN.n11951 VN.t2247 3.904
R1057 VN.n11948 VN.t873 3.904
R1058 VN.n11943 VN.n11942 3.904
R1059 VN.n5445 VN.t1719 3.904
R1060 VN.n6089 VN.n6088 3.904
R1061 VN.n6105 VN.t594 3.904
R1062 VN.n6108 VN.t1753 3.904
R1063 VN.n6086 VN.n6085 3.904
R1064 VN.n6228 VN.n6227 3.904
R1065 VN.n6237 VN.t892 3.904
R1066 VN.n6234 VN.t1144 3.904
R1067 VN.n6225 VN.n6224 3.904
R1068 VN.n7029 VN.n7028 3.904
R1069 VN.n7046 VN.t2518 3.904
R1070 VN.n7043 VN.t1471 3.904
R1071 VN.n7026 VN.n7025 3.904
R1072 VN.n6673 VN.n6672 3.904
R1073 VN.n6682 VN.t468 3.904
R1074 VN.n6679 VN.t565 3.904
R1075 VN.n6670 VN.n6669 3.904
R1076 VN.n7418 VN.n7417 3.904
R1077 VN.n7435 VN.t1944 3.904
R1078 VN.n7432 VN.t999 3.904
R1079 VN.n7415 VN.n7414 3.904
R1080 VN.n7864 VN.n7863 3.904
R1081 VN.n7873 VN.t2395 3.904
R1082 VN.n7870 VN.t2498 3.904
R1083 VN.n7861 VN.n7860 3.904
R1084 VN.n8263 VN.n8262 3.904
R1085 VN.n8280 VN.t1377 3.904
R1086 VN.n8277 VN.t1857 3.904
R1087 VN.n8260 VN.n8259 3.904
R1088 VN.n8713 VN.n8712 3.904
R1089 VN.n8722 VN.t732 3.904
R1090 VN.n8719 VN.t828 3.904
R1091 VN.n8710 VN.n8709 3.904
R1092 VN.n9125 VN.n9124 3.904
R1093 VN.n9142 VN.t2234 3.904
R1094 VN.n9139 VN.t67 3.904
R1095 VN.n9122 VN.n9121 3.904
R1096 VN.n9575 VN.n9574 3.904
R1097 VN.n9584 VN.t1497 3.904
R1098 VN.n9581 VN.t1609 3.904
R1099 VN.n9572 VN.n9571 3.904
R1100 VN.n10007 VN.n10006 3.904
R1101 VN.n10024 VN.t488 3.904
R1102 VN.n10021 VN.t2059 3.904
R1103 VN.n10004 VN.n10003 3.904
R1104 VN.n10450 VN.n10449 3.904
R1105 VN.n10460 VN.t898 3.904
R1106 VN.n10457 VN.t1013 3.904
R1107 VN.n10447 VN.n10446 3.904
R1108 VN.n10886 VN.n10885 3.904
R1109 VN.n10898 VN.t153 3.904
R1110 VN.n10895 VN.t1474 3.904
R1111 VN.n10883 VN.n10882 3.904
R1112 VN.n11252 VN.n11251 3.904
R1113 VN.n11258 VN.t341 3.904
R1114 VN.n11261 VN.t729 3.904
R1115 VN.n11249 VN.n11248 3.904
R1116 VN.n11821 VN.t1407 3.904
R1117 VN.n11963 VN.n11962 3.904
R1118 VN.n11974 VN.t1385 3.904
R1119 VN.n11971 VN.t2532 3.904
R1120 VN.n11966 VN.n11965 3.904
R1121 VN.n4683 VN.t1446 3.904
R1122 VN.n5301 VN.n5300 3.904
R1123 VN.n5316 VN.t307 3.904
R1124 VN.n5319 VN.t1480 3.904
R1125 VN.n5304 VN.n5303 3.904
R1126 VN.n5451 VN.n5450 3.904
R1127 VN.n5462 VN.t344 3.904
R1128 VN.n5459 VN.t846 3.904
R1129 VN.n5454 VN.n5453 3.904
R1130 VN.n5812 VN.n5811 3.904
R1131 VN.n5832 VN.t2249 3.904
R1132 VN.n5829 VN.t879 3.904
R1133 VN.n5815 VN.n5814 3.904
R1134 VN.n6243 VN.n6242 3.904
R1135 VN.n6254 VN.t147 3.904
R1136 VN.n6251 VN.t280 3.904
R1137 VN.n6246 VN.n6245 3.904
R1138 VN.n7055 VN.n7054 3.904
R1139 VN.n7075 VN.t1658 3.904
R1140 VN.n7072 VN.t727 3.904
R1141 VN.n7058 VN.n7057 3.904
R1142 VN.n6688 VN.n6687 3.904
R1143 VN.n6699 VN.t2119 3.904
R1144 VN.n6696 VN.t2225 3.904
R1145 VN.n6691 VN.n6690 3.904
R1146 VN.n7444 VN.n7443 3.904
R1147 VN.n7464 VN.t1074 3.904
R1148 VN.n7461 VN.t118 3.904
R1149 VN.n7447 VN.n7446 3.904
R1150 VN.n7879 VN.n7878 3.904
R1151 VN.n7890 VN.t1527 3.904
R1152 VN.n7887 VN.t1635 3.904
R1153 VN.n7882 VN.n7881 3.904
R1154 VN.n8289 VN.n8288 3.904
R1155 VN.n8309 VN.t512 3.904
R1156 VN.n8306 VN.t2352 3.904
R1157 VN.n8292 VN.n8291 3.904
R1158 VN.n8728 VN.n8727 3.904
R1159 VN.n8739 VN.t1213 3.904
R1160 VN.n8736 VN.t1332 3.904
R1161 VN.n8731 VN.n8730 3.904
R1162 VN.n9151 VN.n9150 3.904
R1163 VN.n9171 VN.t171 3.904
R1164 VN.n9168 VN.t1757 3.904
R1165 VN.n9154 VN.n9153 3.904
R1166 VN.n9590 VN.n9589 3.904
R1167 VN.n9601 VN.t631 3.904
R1168 VN.n9598 VN.t743 3.904
R1169 VN.n9593 VN.n9592 3.904
R1170 VN.n10033 VN.n10032 3.904
R1171 VN.n10053 VN.t2142 3.904
R1172 VN.n10050 VN.t1188 3.904
R1173 VN.n10036 VN.n10035 3.904
R1174 VN.n10466 VN.n10465 3.904
R1175 VN.n10477 VN.t2561 3.904
R1176 VN.n10474 VN.t139 3.904
R1177 VN.n10469 VN.n10468 3.904
R1178 VN.n10907 VN.n10906 3.904
R1179 VN.n10927 VN.t1952 3.904
R1180 VN.n10924 VN.t607 3.904
R1181 VN.n10910 VN.n10909 3.904
R1182 VN.n11234 VN.n11233 3.904
R1183 VN.n11242 VN.t1985 3.904
R1184 VN.n11245 VN.t2505 3.904
R1185 VN.n11237 VN.n11236 3.904
R1186 VN.n6220 VN.t2017 3.904
R1187 VN.n6654 VN.n6653 3.904
R1188 VN.n6665 VN.t1197 3.904
R1189 VN.n6662 VN.t1432 3.904
R1190 VN.n6657 VN.n6656 3.904
R1191 VN.n7381 VN.n7380 3.904
R1192 VN.n7401 VN.t293 3.904
R1193 VN.n7398 VN.t1739 3.904
R1194 VN.n7384 VN.n7383 3.904
R1195 VN.n7845 VN.n7844 3.904
R1196 VN.n7856 VN.t738 3.904
R1197 VN.n7853 VN.t833 3.904
R1198 VN.n7848 VN.n7847 3.904
R1199 VN.n8226 VN.n8225 3.904
R1200 VN.n8246 VN.t2241 3.904
R1201 VN.n8243 VN.t205 3.904
R1202 VN.n8229 VN.n8228 3.904
R1203 VN.n8694 VN.n8693 3.904
R1204 VN.n8705 VN.t1597 3.904
R1205 VN.n8702 VN.t1698 3.904
R1206 VN.n8697 VN.n8696 3.904
R1207 VN.n9088 VN.n9087 3.904
R1208 VN.n9108 VN.t576 3.904
R1209 VN.n9105 VN.t2168 3.904
R1210 VN.n9091 VN.n9090 3.904
R1211 VN.n9556 VN.n9555 3.904
R1212 VN.n9567 VN.t1006 3.904
R1213 VN.n9564 VN.t1121 3.904
R1214 VN.n9559 VN.n9558 3.904
R1215 VN.n9970 VN.n9969 3.904
R1216 VN.n9990 VN.t2509 3.904
R1217 VN.n9987 VN.t410 3.904
R1218 VN.n9973 VN.n9972 3.904
R1219 VN.n10431 VN.n10430 3.904
R1220 VN.n10442 VN.t1770 3.904
R1221 VN.n10439 VN.t1885 3.904
R1222 VN.n10434 VN.n10433 3.904
R1223 VN.n10849 VN.n10848 3.904
R1224 VN.n10869 VN.t1026 3.904
R1225 VN.n10866 VN.t2342 3.904
R1226 VN.n10852 VN.n10851 3.904
R1227 VN.n11267 VN.n11266 3.904
R1228 VN.n11275 VN.t1205 3.904
R1229 VN.n11278 VN.t1594 3.904
R1230 VN.n11270 VN.n11269 3.904
R1231 VN.n11914 VN.n11913 3.904
R1232 VN.n11929 VN.t475 3.904
R1233 VN.n11926 VN.t1744 3.904
R1234 VN.n11917 VN.n11916 3.904
R1235 VN.n11862 VN.t625 3.904
R1236 VN.n11753 VN.t1490 3.904
R1237 VN.n11891 VN.n11890 3.904
R1238 VN.n11902 VN.t1340 3.904
R1239 VN.n11899 VN.t44 3.904
R1240 VN.n11894 VN.n11893 3.904
R1241 VN.n6648 VN.t2304 3.904
R1242 VN.n7721 VN.n7720 3.904
R1243 VN.n7737 VN.t1161 3.904
R1244 VN.n7740 VN.t31 3.904
R1245 VN.n7718 VN.n7717 3.904
R1246 VN.n7830 VN.n7829 3.904
R1247 VN.n7839 VN.t1483 3.904
R1248 VN.n7836 VN.t1705 3.904
R1249 VN.n7827 VN.n7826 3.904
R1250 VN.n8200 VN.n8199 3.904
R1251 VN.n8217 VN.t585 3.904
R1252 VN.n8214 VN.t940 3.904
R1253 VN.n8197 VN.n8196 3.904
R1254 VN.n8679 VN.n8678 3.904
R1255 VN.n8688 VN.t2463 3.904
R1256 VN.n8685 VN.t2569 3.904
R1257 VN.n8676 VN.n8675 3.904
R1258 VN.n9062 VN.n9061 3.904
R1259 VN.n9079 VN.t1445 3.904
R1260 VN.n9076 VN.t517 3.904
R1261 VN.n9059 VN.n9058 3.904
R1262 VN.n9541 VN.n9540 3.904
R1263 VN.n9550 VN.t1875 3.904
R1264 VN.n9547 VN.t1994 3.904
R1265 VN.n9538 VN.n9537 3.904
R1266 VN.n9944 VN.n9943 3.904
R1267 VN.n9961 VN.t845 3.904
R1268 VN.n9958 VN.t2437 3.904
R1269 VN.n9941 VN.n9940 3.904
R1270 VN.n10415 VN.n10414 3.904
R1271 VN.n10425 VN.t1317 3.904
R1272 VN.n10422 VN.t1418 3.904
R1273 VN.n10412 VN.n10411 3.904
R1274 VN.n10828 VN.n10827 3.904
R1275 VN.n10840 VN.t564 3.904
R1276 VN.n10837 VN.t682 3.904
R1277 VN.n10825 VN.n10824 3.904
R1278 VN.n11286 VN.n11285 3.904
R1279 VN.n11291 VN.t2077 3.904
R1280 VN.n11294 VN.t2459 3.904
R1281 VN.n11283 VN.n11282 3.904
R1282 VN.n11764 VN.t1867 3.904
R1283 VN.n11633 VN.n11632 3.904
R1284 VN.n11644 VN.t1703 3.904
R1285 VN.n11641 VN.t504 3.904
R1286 VN.n11636 VN.n11635 3.904
R1287 VN.n8654 VN.t1782 3.904
R1288 VN.n9428 VN.n9427 3.904
R1289 VN.n9444 VN.t655 3.904
R1290 VN.n9447 VN.t2128 3.904
R1291 VN.n9425 VN.n9424 3.904
R1292 VN.n9507 VN.n9506 3.904
R1293 VN.n9516 VN.t962 3.904
R1294 VN.n9513 VN.t1212 3.904
R1295 VN.n9504 VN.n9503 3.904
R1296 VN.n9881 VN.n9880 3.904
R1297 VN.n9898 VN.t2588 3.904
R1298 VN.n9895 VN.t1534 3.904
R1299 VN.n9878 VN.n9877 3.904
R1300 VN.n10380 VN.n10379 3.904
R1301 VN.n10390 VN.t528 3.904
R1302 VN.n10387 VN.t630 3.904
R1303 VN.n10377 VN.n10376 3.904
R1304 VN.n10770 VN.n10769 3.904
R1305 VN.n10782 VN.t2303 3.904
R1306 VN.n10779 VN.t1066 3.904
R1307 VN.n10767 VN.n10766 3.904
R1308 VN.n11319 VN.n11318 3.904
R1309 VN.n11325 VN.t2452 3.904
R1310 VN.n11328 VN.t337 3.904
R1311 VN.n11316 VN.n11315 3.904
R1312 VN.n11810 VN.t2358 3.904
R1313 VN.n11870 VN.n11869 3.904
R1314 VN.n11881 VN.t832 3.904
R1315 VN.n11878 VN.t956 3.904
R1316 VN.n11873 VN.n11872 3.904
R1317 VN.n7822 VN.t2576 3.904
R1318 VN.n8570 VN.n8569 3.904
R1319 VN.n8585 VN.t1454 3.904
R1320 VN.n8588 VN.t1815 3.904
R1321 VN.n8573 VN.n8572 3.904
R1322 VN.n8660 VN.n8659 3.904
R1323 VN.n8671 VN.t686 3.904
R1324 VN.n8668 VN.t906 3.904
R1325 VN.n8663 VN.n8662 3.904
R1326 VN.n9025 VN.n9024 3.904
R1327 VN.n9045 VN.t2315 3.904
R1328 VN.n9042 VN.t1251 3.904
R1329 VN.n9028 VN.n9027 3.904
R1330 VN.n9522 VN.n9521 3.904
R1331 VN.n9533 VN.t227 3.904
R1332 VN.n9530 VN.t351 3.904
R1333 VN.n9525 VN.n9524 3.904
R1334 VN.n9907 VN.n9906 3.904
R1335 VN.n9927 VN.t1718 3.904
R1336 VN.n9924 VN.t784 3.904
R1337 VN.n9910 VN.n9909 3.904
R1338 VN.n10396 VN.n10395 3.904
R1339 VN.n10407 VN.t2183 3.904
R1340 VN.n10404 VN.t2287 3.904
R1341 VN.n10399 VN.n10398 3.904
R1342 VN.n10791 VN.n10790 3.904
R1343 VN.n10811 VN.t1430 3.904
R1344 VN.n10808 VN.t192 3.904
R1345 VN.n10794 VN.n10793 3.904
R1346 VN.n11301 VN.n11300 3.904
R1347 VN.n11309 VN.t1589 3.904
R1348 VN.n11312 VN.t1980 3.904
R1349 VN.n11304 VN.n11303 3.904
R1350 VN.n11773 VN.t1088 3.904
R1351 VN.n11588 VN.n11587 3.904
R1352 VN.n11599 VN.t913 3.904
R1353 VN.n11596 VN.t2114 3.904
R1354 VN.n11591 VN.n11590 3.904
R1355 VN.n10355 VN.t2368 3.904
R1356 VN.n11479 VN.n11478 3.904
R1357 VN.n11491 VN.t1513 3.904
R1358 VN.n11494 VN.t143 3.904
R1359 VN.n11476 VN.n11475 3.904
R1360 VN.n11353 VN.n11352 3.904
R1361 VN.n11359 VN.t1546 3.904
R1362 VN.n11362 VN.t2075 3.904
R1363 VN.n11350 VN.n11349 3.904
R1364 VN.n11799 VN.t216 3.904
R1365 VN.n11611 VN.n11610 3.904
R1366 VN.n11622 VN.t2575 3.904
R1367 VN.n11619 VN.t1370 3.904
R1368 VN.n11614 VN.n11613 3.904
R1369 VN.n9499 VN.t2089 3.904
R1370 VN.n10315 VN.n10314 3.904
R1371 VN.n10330 VN.t925 3.904
R1372 VN.n10333 VN.t2403 3.904
R1373 VN.n10318 VN.n10317 3.904
R1374 VN.n10361 VN.n10360 3.904
R1375 VN.n10372 VN.t1272 3.904
R1376 VN.n10369 VN.t1496 3.904
R1377 VN.n10364 VN.n10363 3.904
R1378 VN.n10733 VN.n10732 3.904
R1379 VN.n10753 VN.t645 3.904
R1380 VN.n10750 VN.t1806 3.904
R1381 VN.n10736 VN.n10735 3.904
R1382 VN.n11335 VN.n11334 3.904
R1383 VN.n11343 VN.t797 3.904
R1384 VN.n11346 VN.t1203 3.904
R1385 VN.n11338 VN.n11337 3.904
R1386 VN.n12176 VN.t1091 3.904
R1387 VN.n12173 VN.t1355 3.904
R1388 VN.n11093 VN.n11092 3.904
R1389 VN.n11105 VN.t214 3.904
R1390 VN.n11102 VN.t2127 3.904
R1391 VN.n11096 VN.n11095 3.904
R1392 VN.n11499 VN.n11498 3.904
R1393 VN.n11508 VN.t976 3.904
R1394 VN.n11511 VN.t1379 3.904
R1395 VN.n11502 VN.n11501 3.904
R1396 VN.n10337 VN.n10336 3.904
R1397 VN.n10652 VN.t242 3.904
R1398 VN.n10655 VN.t484 3.904
R1399 VN.n10658 VN.n10657 3.904
R1400 VN.n10665 VN.n10664 3.904
R1401 VN.n10678 VN.t1860 3.904
R1402 VN.n10681 VN.t1397 3.904
R1403 VN.n10668 VN.n10667 3.904
R1404 VN.n9750 VN.n9749 3.904
R1405 VN.n9759 VN.t273 3.904
R1406 VN.n9762 VN.t511 3.904
R1407 VN.n9753 VN.n9752 3.904
R1408 VN.n9451 VN.n9450 3.904
R1409 VN.n9464 VN.t1887 3.904
R1410 VN.n9467 VN.t1425 3.904
R1411 VN.n9454 VN.n9453 3.904
R1412 VN.n8888 VN.n8887 3.904
R1413 VN.n8897 VN.t298 3.904
R1414 VN.n8900 VN.t532 3.904
R1415 VN.n8891 VN.n8890 3.904
R1416 VN.n8592 VN.n8591 3.904
R1417 VN.n8605 VN.t1716 3.904
R1418 VN.n8608 VN.t1450 3.904
R1419 VN.n8595 VN.n8594 3.904
R1420 VN.n8039 VN.n8038 3.904
R1421 VN.n8048 VN.t226 3.904
R1422 VN.n8051 VN.t348 3.904
R1423 VN.n8042 VN.n8041 3.904
R1424 VN.n7744 VN.n7743 3.904
R1425 VN.n7757 VN.t2313 3.904
R1426 VN.n7760 VN.t1381 3.904
R1427 VN.n7747 VN.n7746 3.904
R1428 VN.n6848 VN.n6847 3.904
R1429 VN.n6857 VN.t807 3.904
R1430 VN.n6860 VN.t905 3.904
R1431 VN.n6851 VN.n6850 3.904
R1432 VN.n6996 VN.n6995 3.904
R1433 VN.n7012 VN.t374 3.904
R1434 VN.n7009 VN.t1813 3.904
R1435 VN.n6999 VN.n6998 3.904
R1436 VN.n6403 VN.n6402 3.904
R1437 VN.n6412 VN.t1283 3.904
R1438 VN.n6415 VN.t1506 3.904
R1439 VN.n6406 VN.n6405 3.904
R1440 VN.n6112 VN.n6111 3.904
R1441 VN.n6125 VN.t934 3.904
R1442 VN.n6128 VN.t2137 3.904
R1443 VN.n6115 VN.n6114 3.904
R1444 VN.n5611 VN.n5610 3.904
R1445 VN.n5620 VN.t1568 3.904
R1446 VN.n5623 VN.t2099 3.904
R1447 VN.n5614 VN.n5613 3.904
R1448 VN.n5323 VN.n5322 3.904
R1449 VN.n5336 VN.t1538 3.904
R1450 VN.n5339 VN.t165 3.904
R1451 VN.n5326 VN.n5325 3.904
R1452 VN.n4832 VN.n4831 3.904
R1453 VN.n4841 VN.t2162 3.904
R1454 VN.n4844 VN.t127 3.904
R1455 VN.n4835 VN.n4834 3.904
R1456 VN.n4545 VN.n4544 3.904
R1457 VN.n4558 VN.t2131 3.904
R1458 VN.n4561 VN.t759 3.904
R1459 VN.n4548 VN.n4547 3.904
R1460 VN.n4075 VN.n4074 3.904
R1461 VN.n4084 VN.t197 3.904
R1462 VN.n4087 VN.t730 3.904
R1463 VN.n4078 VN.n4077 3.904
R1464 VN.n3791 VN.n3790 3.904
R1465 VN.n3804 VN.t154 3.904
R1466 VN.n3807 VN.t1357 3.904
R1467 VN.n3794 VN.n3793 3.904
R1468 VN.n3331 VN.n3330 3.904
R1469 VN.n3340 VN.t789 3.904
R1470 VN.n3343 VN.t1189 3.904
R1471 VN.n3334 VN.n3333 3.904
R1472 VN.n3048 VN.n3047 3.904
R1473 VN.n3061 VN.t632 3.904
R1474 VN.n3064 VN.t1925 3.904
R1475 VN.n3051 VN.n3050 3.904
R1476 VN.n2609 VN.n2608 3.904
R1477 VN.n2618 VN.t1387 3.904
R1478 VN.n2621 VN.t1487 3.904
R1479 VN.n2612 VN.n2611 3.904
R1480 VN.n2329 VN.n2328 3.904
R1481 VN.n2342 VN.t910 3.904
R1482 VN.n2345 VN.t2506 3.904
R1483 VN.n2332 VN.n2331 3.904
R1484 VN.n1900 VN.n1899 3.904
R1485 VN.n1909 VN.t1954 3.904
R1486 VN.n1912 VN.t2072 3.904
R1487 VN.n1903 VN.n1902 3.904
R1488 VN.n1621 VN.n1620 3.904
R1489 VN.n1634 VN.t656 3.904
R1490 VN.n1637 VN.t572 3.904
R1491 VN.n1624 VN.n1623 3.904
R1492 VN.n1210 VN.n1209 3.904
R1493 VN.n1219 VN.t1678 3.904
R1494 VN.n1222 VN.t1783 3.904
R1495 VN.n1213 VN.n1212 3.904
R1496 VN.n934 VN.n933 3.904
R1497 VN.n947 VN.t1240 3.904
R1498 VN.n950 VN.t303 3.904
R1499 VN.n937 VN.n936 3.904
R1500 VN.n535 VN.n534 3.904
R1501 VN.n544 VN.t2267 3.904
R1502 VN.n547 VN.t2376 3.904
R1503 VN.n538 VN.n537 3.904
R1504 VN.n262 VN.n261 3.904
R1505 VN.n275 VN.t1810 3.904
R1506 VN.n278 VN.t864 3.904
R1507 VN.n265 VN.n264 3.904
R1508 VN.n12286 VN.n12285 3.904
R1509 VN.n12289 VN.t328 3.904
R1510 VN.n12292 VN.t454 3.904
R1511 VN.n12295 VN.n12294 3.904
R1512 VN.n12303 VN.n12302 3.904
R1513 VN.n12316 VN.t2406 3.904
R1514 VN.n12319 VN.t1350 3.904
R1515 VN.n12306 VN.n12305 3.904
R1516 VN.n12268 VN.n12267 3.904
R1517 VN.n12271 VN.t781 3.904
R1518 VN.n12274 VN.t1004 3.904
R1519 VN.n12277 VN.n12276 3.904
R1520 VN.n106 VN.t1632 3.904
R1521 VN.n104 VN.t478 3.904
R1522 VN.n11514 VN.t243 3.904
R1523 VN.n11516 VN.t514 3.904
R1524 VN.n10638 VN.n10637 3.904
R1525 VN.n10646 VN.t1890 3.904
R1526 VN.n10649 VN.t2139 3.904
R1527 VN.n10641 VN.n10640 3.904
R1528 VN.n10689 VN.n10688 3.904
R1529 VN.n10693 VN.t991 3.904
R1530 VN.n10696 VN.t535 3.904
R1531 VN.n10686 VN.n10685 3.904
R1532 VN.n110 VN.t761 3.904
R1533 VN.n108 VN.t2133 3.904
R1534 VN.n12628 VN.n12627 3.904
R1535 VN.n12625 VN.t2552 3.904
R1536 VN.n12622 VN.t130 3.904
R1537 VN.n12348 VN.n12347 3.904
R1538 VN.n12327 VN.n12326 3.904
R1539 VN.n12634 VN.t1539 3.904
R1540 VN.n12637 VN.t601 3.904
R1541 VN.n12324 VN.n12323 3.904
R1542 VN.n12341 VN.n12340 3.904
R1543 VN.n12338 VN.t1974 3.904
R1544 VN.n12335 VN.t2102 3.904
R1545 VN.n12332 VN.n12331 3.904
R1546 VN.n286 VN.n285 3.904
R1547 VN.n290 VN.t935 3.904
R1548 VN.n293 VN.t2526 3.904
R1549 VN.n283 VN.n282 3.904
R1550 VN.n555 VN.n554 3.904
R1551 VN.n560 VN.t1403 3.904
R1552 VN.n563 VN.t1509 3.904
R1553 VN.n552 VN.n551 3.904
R1554 VN.n958 VN.n957 3.904
R1555 VN.n962 VN.t375 3.904
R1556 VN.n965 VN.t778 3.904
R1557 VN.n955 VN.n954 3.904
R1558 VN.n1230 VN.n1229 3.904
R1559 VN.n1235 VN.t2176 3.904
R1560 VN.n1238 VN.t2275 3.904
R1561 VN.n1227 VN.n1226 3.904
R1562 VN.n1645 VN.n1644 3.904
R1563 VN.n1649 VN.t1131 3.904
R1564 VN.n1652 VN.t2230 3.904
R1565 VN.n1642 VN.n1641 3.904
R1566 VN.n1920 VN.n1919 3.904
R1567 VN.n1925 VN.t1086 3.904
R1568 VN.n1928 VN.t1201 3.904
R1569 VN.n1917 VN.n1916 3.904
R1570 VN.n2353 VN.n2352 3.904
R1571 VN.n2357 VN.t2572 3.904
R1572 VN.n2360 VN.t1643 3.904
R1573 VN.n2350 VN.n2349 3.904
R1574 VN.n2629 VN.n2628 3.904
R1575 VN.n2634 VN.t521 3.904
R1576 VN.n2637 VN.t620 3.904
R1577 VN.n2626 VN.n2625 3.904
R1578 VN.n3072 VN.n3071 3.904
R1579 VN.n3076 VN.t2408 3.904
R1580 VN.n3079 VN.t1051 3.904
R1581 VN.n3069 VN.n3068 3.904
R1582 VN.n3351 VN.n3350 3.904
R1583 VN.n3356 VN.t2442 3.904
R1584 VN.n3359 VN.t461 3.904
R1585 VN.n3348 VN.n3347 3.904
R1586 VN.n3815 VN.n3814 3.904
R1587 VN.n3819 VN.t1817 3.904
R1588 VN.n3822 VN.t490 3.904
R1589 VN.n3812 VN.n3811 3.904
R1590 VN.n4095 VN.n4094 3.904
R1591 VN.n4100 VN.t1854 3.904
R1592 VN.n4103 VN.t2384 3.904
R1593 VN.n4092 VN.n4091 3.904
R1594 VN.n4569 VN.n4568 3.904
R1595 VN.n4573 VN.t1255 3.904
R1596 VN.n4576 VN.t2412 3.904
R1597 VN.n4566 VN.n4565 3.904
R1598 VN.n4852 VN.n4851 3.904
R1599 VN.n4857 VN.t1294 3.904
R1600 VN.n4860 VN.t1791 3.904
R1601 VN.n4849 VN.n4848 3.904
R1602 VN.n5347 VN.n5346 3.904
R1603 VN.n5351 VN.t667 3.904
R1604 VN.n5354 VN.t1828 3.904
R1605 VN.n5344 VN.n5343 3.904
R1606 VN.n5631 VN.n5630 3.904
R1607 VN.n5636 VN.t698 3.904
R1608 VN.n5639 VN.t1222 3.904
R1609 VN.n5628 VN.n5627 3.904
R1610 VN.n6136 VN.n6135 3.904
R1611 VN.n6140 VN.t11 3.904
R1612 VN.n6143 VN.t1263 3.904
R1613 VN.n6133 VN.n6132 3.904
R1614 VN.n6423 VN.n6422 3.904
R1615 VN.n6428 VN.t538 3.904
R1616 VN.n6431 VN.t639 3.904
R1617 VN.n6420 VN.n6419 3.904
R1618 VN.n6985 VN.n6984 3.904
R1619 VN.n6992 VN.t2027 3.904
R1620 VN.n6989 VN.t1077 3.904
R1621 VN.n6982 VN.n6981 3.904
R1622 VN.n6868 VN.n6867 3.904
R1623 VN.n6873 VN.t2461 3.904
R1624 VN.n6876 VN.t2567 3.904
R1625 VN.n6865 VN.n6864 3.904
R1626 VN.n7768 VN.n7767 3.904
R1627 VN.n7772 VN.t1443 3.904
R1628 VN.n7775 VN.t318 3.904
R1629 VN.n7765 VN.n7764 3.904
R1630 VN.n8059 VN.n8058 3.904
R1631 VN.n8064 VN.t1683 3.904
R1632 VN.n8067 VN.t1910 3.904
R1633 VN.n8056 VN.n8055 3.904
R1634 VN.n8616 VN.n8615 3.904
R1635 VN.n8620 VN.t766 3.904
R1636 VN.n8623 VN.t582 3.904
R1637 VN.n8613 VN.n8612 3.904
R1638 VN.n8908 VN.n8907 3.904
R1639 VN.n8913 VN.t1947 3.904
R1640 VN.n8916 VN.t2186 3.904
R1641 VN.n8905 VN.n8904 3.904
R1642 VN.n9475 VN.n9474 3.904
R1643 VN.n9798 VN.t1015 3.904
R1644 VN.n9801 VN.t559 3.904
R1645 VN.n9472 VN.n9471 3.904
R1646 VN.n9793 VN.n9792 3.904
R1647 VN.n9790 VN.t1923 3.904
R1648 VN.n9787 VN.t2163 3.904
R1649 VN.n9480 VN.n9479 3.904
R1650 VN.n10701 VN.t255 3.904
R1651 VN.n10698 VN.t2190 3.904
R1652 VN.n9767 VN.n9766 3.904
R1653 VN.n9781 VN.t1048 3.904
R1654 VN.n9784 VN.t1296 3.904
R1655 VN.n9770 VN.n9769 3.904
R1656 VN.n9809 VN.n9808 3.904
R1657 VN.n9813 VN.t141 3.904
R1658 VN.n9816 VN.t2218 3.904
R1659 VN.n9806 VN.n9805 3.904
R1660 VN.n114 VN.t2537 3.904
R1661 VN.n112 VN.t1259 3.904
R1662 VN.n12419 VN.n12418 3.904
R1663 VN.n12424 VN.t1684 3.904
R1664 VN.n12427 VN.t1795 3.904
R1665 VN.n12416 VN.n12415 3.904
R1666 VN.n12645 VN.n12644 3.904
R1667 VN.n12665 VN.t669 3.904
R1668 VN.n12668 VN.t2255 3.904
R1669 VN.n12642 VN.n12641 3.904
R1670 VN.n12659 VN.n12658 3.904
R1671 VN.n12656 VN.t1107 3.904
R1672 VN.n12653 VN.t1225 3.904
R1673 VN.n12650 VN.n12649 3.904
R1674 VN.n301 VN.n300 3.904
R1675 VN.n305 VN.t13 3.904
R1676 VN.n308 VN.t507 3.904
R1677 VN.n298 VN.n297 3.904
R1678 VN.n571 VN.n570 3.904
R1679 VN.n576 VN.t1870 3.904
R1680 VN.n579 VN.t1983 3.904
R1681 VN.n568 VN.n567 3.904
R1682 VN.n973 VN.n972 3.904
R1683 VN.n977 VN.t834 3.904
R1684 VN.n980 VN.t2427 3.904
R1685 VN.n970 VN.n969 3.904
R1686 VN.n1246 VN.n1245 3.904
R1687 VN.n1251 VN.t1309 3.904
R1688 VN.n1254 VN.t1406 3.904
R1689 VN.n1243 VN.n1242 3.904
R1690 VN.n1660 VN.n1659 3.904
R1691 VN.n1664 VN.t267 3.904
R1692 VN.n1667 VN.t1365 3.904
R1693 VN.n1657 VN.n1656 3.904
R1694 VN.n1936 VN.n1935 3.904
R1695 VN.n1941 VN.t213 3.904
R1696 VN.n1944 VN.t333 3.904
R1697 VN.n1933 VN.n1932 3.904
R1698 VN.n2368 VN.n2367 3.904
R1699 VN.n2372 VN.t1833 3.904
R1700 VN.n2375 VN.t772 3.904
R1701 VN.n2365 VN.n2364 3.904
R1702 VN.n2645 VN.n2644 3.904
R1703 VN.n2650 VN.t2172 3.904
R1704 VN.n2653 VN.t2400 3.904
R1705 VN.n2642 VN.n2641 3.904
R1706 VN.n3087 VN.n3086 3.904
R1707 VN.n3091 VN.t1541 3.904
R1708 VN.n3094 VN.t180 3.904
R1709 VN.n3084 VN.n3083 3.904
R1710 VN.n3367 VN.n3366 3.904
R1711 VN.n3372 VN.t1579 3.904
R1712 VN.n3375 VN.t2110 3.904
R1713 VN.n3364 VN.n3363 3.904
R1714 VN.n3830 VN.n3829 3.904
R1715 VN.n3834 VN.t944 3.904
R1716 VN.n3837 VN.t2145 3.904
R1717 VN.n3827 VN.n3826 3.904
R1718 VN.n4111 VN.n4110 3.904
R1719 VN.n4116 VN.t985 3.904
R1720 VN.n4119 VN.t1515 3.904
R1721 VN.n4108 VN.n4107 3.904
R1722 VN.n4584 VN.n4583 3.904
R1723 VN.n4588 VN.t385 3.904
R1724 VN.n4591 VN.t1551 3.904
R1725 VN.n4581 VN.n4580 3.904
R1726 VN.n4868 VN.n4867 3.904
R1727 VN.n4873 VN.t429 3.904
R1728 VN.n4876 VN.t916 3.904
R1729 VN.n4865 VN.n4864 3.904
R1730 VN.n5362 VN.n5361 3.904
R1731 VN.n5366 VN.t2327 3.904
R1732 VN.n5369 VN.t951 3.904
R1733 VN.n5359 VN.n5358 3.904
R1734 VN.n5647 VN.n5646 3.904
R1735 VN.n5652 VN.t2475 3.904
R1736 VN.n5655 VN.t358 3.904
R1737 VN.n5644 VN.n5643 3.904
R1738 VN.n6151 VN.n6150 3.904
R1739 VN.n6155 VN.t1728 3.904
R1740 VN.n6158 VN.t525 3.904
R1741 VN.n6148 VN.n6147 3.904
R1742 VN.n6439 VN.n6438 3.904
R1743 VN.n6444 VN.t2193 3.904
R1744 VN.n6447 VN.t2298 3.904
R1745 VN.n6436 VN.n6435 3.904
R1746 VN.n6970 VN.n6969 3.904
R1747 VN.n6977 VN.t1152 3.904
R1748 VN.n6974 VN.t1995 3.904
R1749 VN.n6967 VN.n6966 3.904
R1750 VN.n6884 VN.n6883 3.904
R1751 VN.n6889 VN.t836 3.904
R1752 VN.n6892 VN.t1069 3.904
R1753 VN.n6881 VN.n6880 3.904
R1754 VN.n7783 VN.n7782 3.904
R1755 VN.n7787 VN.t2445 3.904
R1756 VN.n7790 VN.t1967 3.904
R1757 VN.n7780 VN.n7779 3.904
R1758 VN.n8075 VN.n8074 3.904
R1759 VN.n8080 VN.t817 3.904
R1760 VN.n8083 VN.t1035 3.904
R1761 VN.n8072 VN.n8071 3.904
R1762 VN.n8631 VN.n8630 3.904
R1763 VN.n8952 VN.t2420 3.904
R1764 VN.n8955 VN.t2240 3.904
R1765 VN.n8628 VN.n8627 3.904
R1766 VN.n8947 VN.n8946 3.904
R1767 VN.n8944 VN.t1078 3.904
R1768 VN.n8941 VN.t1321 3.904
R1769 VN.n8636 VN.n8635 3.904
R1770 VN.n9821 VN.t1936 3.904
R1771 VN.n9818 VN.t1351 3.904
R1772 VN.n8921 VN.n8920 3.904
R1773 VN.n8935 VN.t203 3.904
R1774 VN.n8938 VN.t459 3.904
R1775 VN.n8924 VN.n8923 3.904
R1776 VN.n8963 VN.n8962 3.904
R1777 VN.n8967 VN.t1558 3.904
R1778 VN.n8970 VN.t1375 3.904
R1779 VN.n8960 VN.n8959 3.904
R1780 VN.n118 VN.t1672 3.904
R1781 VN.n116 VN.t389 3.904
R1782 VN.n12435 VN.n12434 3.904
R1783 VN.n12440 VN.t818 3.904
R1784 VN.n12443 VN.t920 3.904
R1785 VN.n12432 VN.n12431 3.904
R1786 VN.n12676 VN.n12675 3.904
R1787 VN.n12776 VN.t2329 3.904
R1788 VN.n12779 VN.t195 3.904
R1789 VN.n12673 VN.n12672 3.904
R1790 VN.n12770 VN.n12769 3.904
R1791 VN.n12767 VN.t1592 3.904
R1792 VN.n12764 VN.t1691 3.904
R1793 VN.n12681 VN.n12680 3.904
R1794 VN.n316 VN.n315 3.904
R1795 VN.n320 VN.t566 3.904
R1796 VN.n323 VN.t2160 3.904
R1797 VN.n313 VN.n312 3.904
R1798 VN.n587 VN.n586 3.904
R1799 VN.n592 VN.t1000 3.904
R1800 VN.n595 VN.t1110 3.904
R1801 VN.n584 VN.n583 3.904
R1802 VN.n988 VN.n987 3.904
R1803 VN.n992 VN.t2497 3.904
R1804 VN.n995 VN.t1565 3.904
R1805 VN.n985 VN.n984 3.904
R1806 VN.n1262 VN.n1261 3.904
R1807 VN.n1267 VN.t448 3.904
R1808 VN.n1270 VN.t546 3.904
R1809 VN.n1259 VN.n1258 3.904
R1810 VN.n1675 VN.n1674 3.904
R1811 VN.n1679 VN.t2053 3.904
R1812 VN.n1682 VN.t500 3.904
R1813 VN.n1672 VN.n1671 3.904
R1814 VN.n1952 VN.n1951 3.904
R1815 VN.n1957 VN.t1863 3.904
R1816 VN.n1960 VN.t2123 3.904
R1817 VN.n1949 VN.n1948 3.904
R1818 VN.n2383 VN.n2382 3.904
R1819 VN.n2387 VN.t958 3.904
R1820 VN.n2390 VN.t2424 3.904
R1821 VN.n2380 VN.n2379 3.904
R1822 VN.n2661 VN.n2660 3.904
R1823 VN.n2666 VN.t1305 3.904
R1824 VN.n2669 VN.t1531 3.904
R1825 VN.n2658 VN.n2657 3.904
R1826 VN.n3102 VN.n3101 3.904
R1827 VN.n3106 VN.t672 3.904
R1828 VN.n3109 VN.t1838 3.904
R1829 VN.n3099 VN.n3098 3.904
R1830 VN.n3383 VN.n3382 3.904
R1831 VN.n3388 VN.t712 3.904
R1832 VN.n3391 VN.t1233 3.904
R1833 VN.n3380 VN.n3379 3.904
R1834 VN.n3845 VN.n3844 3.904
R1835 VN.n3849 VN.t19 3.904
R1836 VN.n3852 VN.t1275 3.904
R1837 VN.n3842 VN.n3841 3.904
R1838 VN.n4127 VN.n4126 3.904
R1839 VN.n4132 VN.t96 3.904
R1840 VN.n4135 VN.t647 3.904
R1841 VN.n4124 VN.n4123 3.904
R1842 VN.n4599 VN.n4598 3.904
R1843 VN.n4603 VN.t2039 3.904
R1844 VN.n4606 VN.t678 3.904
R1845 VN.n4596 VN.n4595 3.904
R1846 VN.n4884 VN.n4883 3.904
R1847 VN.n4889 VN.t2203 3.904
R1848 VN.n4892 VN.t2579 3.904
R1849 VN.n4881 VN.n4880 3.904
R1850 VN.n5377 VN.n5376 3.904
R1851 VN.n5381 VN.t1462 3.904
R1852 VN.n5384 VN.t220 3.904
R1853 VN.n5374 VN.n5373 3.904
R1854 VN.n5663 VN.n5662 3.904
R1855 VN.n5668 VN.t1614 3.904
R1856 VN.n5671 VN.t2007 3.904
R1857 VN.n5660 VN.n5659 3.904
R1858 VN.n6166 VN.n6165 3.904
R1859 VN.n6170 VN.t852 3.904
R1860 VN.n6173 VN.t2014 3.904
R1861 VN.n6163 VN.n6162 3.904
R1862 VN.n6455 VN.n6454 3.904
R1863 VN.n6460 VN.t2519 3.904
R1864 VN.n6463 VN.t229 3.904
R1865 VN.n6452 VN.n6451 3.904
R1866 VN.n6955 VN.n6954 3.904
R1867 VN.n6962 VN.t1606 3.904
R1868 VN.n6959 VN.t1122 3.904
R1869 VN.n6952 VN.n6951 3.904
R1870 VN.n6900 VN.n6899 3.904
R1871 VN.n6905 VN.t2499 3.904
R1872 VN.n6908 VN.t196 3.904
R1873 VN.n6897 VN.n6896 3.904
R1874 VN.n7798 VN.n7797 3.904
R1875 VN.n8119 VN.t1582 3.904
R1876 VN.n8122 VN.t1100 3.904
R1877 VN.n7795 VN.n7794 3.904
R1878 VN.n8114 VN.n8113 3.904
R1879 VN.n8111 VN.t2474 3.904
R1880 VN.n8108 VN.t163 3.904
R1881 VN.n7803 VN.n7802 3.904
R1882 VN.n8975 VN.t808 3.904
R1883 VN.n8972 VN.t509 3.904
R1884 VN.n8088 VN.n8087 3.904
R1885 VN.n8102 VN.t1613 3.904
R1886 VN.n8105 VN.t1827 3.904
R1887 VN.n8091 VN.n8090 3.904
R1888 VN.n8130 VN.n8129 3.904
R1889 VN.n8134 VN.t717 3.904
R1890 VN.n8137 VN.t233 3.904
R1891 VN.n8127 VN.n8126 3.904
R1892 VN.n122 VN.t2171 3.904
R1893 VN.n120 VN.t2042 3.904
R1894 VN.n12451 VN.n12450 3.904
R1895 VN.n12456 VN.t1320 3.904
R1896 VN.n12459 VN.t1419 3.904
R1897 VN.n12448 VN.n12447 3.904
R1898 VN.n12790 VN.n12789 3.904
R1899 VN.n12810 VN.t281 3.904
R1900 VN.n12787 VN.t1851 3.904
R1901 VN.n12784 VN.n12783 3.904
R1902 VN.n12804 VN.n12803 3.904
R1903 VN.n12801 VN.t726 3.904
R1904 VN.n12798 VN.t822 3.904
R1905 VN.n12795 VN.n12794 3.904
R1906 VN.n331 VN.n330 3.904
R1907 VN.n335 VN.t2226 3.904
R1908 VN.n338 VN.t1292 3.904
R1909 VN.n328 VN.n327 3.904
R1910 VN.n603 VN.n602 3.904
R1911 VN.n608 VN.t119 3.904
R1912 VN.n611 VN.t246 3.904
R1913 VN.n600 VN.n599 3.904
R1914 VN.n1003 VN.n1002 3.904
R1915 VN.n1007 VN.t1752 3.904
R1916 VN.n1010 VN.t695 3.904
R1917 VN.n1000 VN.n999 3.904
R1918 VN.n1278 VN.n1277 3.904
R1919 VN.n1283 VN.t2094 3.904
R1920 VN.n1286 VN.t2323 3.904
R1921 VN.n1275 VN.n1274 3.904
R1922 VN.n1690 VN.n1689 3.904
R1923 VN.n1694 VN.t1184 3.904
R1924 VN.n1697 VN.t2156 3.904
R1925 VN.n1687 VN.n1686 3.904
R1926 VN.n1968 VN.n1967 3.904
R1927 VN.n1973 VN.t993 3.904
R1928 VN.n1976 VN.t1248 3.904
R1929 VN.n1965 VN.n1964 3.904
R1930 VN.n2398 VN.n2397 3.904
R1931 VN.n2402 VN.t50 3.904
R1932 VN.n2405 VN.t1562 3.904
R1933 VN.n2395 VN.n2394 3.904
R1934 VN.n2677 VN.n2676 3.904
R1935 VN.n2682 VN.t441 3.904
R1936 VN.n2685 VN.t660 3.904
R1937 VN.n2674 VN.n2673 3.904
R1938 VN.n3117 VN.n3116 3.904
R1939 VN.n3121 VN.t2331 3.904
R1940 VN.n3124 VN.t966 3.904
R1941 VN.n3114 VN.n3113 3.904
R1942 VN.n3399 VN.n3398 3.904
R1943 VN.n3404 VN.t2367 3.904
R1944 VN.n3407 VN.t369 3.904
R1945 VN.n3396 VN.n3395 3.904
R1946 VN.n3860 VN.n3859 3.904
R1947 VN.n3864 VN.t1734 3.904
R1948 VN.n3867 VN.t405 3.904
R1949 VN.n3857 VN.n3856 3.904
R1950 VN.n4143 VN.n4142 3.904
R1951 VN.n4148 VN.t1896 3.904
R1952 VN.n4151 VN.t2306 3.904
R1953 VN.n4140 VN.n4139 3.904
R1954 VN.n4614 VN.n4613 3.904
R1955 VN.n4618 VN.t1167 3.904
R1956 VN.n4621 VN.t2457 3.904
R1957 VN.n4611 VN.n4610 3.904
R1958 VN.n4900 VN.n4899 3.904
R1959 VN.n4905 VN.t1335 3.904
R1960 VN.n4908 VN.t1709 3.904
R1961 VN.n4897 VN.n4896 3.904
R1962 VN.n5392 VN.n5391 3.904
R1963 VN.n5396 VN.t589 3.904
R1964 VN.n5399 VN.t1173 3.904
R1965 VN.n5389 VN.n5388 3.904
R1966 VN.n5679 VN.n5678 3.904
R1967 VN.n5684 VN.t2531 3.904
R1968 VN.n5687 VN.t1903 3.904
R1969 VN.n5676 VN.n5675 3.904
R1970 VN.n6181 VN.n6180 3.904
R1971 VN.n6185 VN.t758 3.904
R1972 VN.n6188 VN.t1141 3.904
R1973 VN.n6178 VN.n6177 3.904
R1974 VN.n6471 VN.n6470 3.904
R1975 VN.n6476 VN.t1659 3.904
R1976 VN.n6479 VN.t1876 3.904
R1977 VN.n6468 VN.n6467 3.904
R1978 VN.n6625 VN.n6624 3.904
R1979 VN.n6947 VN.t739 3.904
R1980 VN.n6944 VN.t259 3.904
R1981 VN.n6622 VN.n6621 3.904
R1982 VN.n6939 VN.n6938 3.904
R1983 VN.n6936 VN.t1636 3.904
R1984 VN.n6933 VN.t1852 3.904
R1985 VN.n6630 VN.n6629 3.904
R1986 VN.n8142 VN.t2488 3.904
R1987 VN.n8139 VN.t1880 3.904
R1988 VN.n6913 VN.n6912 3.904
R1989 VN.n6927 VN.t764 3.904
R1990 VN.n6930 VN.t981 3.904
R1991 VN.n6916 VN.n6915 3.904
R1992 VN.n6610 VN.n6609 3.904
R1993 VN.n6617 VN.t2396 3.904
R1994 VN.n6614 VN.t1908 3.904
R1995 VN.n6607 VN.n6606 3.904
R1996 VN.n126 VN.t1304 3.904
R1997 VN.n124 VN.t2511 3.904
R1998 VN.n12467 VN.n12466 3.904
R1999 VN.n12472 VN.t457 3.904
R2000 VN.n12475 VN.t555 3.904
R2001 VN.n12464 VN.n12463 3.904
R2002 VN.n12821 VN.n12820 3.904
R2003 VN.n12841 VN.t1932 3.904
R2004 VN.n12818 VN.t980 3.904
R2005 VN.n12815 VN.n12814 3.904
R2006 VN.n12835 VN.n12834 3.904
R2007 VN.n12832 VN.t2379 3.904
R2008 VN.n12829 VN.t2482 3.904
R2009 VN.n12826 VN.n12825 3.904
R2010 VN.n346 VN.n345 3.904
R2011 VN.n350 VN.t1479 3.904
R2012 VN.n353 VN.t425 3.904
R2013 VN.n343 VN.n342 3.904
R2014 VN.n619 VN.n618 3.904
R2015 VN.n624 VN.t1786 3.904
R2016 VN.n627 VN.t2037 3.904
R2017 VN.n616 VN.n615 3.904
R2018 VN.n1018 VN.n1017 3.904
R2019 VN.n1022 VN.t878 3.904
R2020 VN.n1025 VN.t2354 3.904
R2021 VN.n1015 VN.n1014 3.904
R2022 VN.n1294 VN.n1293 3.904
R2023 VN.n1299 VN.t1218 3.904
R2024 VN.n1302 VN.t1457 3.904
R2025 VN.n1291 VN.n1290 3.904
R2026 VN.n1705 VN.n1704 3.904
R2027 VN.n1709 VN.t312 3.904
R2028 VN.n1712 VN.t1288 3.904
R2029 VN.n1702 VN.n1701 3.904
R2030 VN.n1984 VN.n1983 3.904
R2031 VN.n1989 VN.t109 3.904
R2032 VN.n1992 VN.t380 3.904
R2033 VN.n1981 VN.n1980 3.904
R2034 VN.n2413 VN.n2412 3.904
R2035 VN.n2417 VN.t1746 3.904
R2036 VN.n2420 VN.t692 3.904
R2037 VN.n2410 VN.n2409 3.904
R2038 VN.n2693 VN.n2692 3.904
R2039 VN.n2698 VN.t2086 3.904
R2040 VN.n2701 VN.t2320 3.904
R2041 VN.n2690 VN.n2689 3.904
R2042 VN.n3132 VN.n3131 3.904
R2043 VN.n3136 VN.t1467 3.904
R2044 VN.n3139 VN.t62 3.904
R2045 VN.n3129 VN.n3128 3.904
R2046 VN.n3415 VN.n3414 3.904
R2047 VN.n3420 VN.t1620 3.904
R2048 VN.n3423 VN.t2021 3.904
R2049 VN.n3412 VN.n3411 3.904
R2050 VN.n3875 VN.n3874 3.904
R2051 VN.n3879 VN.t860 3.904
R2052 VN.n3882 VN.t2188 3.904
R2053 VN.n3872 VN.n3871 3.904
R2054 VN.n4159 VN.n4158 3.904
R2055 VN.n4164 VN.t1021 3.904
R2056 VN.n4167 VN.t1435 3.904
R2057 VN.n4156 VN.n4155 3.904
R2058 VN.n4629 VN.n4628 3.904
R2059 VN.n4633 VN.t296 3.904
R2060 VN.n4636 VN.t329 3.904
R2061 VN.n4626 VN.n4625 3.904
R2062 VN.n4916 VN.n4915 3.904
R2063 VN.n4921 VN.t1689 3.904
R2064 VN.n4924 VN.t1060 3.904
R2065 VN.n4913 VN.n4912 3.904
R2066 VN.n5407 VN.n5406 3.904
R2067 VN.n5411 VN.t2441 3.904
R2068 VN.n5414 VN.t305 3.904
R2069 VN.n5404 VN.n5403 3.904
R2070 VN.n5695 VN.n5694 3.904
R2071 VN.n5700 VN.t1667 3.904
R2072 VN.n5703 VN.t1029 3.904
R2073 VN.n5692 VN.n5691 3.904
R2074 VN.n6196 VN.n6195 3.904
R2075 VN.n6515 VN.t2414 3.904
R2076 VN.n6518 VN.t276 3.904
R2077 VN.n6193 VN.n6192 3.904
R2078 VN.n6510 VN.n6509 3.904
R2079 VN.n6507 VN.t791 3.904
R2080 VN.n6504 VN.t1007 3.904
R2081 VN.n6201 VN.n6200 3.904
R2082 VN.n7331 VN.t1652 3.904
R2083 VN.n7328 VN.t1033 3.904
R2084 VN.n6484 VN.n6483 3.904
R2085 VN.n6498 VN.t2444 3.904
R2086 VN.n6501 VN.t132 3.904
R2087 VN.n6487 VN.n6486 3.904
R2088 VN.n6526 VN.n6525 3.904
R2089 VN.n6530 VN.t1552 3.904
R2090 VN.n6533 VN.t1926 3.904
R2091 VN.n6523 VN.n6522 3.904
R2092 VN.n130 VN.t440 3.904
R2093 VN.n128 VN.t1648 3.904
R2094 VN.n12483 VN.n12482 3.904
R2095 VN.n12488 VN.t2105 3.904
R2096 VN.n12491 VN.t2213 3.904
R2097 VN.n12480 VN.n12479 3.904
R2098 VN.n12849 VN.n12848 3.904
R2099 VN.n12869 VN.t1194 3.904
R2100 VN.n12872 VN.t89 3.904
R2101 VN.n12846 VN.n12845 3.904
R2102 VN.n12863 VN.n12862 3.904
R2103 VN.n12860 VN.t1511 3.904
R2104 VN.n12857 VN.t1733 3.904
R2105 VN.n12854 VN.n12853 3.904
R2106 VN.n361 VN.n360 3.904
R2107 VN.n365 VN.t611 3.904
R2108 VN.n368 VN.t2071 3.904
R2109 VN.n358 VN.n357 3.904
R2110 VN.n635 VN.n634 3.904
R2111 VN.n640 VN.t909 3.904
R2112 VN.n643 VN.t1164 3.904
R2113 VN.n632 VN.n631 3.904
R2114 VN.n1033 VN.n1032 3.904
R2115 VN.n1037 VN.t2538 3.904
R2116 VN.n1040 VN.t1486 3.904
R2117 VN.n1030 VN.n1029 3.904
R2118 VN.n1310 VN.n1309 3.904
R2119 VN.n1315 VN.t355 3.904
R2120 VN.n1318 VN.t587 3.904
R2121 VN.n1307 VN.n1306 3.904
R2122 VN.n1720 VN.n1719 3.904
R2123 VN.n1724 VN.t1961 3.904
R2124 VN.n1727 VN.t421 3.904
R2125 VN.n1717 VN.n1716 3.904
R2126 VN.n2000 VN.n1999 3.904
R2127 VN.n2005 VN.t1778 3.904
R2128 VN.n2008 VN.t2034 3.904
R2129 VN.n1997 VN.n1996 3.904
R2130 VN.n2428 VN.n2427 3.904
R2131 VN.n2432 VN.t872 3.904
R2132 VN.n2435 VN.t2350 3.904
R2133 VN.n2425 VN.n2424 3.904
R2134 VN.n2709 VN.n2708 3.904
R2135 VN.n2714 VN.t1347 3.904
R2136 VN.n2717 VN.t1452 3.904
R2137 VN.n2706 VN.n2705 3.904
R2138 VN.n3147 VN.n3146 3.904
R2139 VN.n3151 VN.t597 3.904
R2140 VN.n3154 VN.t1882 3.904
R2141 VN.n3144 VN.n3143 3.904
R2142 VN.n3431 VN.n3430 3.904
R2143 VN.n3436 VN.t749 3.904
R2144 VN.n3439 VN.t1146 3.904
R2145 VN.n3428 VN.n3427 3.904
R2146 VN.n3890 VN.n3889 3.904
R2147 VN.n3894 VN.t2522 3.904
R2148 VN.n3897 VN.t2006 3.904
R2149 VN.n3887 VN.n3886 3.904
R2150 VN.n4175 VN.n4174 3.904
R2151 VN.n4180 VN.t843 3.904
R2152 VN.n4183 VN.t221 3.904
R2153 VN.n4172 VN.n4171 3.904
R2154 VN.n4644 VN.n4643 3.904
R2155 VN.n4648 VN.t1600 3.904
R2156 VN.n4651 VN.t1975 3.904
R2157 VN.n4641 VN.n4640 3.904
R2158 VN.n4932 VN.n4931 3.904
R2159 VN.n4937 VN.t821 3.904
R2160 VN.n4940 VN.t186 3.904
R2161 VN.n4929 VN.n4928 3.904
R2162 VN.n5422 VN.n5421 3.904
R2163 VN.n5739 VN.t1577 3.904
R2164 VN.n5742 VN.t1953 3.904
R2165 VN.n5419 VN.n5418 3.904
R2166 VN.n5734 VN.n5733 3.904
R2167 VN.n5731 VN.t802 3.904
R2168 VN.n5728 VN.t159 3.904
R2169 VN.n5427 VN.n5426 3.904
R2170 VN.n6538 VN.t804 3.904
R2171 VN.n6535 VN.t1050 3.904
R2172 VN.n5708 VN.n5707 3.904
R2173 VN.n5722 VN.t2455 3.904
R2174 VN.n5725 VN.t1821 3.904
R2175 VN.n5711 VN.n5710 3.904
R2176 VN.n5750 VN.n5749 3.904
R2177 VN.n5754 VN.t710 3.904
R2178 VN.n5757 VN.t1085 3.904
R2179 VN.n5747 VN.n5746 3.904
R2180 VN.n134 VN.t2085 3.904
R2181 VN.n132 VN.t887 3.904
R2182 VN.n12499 VN.n12498 3.904
R2183 VN.n12504 VN.t1228 3.904
R2184 VN.n12507 VN.t1466 3.904
R2185 VN.n12496 VN.n12495 3.904
R2186 VN.n12880 VN.n12879 3.904
R2187 VN.n12900 VN.t325 3.904
R2188 VN.n12903 VN.t1767 3.904
R2189 VN.n12877 VN.n12876 3.904
R2190 VN.n12894 VN.n12893 3.904
R2191 VN.n12891 VN.t642 3.904
R2192 VN.n12888 VN.t858 3.904
R2193 VN.n12885 VN.n12884 3.904
R2194 VN.n376 VN.n375 3.904
R2195 VN.n380 VN.t2263 3.904
R2196 VN.n383 VN.t1200 3.904
R2197 VN.n373 VN.n372 3.904
R2198 VN.n651 VN.n650 3.904
R2199 VN.n656 VN.t2571 3.904
R2200 VN.n659 VN.t295 3.904
R2201 VN.n648 VN.n647 3.904
R2202 VN.n1048 VN.n1047 3.904
R2203 VN.n1052 VN.t1673 3.904
R2204 VN.n1055 VN.t619 3.904
R2205 VN.n1045 VN.n1044 3.904
R2206 VN.n1326 VN.n1325 3.904
R2207 VN.n1331 VN.t2000 3.904
R2208 VN.n1334 VN.t2243 3.904
R2209 VN.n1323 VN.n1322 3.904
R2210 VN.n1735 VN.n1734 3.904
R2211 VN.n1739 VN.t1094 3.904
R2212 VN.n1742 VN.t2068 3.904
R2213 VN.n1732 VN.n1731 3.904
R2214 VN.n2016 VN.n2015 3.904
R2215 VN.n2021 VN.t1036 3.904
R2216 VN.n2024 VN.t1159 3.904
R2217 VN.n2013 VN.n2012 3.904
R2218 VN.n2443 VN.n2442 3.904
R2219 VN.n2447 VN.t2534 3.904
R2220 VN.n2450 VN.t1603 3.904
R2221 VN.n2440 VN.n2439 3.904
R2222 VN.n2725 VN.n2724 3.904
R2223 VN.n2730 VN.t481 3.904
R2224 VN.n2733 VN.t583 3.904
R2225 VN.n2722 VN.n2721 3.904
R2226 VN.n3162 VN.n3161 3.904
R2227 VN.n3166 VN.t2252 3.904
R2228 VN.n3169 VN.t1163 3.904
R2229 VN.n3159 VN.n3158 3.904
R2230 VN.n3447 VN.n3446 3.904
R2231 VN.n3452 VN.t2528 3.904
R2232 VN.n3455 VN.t1898 3.904
R2233 VN.n3444 VN.n3443 3.904
R2234 VN.n3905 VN.n3904 3.904
R2235 VN.n3909 VN.t754 3.904
R2236 VN.n3912 VN.t1133 3.904
R2237 VN.n3902 VN.n3901 3.904
R2238 VN.n4191 VN.n4190 3.904
R2239 VN.n4196 VN.t2507 3.904
R2240 VN.n4199 VN.t1871 3.904
R2241 VN.n4188 VN.n4187 3.904
R2242 VN.n4659 VN.n4658 3.904
R2243 VN.n4976 VN.t734 3.904
R2244 VN.n4979 VN.t1108 3.904
R2245 VN.n4656 VN.n4655 3.904
R2246 VN.n4971 VN.n4970 3.904
R2247 VN.n4968 VN.t2481 3.904
R2248 VN.n4965 VN.t1843 3.904
R2249 VN.n4664 VN.n4663 3.904
R2250 VN.n5762 VN.t2484 3.904
R2251 VN.n5759 VN.t212 3.904
R2252 VN.n4945 VN.n4944 3.904
R2253 VN.n4959 VN.t1618 3.904
R2254 VN.n4962 VN.t971 3.904
R2255 VN.n4948 VN.n4947 3.904
R2256 VN.n4987 VN.n4986 3.904
R2257 VN.n4991 VN.t2389 3.904
R2258 VN.n4994 VN.t240 3.904
R2259 VN.n4984 VN.n4983 3.904
R2260 VN.n138 VN.t1210 3.904
R2261 VN.n136 VN.t2548 3.904
R2262 VN.n12515 VN.n12514 3.904
R2263 VN.n12520 VN.t362 3.904
R2264 VN.n12523 VN.t595 3.904
R2265 VN.n12512 VN.n12511 3.904
R2266 VN.n12911 VN.n12910 3.904
R2267 VN.n12931 VN.t1971 3.904
R2268 VN.n12934 VN.t896 3.904
R2269 VN.n12908 VN.n12907 3.904
R2270 VN.n12925 VN.n12924 3.904
R2271 VN.n12922 VN.t2301 3.904
R2272 VN.n12919 VN.t2520 3.904
R2273 VN.n12916 VN.n12915 3.904
R2274 VN.n391 VN.n390 3.904
R2275 VN.n395 VN.t1398 3.904
R2276 VN.n398 VN.t332 3.904
R2277 VN.n388 VN.n387 3.904
R2278 VN.n667 VN.n666 3.904
R2279 VN.n672 VN.t1700 3.904
R2280 VN.n675 VN.t1946 3.904
R2281 VN.n664 VN.n663 3.904
R2282 VN.n1063 VN.n1062 3.904
R2283 VN.n1067 VN.t806 3.904
R2284 VN.n1070 VN.t2271 3.904
R2285 VN.n1060 VN.n1059 3.904
R2286 VN.n1342 VN.n1341 3.904
R2287 VN.n1347 VN.t1268 3.904
R2288 VN.n1350 VN.t1380 3.904
R2289 VN.n1339 VN.n1338 3.904
R2290 VN.n1750 VN.n1749 3.904
R2291 VN.n1754 VN.t225 3.904
R2292 VN.n1757 VN.t1329 3.904
R2293 VN.n1747 VN.n1746 3.904
R2294 VN.n2032 VN.n2031 3.904
R2295 VN.n2037 VN.t164 3.904
R2296 VN.n2040 VN.t292 3.904
R2297 VN.n2029 VN.n2028 3.904
R2298 VN.n2458 VN.n2457 3.904
R2299 VN.n2462 VN.t1670 3.904
R2300 VN.n2465 VN.t323 3.904
R2301 VN.n2455 VN.n2454 3.904
R2302 VN.n2741 VN.n2740 3.904
R2303 VN.n2746 VN.t1686 3.904
R2304 VN.n2749 VN.t1915 3.904
R2305 VN.n2738 VN.n2737 3.904
R2306 VN.n3177 VN.n3176 3.904
R2307 VN.n3181 VN.t2434 3.904
R2308 VN.n3184 VN.t294 3.904
R2309 VN.n3174 VN.n3173 3.904
R2310 VN.n3463 VN.n3462 3.904
R2311 VN.n3468 VN.t1664 3.904
R2312 VN.n3471 VN.t1023 3.904
R2313 VN.n3460 VN.n3459 3.904
R2314 VN.n3920 VN.n3919 3.904
R2315 VN.n4235 VN.t2411 3.904
R2316 VN.n4238 VN.t270 3.904
R2317 VN.n3917 VN.n3916 3.904
R2318 VN.n4230 VN.n4229 3.904
R2319 VN.n4227 VN.t1644 3.904
R2320 VN.n4224 VN.t1001 3.904
R2321 VN.n3925 VN.n3924 3.904
R2322 VN.n4999 VN.t1649 3.904
R2323 VN.n4996 VN.t1889 3.904
R2324 VN.n4204 VN.n4203 3.904
R2325 VN.n4218 VN.t773 3.904
R2326 VN.n4221 VN.t123 3.904
R2327 VN.n4207 VN.n4206 3.904
R2328 VN.n4246 VN.n4245 3.904
R2329 VN.n4250 VN.t1548 3.904
R2330 VN.n4253 VN.t1920 3.904
R2331 VN.n4243 VN.n4242 3.904
R2332 VN.n142 VN.t347 3.904
R2333 VN.n140 VN.t1680 3.904
R2334 VN.n12531 VN.n12530 3.904
R2335 VN.n12536 VN.t2012 3.904
R2336 VN.n12539 VN.t2250 3.904
R2337 VN.n12528 VN.n12527 3.904
R2338 VN.n12942 VN.n12941 3.904
R2339 VN.n12962 VN.t1103 3.904
R2340 VN.n12965 VN.t2558 3.904
R2341 VN.n12939 VN.n12938 3.904
R2342 VN.n12956 VN.n12955 3.904
R2343 VN.n12953 VN.t1428 3.904
R2344 VN.n12950 VN.t1660 3.904
R2345 VN.n12947 VN.n12946 3.904
R2346 VN.n406 VN.n405 3.904
R2347 VN.n410 VN.t537 3.904
R2348 VN.n413 VN.t1978 3.904
R2349 VN.n403 VN.n402 3.904
R2350 VN.n683 VN.n682 3.904
R2351 VN.n688 VN.t955 3.904
R2352 VN.n691 VN.t1076 3.904
R2353 VN.n680 VN.n679 3.904
R2354 VN.n1078 VN.n1077 3.904
R2355 VN.n1082 VN.t2460 3.904
R2356 VN.n1085 VN.t1530 3.904
R2357 VN.n1075 VN.n1074 3.904
R2358 VN.n1358 VN.n1357 3.904
R2359 VN.n1363 VN.t399 3.904
R2360 VN.n1366 VN.t515 3.904
R2361 VN.n1355 VN.n1354 3.904
R2362 VN.n1765 VN.n1764 3.904
R2363 VN.n1769 VN.t1873 3.904
R2364 VN.n1772 VN.t2003 3.904
R2365 VN.n1762 VN.n1761 3.904
R2366 VN.n2048 VN.n2047 3.904
R2367 VN.n2053 VN.t840 3.904
R2368 VN.n2056 VN.t1073 3.904
R2369 VN.n2045 VN.n2044 3.904
R2370 VN.n2473 VN.n2472 3.904
R2371 VN.n2477 VN.t2447 3.904
R2372 VN.n2480 VN.t1970 3.904
R2373 VN.n2470 VN.n2469 3.904
R2374 VN.n2757 VN.n2756 3.904
R2375 VN.n2762 VN.t820 3.904
R2376 VN.n2765 VN.t1040 3.904
R2377 VN.n2754 VN.n2753 3.904
R2378 VN.n3192 VN.n3191 3.904
R2379 VN.n3507 VN.t1574 3.904
R2380 VN.n3510 VN.t1945 3.904
R2381 VN.n3189 VN.n3188 3.904
R2382 VN.n3502 VN.n3501 3.904
R2383 VN.n3499 VN.t796 3.904
R2384 VN.n3496 VN.t151 3.904
R2385 VN.n3197 VN.n3196 3.904
R2386 VN.n4258 VN.t800 3.904
R2387 VN.n4255 VN.t1045 3.904
R2388 VN.n3476 VN.n3475 3.904
R2389 VN.n3490 VN.t2450 3.904
R2390 VN.n3493 VN.t1814 3.904
R2391 VN.n3479 VN.n3478 3.904
R2392 VN.n3518 VN.n3517 3.904
R2393 VN.n3522 VN.t705 3.904
R2394 VN.n3525 VN.t1075 3.904
R2395 VN.n3515 VN.n3514 3.904
R2396 VN.n146 VN.t1990 3.904
R2397 VN.n144 VN.t814 3.904
R2398 VN.n12547 VN.n12546 3.904
R2399 VN.n12552 VN.t1139 3.904
R2400 VN.n12555 VN.t1389 3.904
R2401 VN.n12544 VN.n12543 3.904
R2402 VN.n12973 VN.n12972 3.904
R2403 VN.n12993 VN.t237 3.904
R2404 VN.n12996 VN.t1688 3.904
R2405 VN.n12970 VN.n12969 3.904
R2406 VN.n12987 VN.n12986 3.904
R2407 VN.n12984 VN.t681 3.904
R2408 VN.n12981 VN.t792 3.904
R2409 VN.n12978 VN.n12977 3.904
R2410 VN.n421 VN.n420 3.904
R2411 VN.n425 VN.t2192 3.904
R2412 VN.n428 VN.t1247 3.904
R2413 VN.n418 VN.n417 3.904
R2414 VN.n699 VN.n698 3.904
R2415 VN.n704 VN.t42 3.904
R2416 VN.n707 VN.t202 3.904
R2417 VN.n696 VN.n695 3.904
R2418 VN.n1093 VN.n1092 3.904
R2419 VN.n1097 VN.t1595 3.904
R2420 VN.n1100 VN.t677 3.904
R2421 VN.n1090 VN.n1089 3.904
R2422 VN.n1374 VN.n1373 3.904
R2423 VN.n1379 VN.t2064 3.904
R2424 VN.n1382 VN.t2284 3.904
R2425 VN.n1371 VN.n1370 3.904
R2426 VN.n1780 VN.n1779 3.904
R2427 VN.n1784 VN.t1130 3.904
R2428 VN.n1787 VN.t1129 3.904
R2429 VN.n1777 VN.n1776 3.904
R2430 VN.n2064 VN.n2063 3.904
R2431 VN.n2069 VN.t2503 3.904
R2432 VN.n2072 VN.t198 3.904
R2433 VN.n2061 VN.n2060 3.904
R2434 VN.n2488 VN.n2487 3.904
R2435 VN.n2801 VN.t1584 3.904
R2436 VN.n2804 VN.t1102 3.904
R2437 VN.n2485 VN.n2484 3.904
R2438 VN.n2796 VN.n2795 3.904
R2439 VN.n2793 VN.t2477 3.904
R2440 VN.n2790 VN.t168 3.904
R2441 VN.n2493 VN.n2492 3.904
R2442 VN.n3530 VN.t2478 3.904
R2443 VN.n3527 VN.t200 3.904
R2444 VN.n2770 VN.n2769 3.904
R2445 VN.n2784 VN.t1616 3.904
R2446 VN.n2787 VN.t1829 3.904
R2447 VN.n2773 VN.n2772 3.904
R2448 VN.n2812 VN.n2811 3.904
R2449 VN.n2816 VN.t720 3.904
R2450 VN.n2819 VN.t235 3.904
R2451 VN.n2809 VN.n2808 3.904
R2452 VN.n150 VN.t1116 3.904
R2453 VN.n148 VN.t2471 3.904
R2454 VN.n12563 VN.n12562 3.904
R2455 VN.n12568 VN.t409 3.904
R2456 VN.n12571 VN.t523 3.904
R2457 VN.n12560 VN.n12559 3.904
R2458 VN.n13004 VN.n13003 3.904
R2459 VN.n13024 VN.t1884 3.904
R2460 VN.n13027 VN.t939 3.904
R2461 VN.n13001 VN.n13000 3.904
R2462 VN.n13018 VN.n13017 3.904
R2463 VN.n13015 VN.t2341 3.904
R2464 VN.n13012 VN.t2446 3.904
R2465 VN.n13009 VN.n13008 3.904
R2466 VN.n436 VN.n435 3.904
R2467 VN.n440 VN.t1323 3.904
R2468 VN.n443 VN.t2365 3.904
R2469 VN.n433 VN.n432 3.904
R2470 VN.n715 VN.n714 3.904
R2471 VN.n720 VN.t1220 3.904
R2472 VN.n723 VN.t1441 3.904
R2473 VN.n712 VN.n711 3.904
R2474 VN.n1108 VN.n1107 3.904
R2475 VN.n1112 VN.t291 3.904
R2476 VN.n1115 VN.t2338 3.904
R2477 VN.n1105 VN.n1104 3.904
R2478 VN.n1390 VN.n1389 3.904
R2479 VN.n1395 VN.t1192 3.904
R2480 VN.n1398 VN.t1415 3.904
R2481 VN.n1387 VN.n1386 3.904
R2482 VN.n1795 VN.n1794 3.904
R2483 VN.n2108 VN.t264 3.904
R2484 VN.n2111 VN.t263 3.904
R2485 VN.n1792 VN.n1791 3.904
R2486 VN.n2103 VN.n2102 3.904
R2487 VN.n2100 VN.t1641 3.904
R2488 VN.n2097 VN.t1855 3.904
R2489 VN.n1800 VN.n1799 3.904
R2490 VN.n2824 VN.t2491 3.904
R2491 VN.n2821 VN.t1883 3.904
R2492 VN.n2077 VN.n2076 3.904
R2493 VN.n2091 VN.t769 3.904
R2494 VN.n2094 VN.t986 3.904
R2495 VN.n2080 VN.n2079 3.904
R2496 VN.n2119 VN.n2118 3.904
R2497 VN.n2123 VN.t1914 3.904
R2498 VN.n2126 VN.t1913 3.904
R2499 VN.n2116 VN.n2115 3.904
R2500 VN.n154 VN.t395 3.904
R2501 VN.n152 VN.t1608 3.904
R2502 VN.n12579 VN.n12578 3.904
R2503 VN.n12584 VN.t2058 3.904
R2504 VN.n12587 VN.t2177 3.904
R2505 VN.n12576 VN.n12575 3.904
R2506 VN.n13035 VN.n13034 3.904
R2507 VN.n13055 VN.t1012 3.904
R2508 VN.n13058 VN.t1519 3.904
R2509 VN.n13032 VN.n13031 3.904
R2510 VN.n13049 VN.n13048 3.904
R2511 VN.n13046 VN.t379 3.904
R2512 VN.n13043 VN.t602 3.904
R2513 VN.n13040 VN.n13039 3.904
R2514 VN.n451 VN.n450 3.904
R2515 VN.n455 VN.t1966 3.904
R2516 VN.n458 VN.t1495 3.904
R2517 VN.n448 VN.n447 3.904
R2518 VN.n731 VN.n730 3.904
R2519 VN.n736 VN.t357 3.904
R2520 VN.n739 VN.t573 3.904
R2521 VN.n728 VN.n727 3.904
R2522 VN.n1123 VN.n1122 3.904
R2523 VN.n1434 VN.t1943 3.904
R2524 VN.n1437 VN.t1473 3.904
R2525 VN.n1120 VN.n1119 3.904
R2526 VN.n1429 VN.n1428 3.904
R2527 VN.n1426 VN.t322 3.904
R2528 VN.n1423 VN.t553 3.904
R2529 VN.n1128 VN.n1127 3.904
R2530 VN.n2131 VN.t1182 3.904
R2531 VN.n2128 VN.t1039 3.904
R2532 VN.n1403 VN.n1402 3.904
R2533 VN.n1417 VN.t1969 3.904
R2534 VN.n1420 VN.t2209 3.904
R2535 VN.n1406 VN.n1405 3.904
R2536 VN.n1445 VN.n1444 3.904
R2537 VN.n1449 VN.t1072 3.904
R2538 VN.n1452 VN.t606 3.904
R2539 VN.n1442 VN.n1441 3.904
R2540 VN.n158 VN.t1537 3.904
R2541 VN.n156 VN.t742 3.904
R2542 VN.n12595 VN.n12594 3.904
R2543 VN.n12600 VN.t2055 3.904
R2544 VN.n12603 VN.t2280 3.904
R2545 VN.n12592 VN.n12591 3.904
R2546 VN.n13066 VN.n13065 3.904
R2547 VN.n13086 VN.t1119 3.904
R2548 VN.n13089 VN.t650 3.904
R2549 VN.n13063 VN.n13062 3.904
R2550 VN.n13080 VN.n13079 3.904
R2551 VN.n13077 VN.t2033 3.904
R2552 VN.n13074 VN.t2256 3.904
R2553 VN.n13071 VN.n13070 3.904
R2554 VN.n466 VN.n465 3.904
R2555 VN.n774 VN.t1099 3.904
R2556 VN.n777 VN.t628 3.904
R2557 VN.n463 VN.n462 3.904
R2558 VN.n769 VN.n768 3.904
R2559 VN.n766 VN.t2002 3.904
R2560 VN.n763 VN.t2231 3.904
R2561 VN.n471 VN.n470 3.904
R2562 VN.n1457 VN.t343 3.904
R2563 VN.n1454 VN.t2258 3.904
R2564 VN.n742 VN.n741 3.904
R2565 VN.n757 VN.t1128 3.904
R2566 VN.n760 VN.t1366 3.904
R2567 VN.n745 VN.n744 3.904
R2568 VN.n787 VN.n786 3.904
R2569 VN.n796 VN.t232 3.904
R2570 VN.n799 VN.t2282 3.904
R2571 VN.n790 VN.n789 3.904
R2572 VN.n162 VN.t665 3.904
R2573 VN.n160 VN.t285 3.904
R2574 VN.n12608 VN.n12607 3.904
R2575 VN.n12616 VN.t1187 3.904
R2576 VN.n12619 VN.t1410 3.904
R2577 VN.n12611 VN.n12610 3.904
R2578 VN.n13098 VN.n13097 3.904
R2579 VN.n13106 VN.t256 3.904
R2580 VN.n13109 VN.t2309 3.904
R2581 VN.n13101 VN.n13100 3.904
R2582 VN.n12750 VN.n12749 3.904
R2583 VN.n12758 VN.t1157 3.904
R2584 VN.n12761 VN.t1391 3.904
R2585 VN.n12753 VN.n12752 3.904
R2586 VN.n804 VN.t2019 3.904
R2587 VN.n801 VN.t1413 3.904
R2588 VN.n166 VN.t2325 3.904
R2589 VN.n164 VN.t1937 3.904
R2590 VN.n12379 VN.n12378 3.904
R2591 VN.n12390 VN.t316 3.904
R2592 VN.n12387 VN.t550 3.904
R2593 VN.n12382 VN.n12381 3.904
R2594 VN.n12227 VN.n12226 3.904
R2595 VN.n12235 VN.t1907 3.904
R2596 VN.n12218 VN.t1439 3.904
R2597 VN.n12230 VN.n12229 3.904
R2598 VN.n12724 VN.n12723 3.904
R2599 VN.n12742 VN.t289 3.904
R2600 VN.n12739 VN.t526 3.904
R2601 VN.n12727 VN.n12726 3.904
R2602 VN.n12400 VN.n12399 3.904
R2603 VN.n12403 VN.t2207 3.904
R2604 VN.n6584 VN.t2336 3.904
R2605 VN.n6582 VN.n6581 3.904
R2606 VN.n6603 VN.n6602 3.643
R2607 VN.n7327 VN.t1219 3.643
R2608 VN.n11382 VN.t2348 3.643
R2609 VN.n11366 VN.t945 3.643
R2610 VN.n11666 VN.t387 3.643
R2611 VN.n11667 VN.t1754 3.643
R2612 VN.n11574 VN.t987 3.643
R2613 VN.n11577 VN.n11576 3.643
R2614 VN.n11569 VN.t2148 3.643
R2615 VN.n11547 VN.n11546 3.643
R2616 VN.n11777 VN.t60 3.643
R2617 VN.n11790 VN.t1256 3.643
R2618 VN.n12407 VN.t1891 3.643
R2619 VN.n12410 VN.n12409 3.643
R2620 VN.n13116 VN.t1521 3.643
R2621 VN.n84 VN.t408 3.643
R2622 VN.n11676 VN.t2020 3.643
R2623 VN.n11677 VN.t983 3.643
R2624 VN.n12157 VN.t1158 3.643
R2625 VN.n12170 VN.n12169 3.643
R2626 VN.n12167 VN.n12166 3.643
R2627 VN.n12154 VN.t2310 3.643
R2628 VN.n12369 VN.t1581 3.643
R2629 VN.n12350 VN.t2428 3.643
R2630 VN.n12244 VN.t2466 3.643
R2631 VN.n12261 VN.n12260 3.643
R2632 VN.n12264 VN.n12263 3.643
R2633 VN.n12241 VN.t1084 3.643
R2634 VN.n12709 VN.t989 3.643
R2635 VN.n12718 VN.n12717 3.643
R2636 VN.n12715 VN.n12714 3.643
R2637 VN.n12706 VN.t2150 3.643
R2638 VN.n215 VN.t2018 3.643
R2639 VN.n232 VN.n231 3.643
R2640 VN.n229 VN.n228 3.643
R2641 VN.n212 VN.t520 3.643
R2642 VN.n520 VN.t433 3.643
R2643 VN.n529 VN.n528 3.643
R2644 VN.n526 VN.n525 3.643
R2645 VN.n517 VN.t1556 3.643
R2646 VN.n886 VN.t1433 3.643
R2647 VN.n903 VN.n902 3.643
R2648 VN.n900 VN.n899 3.643
R2649 VN.n883 VN.t2562 3.643
R2650 VN.n1195 VN.t2361 3.643
R2651 VN.n1204 VN.n1203 3.643
R2652 VN.n1201 VN.n1200 3.643
R2653 VN.n1192 VN.t961 3.643
R2654 VN.n1569 VN.t835 3.643
R2655 VN.n1586 VN.n1585 3.643
R2656 VN.n1583 VN.n1582 3.643
R2657 VN.n1566 VN.t1984 3.643
R2658 VN.n1885 VN.t1295 3.643
R2659 VN.n1894 VN.n1893 3.643
R2660 VN.n1891 VN.n1890 3.643
R2661 VN.n1882 VN.t2413 3.643
R2662 VN.n2277 VN.t1113 3.643
R2663 VN.n2294 VN.n2293 3.643
R2664 VN.n2291 VN.n2290 3.643
R2665 VN.n2274 VN.t2261 3.643
R2666 VN.n2594 VN.t2051 3.643
R2667 VN.n2603 VN.n2602 3.643
R2668 VN.n2600 VN.n2599 3.643
R2669 VN.n2591 VN.t662 3.643
R2670 VN.n2999 VN.t816 3.643
R2671 VN.n3016 VN.n3015 3.643
R2672 VN.n3013 VN.n3012 3.643
R2673 VN.n2996 VN.t1671 3.643
R2674 VN.n3316 VN.t1470 3.643
R2675 VN.n3325 VN.n3324 3.643
R2676 VN.n3322 VN.n3321 3.643
R2677 VN.n3313 VN.t5 3.643
R2678 VN.n3739 VN.t238 3.643
R2679 VN.n3756 VN.n3755 3.643
R2680 VN.n3753 VN.n3752 3.643
R2681 VN.n3736 VN.t1390 3.643
R2682 VN.n4060 VN.t998 3.643
R2683 VN.n4069 VN.n4068 3.643
R2684 VN.n4066 VN.n4065 3.643
R2685 VN.n4057 VN.t2024 3.643
R2686 VN.n4496 VN.t2195 3.643
R2687 VN.n4513 VN.n4512 3.643
R2688 VN.n4510 VN.n4509 3.643
R2689 VN.n4493 VN.t793 3.643
R2690 VN.n4817 VN.t447 3.643
R2691 VN.n4826 VN.n4825 3.643
R2692 VN.n4823 VN.n4822 3.643
R2693 VN.n4814 VN.t1564 3.643
R2694 VN.n5271 VN.t1598 3.643
R2695 VN.n5288 VN.n5287 3.643
R2696 VN.n5285 VN.n5284 3.643
R2697 VN.n5268 VN.t206 3.643
R2698 VN.n5596 VN.t2370 3.643
R2699 VN.n5605 VN.n5604 3.643
R2700 VN.n5602 VN.n5601 3.643
R2701 VN.n5593 VN.t969 3.643
R2702 VN.n6063 VN.t1008 3.643
R2703 VN.n6080 VN.n6079 3.643
R2704 VN.n6077 VN.n6076 3.643
R2705 VN.n6060 VN.t2169 3.643
R2706 VN.n6388 VN.t2076 3.643
R2707 VN.n6397 VN.n6396 3.643
R2708 VN.n6394 VN.n6393 3.643
R2709 VN.n6385 VN.t413 3.643
R2710 VN.n7306 VN.t456 3.643
R2711 VN.n7323 VN.n7322 3.643
R2712 VN.n7320 VN.n7319 3.643
R2713 VN.n7303 VN.t1576 3.643
R2714 VN.n6833 VN.t1489 3.643
R2715 VN.n6842 VN.n6841 3.643
R2716 VN.n6839 VN.n6838 3.643
R2717 VN.n6830 VN.t38 3.643
R2718 VN.n7695 VN.t2496 3.643
R2719 VN.n7712 VN.n7711 3.643
R2720 VN.n7709 VN.n7708 3.643
R2721 VN.n7692 VN.t978 3.643
R2722 VN.n8024 VN.t889 3.643
R2723 VN.n8033 VN.n8032 3.643
R2724 VN.n8030 VN.n8029 3.643
R2725 VN.n8021 VN.t2047 3.643
R2726 VN.n8540 VN.t1917 3.643
R2727 VN.n8557 VN.n8556 3.643
R2728 VN.n8554 VN.n8553 3.643
R2729 VN.n8537 VN.t545 3.643
R2730 VN.n8873 VN.t1756 3.643
R2731 VN.n8882 VN.n8881 3.643
R2732 VN.n8879 VN.n8878 3.643
R2733 VN.n8870 VN.t392 3.643
R2734 VN.n9402 VN.t2103 3.643
R2735 VN.n9419 VN.n9418 3.643
R2736 VN.n9416 VN.n9415 3.643
R2737 VN.n9399 VN.t718 3.643
R2738 VN.n9735 VN.t928 3.643
R2739 VN.n9744 VN.n9743 3.643
R2740 VN.n9741 VN.n9740 3.643
R2741 VN.n9732 VN.t2107 3.643
R2742 VN.n10285 VN.t2070 3.643
R2743 VN.n10302 VN.n10301 3.643
R2744 VN.n10299 VN.n10298 3.643
R2745 VN.n10282 VN.t688 3.643
R2746 VN.n10622 VN.t903 3.643
R2747 VN.n10632 VN.n10631 3.643
R2748 VN.n10629 VN.n10628 3.643
R2749 VN.n10619 VN.t2074 3.643
R2750 VN.n11454 VN.t1186 3.643
R2751 VN.n11470 VN.n11469 3.643
R2752 VN.n11467 VN.n11466 3.643
R2753 VN.n11451 VN.t664 3.643
R2754 VN.n11114 VN.t877 3.643
R2755 VN.n11120 VN.n11119 3.643
R2756 VN.n11123 VN.n11122 3.643
R2757 VN.n11111 VN.t2046 3.643
R2758 VN.n11722 VN.t2398 3.643
R2759 VN.n11723 VN.t1266 3.643
R2760 VN.n12030 VN.t621 3.643
R2761 VN.n12041 VN.n12040 3.643
R2762 VN.n12038 VN.n12037 3.643
R2763 VN.n12033 VN.t1625 3.643
R2764 VN.n2510 VN.t2514 3.643
R2765 VN.n2495 VN.t1127 3.643
R2766 VN.n3025 VN.t1174 3.643
R2767 VN.n3041 VN.n3040 3.643
R2768 VN.n3044 VN.n3043 3.643
R2769 VN.n3022 VN.t2025 3.643
R2770 VN.n3224 VN.t1933 3.643
R2771 VN.n3233 VN.n3232 3.643
R2772 VN.n3230 VN.n3229 3.643
R2773 VN.n3221 VN.t557 3.643
R2774 VN.n3588 VN.t714 3.643
R2775 VN.n3605 VN.n3604 3.643
R2776 VN.n3602 VN.n3601 3.643
R2777 VN.n3585 VN.t1714 3.643
R2778 VN.n3968 VN.t1362 3.643
R2779 VN.n3977 VN.n3976 3.643
R2780 VN.n3974 VN.n3973 3.643
R2781 VN.n3965 VN.t2485 3.643
R2782 VN.n4345 VN.t100 3.643
R2783 VN.n4362 VN.n4361 3.643
R2784 VN.n4359 VN.n4358 3.643
R2785 VN.n4342 VN.t1279 3.643
R2786 VN.n4725 VN.t767 3.643
R2787 VN.n4734 VN.n4733 3.643
R2788 VN.n4731 VN.n4730 3.643
R2789 VN.n4722 VN.t1900 3.643
R2790 VN.n5120 VN.t2079 3.643
R2791 VN.n5137 VN.n5136 3.643
R2792 VN.n5134 VN.n5133 3.643
R2793 VN.n5117 VN.t684 3.643
R2794 VN.n5504 VN.t177 3.643
R2795 VN.n5513 VN.n5512 3.643
R2796 VN.n5510 VN.n5509 3.643
R2797 VN.n5501 VN.t1339 3.643
R2798 VN.n5912 VN.t313 3.643
R2799 VN.n5929 VN.n5928 3.643
R2800 VN.n5926 VN.n5925 3.643
R2801 VN.n5909 VN.t1464 3.643
R2802 VN.n6296 VN.t1242 3.643
R2803 VN.n6305 VN.n6304 3.643
R2804 VN.n6302 VN.n6301 3.643
R2805 VN.n6293 VN.t2106 3.643
R2806 VN.n7155 VN.t2257 3.643
R2807 VN.n7172 VN.n7171 3.643
R2808 VN.n7169 VN.n7168 3.643
R2809 VN.n7152 VN.t854 3.643
R2810 VN.n6741 VN.t658 3.643
R2811 VN.n6750 VN.n6749 3.643
R2812 VN.n6747 VN.n6746 3.643
R2813 VN.n6738 VN.t1784 3.643
R2814 VN.n7544 VN.t1666 3.643
R2815 VN.n7561 VN.n7560 3.643
R2816 VN.n7558 VN.n7557 3.643
R2817 VN.n7541 VN.t287 3.643
R2818 VN.n7932 VN.t185 3.643
R2819 VN.n7941 VN.n7940 3.643
R2820 VN.n7938 VN.n7937 3.643
R2821 VN.n7929 VN.t1217 3.643
R2822 VN.n8389 VN.t1089 3.643
R2823 VN.n8406 VN.n8405 3.643
R2824 VN.n8403 VN.n8402 3.643
R2825 VN.n8386 VN.t2235 3.643
R2826 VN.n8781 VN.t1052 3.643
R2827 VN.n8790 VN.n8789 3.643
R2828 VN.n8787 VN.n8786 3.643
R2829 VN.n8778 VN.t2210 3.643
R2830 VN.n9251 VN.t1948 3.643
R2831 VN.n9268 VN.n9267 3.643
R2832 VN.n9265 VN.n9264 3.643
R2833 VN.n9248 VN.t570 3.643
R2834 VN.n9643 VN.t491 3.643
R2835 VN.n9652 VN.n9651 3.643
R2836 VN.n9649 VN.n9648 3.643
R2837 VN.n9640 VN.t1617 3.643
R2838 VN.n10133 VN.t1382 3.643
R2839 VN.n10150 VN.n10149 3.643
R2840 VN.n10147 VN.n10146 3.643
R2841 VN.n10130 VN.t2502 3.643
R2842 VN.n10520 VN.t2416 3.643
R2843 VN.n10530 VN.n10529 3.643
R2844 VN.n10527 VN.n10526 3.643
R2845 VN.n10517 VN.t1019 3.643
R2846 VN.n11002 VN.t1062 3.643
R2847 VN.n11014 VN.n11013 3.643
R2848 VN.n11011 VN.n11010 3.643
R2849 VN.n10999 VN.t1922 3.643
R2850 VN.n11184 VN.t1830 3.643
R2851 VN.n11190 VN.n11189 3.643
R2852 VN.n11193 VN.n11192 3.643
R2853 VN.n11181 VN.t469 3.643
R2854 VN.n11858 VN.t1529 3.643
R2855 VN.n11859 VN.t397 3.643
R2856 VN.n12053 VN.t2272 3.643
R2857 VN.n12064 VN.n12063 3.643
R2858 VN.n12061 VN.n12060 3.643
R2859 VN.n12056 VN.t867 3.643
R2860 VN.n1818 VN.t2239 3.643
R2861 VN.n1802 VN.t831 3.643
R2862 VN.n2307 VN.t603 3.643
R2863 VN.n2322 VN.n2321 3.643
R2864 VN.n2325 VN.n2324 3.643
R2865 VN.n2310 VN.t1726 3.643
R2866 VN.n2517 VN.t1651 3.643
R2867 VN.n2528 VN.n2527 3.643
R2868 VN.n2525 VN.n2524 3.643
R2869 VN.n2520 VN.t261 3.643
R2870 VN.n2874 VN.t446 3.643
R2871 VN.n2894 VN.n2893 3.643
R2872 VN.n2891 VN.n2890 3.643
R2873 VN.n2877 VN.t1150 3.643
R2874 VN.n3239 VN.t1058 3.643
R2875 VN.n3250 VN.n3249 3.643
R2876 VN.n3247 VN.n3246 3.643
R2877 VN.n3242 VN.t2216 3.643
R2878 VN.n3614 VN.t2369 3.643
R2879 VN.n3634 VN.n3633 3.643
R2880 VN.n3631 VN.n3630 3.643
R2881 VN.n3617 VN.t968 3.643
R2882 VN.n3983 VN.t495 3.643
R2883 VN.n3994 VN.n3993 3.643
R2884 VN.n3991 VN.n3990 3.643
R2885 VN.n3986 VN.t1621 3.643
R2886 VN.n4371 VN.t1772 3.643
R2887 VN.n4391 VN.n4390 3.643
R2888 VN.n4388 VN.n4387 3.643
R2889 VN.n4374 VN.t412 3.643
R2890 VN.n4740 VN.t2421 3.643
R2891 VN.n4751 VN.n4750 3.643
R2892 VN.n4748 VN.n4747 3.643
R2893 VN.n4743 VN.t1025 3.643
R2894 VN.n5146 VN.t2540 3.643
R2895 VN.n5166 VN.n5165 3.643
R2896 VN.n5163 VN.n5162 3.643
R2897 VN.n5149 VN.t1170 3.643
R2898 VN.n5519 VN.t670 3.643
R2899 VN.n5530 VN.n5529 3.643
R2900 VN.n5527 VN.n5526 3.643
R2901 VN.n5522 VN.t1797 3.643
R2902 VN.n5938 VN.t1962 3.643
R2903 VN.n5958 VN.n5957 3.643
R2904 VN.n5955 VN.n5954 3.643
R2905 VN.n5941 VN.t592 3.643
R2906 VN.n6311 VN.t377 3.643
R2907 VN.n6322 VN.n6321 3.643
R2908 VN.n6319 VN.n6318 3.643
R2909 VN.n6314 VN.t1229 3.643
R2910 VN.n7181 VN.t1394 3.643
R2911 VN.n7201 VN.n7200 3.643
R2912 VN.n7198 VN.n7197 3.643
R2913 VN.n7184 VN.t2516 3.643
R2914 VN.n6756 VN.t2431 3.643
R2915 VN.n6767 VN.n6766 3.643
R2916 VN.n6764 VN.n6763 3.643
R2917 VN.n6759 VN.t908 3.643
R2918 VN.n7570 VN.t798 3.643
R2919 VN.n7590 VN.n7589 3.643
R2920 VN.n7587 VN.n7586 3.643
R2921 VN.n7573 VN.t1939 3.643
R2922 VN.n7947 VN.t1842 3.643
R2923 VN.n7958 VN.n7957 3.643
R2924 VN.n7955 VN.n7954 3.643
R2925 VN.n7950 VN.t487 3.643
R2926 VN.n8415 VN.t219 3.643
R2927 VN.n8435 VN.n8434 3.643
R2928 VN.n8432 VN.n8431 3.643
R2929 VN.n8418 VN.t1372 3.643
R2930 VN.n8796 VN.t181 3.643
R2931 VN.n8807 VN.n8806 3.643
R2932 VN.n8804 VN.n8803 3.643
R2933 VN.n8799 VN.t1344 3.643
R2934 VN.n9277 VN.t1079 3.643
R2935 VN.n9297 VN.n9296 3.643
R2936 VN.n9294 VN.n9293 3.643
R2937 VN.n9280 VN.t2229 3.643
R2938 VN.n9658 VN.t2146 3.643
R2939 VN.n9669 VN.n9668 3.643
R2940 VN.n9666 VN.n9665 3.643
R2941 VN.n9661 VN.t748 3.643
R2942 VN.n10159 VN.t516 3.643
R2943 VN.n10179 VN.n10178 3.643
R2944 VN.n10176 VN.n10175 3.643
R2945 VN.n10162 VN.t1640 3.643
R2946 VN.n10536 VN.t1554 3.643
R2947 VN.n10550 VN.n10549 3.643
R2948 VN.n10547 VN.n10546 3.643
R2949 VN.n10539 VN.t149 3.643
R2950 VN.n10557 VN.t680 3.643
R2951 VN.n10571 VN.n10570 3.643
R2952 VN.n10568 VN.n10567 3.643
R2953 VN.n10560 VN.t1812 3.643
R2954 VN.n11050 VN.t1979 3.643
R2955 VN.n11074 VN.n11073 3.643
R2956 VN.n11071 VN.n11070 3.643
R2957 VN.n11053 VN.t315 3.643
R2958 VN.n11148 VN.t36 3.643
R2959 VN.n11156 VN.n11155 3.643
R2960 VN.n11159 VN.n11158 3.643
R2961 VN.n11151 VN.t1244 3.643
R2962 VN.n12070 VN.t1245 3.643
R2963 VN.n12086 VN.n12085 3.643
R2964 VN.n12083 VN.n12082 3.643
R2965 VN.n12073 VN.t2387 3.643
R2966 VN.n11711 VN.t2109 3.643
R2967 VN.n11712 VN.t933 3.643
R2968 VN.n10197 VN.t2285 3.643
R2969 VN.n10214 VN.n10213 3.643
R2970 VN.n10211 VN.n10210 3.643
R2971 VN.n10194 VN.t768 3.643
R2972 VN.n9314 VN.t204 3.643
R2973 VN.n9331 VN.n9330 3.643
R2974 VN.n9328 VN.n9327 3.643
R2975 VN.n9311 VN.t1364 3.643
R2976 VN.n8452 VN.t1869 3.643
R2977 VN.n8469 VN.n8468 3.643
R2978 VN.n8466 VN.n8465 3.643
R2979 VN.n8449 VN.t505 3.643
R2980 VN.n7607 VN.t2453 3.643
R2981 VN.n7624 VN.n7623 3.643
R2982 VN.n7621 VN.n7620 3.643
R2983 VN.n7604 VN.t1068 3.643
R2984 VN.n7218 VN.t529 3.643
R2985 VN.n7235 VN.n7234 3.643
R2986 VN.n7232 VN.n7231 3.643
R2987 VN.n7215 VN.t1654 3.643
R2988 VN.n5975 VN.t1097 3.643
R2989 VN.n5992 VN.n5991 3.643
R2990 VN.n5989 VN.n5988 3.643
R2991 VN.n5972 VN.t2245 3.643
R2992 VN.n5183 VN.t1675 3.643
R2993 VN.n5200 VN.n5199 3.643
R2994 VN.n5197 VN.n5196 3.643
R2995 VN.n5180 VN.t301 3.643
R2996 VN.n4408 VN.t2265 3.643
R2997 VN.n4425 VN.n4424 3.643
R2998 VN.n4422 VN.n4421 3.643
R2999 VN.n4405 VN.t862 3.643
R3000 VN.n3651 VN.t1500 3.643
R3001 VN.n3668 VN.n3667 3.643
R3002 VN.n3665 VN.n3664 3.643
R3003 VN.n3648 VN.t69 3.643
R3004 VN.n2911 VN.t2090 3.643
R3005 VN.n2928 VN.n2927 3.643
R3006 VN.n2925 VN.n2924 3.643
R3007 VN.n2908 VN.t427 3.643
R3008 VN.n2189 VN.t2381 3.643
R3009 VN.n2206 VN.n2205 3.643
R3010 VN.n2203 VN.n2202 3.643
R3011 VN.n2186 VN.t851 3.643
R3012 VN.n1598 VN.t801 3.643
R3013 VN.n1614 VN.n1613 3.643
R3014 VN.n1617 VN.n1616 3.643
R3015 VN.n1595 VN.t1941 3.643
R3016 VN.n1145 VN.t2432 3.643
R3017 VN.n1130 VN.t1043 3.643
R3018 VN.n1827 VN.t1374 3.643
R3019 VN.n1836 VN.n1835 3.643
R3020 VN.n1833 VN.n1832 3.643
R3021 VN.n1824 VN.t2494 3.643
R3022 VN.n2536 VN.t779 3.643
R3023 VN.n2545 VN.n2544 3.643
R3024 VN.n2542 VN.n2541 3.643
R3025 VN.n2533 VN.t1911 3.643
R3026 VN.n3258 VN.t184 3.643
R3027 VN.n3267 VN.n3266 3.643
R3028 VN.n3264 VN.n3263 3.643
R3029 VN.n3255 VN.t1349 3.643
R3030 VN.n4002 VN.t2152 3.643
R3031 VN.n4011 VN.n4010 3.643
R3032 VN.n4008 VN.n4007 3.643
R3033 VN.n3999 VN.t750 3.643
R3034 VN.n4759 VN.t391 3.643
R3035 VN.n4768 VN.n4767 3.643
R3036 VN.n4765 VN.n4764 3.643
R3037 VN.n4756 VN.t1520 3.643
R3038 VN.n5538 VN.t2330 3.643
R3039 VN.n5547 VN.n5546 3.643
R3040 VN.n5544 VN.n5543 3.643
R3041 VN.n5535 VN.t922 3.643
R3042 VN.n6330 VN.t2164 3.643
R3043 VN.n6339 VN.n6338 3.643
R3044 VN.n6336 VN.n6335 3.643
R3045 VN.n6327 VN.t364 3.643
R3046 VN.n6775 VN.t1570 3.643
R3047 VN.n6784 VN.n6783 3.643
R3048 VN.n6781 VN.n6780 3.643
R3049 VN.n6772 VN.t170 3.643
R3050 VN.n7966 VN.t970 3.643
R3051 VN.n7975 VN.n7974 3.643
R3052 VN.n7972 VN.n7971 3.643
R3053 VN.n7963 VN.t2141 3.643
R3054 VN.n8815 VN.t1839 3.643
R3055 VN.n8824 VN.n8823 3.643
R3056 VN.n8821 VN.n8820 3.643
R3057 VN.n8812 VN.t480 3.643
R3058 VN.n9677 VN.t1276 3.643
R3059 VN.n9686 VN.n9685 3.643
R3060 VN.n9683 VN.n9682 3.643
R3061 VN.n9674 VN.t2407 3.643
R3062 VN.n11401 VN.t406 3.643
R3063 VN.n11419 VN.n11418 3.643
R3064 VN.n11416 VN.n11415 3.643
R3065 VN.n11404 VN.t2404 3.643
R3066 VN.n11089 VN.t59 3.643
R3067 VN.n11384 VN.n11383 3.643
R3068 VN.n11387 VN.n11386 3.643
R3069 VN.n11390 VN.t1264 3.643
R3070 VN.n12104 VN.t378 3.643
R3071 VN.n12120 VN.n12119 3.643
R3072 VN.n12117 VN.n12116 3.643
R3073 VN.n12107 VN.t1518 3.643
R3074 VN.n11698 VN.t1232 3.643
R3075 VN.n11699 VN.t9 3.643
R3076 VN.n492 VN.t2165 3.643
R3077 VN.n473 VN.t763 3.643
R3078 VN.n919 VN.t531 3.643
R3079 VN.n927 VN.n926 3.643
R3080 VN.n930 VN.n929 3.643
R3081 VN.n916 VN.t1656 3.643
R3082 VN.n1160 VN.t1572 3.643
R3083 VN.n1168 VN.n1167 3.643
R3084 VN.n1165 VN.n1164 3.643
R3085 VN.n1157 VN.t174 3.643
R3086 VN.n1513 VN.t2577 3.643
R3087 VN.n1531 VN.n1530 3.643
R3088 VN.n1528 VN.n1527 3.643
R3089 VN.n1510 VN.t1070 3.643
R3090 VN.n1850 VN.t508 3.643
R3091 VN.n1858 VN.n1857 3.643
R3092 VN.n1855 VN.n1854 3.643
R3093 VN.n1847 VN.t1628 3.643
R3094 VN.n2221 VN.t1512 3.643
R3095 VN.n2239 VN.n2238 3.643
R3096 VN.n2236 VN.n2235 3.643
R3097 VN.n2218 VN.t93 3.643
R3098 VN.n2559 VN.t2430 3.643
R3099 VN.n2567 VN.n2566 3.643
R3100 VN.n2564 VN.n2563 3.643
R3101 VN.n2556 VN.t1038 3.643
R3102 VN.n2943 VN.t1214 3.643
R3103 VN.n2961 VN.n2960 3.643
R3104 VN.n2958 VN.n2957 3.643
R3105 VN.n2940 VN.t2073 3.643
R3106 VN.n3281 VN.t1841 3.643
R3107 VN.n3289 VN.n3288 3.643
R3108 VN.n3286 VN.n3285 3.643
R3109 VN.n3278 VN.t482 3.643
R3110 VN.n3683 VN.t1973 3.643
R3111 VN.n3701 VN.n3700 3.643
R3112 VN.n3698 VN.n3697 3.643
R3113 VN.n3680 VN.t599 3.643
R3114 VN.n4025 VN.t29 3.643
R3115 VN.n4033 VN.n4032 3.643
R3116 VN.n4030 VN.n4029 3.643
R3117 VN.n4022 VN.t1236 3.643
R3118 VN.n4440 VN.t1400 3.643
R3119 VN.n4458 VN.n4457 3.643
R3120 VN.n4455 VN.n4454 3.643
R3121 VN.n4437 VN.t2524 3.643
R3122 VN.n4782 VN.t2044 3.643
R3123 VN.n4790 VN.n4789 3.643
R3124 VN.n4787 VN.n4786 3.643
R3125 VN.n4779 VN.t652 3.643
R3126 VN.n5215 VN.t809 3.643
R3127 VN.n5233 VN.n5232 3.643
R3128 VN.n5230 VN.n5229 3.643
R3129 VN.n5212 VN.t1949 3.643
R3130 VN.n5561 VN.t1580 3.643
R3131 VN.n5569 VN.n5568 3.643
R3132 VN.n5566 VN.n5565 3.643
R3133 VN.n5558 VN.t2584 3.643
R3134 VN.n6007 VN.t230 3.643
R3135 VN.n6025 VN.n6024 3.643
R3136 VN.n6022 VN.n6021 3.643
R3137 VN.n6004 VN.t1383 3.643
R3138 VN.n6353 VN.t1297 3.643
R3139 VN.n6361 VN.n6360 3.643
R3140 VN.n6358 VN.n6357 3.643
R3141 VN.n6350 VN.t2149 3.643
R3142 VN.n7250 VN.t2184 3.643
R3143 VN.n7268 VN.n7267 3.643
R3144 VN.n7265 VN.n7264 3.643
R3145 VN.n7247 VN.t785 3.643
R3146 VN.n6798 VN.t700 3.643
R3147 VN.n6806 VN.n6805 3.643
R3148 VN.n6803 VN.n6802 3.643
R3149 VN.n6795 VN.t1831 3.643
R3150 VN.n7639 VN.t1591 3.643
R3151 VN.n7657 VN.n7656 3.643
R3152 VN.n7654 VN.n7653 3.643
R3153 VN.n7636 VN.t194 3.643
R3154 VN.n7989 VN.t74 3.643
R3155 VN.n7997 VN.n7996 3.643
R3156 VN.n7994 VN.n7993 3.643
R3157 VN.n7986 VN.t1267 3.643
R3158 VN.n8484 VN.t997 3.643
R3159 VN.n8502 VN.n8501 3.643
R3160 VN.n8499 VN.n8498 3.643
R3161 VN.n8481 VN.t2159 3.643
R3162 VN.n8838 VN.t967 3.643
R3163 VN.n8846 VN.n8845 3.643
R3164 VN.n8843 VN.n8842 3.643
R3165 VN.n8835 VN.t2135 3.643
R3166 VN.n9346 VN.t1992 3.643
R3167 VN.n9364 VN.n9363 3.643
R3168 VN.n9361 VN.n9360 3.643
R3169 VN.n9343 VN.t497 3.643
R3170 VN.n9700 VN.t407 3.643
R3171 VN.n9708 VN.n9707 3.643
R3172 VN.n9705 VN.n9704 3.643
R3173 VN.n9697 VN.t1540 3.643
R3174 VN.n10229 VN.t1416 3.643
R3175 VN.n10247 VN.n10246 3.643
R3176 VN.n10244 VN.n10243 3.643
R3177 VN.n10226 VN.t2543 3.643
R3178 VN.n10585 VN.t2340 3.643
R3179 VN.n10593 VN.n10592 3.643
R3180 VN.n10590 VN.n10589 3.643
R3181 VN.n10582 VN.t937 3.643
R3182 VN.n11428 VN.t2056 3.643
R3183 VN.n11446 VN.n11445 3.643
R3184 VN.n11443 VN.n11442 3.643
R3185 VN.n11431 VN.t1536 3.643
R3186 VN.n11129 VN.t1751 3.643
R3187 VN.n11140 VN.n11139 3.643
R3188 VN.n11143 VN.n11142 3.643
R3189 VN.n11132 VN.t396 3.643
R3190 VN.n10605 VN.t1776 3.643
R3191 VN.n10614 VN.n10613 3.643
R3192 VN.n10611 VN.n10610 3.643
R3193 VN.n10602 VN.t428 3.643
R3194 VN.n10256 VN.t423 3.643
R3195 VN.n10268 VN.n10267 3.643
R3196 VN.n10265 VN.n10264 3.643
R3197 VN.n10259 VN.t1559 3.643
R3198 VN.n9714 VN.t2057 3.643
R3199 VN.n9727 VN.n9726 3.643
R3200 VN.n9724 VN.n9723 3.643
R3201 VN.n9717 VN.t671 3.643
R3202 VN.n9373 VN.t1118 3.643
R3203 VN.n9385 VN.n9384 3.643
R3204 VN.n9382 VN.n9381 3.643
R3205 VN.n9376 VN.t2268 3.643
R3206 VN.n8852 VN.t65 3.643
R3207 VN.n8865 VN.n8864 3.643
R3208 VN.n8862 VN.n8861 3.643
R3209 VN.n8855 VN.t1260 3.643
R3210 VN.n8511 VN.t266 3.643
R3211 VN.n8523 VN.n8522 3.643
R3212 VN.n8520 VN.n8519 3.643
R3213 VN.n8514 VN.t1290 3.643
R3214 VN.n8003 VN.t1760 3.643
R3215 VN.n8016 VN.n8015 3.643
R3216 VN.n8013 VN.n8012 3.643
R3217 VN.n8006 VN.t398 3.643
R3218 VN.n7666 VN.t724 3.643
R3219 VN.n7678 VN.n7677 3.643
R3220 VN.n7675 VN.n7674 3.643
R3221 VN.n7669 VN.t1850 3.643
R3222 VN.n6812 VN.t2357 3.643
R3223 VN.n6825 VN.n6824 3.643
R3224 VN.n6822 VN.n6821 3.643
R3225 VN.n6815 VN.t954 3.643
R3226 VN.n7277 VN.t1319 3.643
R3227 VN.n7289 VN.n7288 3.643
R3228 VN.n7286 VN.n7285 3.643
R3229 VN.n7280 VN.t2439 3.643
R3230 VN.n6367 VN.t431 3.643
R3231 VN.n6380 VN.n6379 3.643
R3232 VN.n6377 VN.n6376 3.643
R3233 VN.n6370 VN.t1280 3.643
R3234 VN.n6034 VN.t1877 3.643
R3235 VN.n6046 VN.n6045 3.643
R3236 VN.n6043 VN.n6042 3.643
R3237 VN.n6037 VN.t518 3.643
R3238 VN.n5575 VN.t715 3.643
R3239 VN.n5588 VN.n5587 3.643
R3240 VN.n5585 VN.n5584 3.643
R3241 VN.n5578 VN.t1840 3.643
R3242 VN.n5242 VN.t2464 3.643
R3243 VN.n5254 VN.n5253 3.643
R3244 VN.n5251 VN.n5250 3.643
R3245 VN.n5245 VN.t1080 3.643
R3246 VN.n4796 VN.t1308 3.643
R3247 VN.n4809 VN.n4808 3.643
R3248 VN.n4806 VN.n4805 3.643
R3249 VN.n4799 VN.t2311 3.643
R3250 VN.n4467 VN.t539 3.643
R3251 VN.n4479 VN.n4478 3.643
R3252 VN.n4476 VN.n4475 3.643
R3253 VN.n4470 VN.t1661 3.643
R3254 VN.n4039 VN.t1738 3.643
R3255 VN.n4052 VN.n4051 3.643
R3256 VN.n4049 VN.n4048 3.643
R3257 VN.n4042 VN.t372 3.643
R3258 VN.n3710 VN.t1105 3.643
R3259 VN.n3722 VN.n3721 3.643
R3260 VN.n3719 VN.n3718 3.643
R3261 VN.n3713 VN.t2254 3.643
R3262 VN.n3295 VN.t2335 3.643
R3263 VN.n3308 VN.n3307 3.643
R3264 VN.n3305 VN.n3304 3.643
R3265 VN.n3298 VN.t930 3.643
R3266 VN.n2970 VN.t1682 3.643
R3267 VN.n2982 VN.n2981 3.643
R3268 VN.n2979 VN.n2978 3.643
R3269 VN.n2973 VN.t2536 3.643
R3270 VN.n2573 VN.t1569 3.643
R3271 VN.n2586 VN.n2585 3.643
R3272 VN.n2583 VN.n2582 3.643
R3273 VN.n2576 VN.t166 3.643
R3274 VN.n2248 VN.t644 3.643
R3275 VN.n2260 VN.n2259 3.643
R3276 VN.n2257 VN.n2256 3.643
R3277 VN.n2251 VN.t1768 3.643
R3278 VN.n1864 VN.t2161 3.643
R3279 VN.n1877 VN.n1876 3.643
R3280 VN.n1874 VN.n1873 3.643
R3281 VN.n1867 VN.t756 3.643
R3282 VN.n1543 VN.t1706 3.643
R3283 VN.n1552 VN.n1551 3.643
R3284 VN.n1534 VN.n1533 3.643
R3285 VN.n1546 VN.t340 3.643
R3286 VN.n1174 VN.t702 3.643
R3287 VN.n1187 VN.n1186 3.643
R3288 VN.n1184 VN.n1183 3.643
R3289 VN.n1177 VN.t1836 3.643
R3290 VN.n857 VN.t2305 3.643
R3291 VN.n869 VN.n868 3.643
R3292 VN.n866 VN.n865 3.643
R3293 VN.n860 VN.t787 3.643
R3294 VN.n499 VN.t1299 3.643
R3295 VN.n512 VN.n511 3.643
R3296 VN.n509 VN.n508 3.643
R3297 VN.n502 VN.t2418 3.643
R3298 VN.n246 VN.t231 3.643
R3299 VN.n255 VN.n254 3.643
R3300 VN.n258 VN.n257 3.643
R3301 VN.n249 VN.t1386 3.643
R3302 VN.n12700 VN.t1856 3.643
R3303 VN.n12683 VN.t493 3.643
R3304 VN.n11685 VN.t367 3.643
R3305 VN.n11686 VN.t1727 3.643
R3306 VN.n12130 VN.t2032 3.643
R3307 VN.n12149 VN.n12148 3.643
R3308 VN.n12146 VN.n12145 3.643
R3309 VN.n12133 VN.t651 3.643
R3310 VN.n11023 VN.t334 3.643
R3311 VN.n11041 VN.n11040 3.643
R3312 VN.n11038 VN.n11037 3.643
R3313 VN.n11026 VN.t1047 3.643
R3314 VN.n11166 VN.t953 3.643
R3315 VN.n11174 VN.n11173 3.643
R3316 VN.n11177 VN.n11176 3.643
R3317 VN.n11169 VN.t2120 3.643
R3318 VN.n11733 VN.t1607 3.643
R3319 VN.n11734 VN.t486 3.643
R3320 VN.n11985 VN.t2232 3.643
R3321 VN.n11996 VN.n11995 3.643
R3322 VN.n11993 VN.n11992 3.643
R3323 VN.n11988 VN.t826 3.643
R3324 VN.n3942 VN.t569 3.643
R3325 VN.n3927 VN.t1694 3.643
R3326 VN.n4522 VN.t1730 3.643
R3327 VN.n4538 VN.n4537 3.643
R3328 VN.n4541 VN.n4540 3.643
R3329 VN.n4519 VN.t363 3.643
R3330 VN.n4691 VN.t2501 3.643
R3331 VN.n4700 VN.n4699 3.643
R3332 VN.n4697 VN.n4696 3.643
R3333 VN.n4688 VN.t1114 3.643
R3334 VN.n5057 VN.t1298 3.643
R3335 VN.n5074 VN.n5073 3.643
R3336 VN.n5071 VN.n5070 3.643
R3337 VN.n5054 VN.t2302 3.643
R3338 VN.n5470 VN.t1921 3.643
R3339 VN.n5479 VN.n5478 3.643
R3340 VN.n5476 VN.n5475 3.643
R3341 VN.n5467 VN.t551 3.643
R3342 VN.n5849 VN.t701 3.643
R3343 VN.n5866 VN.n5865 3.643
R3344 VN.n5863 VN.n5862 3.643
R3345 VN.n5846 VN.t1835 3.643
R3346 VN.n6262 VN.t1624 3.643
R3347 VN.n6271 VN.n6270 3.643
R3348 VN.n6268 VN.n6267 3.643
R3349 VN.n6259 VN.t2476 3.643
R3350 VN.n7092 VN.t77 3.643
R3351 VN.n7109 VN.n7108 3.643
R3352 VN.n7106 VN.n7105 3.643
R3353 VN.n7089 VN.t1270 3.643
R3354 VN.n6707 VN.t1030 3.643
R3355 VN.n6716 VN.n6715 3.643
R3356 VN.n6713 VN.n6712 3.643
R3357 VN.n6704 VN.t2196 3.643
R3358 VN.n7481 VN.t866 3.643
R3359 VN.n7498 VN.n7497 3.643
R3360 VN.n7495 VN.n7494 3.643
R3361 VN.n7478 VN.t2029 3.643
R3362 VN.n7898 VN.t1802 3.643
R3363 VN.n7907 VN.n7906 3.643
R3364 VN.n7904 VN.n7903 3.643
R3365 VN.n7895 VN.t444 3.643
R3366 VN.n8326 VN.t308 3.643
R3367 VN.n8343 VN.n8342 3.643
R3368 VN.n8340 VN.n8339 3.643
R3369 VN.n8323 VN.t1447 3.643
R3370 VN.n8747 VN.t128 3.643
R3371 VN.n8756 VN.n8755 3.643
R3372 VN.n8753 VN.n8752 3.643
R3373 VN.n8744 VN.t1301 3.643
R3374 VN.n9188 VN.t1168 3.643
R3375 VN.n9205 VN.n9204 3.643
R3376 VN.n9202 VN.n9201 3.643
R3377 VN.n9185 VN.t2307 3.643
R3378 VN.n9609 VN.t2223 3.643
R3379 VN.n9618 VN.n9617 3.643
R3380 VN.n9615 VN.n9614 3.643
R3381 VN.n9606 VN.t706 3.643
R3382 VN.n10070 VN.t591 3.643
R3383 VN.n10087 VN.n10086 3.643
R3384 VN.n10084 VN.n10083 3.643
R3385 VN.n10067 VN.t1711 3.643
R3386 VN.n10485 VN.t1631 3.643
R3387 VN.n10495 VN.n10494 3.643
R3388 VN.n10492 VN.n10491 3.643
R3389 VN.n10482 VN.t244 3.643
R3390 VN.n10944 VN.t284 3.643
R3391 VN.n10956 VN.n10955 3.643
R3392 VN.n10953 VN.n10952 3.643
R3393 VN.n10941 VN.t1135 3.643
R3394 VN.n11218 VN.t1041 3.643
R3395 VN.n11224 VN.n11223 3.643
R3396 VN.n11227 VN.n11226 3.643
R3397 VN.n11215 VN.t2200 3.643
R3398 VN.n11834 VN.t741 3.643
R3399 VN.n11835 VN.t2140 3.643
R3400 VN.n12008 VN.t1367 3.643
R3401 VN.n12019 VN.n12018 3.643
R3402 VN.n12016 VN.n12015 3.643
R3403 VN.n12011 VN.t2490 3.643
R3404 VN.n3215 VN.t283 3.643
R3405 VN.n3199 VN.t1424 3.643
R3406 VN.n3769 VN.t1465 3.643
R3407 VN.n3784 VN.n3783 3.643
R3408 VN.n3787 VN.n3786 3.643
R3409 VN.n3772 VN.t2583 3.643
R3410 VN.n3949 VN.t2228 3.643
R3411 VN.n3960 VN.n3959 3.643
R3412 VN.n3957 VN.n3956 3.643
R3413 VN.n3952 VN.t824 3.643
R3414 VN.n4308 VN.t988 3.643
R3415 VN.n4328 VN.n4327 3.643
R3416 VN.n4325 VN.n4324 3.643
R3417 VN.n4311 VN.t2013 3.643
R3418 VN.n4706 VN.t1638 3.643
R3419 VN.n4717 VN.n4716 3.643
R3420 VN.n4714 VN.n4713 3.643
R3421 VN.n4709 VN.t250 3.643
R3422 VN.n5083 VN.t432 3.643
R3423 VN.n5103 VN.n5102 3.643
R3424 VN.n5100 VN.n5099 3.643
R3425 VN.n5086 VN.t1555 3.643
R3426 VN.n5485 VN.t1046 3.643
R3427 VN.n5496 VN.n5495 3.643
R3428 VN.n5493 VN.n5492 3.643
R3429 VN.n5488 VN.t2206 3.643
R3430 VN.n5875 VN.t2360 3.643
R3431 VN.n5895 VN.n5894 3.643
R3432 VN.n5892 VN.n5891 3.643
R3433 VN.n5878 VN.t959 3.643
R3434 VN.n6277 VN.t753 3.643
R3435 VN.n6288 VN.n6287 3.643
R3436 VN.n6285 VN.n6284 3.643
R3437 VN.n6280 VN.t1615 3.643
R3438 VN.n7118 VN.t604 3.643
R3439 VN.n7138 VN.n7137 3.643
R3440 VN.n7135 VN.n7134 3.643
R3441 VN.n7121 VN.t1729 3.643
R3442 VN.n6722 VN.t1526 3.643
R3443 VN.n6733 VN.n6732 3.643
R3444 VN.n6730 VN.n6729 3.643
R3445 VN.n6725 VN.t116 3.643
R3446 VN.n7507 VN.t2530 3.643
R3447 VN.n7527 VN.n7526 3.643
R3448 VN.n7524 VN.n7523 3.643
R3449 VN.n7510 VN.t1155 3.643
R3450 VN.n7913 VN.t926 3.643
R3451 VN.n7924 VN.n7923 3.643
R3452 VN.n7921 VN.n7920 3.643
R3453 VN.n7916 VN.t2091 3.643
R3454 VN.n8352 VN.t1956 3.643
R3455 VN.n8372 VN.n8371 3.643
R3456 VN.n8369 VN.n8368 3.643
R3457 VN.n8355 VN.t577 3.643
R3458 VN.n8762 VN.t1927 3.643
R3459 VN.n8773 VN.n8772 3.643
R3460 VN.n8770 VN.n8769 3.643
R3461 VN.n8765 VN.t435 3.643
R3462 VN.n9214 VN.t299 3.643
R3463 VN.n9234 VN.n9233 3.643
R3464 VN.n9231 VN.n9230 3.643
R3465 VN.n9217 VN.t1437 3.643
R3466 VN.n9624 VN.t1358 3.643
R3467 VN.n9635 VN.n9634 3.643
R3468 VN.n9632 VN.n9631 3.643
R3469 VN.n9627 VN.t2479 3.643
R3470 VN.n10096 VN.t2244 3.643
R3471 VN.n10116 VN.n10115 3.643
R3472 VN.n10113 VN.n10112 3.643
R3473 VN.n10099 VN.t839 3.643
R3474 VN.n10501 VN.t760 3.643
R3475 VN.n10512 VN.n10511 3.643
R3476 VN.n10509 VN.n10508 3.643
R3477 VN.n10504 VN.t1892 3.643
R3478 VN.n10965 VN.t1935 3.643
R3479 VN.n10985 VN.n10984 3.643
R3480 VN.n10982 VN.n10981 3.643
R3481 VN.n10968 VN.t272 3.643
R3482 VN.n11200 VN.t169 3.643
R3483 VN.n11208 VN.n11207 3.643
R3484 VN.n11211 VN.n11210 3.643
R3485 VN.n11203 VN.t1331 3.643
R3486 VN.n11744 VN.t813 3.643
R3487 VN.n11745 VN.t2219 3.643
R3488 VN.n11940 VN.t1442 3.643
R3489 VN.n11951 VN.n11950 3.643
R3490 VN.n11948 VN.n11947 3.643
R3491 VN.n11943 VN.t2566 3.643
R3492 VN.n5444 VN.t1134 3.643
R3493 VN.n5429 VN.t2279 3.643
R3494 VN.n6089 VN.t2318 3.643
R3495 VN.n6105 VN.n6104 3.643
R3496 VN.n6108 VN.n6107 3.643
R3497 VN.n6086 VN.t911 3.643
R3498 VN.n6228 VN.t825 3.643
R3499 VN.n6237 VN.n6236 3.643
R3500 VN.n6234 VN.n6233 3.643
R3501 VN.n6225 VN.t1685 3.643
R3502 VN.n7029 VN.t1844 3.643
R3503 VN.n7046 VN.n7045 3.643
R3504 VN.n7043 VN.n7042 3.643
R3505 VN.n7026 VN.t356 3.643
R3506 VN.n6673 VN.t254 3.643
R3507 VN.n6682 VN.n6681 3.643
R3508 VN.n6679 VN.n6678 3.643
R3509 VN.n6670 VN.t1401 3.643
R3510 VN.n7418 VN.t1287 3.643
R3511 VN.n7435 VN.n7434 3.643
R3512 VN.n7432 VN.n7431 3.643
R3513 VN.n7415 VN.t2409 3.643
R3514 VN.n7864 VN.t2208 3.643
R3515 VN.n7873 VN.n7872 3.643
R3516 VN.n7870 VN.n7869 3.643
R3517 VN.n7861 VN.t810 3.643
R3518 VN.n8263 VN.t691 3.643
R3519 VN.n8280 VN.n8279 3.643
R3520 VN.n8277 VN.n8276 3.643
R3521 VN.n8260 VN.t1819 3.643
R3522 VN.n8713 VN.t548 3.643
R3523 VN.n8722 VN.n8721 3.643
R3524 VN.n8719 VN.n8718 3.643
R3525 VN.n8710 VN.t1669 3.643
R3526 VN.n9125 VN.t386 3.643
R3527 VN.n9142 VN.n9141 3.643
R3528 VN.n9139 VN.n9138 3.643
R3529 VN.n9122 VN.t1516 3.643
R3530 VN.n9575 VN.t1315 3.643
R3531 VN.n9584 VN.n9583 3.643
R3532 VN.n9581 VN.n9580 3.643
R3533 VN.n9572 VN.t2436 3.643
R3534 VN.n10007 VN.t2328 3.643
R3535 VN.n10024 VN.n10023 3.643
R3536 VN.n10021 VN.n10020 3.643
R3537 VN.n10004 VN.t918 3.643
R3538 VN.n10450 VN.t723 3.643
R3539 VN.n10460 VN.n10459 3.643
R3540 VN.n10457 VN.n10456 3.643
R3541 VN.n10447 VN.t1849 3.643
R3542 VN.n10886 VN.t2026 3.643
R3543 VN.n10898 VN.n10897 3.643
R3544 VN.n10895 VN.n10894 3.643
R3545 VN.n10883 VN.t359 3.643
R3546 VN.n11252 VN.t265 3.643
R3547 VN.n11258 VN.n11257 3.643
R3548 VN.n11261 VN.n11260 3.643
R3549 VN.n11249 VN.t1289 3.643
R3550 VN.n11823 VN.t2470 3.643
R3551 VN.n11824 VN.t1354 3.643
R3552 VN.n11963 VN.t574 3.643
R3553 VN.n11974 VN.n11973 3.643
R3554 VN.n11971 VN.n11970 3.643
R3555 VN.n11966 VN.t1696 3.643
R3556 VN.n4682 VN.t838 3.643
R3557 VN.n4666 VN.t1987 3.643
R3558 VN.n5301 VN.t2031 3.643
R3559 VN.n5316 VN.n5315 3.643
R3560 VN.n5319 VN.n5318 3.643
R3561 VN.n5304 VN.t643 3.643
R3562 VN.n5451 VN.t271 3.643
R3563 VN.n5462 VN.n5461 3.643
R3564 VN.n5459 VN.n5458 3.643
R3565 VN.n5454 VN.t1411 3.643
R3566 VN.n5812 VN.t1571 3.643
R3567 VN.n5832 VN.n5831 3.643
R3568 VN.n5829 VN.n5828 3.643
R3569 VN.n5815 VN.t2573 3.643
R3570 VN.n6243 VN.t2489 3.643
R3571 VN.n6254 VN.n6253 3.643
R3572 VN.n6251 VN.n6250 3.643
R3573 VN.n6246 VN.t819 3.643
R3574 VN.n7055 VN.t972 3.643
R3575 VN.n7075 VN.n7074 3.643
R3576 VN.n7072 VN.n7071 3.643
R3577 VN.n7058 VN.t2144 3.643
R3578 VN.n6688 VN.t1904 3.643
R3579 VN.n6699 VN.n6698 3.643
R3580 VN.n6696 VN.n6695 3.643
R3581 VN.n6691 VN.t540 3.643
R3582 VN.n7444 VN.t420 3.643
R3583 VN.n7464 VN.n7463 3.643
R3584 VN.n7461 VN.n7460 3.643
R3585 VN.n7447 VN.t1544 3.643
R3586 VN.n7879 VN.t1343 3.643
R3587 VN.n7890 VN.n7889 3.643
R3588 VN.n7887 VN.n7886 3.643
R3589 VN.n7882 VN.t2465 3.643
R3590 VN.n8289 VN.t1176 3.643
R3591 VN.n8309 VN.n8308 3.643
R3592 VN.n8306 VN.n8305 3.643
R3593 VN.n8292 VN.t2316 3.643
R3594 VN.n8728 VN.t1005 3.643
R3595 VN.n8739 VN.n8738 3.643
R3596 VN.n8736 VN.n8735 3.643
R3597 VN.n8731 VN.t2167 3.643
R3598 VN.n9151 VN.t2040 3.643
R3599 VN.n9171 VN.n9170 3.643
R3600 VN.n9168 VN.n9167 3.643
R3601 VN.n9154 VN.t648 3.643
R3602 VN.n9590 VN.t455 3.643
R3603 VN.n9601 VN.n9600 3.643
R3604 VN.n9598 VN.n9597 3.643
R3605 VN.n9593 VN.t1575 3.643
R3606 VN.n10033 VN.t1463 3.643
R3607 VN.n10053 VN.n10052 3.643
R3608 VN.n10050 VN.n10049 3.643
R3609 VN.n10036 VN.t2580 3.643
R3610 VN.n10466 VN.t2495 3.643
R3611 VN.n10477 VN.n10476 3.643
R3612 VN.n10474 VN.n10473 3.643
R3613 VN.n10469 VN.t977 3.643
R3614 VN.n10907 VN.t1151 3.643
R3615 VN.n10927 VN.n10926 3.643
R3616 VN.n10924 VN.n10923 3.643
R3617 VN.n10910 VN.t2008 3.643
R3618 VN.n11234 VN.t1916 3.643
R3619 VN.n11242 VN.n11241 3.643
R3620 VN.n11245 VN.n11244 3.643
R3621 VN.n11237 VN.t544 3.643
R3622 VN.n6219 VN.t1695 3.643
R3623 VN.n6203 VN.t2554 3.643
R3624 VN.n6654 VN.t1117 3.643
R3625 VN.n6665 VN.n6664 3.643
R3626 VN.n6662 VN.n6661 3.643
R3627 VN.n6657 VN.t2266 3.643
R3628 VN.n7381 VN.t2155 3.643
R3629 VN.n7401 VN.n7400 3.643
R3630 VN.n7398 VN.n7397 3.643
R3631 VN.n7384 VN.t636 3.643
R3632 VN.n7845 VN.t552 3.643
R3633 VN.n7856 VN.n7855 3.643
R3634 VN.n7853 VN.n7852 3.643
R3635 VN.n7848 VN.t1676 3.643
R3636 VN.n8226 VN.t1561 3.643
R3637 VN.n8246 VN.n8245 3.643
R3638 VN.n8243 VN.n8242 3.643
R3639 VN.n8229 VN.t156 3.643
R3640 VN.n8694 VN.t1408 3.643
R3641 VN.n8705 VN.n8704 3.643
R3642 VN.n8702 VN.n8701 3.643
R3643 VN.n8697 VN.t2533 3.643
R3644 VN.n9088 VN.t2417 3.643
R3645 VN.n9108 VN.n9107 3.643
R3646 VN.n9105 VN.n9104 3.643
R3647 VN.n9091 VN.t1020 3.643
R3648 VN.n9556 VN.t815 3.643
R3649 VN.n9567 VN.n9566 3.643
R3650 VN.n9564 VN.n9563 3.643
R3651 VN.n9559 VN.t1959 3.643
R3652 VN.n9970 VN.t668 3.643
R3653 VN.n9990 VN.n9989 3.643
R3654 VN.n9987 VN.n9986 3.643
R3655 VN.n9973 VN.t1793 3.643
R3656 VN.n10431 VN.t1588 3.643
R3657 VN.n10442 VN.n10441 3.643
R3658 VN.n10439 VN.n10438 3.643
R3659 VN.n10434 VN.t191 3.643
R3660 VN.n10849 VN.t373 3.643
R3661 VN.n10869 VN.n10868 3.643
R3662 VN.n10866 VN.n10865 3.643
R3663 VN.n10852 VN.t1224 3.643
R3664 VN.n11267 VN.t996 3.643
R3665 VN.n11275 VN.n11274 3.643
R3666 VN.n11278 VN.n11277 3.643
R3667 VN.n11270 VN.t2158 3.643
R3668 VN.n11914 VN.t2312 3.643
R3669 VN.n11929 VN.n11928 3.643
R3670 VN.n11926 VN.n11925 3.643
R3671 VN.n11917 VN.t904 3.643
R3672 VN.n11861 VN.t1563 3.643
R3673 VN.n11863 VN.t560 3.643
R3674 VN.n11755 VN.t2426 3.643
R3675 VN.n11756 VN.t1307 3.643
R3676 VN.n11891 VN.t653 3.643
R3677 VN.n11902 VN.n11901 3.643
R3678 VN.n11899 VN.n11898 3.643
R3679 VN.n11894 VN.t1779 3.643
R3680 VN.n6647 VN.t1991 3.643
R3681 VN.n6632 VN.t614 3.643
R3682 VN.n7721 VN.t368 3.643
R3683 VN.n7737 VN.n7736 3.643
R3684 VN.n7740 VN.n7739 3.643
R3685 VN.n7718 VN.t1503 3.643
R3686 VN.n7830 VN.t1414 3.643
R3687 VN.n7839 VN.n7838 3.643
R3688 VN.n7836 VN.n7835 3.643
R3689 VN.n7827 VN.t2541 3.643
R3690 VN.n8200 VN.t2423 3.643
R3691 VN.n8217 VN.n8216 3.643
R3692 VN.n8214 VN.n8213 3.643
R3693 VN.n8197 VN.t902 3.643
R3694 VN.n8679 VN.t2276 3.643
R3695 VN.n8688 VN.n8687 3.643
R3696 VN.n8685 VN.n8684 3.643
R3697 VN.n8676 VN.t871 3.643
R3698 VN.n9062 VN.t762 3.643
R3699 VN.n9079 VN.n9078 3.643
R3700 VN.n9076 VN.n9075 3.643
R3701 VN.n9059 VN.t1893 3.643
R3702 VN.n9541 VN.t1681 3.643
R3703 VN.n9550 VN.n9549 3.643
R3704 VN.n9547 VN.n9546 3.643
R3705 VN.n9538 VN.t310 3.643
R3706 VN.n9944 VN.t172 3.643
R3707 VN.n9961 VN.n9960 3.643
R3708 VN.n9958 VN.n9957 3.643
R3709 VN.n9941 VN.t1334 3.643
R3710 VN.n10415 VN.t1104 3.643
R3711 VN.n10425 VN.n10424 3.643
R3712 VN.n10422 VN.n10421 3.643
R3713 VN.n10412 VN.t2253 3.643
R3714 VN.n10828 VN.t1238 3.643
R3715 VN.n10840 VN.n10839 3.643
R3716 VN.n10837 VN.n10836 3.643
R3717 VN.n10825 VN.t2101 3.643
R3718 VN.n11286 VN.t1866 3.643
R3719 VN.n11291 VN.n11290 3.643
R3720 VN.n11294 VN.n11293 3.643
R3721 VN.n11283 VN.t503 3.643
R3722 VN.n11766 VN.t300 3.643
R3723 VN.n11767 VN.t1674 3.643
R3724 VN.n11633 VN.t1027 3.643
R3725 VN.n11644 VN.n11643 3.643
R3726 VN.n11641 VN.n11640 3.643
R3727 VN.n11636 VN.t2191 3.643
R3728 VN.n8653 VN.t1491 3.643
R3729 VN.n8638 VN.t46 3.643
R3730 VN.n9428 VN.t2380 3.643
R3731 VN.n9444 VN.n9443 3.643
R3732 VN.n9447 VN.n9446 3.643
R3733 VN.n9425 VN.t982 3.643
R3734 VN.n9507 VN.t890 3.643
R3735 VN.n9516 VN.n9515 3.643
R3736 VN.n9513 VN.n9512 3.643
R3737 VN.n9504 VN.t2048 3.643
R3738 VN.n9881 VN.t1918 3.643
R3739 VN.n9898 VN.n9897 3.643
R3740 VN.n9895 VN.n9894 3.643
R3741 VN.n9878 VN.t426 3.643
R3742 VN.n10380 VN.t327 3.643
R3743 VN.n10390 VN.n10389 3.643
R3744 VN.n10387 VN.n10386 3.643
R3745 VN.n10377 VN.t1468 3.643
R3746 VN.n10770 VN.t1623 3.643
R3747 VN.n10782 VN.n10781 3.643
R3748 VN.n10779 VN.n10778 3.643
R3749 VN.n10767 VN.t2472 3.643
R3750 VN.n11319 VN.t2264 3.643
R3751 VN.n11325 VN.n11324 3.643
R3752 VN.n11328 VN.n11327 3.643
R3753 VN.n11316 VN.t861 3.643
R3754 VN.n11812 VN.t776 3.643
R3755 VN.n11813 VN.t2174 3.643
R3756 VN.n11870 VN.t1523 3.643
R3757 VN.n11881 VN.n11880 3.643
R3758 VN.n11878 VN.n11877 3.643
R3759 VN.n11873 VN.t111 3.643
R3760 VN.n7821 VN.t2283 3.643
R3761 VN.n7805 VN.t881 3.643
R3762 VN.n8570 VN.t646 3.643
R3763 VN.n8585 VN.n8584 3.643
R3764 VN.n8588 VN.n8587 3.643
R3765 VN.n8573 VN.t1774 3.643
R3766 VN.n8660 VN.t624 3.643
R3767 VN.n8671 VN.n8670 3.643
R3768 VN.n8668 VN.n8667 3.643
R3769 VN.n8663 VN.t1743 3.643
R3770 VN.n9025 VN.t1634 3.643
R3771 VN.n9045 VN.n9044 3.643
R3772 VN.n9042 VN.n9041 3.643
R3773 VN.n9028 VN.t91 3.643
R3774 VN.n9522 VN.t2551 3.643
R3775 VN.n9533 VN.n9532 3.643
R3776 VN.n9530 VN.n9529 3.643
R3777 VN.n9525 VN.t1180 3.643
R3778 VN.n9907 VN.t1042 3.643
R3779 VN.n9927 VN.n9926 3.643
R3780 VN.n9924 VN.n9923 3.643
R3781 VN.n9910 VN.t2201 3.643
R3782 VN.n10396 VN.t1972 3.643
R3783 VN.n10407 VN.n10406 3.643
R3784 VN.n10404 VN.n10403 3.643
R3785 VN.n10399 VN.t598 3.643
R3786 VN.n10791 VN.t751 3.643
R3787 VN.n10811 VN.n10810 3.643
R3788 VN.n10808 VN.n10807 3.643
R3789 VN.n10794 VN.t1610 3.643
R3790 VN.n11301 VN.t1399 3.643
R3791 VN.n11309 VN.n11308 3.643
R3792 VN.n11312 VN.n11311 3.643
R3793 VN.n11304 VN.t2523 3.643
R3794 VN.n11775 VN.t2041 3.643
R3795 VN.n11776 VN.t880 3.643
R3796 VN.n11588 VN.t252 3.643
R3797 VN.n11599 VN.n11598 3.643
R3798 VN.n11596 VN.n11595 3.643
R3799 VN.n11591 VN.t1278 3.643
R3800 VN.n10354 VN.t2066 3.643
R3801 VN.n10339 VN.t673 3.643
R3802 VN.n11479 VN.t713 3.643
R3803 VN.n11491 VN.n11490 3.643
R3804 VN.n11494 VN.n11493 3.643
R3805 VN.n11476 VN.t1566 3.643
R3806 VN.n11353 VN.t1481 3.643
R3807 VN.n11359 VN.n11358 3.643
R3808 VN.n11362 VN.n11361 3.643
R3809 VN.n11350 VN.t21 3.643
R3810 VN.n11801 VN.t1169 3.643
R3811 VN.n11802 VN.t2539 3.643
R3812 VN.n11611 VN.t1902 3.643
R3813 VN.n11622 VN.n11621 3.643
R3814 VN.n11619 VN.n11618 3.643
R3815 VN.n11614 VN.t536 3.643
R3816 VN.n9498 VN.t1761 3.643
R3817 VN.n9482 VN.t400 3.643
R3818 VN.n10315 VN.t121 3.643
R3819 VN.n10330 VN.n10329 3.643
R3820 VN.n10333 VN.n10332 3.643
R3821 VN.n10318 VN.t1293 3.643
R3822 VN.n10361 VN.t1196 3.643
R3823 VN.n10372 VN.n10371 3.643
R3824 VN.n10369 VN.n10368 3.643
R3825 VN.n10364 VN.t2332 3.643
R3826 VN.n10733 VN.t2487 3.643
R3827 VN.n10753 VN.n10752 3.643
R3828 VN.n10750 VN.n10749 3.643
R3829 VN.n10736 VN.t696 3.643
R3830 VN.n11335 VN.t613 3.643
R3831 VN.n11343 VN.n11342 3.643
R3832 VN.n11346 VN.n11345 3.643
R3833 VN.n11338 VN.t1735 3.643
R3834 VN.n11544 VN.t1440 3.643
R3835 VN.n11093 VN.t135 3.643
R3836 VN.n11105 VN.n11104 3.643
R3837 VN.n11102 VN.n11101 3.643
R3838 VN.n11096 VN.t1178 3.643
R3839 VN.n11499 VN.t317 3.643
R3840 VN.n11508 VN.n11507 3.643
R3841 VN.n11511 VN.n11510 3.643
R3842 VN.n11502 VN.t2326 3.643
R3843 VN.n10337 VN.t2564 3.643
R3844 VN.n10652 VN.n10651 3.643
R3845 VN.n10655 VN.n10654 3.643
R3846 VN.n10658 VN.t1202 3.643
R3847 VN.n10665 VN.t1198 3.643
R3848 VN.n10678 VN.n10677 3.643
R3849 VN.n10681 VN.n10680 3.643
R3850 VN.n10668 VN.t2346 3.643
R3851 VN.n9750 VN.t1 3.643
R3852 VN.n9759 VN.n9758 3.643
R3853 VN.n9762 VN.n9761 3.643
R3854 VN.n9753 VN.t1230 3.643
R3855 VN.n9451 VN.t1226 3.643
R3856 VN.n9464 VN.n9463 3.643
R3857 VN.n9467 VN.n9466 3.643
R3858 VN.n9454 VN.t2372 3.643
R3859 VN.n8888 VN.t40 3.643
R3860 VN.n8897 VN.n8896 3.643
R3861 VN.n8900 VN.n8899 3.643
R3862 VN.n8891 VN.t1261 3.643
R3863 VN.n8592 VN.t948 3.643
R3864 VN.n8605 VN.n8604 3.643
R3865 VN.n8608 VN.n8607 3.643
R3866 VN.n8595 VN.t2124 3.643
R3867 VN.n8039 VN.t2550 3.643
R3868 VN.n8048 VN.n8047 3.643
R3869 VN.n8051 VN.n8050 3.643
R3870 VN.n8042 VN.t1179 3.643
R3871 VN.n7744 VN.t1633 3.643
R3872 VN.n7757 VN.n7756 3.643
R3873 VN.n7760 VN.n7759 3.643
R3874 VN.n7747 VN.t245 3.643
R3875 VN.n6848 VN.t623 3.643
R3876 VN.n6857 VN.n6856 3.643
R3877 VN.n6860 VN.n6859 3.643
R3878 VN.n6851 VN.t1741 3.643
R3879 VN.n6996 VN.t2224 3.643
R3880 VN.n7012 VN.n7011 3.643
R3881 VN.n7009 VN.n7008 3.643
R3882 VN.n6999 VN.t707 3.643
R3883 VN.n6403 VN.t1204 3.643
R3884 VN.n6412 VN.n6411 3.643
R3885 VN.n6415 VN.n6414 3.643
R3886 VN.n6406 VN.t2061 3.643
R3887 VN.n6112 VN.t133 3.643
R3888 VN.n6125 VN.n6124 3.643
R3889 VN.n6128 VN.n6127 3.643
R3890 VN.n6115 VN.t1302 3.643
R3891 VN.n5611 VN.t1501 3.643
R3892 VN.n5620 VN.n5619 3.643
R3893 VN.n5623 VN.n5622 3.643
R3894 VN.n5614 VN.t70 3.643
R3895 VN.n5323 VN.t733 3.643
R3896 VN.n5336 VN.n5335 3.643
R3897 VN.n5339 VN.n5338 3.643
R3898 VN.n5326 VN.t1859 3.643
R3899 VN.n4832 VN.t2093 3.643
R3900 VN.n4841 VN.n4840 3.643
R3901 VN.n4844 VN.n4843 3.643
R3902 VN.n4835 VN.t694 3.643
R3903 VN.n4545 VN.t1325 3.643
R3904 VN.n4558 VN.n4557 3.643
R3905 VN.n4561 VN.n4560 3.643
R3906 VN.n4548 VN.t2448 3.643
R3907 VN.n4075 VN.t117 3.643
R3908 VN.n4084 VN.n4083 3.643
R3909 VN.n4087 VN.n4086 3.643
R3910 VN.n4078 VN.t1291 3.643
R3911 VN.n3791 VN.t1888 3.643
R3912 VN.n3804 VN.n3803 3.643
R3913 VN.n3807 VN.n3806 3.643
R3914 VN.n3794 VN.t524 3.643
R3915 VN.n3331 VN.t725 3.643
R3916 VN.n3340 VN.n3339 3.643
R3917 VN.n3343 VN.n3342 3.643
R3918 VN.n3334 VN.t1725 3.643
R3919 VN.n3048 VN.t2473 3.643
R3920 VN.n3061 VN.n3060 3.643
R3921 VN.n3064 VN.n3063 3.643
R3922 VN.n3051 VN.t805 3.643
R3923 VN.n2609 VN.t1183 3.643
R3924 VN.n2618 VN.n2617 3.643
R3925 VN.n2621 VN.n2620 3.643
R3926 VN.n2612 VN.t2322 3.643
R3927 VN.n2329 VN.t249 3.643
R3928 VN.n2342 VN.n2341 3.643
R3929 VN.n2345 VN.n2344 3.643
R3930 VN.n2332 VN.t1396 3.643
R3931 VN.n1900 VN.t1749 3.643
R3932 VN.n1909 VN.n1908 3.643
R3933 VN.n1912 VN.n1911 3.643
R3934 VN.n1903 VN.t382 3.643
R3935 VN.n1621 VN.t1342 3.643
R3936 VN.n1634 VN.n1633 3.643
R3937 VN.n1637 VN.n1636 3.643
R3938 VN.n1624 VN.t2462 3.643
R3939 VN.n1210 VN.t1493 3.643
R3940 VN.n1219 VN.n1218 3.643
R3941 VN.n1222 VN.n1221 3.643
R3942 VN.n1213 VN.t54 3.643
R3943 VN.n934 VN.t567 3.643
R3944 VN.n947 VN.n946 3.643
R3945 VN.n950 VN.n949 3.643
R3946 VN.n937 VN.t1692 3.643
R3947 VN.n535 VN.t2080 3.643
R3948 VN.n544 VN.n543 3.643
R3949 VN.n547 VN.n546 3.643
R3950 VN.n538 VN.t685 3.643
R3951 VN.n262 VN.t1145 3.643
R3952 VN.n275 VN.n274 3.643
R3953 VN.n278 VN.n277 3.643
R3954 VN.n265 VN.t2289 3.643
R3955 VN.n12286 VN.t102 3.643
R3956 VN.n12289 VN.n12288 3.643
R3957 VN.n12292 VN.n12291 3.643
R3958 VN.n12295 VN.t1282 3.643
R3959 VN.n12303 VN.t1720 3.643
R3960 VN.n12316 VN.n12315 3.643
R3961 VN.n12319 VN.n12318 3.643
R3962 VN.n12306 VN.t211 3.643
R3963 VN.n12268 VN.t716 3.643
R3964 VN.n12271 VN.n12270 3.643
R3965 VN.n12274 VN.n12273 3.643
R3966 VN.n12277 VN.t1567 3.643
R3967 VN.n107 VN.t2198 3.643
R3968 VN.n11518 VN.t1460 3.643
R3969 VN.n10638 VN.t1822 3.643
R3970 VN.n10646 VN.n10645 3.643
R3971 VN.n10649 VN.n10648 3.643
R3972 VN.n10641 VN.t336 3.643
R3973 VN.n10689 VN.t330 3.643
R3974 VN.n10693 VN.n10692 3.643
R3975 VN.n10696 VN.n10695 3.643
R3976 VN.n10686 VN.t1478 3.643
R3977 VN.n111 VN.t1448 3.643
R3978 VN.n12628 VN.t2371 3.643
R3979 VN.n12625 VN.n12624 3.643
R3980 VN.n12622 VN.n12621 3.643
R3981 VN.n12348 VN.t697 3.643
R3982 VN.n12327 VN.t847 3.643
R3983 VN.n12634 VN.n12633 3.643
R3984 VN.n12637 VN.n12636 3.643
R3985 VN.n12324 VN.t1996 3.643
R3986 VN.n12341 VN.t1773 3.643
R3987 VN.n12338 VN.n12337 3.643
R3988 VN.n12335 VN.n12334 3.643
R3989 VN.n12332 VN.t414 3.643
R3990 VN.n286 VN.t282 3.643
R3991 VN.n290 VN.n289 3.643
R3992 VN.n293 VN.n292 3.643
R3993 VN.n283 VN.t1420 3.643
R3994 VN.n555 VN.t1207 3.643
R3995 VN.n560 VN.n559 3.643
R3996 VN.n563 VN.n562 3.643
R3997 VN.n552 VN.t2344 3.643
R3998 VN.n958 VN.t1028 3.643
R3999 VN.n962 VN.n961 3.643
R4000 VN.n965 VN.n964 3.643
R4001 VN.n955 VN.t2194 3.643
R4002 VN.n1230 VN.t1964 3.643
R4003 VN.n1235 VN.n1234 3.643
R4004 VN.n1238 VN.n1237 3.643
R4005 VN.n1227 VN.t593 3.643
R4006 VN.n1645 VN.t479 3.643
R4007 VN.n1649 VN.n1648 3.643
R4008 VN.n1652 VN.n1651 3.643
R4009 VN.n1642 VN.t1596 3.643
R4010 VN.n1920 VN.t876 3.643
R4011 VN.n1925 VN.n1924 3.643
R4012 VN.n1928 VN.n1927 3.643
R4013 VN.n1917 VN.t2036 3.643
R4014 VN.n2353 VN.t1899 3.643
R4015 VN.n2357 VN.n2356 3.643
R4016 VN.n2360 VN.n2359 3.643
R4017 VN.n2350 VN.t534 3.643
R4018 VN.n2629 VN.t458 3.643
R4019 VN.n2634 VN.n2633 3.643
R4020 VN.n2637 VN.n2636 3.643
R4021 VN.n2626 VN.t1455 3.643
R4022 VN.n3072 VN.t1612 3.643
R4023 VN.n3076 VN.n3075 3.643
R4024 VN.n3079 VN.n3078 3.643
R4025 VN.n3069 VN.t2458 3.643
R4026 VN.n3351 VN.t2377 3.643
R4027 VN.n3356 VN.n3355 3.643
R4028 VN.n3359 VN.n3358 3.643
R4029 VN.n3348 VN.t979 3.643
R4030 VN.n3815 VN.t1016 3.643
R4031 VN.n3819 VN.n3818 3.643
R4032 VN.n3822 VN.n3821 3.643
R4033 VN.n3812 VN.t2179 3.643
R4034 VN.n4095 VN.t1785 3.643
R4035 VN.n4100 VN.n4099 3.643
R4036 VN.n4103 VN.n4102 3.643
R4037 VN.n4092 VN.t424 3.643
R4038 VN.n4569 VN.t463 3.643
R4039 VN.n4573 VN.n4572 3.643
R4040 VN.n4576 VN.n4575 3.643
R4041 VN.n4566 VN.t1583 3.643
R4042 VN.n4852 VN.t1216 3.643
R4043 VN.n4857 VN.n4856 3.643
R4044 VN.n4860 VN.n4859 3.643
R4045 VN.n4849 VN.t2353 3.643
R4046 VN.n5347 VN.t2386 3.643
R4047 VN.n5351 VN.n5350 3.643
R4048 VN.n5354 VN.n5353 3.643
R4049 VN.n5344 VN.t990 3.643
R4050 VN.n5631 VN.t634 3.643
R4051 VN.n5636 VN.n5635 3.643
R4052 VN.n5639 VN.n5638 3.643
R4053 VN.n5628 VN.t1758 3.643
R4054 VN.n6136 VN.t1929 3.643
R4055 VN.n6140 VN.n6139 3.643
R4056 VN.n6143 VN.n6142 3.643
R4057 VN.n6133 VN.t436 3.643
R4058 VN.n6423 VN.t339 3.643
R4059 VN.n6428 VN.n6427 3.643
R4060 VN.n6431 VN.n6430 3.643
R4061 VN.n6420 VN.t1190 3.643
R4062 VN.n6985 VN.t1359 3.643
R4063 VN.n6992 VN.n6991 3.643
R4064 VN.n6989 VN.n6988 3.643
R4065 VN.n6982 VN.t2480 3.643
R4066 VN.n6868 VN.t2274 3.643
R4067 VN.n6873 VN.n6872 3.643
R4068 VN.n6876 VN.n6875 3.643
R4069 VN.n6865 VN.t869 3.643
R4070 VN.n7768 VN.t81 3.643
R4071 VN.n7772 VN.n7771 3.643
R4072 VN.n7775 VN.n7774 3.643
R4073 VN.n7765 VN.t1281 3.643
R4074 VN.n8059 VN.t1499 3.643
R4075 VN.n8064 VN.n8063 3.643
R4076 VN.n8067 VN.n8066 3.643
R4077 VN.n8056 VN.t85 3.643
R4078 VN.n8616 VN.t27 3.643
R4079 VN.n8620 VN.n8619 3.643
R4080 VN.n8623 VN.n8622 3.643
R4081 VN.n8613 VN.t1249 3.643
R4082 VN.n8908 VN.t1742 3.643
R4083 VN.n8913 VN.n8912 3.643
R4084 VN.n8916 VN.n8915 3.643
R4085 VN.n8905 VN.t393 3.643
R4086 VN.n9475 VN.t360 3.643
R4087 VN.n9798 VN.n9797 3.643
R4088 VN.n9801 VN.n9800 3.643
R4089 VN.n9472 VN.t1504 3.643
R4090 VN.n9793 VN.t1722 3.643
R4091 VN.n9790 VN.n9789 3.643
R4092 VN.n9787 VN.n9786 3.643
R4093 VN.n9480 VN.t365 3.643
R4094 VN.n9864 VN.t610 3.643
R4095 VN.n9767 VN.t974 3.643
R4096 VN.n9781 VN.n9780 3.643
R4097 VN.n9784 VN.n9783 3.643
R4098 VN.n9770 VN.t2015 3.643
R4099 VN.n9809 VN.t2009 3.643
R4100 VN.n9813 VN.n9812 3.643
R4101 VN.n9816 VN.n9815 3.643
R4102 VN.n9806 VN.t638 3.643
R4103 VN.n115 VN.t579 3.643
R4104 VN.n12419 VN.t1502 3.643
R4105 VN.n12424 VN.n12423 3.643
R4106 VN.n12427 VN.n12426 3.643
R4107 VN.n12416 VN.t2356 3.643
R4108 VN.n12645 VN.t2512 3.643
R4109 VN.n12665 VN.n12664 3.643
R4110 VN.n12668 VN.n12667 3.643
R4111 VN.n12642 VN.t1124 3.643
R4112 VN.n12659 VN.t900 3.643
R4113 VN.n12656 VN.n12655 3.643
R4114 VN.n12653 VN.n12652 3.643
R4115 VN.n12650 VN.t2062 3.643
R4116 VN.n301 VN.t752 3.643
R4117 VN.n305 VN.n304 3.643
R4118 VN.n308 VN.n307 3.643
R4119 VN.n298 VN.t1886 3.643
R4120 VN.n571 VN.t1677 3.643
R4121 VN.n576 VN.n575 3.643
R4122 VN.n579 VN.n578 3.643
R4123 VN.n568 VN.t302 3.643
R4124 VN.n973 VN.t157 3.643
R4125 VN.n977 VN.n976 3.643
R4126 VN.n980 VN.n979 3.643
R4127 VN.n970 VN.t1324 3.643
R4128 VN.n1246 VN.t1098 3.643
R4129 VN.n1251 VN.n1250 3.643
R4130 VN.n1254 VN.n1253 3.643
R4131 VN.n1243 VN.t2246 3.643
R4132 VN.n1660 VN.t2134 3.643
R4133 VN.n1664 VN.n1663 3.643
R4134 VN.n1667 VN.n1666 3.643
R4135 VN.n1657 VN.t731 3.643
R4136 VN.n1936 VN.t134 3.643
R4137 VN.n1941 VN.n1940 3.643
R4138 VN.n1944 VN.n1943 3.643
R4139 VN.n1933 VN.t1162 3.643
R4140 VN.n2368 VN.t1024 3.643
R4141 VN.n2372 VN.n2371 3.643
R4142 VN.n2375 VN.n2374 3.643
R4143 VN.n2365 VN.t2189 3.643
R4144 VN.n2645 VN.t2104 3.643
R4145 VN.n2650 VN.n2649 3.643
R4146 VN.n2653 VN.n2652 3.643
R4147 VN.n2642 VN.t708 3.643
R4148 VN.n3087 VN.t745 3.643
R4149 VN.n3091 VN.n3090 3.643
R4150 VN.n3094 VN.n3093 3.643
R4151 VN.n3084 VN.t1593 3.643
R4152 VN.n3367 VN.t1510 3.643
R4153 VN.n3372 VN.n3371 3.643
R4154 VN.n3375 VN.n3374 3.643
R4155 VN.n3364 VN.t87 3.643
R4156 VN.n3830 VN.t142 3.643
R4157 VN.n3834 VN.n3833 3.643
R4158 VN.n3837 VN.n3836 3.643
R4159 VN.n3827 VN.t1311 3.643
R4160 VN.n4111 VN.t907 3.643
R4161 VN.n4116 VN.n4115 3.643
R4162 VN.n4119 VN.n4118 3.643
R4163 VN.n4108 VN.t2069 3.643
R4164 VN.n4584 VN.t2112 3.643
R4165 VN.n4588 VN.n4587 3.643
R4166 VN.n4591 VN.n4590 3.643
R4167 VN.n4581 VN.t719 3.643
R4168 VN.n4868 VN.t354 3.643
R4169 VN.n4873 VN.n4872 3.643
R4170 VN.n4876 VN.n4875 3.643
R4171 VN.n4865 VN.t1485 3.643
R4172 VN.n5362 VN.t1645 3.643
R4173 VN.n5366 VN.n5365 3.643
R4174 VN.n5369 VN.n5368 3.643
R4175 VN.n5359 VN.t105 3.643
R4176 VN.n5647 VN.t2291 3.643
R4177 VN.n5652 VN.n5651 3.643
R4178 VN.n5655 VN.n5654 3.643
R4179 VN.n5644 VN.t885 3.643
R4180 VN.n6151 VN.t1054 3.643
R4181 VN.n6155 VN.n6154 3.643
R4182 VN.n6158 VN.n6157 3.643
R4183 VN.n6148 VN.t2211 3.643
R4184 VN.n6439 VN.t1982 3.643
R4185 VN.n6444 VN.n6443 3.643
R4186 VN.n6447 VN.n6446 3.643
R4187 VN.n6436 VN.t320 3.643
R4188 VN.n6970 VN.t1789 3.643
R4189 VN.n6977 VN.n6976 3.643
R4190 VN.n6974 VN.n6973 3.643
R4191 VN.n6967 VN.t445 3.643
R4192 VN.n6884 VN.t657 3.643
R4193 VN.n6889 VN.n6888 3.643
R4194 VN.n6892 VN.n6891 3.643
R4195 VN.n6881 VN.t1794 3.643
R4196 VN.n7783 VN.t1763 3.643
R4197 VN.n7787 VN.n7786 3.643
R4198 VN.n7790 VN.n7789 3.643
R4199 VN.n7780 VN.t415 3.643
R4200 VN.n8075 VN.t633 3.643
R4201 VN.n8080 VN.n8079 3.643
R4202 VN.n8083 VN.n8082 3.643
R4203 VN.n8072 VN.t1764 3.643
R4204 VN.n8631 VN.t1737 3.643
R4205 VN.n8952 VN.n8951 3.643
R4206 VN.n8955 VN.n8954 3.643
R4207 VN.n8628 VN.t381 3.643
R4208 VN.n8947 VN.t870 3.643
R4209 VN.n8944 VN.n8943 3.643
R4210 VN.n8941 VN.n8940 3.643
R4211 VN.n8636 VN.t2045 3.643
R4212 VN.n9016 VN.t2295 3.643
R4213 VN.n8921 VN.t124 3.643
R4214 VN.n8935 VN.n8934 3.643
R4215 VN.n8938 VN.n8937 3.643
R4216 VN.n8924 VN.t1175 3.643
R4217 VN.n8963 VN.t865 3.643
R4218 VN.n8967 VN.n8966 3.643
R4219 VN.n8970 VN.n8969 3.643
R4220 VN.n8960 VN.t2035 3.643
R4221 VN.n119 VN.t2237 3.643
R4222 VN.n12435 VN.t635 3.643
R4223 VN.n12440 VN.n12439 3.643
R4224 VN.n12443 VN.n12442 3.643
R4225 VN.n12432 VN.t1488 3.643
R4226 VN.n12676 VN.t489 3.643
R4227 VN.n12776 VN.n12775 3.643
R4228 VN.n12779 VN.n12778 3.643
R4229 VN.n12673 VN.t1611 3.643
R4230 VN.n12770 VN.t1402 3.643
R4231 VN.n12767 VN.n12766 3.643
R4232 VN.n12764 VN.n12763 3.643
R4233 VN.n12681 VN.t2525 3.643
R4234 VN.n316 VN.t2410 3.643
R4235 VN.n320 VN.n319 3.643
R4236 VN.n323 VN.n322 3.643
R4237 VN.n313 VN.t1014 3.643
R4238 VN.n587 VN.t811 3.643
R4239 VN.n592 VN.n591 3.643
R4240 VN.n595 VN.n594 3.643
R4241 VN.n584 VN.t1950 3.643
R4242 VN.n988 VN.t1820 3.643
R4243 VN.n992 VN.n991 3.643
R4244 VN.n995 VN.n994 3.643
R4245 VN.n985 VN.t462 3.643
R4246 VN.n1262 VN.t366 3.643
R4247 VN.n1267 VN.n1266 3.643
R4248 VN.n1270 VN.n1269 3.643
R4249 VN.n1259 VN.t1384 3.643
R4250 VN.n1675 VN.t1258 3.643
R4251 VN.n1679 VN.n1678 3.643
R4252 VN.n1682 VN.n1681 3.643
R4253 VN.n1672 VN.t2385 3.643
R4254 VN.n1952 VN.t1796 3.643
R4255 VN.n1957 VN.n1956 3.643
R4256 VN.n1960 VN.n1959 3.643
R4257 VN.n1949 VN.t437 3.643
R4258 VN.n2383 VN.t152 3.643
R4259 VN.n2387 VN.n2386 3.643
R4260 VN.n2390 VN.n2389 3.643
R4261 VN.n2380 VN.t1322 3.643
R4262 VN.n2661 VN.t1227 3.643
R4263 VN.n2666 VN.n2665 3.643
R4264 VN.n2669 VN.n2668 3.643
R4265 VN.n2658 VN.t2364 3.643
R4266 VN.n3102 VN.t2402 3.643
R4267 VN.n3106 VN.n3105 3.643
R4268 VN.n3109 VN.n3108 3.643
R4269 VN.n3099 VN.t728 3.643
R4270 VN.n3383 VN.t641 3.643
R4271 VN.n3388 VN.n3387 3.643
R4272 VN.n3391 VN.n3390 3.643
R4273 VN.n3380 VN.t1765 3.643
R4274 VN.n3845 VN.t1805 3.643
R4275 VN.n3849 VN.n3848 3.643
R4276 VN.n3852 VN.n3851 3.643
R4277 VN.n3842 VN.t450 3.643
R4278 VN.n4127 VN.t2570 3.643
R4279 VN.n4132 VN.n4131 3.643
R4280 VN.n4135 VN.n4134 3.643
R4281 VN.n4124 VN.t1199 3.643
R4282 VN.n4599 VN.t1368 3.643
R4283 VN.n4603 VN.n4602 3.643
R4284 VN.n4606 VN.n4605 3.643
R4285 VN.n4596 VN.t2373 3.643
R4286 VN.n4884 VN.t1999 3.643
R4287 VN.n4889 VN.n4888 3.643
R4288 VN.n4892 VN.n4891 3.643
R4289 VN.n4881 VN.t618 3.643
R4290 VN.n5377 VN.t774 3.643
R4291 VN.n5381 VN.n5380 3.643
R4292 VN.n5384 VN.n5383 3.643
R4293 VN.n5374 VN.t1905 3.643
R4294 VN.n5663 VN.t1422 3.643
R4295 VN.n5668 VN.n5667 3.643
R4296 VN.n5671 VN.n5670 3.643
R4297 VN.n5660 VN.t2546 3.643
R4298 VN.n6166 VN.t943 3.643
R4299 VN.n6170 VN.n6169 3.643
R4300 VN.n6173 VN.n6172 3.643
R4301 VN.n6163 VN.t2118 3.643
R4302 VN.n6455 VN.t2339 3.643
R4303 VN.n6460 VN.n6459 3.643
R4304 VN.n6463 VN.n6462 3.643
R4305 VN.n6452 VN.t1807 3.643
R4306 VN.n6955 VN.t914 3.643
R4307 VN.n6962 VN.n6961 3.643
R4308 VN.n6959 VN.n6958 3.643
R4309 VN.n6952 VN.t2092 3.643
R4310 VN.n6900 VN.t2317 3.643
R4311 VN.n6905 VN.n6904 3.643
R4312 VN.n6908 VN.n6907 3.643
R4313 VN.n6897 VN.t919 3.643
R4314 VN.n7798 VN.t891 3.643
R4315 VN.n8119 VN.n8118 3.643
R4316 VN.n8122 VN.n8121 3.643
R4317 VN.n7795 VN.t2063 3.643
R4318 VN.n8114 VN.t2290 3.643
R4319 VN.n8111 VN.n8110 3.643
R4320 VN.n8108 VN.n8107 3.643
R4321 VN.n7803 VN.t893 3.643
R4322 VN.n8183 VN.t1160 3.643
R4323 VN.n8088 VN.t1542 3.643
R4324 VN.n8102 VN.n8101 3.643
R4325 VN.n8105 VN.n8104 3.643
R4326 VN.n8091 VN.t2555 3.643
R4327 VN.n8130 VN.t2553 3.643
R4328 VN.n8134 VN.n8133 3.643
R4329 VN.n8137 VN.n8136 3.643
R4330 VN.n8127 VN.t1191 3.643
R4331 VN.n123 VN.t173 3.643
R4332 VN.n12451 VN.t1106 3.643
R4333 VN.n12456 VN.n12455 3.643
R4334 VN.n12459 VN.n12458 3.643
R4335 VN.n12448 VN.t1960 3.643
R4336 VN.n12790 VN.t2143 3.643
R4337 VN.n12810 VN.n12809 3.643
R4338 VN.n12787 VN.n12786 3.643
R4339 VN.n12784 VN.t744 3.643
R4340 VN.n12804 VN.t541 3.643
R4341 VN.n12801 VN.n12800 3.643
R4342 VN.n12798 VN.n12797 3.643
R4343 VN.n12795 VN.t1662 3.643
R4344 VN.n331 VN.t1545 3.643
R4345 VN.n335 VN.n334 3.643
R4346 VN.n338 VN.n337 3.643
R4347 VN.n328 VN.t140 3.643
R4348 VN.n603 VN.t2587 3.643
R4349 VN.n608 VN.n607 3.643
R4350 VN.n611 VN.n610 3.643
R4351 VN.n600 VN.t1081 3.643
R4352 VN.n1003 VN.t947 3.643
R4353 VN.n1007 VN.n1006 3.643
R4354 VN.n1010 VN.n1009 3.643
R4355 VN.n1000 VN.t2111 3.643
R4356 VN.n1278 VN.t2016 3.643
R4357 VN.n1283 VN.n1282 3.643
R4358 VN.n1286 VN.n1285 3.643
R4359 VN.n1275 VN.t629 3.643
R4360 VN.n1690 VN.t390 3.643
R4361 VN.n1694 VN.n1693 3.643
R4362 VN.n1697 VN.n1696 3.643
R4363 VN.n1687 VN.t1517 3.643
R4364 VN.n1968 VN.t921 3.643
R4365 VN.n1973 VN.n1972 3.643
R4366 VN.n1976 VN.n1975 3.643
R4367 VN.n1965 VN.t2082 3.643
R4368 VN.n2398 VN.t1816 3.643
R4369 VN.n2402 VN.n2401 3.643
R4370 VN.n2405 VN.n2404 3.643
R4371 VN.n2395 VN.t460 3.643
R4372 VN.n2677 VN.t361 3.643
R4373 VN.n2682 VN.n2681 3.643
R4374 VN.n2685 VN.n2684 3.643
R4375 VN.n2674 VN.t1494 3.643
R4376 VN.n3117 VN.t1533 3.643
R4377 VN.n3121 VN.n3120 3.643
R4378 VN.n3124 VN.n3123 3.643
R4379 VN.n3114 VN.t2383 3.643
R4380 VN.n3399 VN.t2300 3.643
R4381 VN.n3404 VN.n3403 3.643
R4382 VN.n3407 VN.n3406 3.643
R4383 VN.n3396 VN.t894 3.643
R4384 VN.n3860 VN.t1063 3.643
R4385 VN.n3864 VN.n3863 3.643
R4386 VN.n3867 VN.n3866 3.643
R4387 VN.n3857 VN.t2096 3.643
R4388 VN.n4143 VN.t1699 3.643
R4389 VN.n4148 VN.n4147 3.643
R4390 VN.n4151 VN.n4150 3.643
R4391 VN.n4140 VN.t331 3.643
R4392 VN.n4614 VN.t501 3.643
R4393 VN.n4618 VN.n4617 3.643
R4394 VN.n4621 VN.n4620 3.643
R4395 VN.n4611 VN.t1626 3.643
R4396 VN.n4900 VN.t1125 3.643
R4397 VN.n4905 VN.n4904 3.643
R4398 VN.n4908 VN.n4907 3.643
R4399 VN.n4897 VN.t2270 3.643
R4400 VN.n5392 VN.t72 3.643
R4401 VN.n5396 VN.n5395 3.643
R4402 VN.n5399 VN.n5398 3.643
R4403 VN.n5389 VN.t1274 3.643
R4404 VN.n5679 VN.t2351 3.643
R4405 VN.n5684 VN.n5683 3.643
R4406 VN.n5687 VN.n5686 3.643
R4407 VN.n5676 VN.t963 3.643
R4408 VN.n6181 VN.t18 3.643
R4409 VN.n6185 VN.n6184 3.643
R4410 VN.n6188 VN.n6187 3.643
R4411 VN.n6178 VN.t1241 3.643
R4412 VN.n6471 VN.t1472 3.643
R4413 VN.n6476 VN.n6475 3.643
R4414 VN.n6479 VN.n6478 3.643
R4415 VN.n6468 VN.t931 3.643
R4416 VN.n6625 VN.t2578 3.643
R4417 VN.n6947 VN.n6946 3.643
R4418 VN.n6944 VN.n6943 3.643
R4419 VN.n6622 VN.t1215 3.643
R4420 VN.n6939 VN.t1449 3.643
R4421 VN.n6936 VN.n6935 3.643
R4422 VN.n6933 VN.n6932 3.643
R4423 VN.n6630 VN.t2581 3.643
R4424 VN.n7372 VN.t321 3.643
R4425 VN.n6913 VN.t699 3.643
R4426 VN.n6927 VN.n6926 3.643
R4427 VN.n6930 VN.n6929 3.643
R4428 VN.n6916 VN.t1712 3.643
R4429 VN.n6610 VN.t1708 3.643
R4430 VN.n6617 VN.n6616 3.643
R4431 VN.n6614 VN.n6613 3.643
R4432 VN.n6607 VN.t353 3.643
R4433 VN.n127 VN.t1834 3.643
R4434 VN.n12467 VN.t239 3.643
R4435 VN.n12472 VN.n12471 3.643
R4436 VN.n12475 VN.n12474 3.643
R4437 VN.n12464 VN.t1092 3.643
R4438 VN.n12821 VN.t1271 3.643
R4439 VN.n12841 VN.n12840 3.643
R4440 VN.n12818 VN.n12817 3.643
R4441 VN.n12815 VN.t2401 3.643
R4442 VN.n12835 VN.t2314 3.643
R4443 VN.n12832 VN.n12831 3.643
R4444 VN.n12829 VN.n12828 3.643
R4445 VN.n12826 VN.t794 3.643
R4446 VN.n346 VN.t675 3.643
R4447 VN.n350 VN.n349 3.643
R4448 VN.n353 VN.n352 3.643
R4449 VN.n343 VN.t1804 3.643
R4450 VN.n619 VN.t1717 3.643
R4451 VN.n624 VN.n623 3.643
R4452 VN.n627 VN.n626 3.643
R4453 VN.n616 VN.t349 3.643
R4454 VN.n1018 VN.t25 3.643
R4455 VN.n1022 VN.n1021 3.643
R4456 VN.n1025 VN.n1024 3.643
R4457 VN.n1015 VN.t1234 3.643
R4458 VN.n1294 VN.t1143 3.643
R4459 VN.n1299 VN.n1298 3.643
R4460 VN.n1302 VN.n1301 3.643
R4461 VN.n1291 VN.t2286 3.643
R4462 VN.n1705 VN.t2043 3.643
R4463 VN.n1709 VN.n1708 3.643
R4464 VN.n1712 VN.n1711 3.643
R4465 VN.n1702 VN.t649 3.643
R4466 VN.n1984 VN.t2582 3.643
R4467 VN.n1989 VN.n1988 3.643
R4468 VN.n1992 VN.n1991 3.643
R4469 VN.n1981 VN.t1208 3.643
R4470 VN.n2413 VN.t941 3.643
R4471 VN.n2417 VN.n2416 3.643
R4472 VN.n2420 VN.n2419 3.643
R4473 VN.n2410 VN.t2108 3.643
R4474 VN.n2693 VN.t2011 3.643
R4475 VN.n2698 VN.n2697 3.643
R4476 VN.n2701 VN.n2700 3.643
R4477 VN.n2690 VN.t627 3.643
R4478 VN.n3132 VN.t783 3.643
R4479 VN.n3136 VN.n3135 3.643
R4480 VN.n3139 VN.n3138 3.643
R4481 VN.n3129 VN.t1514 3.643
R4482 VN.n3415 VN.t1427 3.643
R4483 VN.n3420 VN.n3419 3.643
R4484 VN.n3423 VN.n3422 3.643
R4485 VN.n3412 VN.t2557 3.643
R4486 VN.n3875 VN.t189 3.643
R4487 VN.n3879 VN.n3878 3.643
R4488 VN.n3882 VN.n3881 3.643
R4489 VN.n3872 VN.t1356 3.643
R4490 VN.n4159 VN.t829 3.643
R4491 VN.n4164 VN.n4163 3.643
R4492 VN.n4167 VN.n4166 3.643
R4493 VN.n4156 VN.t1977 3.643
R4494 VN.n4629 VN.t1787 3.643
R4495 VN.n4633 VN.n4632 3.643
R4496 VN.n4636 VN.n4635 3.643
R4497 VN.n4626 VN.t438 3.643
R4498 VN.n4916 VN.t1507 3.643
R4499 VN.n4921 VN.n4920 3.643
R4500 VN.n4924 VN.n4923 3.643
R4501 VN.n4913 VN.t104 3.643
R4502 VN.n5407 VN.t1759 3.643
R4503 VN.n5411 VN.n5410 3.643
R4504 VN.n5414 VN.n5413 3.643
R4505 VN.n5404 VN.t404 3.643
R4506 VN.n5695 VN.t1482 3.643
R4507 VN.n5700 VN.n5699 3.643
R4508 VN.n5703 VN.n5702 3.643
R4509 VN.n5692 VN.t56 3.643
R4510 VN.n6196 VN.t1732 3.643
R4511 VN.n6515 VN.n6514 3.643
R4512 VN.n6518 VN.n6517 3.643
R4513 VN.n6193 VN.t376 3.643
R4514 VN.n6510 VN.t605 3.643
R4515 VN.n6507 VN.n6506 3.643
R4516 VN.n6504 VN.n6503 3.643
R4517 VN.n6201 VN.t7 3.643
R4518 VN.n6579 VN.t1998 3.643
R4519 VN.n6484 VN.t2382 3.643
R4520 VN.n6498 VN.n6497 3.643
R4521 VN.n6501 VN.n6500 3.643
R4522 VN.n6487 VN.t1724 3.643
R4523 VN.n6526 VN.t857 3.643
R4524 VN.n6530 VN.n6529 3.643
R4525 VN.n6533 VN.n6532 3.643
R4526 VN.n6523 VN.t2030 3.643
R4527 VN.n131 VN.t960 3.643
R4528 VN.n12483 VN.t2028 3.643
R4529 VN.n12488 VN.n12487 3.643
R4530 VN.n12491 VN.n12490 3.643
R4531 VN.n12480 VN.t222 3.643
R4532 VN.n12849 VN.t402 3.643
R4533 VN.n12869 VN.n12868 3.643
R4534 VN.n12872 VN.n12871 3.643
R4535 VN.n12846 VN.t1532 3.643
R4536 VN.n12863 VN.t1444 3.643
R4537 VN.n12860 VN.n12859 3.643
R4538 VN.n12857 VN.n12856 3.643
R4539 VN.n12854 VN.t2568 3.643
R4540 VN.n361 VN.t2334 3.643
R4541 VN.n365 VN.n364 3.643
R4542 VN.n368 VN.n367 3.643
R4543 VN.n358 VN.t929 3.643
R4544 VN.n635 VN.t844 3.643
R4545 VN.n640 VN.n639 3.643
R4546 VN.n643 VN.n642 3.643
R4547 VN.n632 VN.t1993 3.643
R4548 VN.n1033 VN.t1736 3.643
R4549 VN.n1037 VN.n1036 3.643
R4550 VN.n1040 VN.n1039 3.643
R4551 VN.n1030 VN.t370 3.643
R4552 VN.n1310 VN.t279 3.643
R4553 VN.n1315 VN.n1314 3.643
R4554 VN.n1318 VN.n1317 3.643
R4555 VN.n1307 VN.t1417 3.643
R4556 VN.n1720 VN.t1171 3.643
R4557 VN.n1724 VN.n1723 3.643
R4558 VN.n1727 VN.n1726 3.643
R4559 VN.n1717 VN.t2308 3.643
R4560 VN.n2000 VN.t1713 3.643
R4561 VN.n2005 VN.n2004 3.643
R4562 VN.n2008 VN.n2007 3.643
R4563 VN.n1997 VN.t345 3.643
R4564 VN.n2428 VN.t208 3.643
R4565 VN.n2432 VN.n2431 3.643
R4566 VN.n2435 VN.n2434 3.643
R4567 VN.n2425 VN.t1231 3.643
R4568 VN.n2709 VN.t1138 3.643
R4569 VN.n2714 VN.n2713 3.643
R4570 VN.n2717 VN.n2716 3.643
R4571 VN.n2706 VN.t2281 3.643
R4572 VN.n3147 VN.t2435 3.643
R4573 VN.n3151 VN.n3150 3.643
R4574 VN.n3154 VN.n3153 3.643
R4575 VN.n3144 VN.t770 3.643
R4576 VN.n3431 VN.t562 3.643
R4577 VN.n3436 VN.n3435 3.643
R4578 VN.n3439 VN.n3438 3.643
R4579 VN.n3428 VN.t1687 3.643
R4580 VN.n3890 VN.t938 3.643
R4581 VN.n3894 VN.n3893 3.643
R4582 VN.n3897 VN.n3896 3.643
R4583 VN.n3887 VN.t2113 3.643
R4584 VN.n4175 VN.t666 3.643
R4585 VN.n4180 VN.n4179 3.643
R4586 VN.n4183 VN.n4182 3.643
R4587 VN.n4172 VN.t1803 3.643
R4588 VN.n4644 VN.t912 3.643
R4589 VN.n4648 VN.n4647 3.643
R4590 VN.n4651 VN.n4650 3.643
R4591 VN.n4641 VN.t2083 3.643
R4592 VN.n4932 VN.t640 3.643
R4593 VN.n4937 VN.n4936 3.643
R4594 VN.n4940 VN.n4939 3.643
R4595 VN.n4929 VN.t1775 3.643
R4596 VN.n5422 VN.t886 3.643
R4597 VN.n5739 VN.n5738 3.643
R4598 VN.n5742 VN.n5741 3.643
R4599 VN.n5419 VN.t2054 3.643
R4600 VN.n5734 VN.t616 3.643
R4601 VN.n5731 VN.n5730 3.643
R4602 VN.n5728 VN.n5727 3.643
R4603 VN.n5427 VN.t1748 3.643
R4604 VN.n5803 VN.t1156 3.643
R4605 VN.n5708 VN.t2394 3.643
R4606 VN.n5722 VN.n5721 3.643
R4607 VN.n5725 VN.n5724 3.643
R4608 VN.n5711 VN.t875 3.643
R4609 VN.n5750 VN.t2547 3.643
R4610 VN.n5754 VN.n5753 3.643
R4611 VN.n5757 VN.n5756 3.643
R4612 VN.n5747 VN.t1185 3.643
R4613 VN.n135 VN.t52 3.643
R4614 VN.n12499 VN.t1153 3.643
R4615 VN.n12504 VN.n12503 3.643
R4616 VN.n12507 VN.n12506 3.643
R4617 VN.n12496 VN.t2010 3.643
R4618 VN.n12880 VN.t2050 3.643
R4619 VN.n12900 VN.n12899 3.643
R4620 VN.n12903 VN.n12902 3.643
R4621 VN.n12877 VN.t661 3.643
R4622 VN.n12894 VN.t575 3.643
R4623 VN.n12891 VN.n12890 3.643
R4624 VN.n12888 VN.n12887 3.643
R4625 VN.n12885 VN.t1697 3.643
R4626 VN.n376 VN.t1469 3.643
R4627 VN.n380 VN.n379 3.643
R4628 VN.n383 VN.n382 3.643
R4629 VN.n373 VN.t3 3.643
R4630 VN.n651 VN.t2508 3.643
R4631 VN.n656 VN.n655 3.643
R4632 VN.n659 VN.n658 3.643
R4633 VN.n648 VN.t1120 3.643
R4634 VN.n1048 VN.t863 3.643
R4635 VN.n1052 VN.n1051 3.643
R4636 VN.n1055 VN.n1054 3.643
R4637 VN.n1045 VN.t2022 3.643
R4638 VN.n1326 VN.t1930 3.643
R4639 VN.n1331 VN.n1330 3.643
R4640 VN.n1334 VN.n1333 3.643
R4641 VN.n1323 VN.t554 3.643
R4642 VN.n1735 VN.t443 3.643
R4643 VN.n1739 VN.n1738 3.643
R4644 VN.n1742 VN.n1741 3.643
R4645 VN.n1732 VN.t1438 3.643
R4646 VN.n2016 VN.t841 3.643
R4647 VN.n2021 VN.n2020 3.643
R4648 VN.n2024 VN.n2023 3.643
R4649 VN.n2013 VN.t1988 3.643
R4650 VN.n2443 VN.t1858 3.643
R4651 VN.n2447 VN.n2446 3.643
R4652 VN.n2450 VN.n2449 3.643
R4653 VN.n2440 VN.t498 3.643
R4654 VN.n2725 VN.t275 3.643
R4655 VN.n2730 VN.n2729 3.643
R4656 VN.n2733 VN.n2732 3.643
R4657 VN.n2722 VN.t1412 3.643
R4658 VN.n3162 VN.t64 3.643
R4659 VN.n3166 VN.n3165 3.643
R4660 VN.n3169 VN.n3168 3.643
R4661 VN.n3159 VN.t2130 3.643
R4662 VN.n3447 VN.t2347 3.643
R4663 VN.n3452 VN.n3451 3.643
R4664 VN.n3455 VN.n3454 3.643
R4665 VN.n3444 VN.t952 3.643
R4666 VN.n3905 VN.t15 3.643
R4667 VN.n3909 VN.n3908 3.643
R4668 VN.n3912 VN.n3911 3.643
R4669 VN.n3902 VN.t1235 3.643
R4670 VN.n4191 VN.t2324 3.643
R4671 VN.n4196 VN.n4195 3.643
R4672 VN.n4199 VN.n4198 3.643
R4673 VN.n4188 VN.t927 3.643
R4674 VN.n4659 VN.t2574 3.643
R4675 VN.n4976 VN.n4975 3.643
R4676 VN.n4979 VN.n4978 3.643
R4677 VN.n4656 VN.t1209 3.643
R4678 VN.n4971 VN.t2299 3.643
R4679 VN.n4968 VN.n4967 3.643
R4680 VN.n4965 VN.n4964 3.643
R4681 VN.n4664 VN.t901 3.643
R4682 VN.n5040 VN.t314 3.643
R4683 VN.n4945 VN.t1550 3.643
R4684 VN.n4959 VN.n4958 3.643
R4685 VN.n4962 VN.n4961 3.643
R4686 VN.n4948 VN.t2563 3.643
R4687 VN.n4987 VN.t1702 3.643
R4688 VN.n4991 VN.n4990 3.643
R4689 VN.n4994 VN.n4993 3.643
R4690 VN.n4984 VN.t346 3.643
R4691 VN.n139 VN.t1747 3.643
R4692 VN.n12515 VN.t286 3.643
R4693 VN.n12520 VN.n12519 3.643
R4694 VN.n12523 VN.n12522 3.643
R4695 VN.n12512 VN.t1137 3.643
R4696 VN.n12911 VN.t1181 3.643
R4697 VN.n12931 VN.n12930 3.643
R4698 VN.n12934 VN.n12933 3.643
R4699 VN.n12908 VN.t2321 3.643
R4700 VN.n12925 VN.t2233 3.643
R4701 VN.n12922 VN.n12921 3.643
R4702 VN.n12919 VN.n12918 3.643
R4703 VN.n12916 VN.t827 3.643
R4704 VN.n391 VN.t600 3.643
R4705 VN.n395 VN.n394 3.643
R4706 VN.n398 VN.n397 3.643
R4707 VN.n388 VN.t1723 3.643
R4708 VN.n667 VN.t1646 3.643
R4709 VN.n672 VN.n671 3.643
R4710 VN.n675 VN.n674 3.643
R4711 VN.n664 VN.t258 3.643
R4712 VN.n1063 VN.t113 3.643
R4713 VN.n1067 VN.n1066 3.643
R4714 VN.n1070 VN.n1069 3.643
R4715 VN.n1060 VN.t1148 3.643
R4716 VN.n1342 VN.t1055 3.643
R4717 VN.n1347 VN.n1346 3.643
R4718 VN.n1350 VN.n1349 3.643
R4719 VN.n1339 VN.t2212 3.643
R4720 VN.n1750 VN.t2088 3.643
R4721 VN.n1754 VN.n1753 3.643
R4722 VN.n1757 VN.n1756 3.643
R4723 VN.n1747 VN.t693 3.643
R4724 VN.n2032 VN.t2504 3.643
R4725 VN.n2037 VN.n2036 3.643
R4726 VN.n2040 VN.n2039 3.643
R4727 VN.n2029 VN.t1115 3.643
R4728 VN.n2458 VN.t86 3.643
R4729 VN.n2462 VN.n2461 3.643
R4730 VN.n2465 VN.n2464 3.643
R4731 VN.n2455 VN.t1285 3.643
R4732 VN.n2741 VN.t1505 3.643
R4733 VN.n2746 VN.n2745 3.643
R4734 VN.n2749 VN.n2748 3.643
R4735 VN.n2738 VN.t98 3.643
R4736 VN.n3177 VN.t1755 3.643
R4737 VN.n3181 VN.n3180 3.643
R4738 VN.n3184 VN.n3183 3.643
R4739 VN.n3174 VN.t1254 3.643
R4740 VN.n3463 VN.t1477 3.643
R4741 VN.n3468 VN.n3467 3.643
R4742 VN.n3471 VN.n3470 3.643
R4743 VN.n3460 VN.t34 3.643
R4744 VN.n3920 VN.t1731 3.643
R4745 VN.n4235 VN.n4234 3.643
R4746 VN.n4238 VN.n4237 3.643
R4747 VN.n3917 VN.t371 3.643
R4748 VN.n4230 VN.t1458 3.643
R4749 VN.n4227 VN.n4226 3.643
R4750 VN.n4224 VN.n4223 3.643
R4751 VN.n3925 VN.t2589 3.643
R4752 VN.n4299 VN.t1989 3.643
R4753 VN.n4204 VN.t709 3.643
R4754 VN.n4218 VN.n4217 3.643
R4755 VN.n4221 VN.n4220 3.643
R4756 VN.n4207 VN.t1721 3.643
R4757 VN.n4246 VN.t855 3.643
R4758 VN.n4250 VN.n4249 3.643
R4759 VN.n4253 VN.n4252 3.643
R4760 VN.n4243 VN.t2023 3.643
R4761 VN.n143 VN.t874 3.643
R4762 VN.n12531 VN.t1938 3.643
R4763 VN.n12536 VN.n12535 3.643
R4764 VN.n12539 VN.n12538 3.643
R4765 VN.n12528 VN.t274 3.643
R4766 VN.n12942 VN.t311 3.643
R4767 VN.n12962 VN.n12961 3.643
R4768 VN.n12965 VN.n12964 3.643
R4769 VN.n12939 VN.t1453 3.643
R4770 VN.n12956 VN.t1369 3.643
R4771 VN.n12953 VN.n12952 3.643
R4772 VN.n12950 VN.n12949 3.643
R4773 VN.n12947 VN.t2492 3.643
R4774 VN.n406 VN.t2375 3.643
R4775 VN.n410 VN.n409 3.643
R4776 VN.n413 VN.n412 3.643
R4777 VN.n403 VN.t850 3.643
R4778 VN.n683 VN.t775 3.643
R4779 VN.n688 VN.n687 3.643
R4780 VN.n691 VN.n690 3.643
R4781 VN.n680 VN.t1906 3.643
R4782 VN.n1078 VN.t1781 3.643
R4783 VN.n1082 VN.n1081 3.643
R4784 VN.n1085 VN.n1084 3.643
R4785 VN.n1075 VN.t422 3.643
R4786 VN.n1358 VN.t182 3.643
R4787 VN.n1363 VN.n1362 3.643
R4788 VN.n1366 VN.n1365 3.643
R4789 VN.n1355 VN.t1345 3.643
R4790 VN.n1765 VN.t1341 3.643
R4791 VN.n1769 VN.n1768 3.643
R4792 VN.n1772 VN.n1771 3.643
R4793 VN.n1762 VN.t2469 3.643
R4794 VN.n2048 VN.t659 3.643
R4795 VN.n2053 VN.n2052 3.643
R4796 VN.n2056 VN.n2055 3.643
R4797 VN.n2045 VN.t1800 3.643
R4798 VN.n2473 VN.t1766 3.643
R4799 VN.n2477 VN.n2476 3.643
R4800 VN.n2480 VN.n2479 3.643
R4801 VN.n2470 VN.t417 3.643
R4802 VN.n2757 VN.t637 3.643
R4803 VN.n2762 VN.n2761 3.643
R4804 VN.n2765 VN.n2764 3.643
R4805 VN.n2754 VN.t1769 3.643
R4806 VN.n3192 VN.t883 3.643
R4807 VN.n3507 VN.n3506 3.643
R4808 VN.n3510 VN.n3509 3.643
R4809 VN.n3189 VN.t384 3.643
R4810 VN.n3502 VN.t609 3.643
R4811 VN.n3499 VN.n3498 3.643
R4812 VN.n3496 VN.n3495 3.643
R4813 VN.n3197 VN.t1740 3.643
R4814 VN.n3571 VN.t1149 3.643
R4815 VN.n3476 VN.t2388 3.643
R4816 VN.n3490 VN.n3489 3.643
R4817 VN.n3493 VN.n3492 3.643
R4818 VN.n3479 VN.t868 3.643
R4819 VN.n3518 VN.t2544 3.643
R4820 VN.n3522 VN.n3521 3.643
R4821 VN.n3525 VN.n3524 3.643
R4822 VN.n3515 VN.t2038 3.643
R4823 VN.n147 VN.t2535 3.643
R4824 VN.n12547 VN.t1065 3.643
R4825 VN.n12552 VN.n12551 3.643
R4826 VN.n12555 VN.n12554 3.643
R4827 VN.n12544 VN.t1924 3.643
R4828 VN.n12973 VN.t2100 3.643
R4829 VN.n12993 VN.n12992 3.643
R4830 VN.n12996 VN.n12995 3.643
R4831 VN.n12970 VN.t584 3.643
R4832 VN.n12987 VN.t502 3.643
R4833 VN.n12984 VN.n12983 3.643
R4834 VN.n12981 VN.n12980 3.643
R4835 VN.n12978 VN.t1627 3.643
R4836 VN.n421 VN.t1508 3.643
R4837 VN.n425 VN.n424 3.643
R4838 VN.n428 VN.n427 3.643
R4839 VN.n418 VN.t84 3.643
R4840 VN.n699 VN.t2425 3.643
R4841 VN.n704 VN.n703 3.643
R4842 VN.n707 VN.n706 3.643
R4843 VN.n696 VN.t1032 3.643
R4844 VN.n1093 VN.t496 3.643
R4845 VN.n1097 VN.n1096 3.643
R4846 VN.n1100 VN.n1099 3.643
R4847 VN.n1090 VN.t1630 3.643
R4848 VN.n1374 VN.t1853 3.643
R4849 VN.n1379 VN.n1378 3.643
R4850 VN.n1382 VN.n1381 3.643
R4851 VN.n1371 VN.t499 3.643
R4852 VN.n1780 VN.t476 3.643
R4853 VN.n1784 VN.n1783 3.643
R4854 VN.n1787 VN.n1786 3.643
R4855 VN.n1777 VN.t1605 3.643
R4856 VN.n2064 VN.t2319 3.643
R4857 VN.n2069 VN.n2068 3.643
R4858 VN.n2072 VN.n2071 3.643
R4859 VN.n2061 VN.t923 3.643
R4860 VN.n2488 VN.t895 3.643
R4861 VN.n2801 VN.n2800 3.643
R4862 VN.n2804 VN.n2803 3.643
R4863 VN.n2485 VN.t2065 3.643
R4864 VN.n2796 VN.t2294 3.643
R4865 VN.n2793 VN.n2792 3.643
R4866 VN.n2790 VN.n2789 3.643
R4867 VN.n2493 VN.t897 3.643
R4868 VN.n2865 VN.t1165 3.643
R4869 VN.n2770 VN.t1547 3.643
R4870 VN.n2784 VN.n2783 3.643
R4871 VN.n2787 VN.n2786 3.643
R4872 VN.n2773 VN.t2559 3.643
R4873 VN.n2812 VN.t2556 3.643
R4874 VN.n2816 VN.n2815 3.643
R4875 VN.n2819 VN.n2818 3.643
R4876 VN.n2809 VN.t1193 3.643
R4877 VN.n151 VN.t1792 3.643
R4878 VN.n12563 VN.t190 3.643
R4879 VN.n12568 VN.n12567 3.643
R4880 VN.n12571 VN.n12570 3.643
R4881 VN.n12560 VN.t1049 3.643
R4882 VN.n13004 VN.t1223 3.643
R4883 VN.n13024 VN.n13023 3.643
R4884 VN.n13027 VN.n13026 3.643
R4885 VN.n13001 VN.t2363 3.643
R4886 VN.n13018 VN.t2157 3.643
R4887 VN.n13015 VN.n13014 3.643
R4888 VN.n13012 VN.n13011 3.643
R4889 VN.n13009 VN.t755 3.643
R4890 VN.n436 VN.t2178 3.643
R4891 VN.n440 VN.n439 3.643
R4892 VN.n443 VN.n442 3.643
R4893 VN.n433 VN.t788 3.643
R4894 VN.n715 VN.t1010 3.643
R4895 VN.n720 VN.n719 3.643
R4896 VN.n723 VN.n722 3.643
R4897 VN.n712 VN.t2180 3.643
R4898 VN.n1108 VN.t2153 3.643
R4899 VN.n1112 VN.n1111 3.643
R4900 VN.n1115 VN.n1114 3.643
R4901 VN.n1105 VN.t757 3.643
R4902 VN.n1390 VN.t984 3.643
R4903 VN.n1395 VN.n1394 3.643
R4904 VN.n1398 VN.n1397 3.643
R4905 VN.n1387 VN.t2154 3.643
R4906 VN.n1795 VN.t2129 3.643
R4907 VN.n2108 VN.n2107 3.643
R4908 VN.n2111 VN.n2110 3.643
R4909 VN.n1792 VN.t740 3.643
R4910 VN.n2103 VN.t1451 3.643
R4911 VN.n2100 VN.n2099 3.643
R4912 VN.n2097 VN.n2096 3.643
R4913 VN.n1800 VN.t2585 3.643
R4914 VN.n2172 VN.t324 3.643
R4915 VN.n2077 VN.t704 3.643
R4916 VN.n2091 VN.n2090 3.643
R4917 VN.n2094 VN.n2093 3.643
R4918 VN.n2080 VN.t1715 3.643
R4919 VN.n2119 VN.t1253 3.643
R4920 VN.n2123 VN.n2122 3.643
R4921 VN.n2126 VN.n2125 3.643
R4922 VN.n2116 VN.t2397 3.643
R4923 VN.n155 VN.t917 3.643
R4924 VN.n12579 VN.t1848 3.643
R4925 VN.n12584 VN.n12583 3.643
R4926 VN.n12587 VN.n12586 3.643
R4927 VN.n12576 VN.t179 3.643
R4928 VN.n13035 VN.t1333 3.643
R4929 VN.n13055 VN.n13054 3.643
R4930 VN.n13058 VN.n13057 3.643
R4931 VN.n13032 VN.t2467 3.643
R4932 VN.n13049 VN.t162 3.643
R4933 VN.n13046 VN.n13045 3.643
R4934 VN.n13043 VN.n13042 3.643
R4935 VN.n13040 VN.t1338 3.643
R4936 VN.n451 VN.t1310 3.643
R4937 VN.n455 VN.n454 3.643
R4938 VN.n458 VN.n457 3.643
R4939 VN.n448 VN.t2440 3.643
R4940 VN.n731 VN.t136 3.643
R4941 VN.n736 VN.n735 3.643
R4942 VN.n739 VN.n738 3.643
R4943 VN.n728 VN.t1312 3.643
R4944 VN.n1123 VN.t1284 3.643
R4945 VN.n1434 VN.n1433 3.643
R4946 VN.n1437 VN.n1436 3.643
R4947 VN.n1120 VN.t2415 3.643
R4948 VN.n1429 VN.t95 3.643
R4949 VN.n1426 VN.n1425 3.643
R4950 VN.n1423 VN.n1422 3.643
R4951 VN.n1128 VN.t1286 3.643
R4952 VN.n1498 VN.t1528 3.643
R4953 VN.n1403 VN.t1895 3.643
R4954 VN.n1417 VN.n1416 3.643
R4955 VN.n1420 VN.n1419 3.643
R4956 VN.n1406 VN.t419 3.643
R4957 VN.n1445 VN.t416 3.643
R4958 VN.n1449 VN.n1448 3.643
R4959 VN.n1452 VN.n1451 3.643
R4960 VN.n1442 VN.t1553 3.643
R4961 VN.n159 VN.t492 3.643
R4962 VN.n12595 VN.t1847 3.643
R4963 VN.n12600 VN.n12599 3.643
R4964 VN.n12603 VN.n12602 3.643
R4965 VN.n12592 VN.t1353 3.643
R4966 VN.n13066 VN.t471 3.643
R4967 VN.n13086 VN.n13085 3.643
R4968 VN.n13089 VN.n13088 3.643
R4969 VN.n13063 VN.t1599 3.643
R4970 VN.n13080 VN.t1824 3.643
R4971 VN.n13077 VN.n13076 3.643
R4972 VN.n13074 VN.n13073 3.643
R4973 VN.n13071 VN.t474 3.643
R4974 VN.n466 VN.t449 3.643
R4975 VN.n774 VN.n773 3.643
R4976 VN.n777 VN.n776 3.643
R4977 VN.n463 VN.t1578 3.643
R4978 VN.n769 VN.t1799 3.643
R4979 VN.n766 VN.n765 3.643
R4980 VN.n763 VN.n762 3.643
R4981 VN.n471 VN.t451 3.643
R4982 VN.n848 VN.t679 3.643
R4983 VN.n742 VN.t1057 3.643
R4984 VN.n757 VN.n756 3.643
R4985 VN.n760 VN.n759 3.643
R4986 VN.n745 VN.t2097 3.643
R4987 VN.n787 VN.t2095 3.643
R4988 VN.n796 VN.n795 3.643
R4989 VN.n799 VN.n798 3.643
R4990 VN.n790 VN.t711 3.643
R4991 VN.n163 VN.t2147 3.643
R4992 VN.n12608 VN.t975 3.643
R4993 VN.n12616 VN.n12615 3.643
R4994 VN.n12619 VN.n12618 3.643
R4995 VN.n12611 VN.t485 3.643
R4996 VN.n13098 VN.t2121 3.643
R4997 VN.n13106 VN.n13105 3.643
R4998 VN.n13109 VN.n13108 3.643
R4999 VN.n13101 VN.t735 3.643
R5000 VN.n12750 VN.t949 3.643
R5001 VN.n12758 VN.n12757 3.643
R5002 VN.n12761 VN.n12760 3.643
R5003 VN.n12753 VN.t2126 3.643
R5004 VN.n198 VN.t2366 3.643
R5005 VN.n167 VN.t1277 3.643
R5006 VN.n12379 VN.t83 3.643
R5007 VN.n12390 VN.n12389 3.643
R5008 VN.n12387 VN.n12386 3.643
R5009 VN.n12382 VN.t2138 3.643
R5010 VN.n12227 VN.t1246 3.643
R5011 VN.n12235 VN.n12234 3.643
R5012 VN.n12218 VN.n12217 3.643
R5013 VN.n12230 VN.t2390 3.643
R5014 VN.n12724 VN.t218 3.643
R5015 VN.n12742 VN.n12741 3.643
R5016 VN.n12739 VN.n12738 3.643
R5017 VN.n12727 VN.t1250 3.643
R5018 VN.n12400 VN.t1265 3.643
R5019 VN.n12403 VN.n12402 3.643
R5020 VN.n6584 VN.n6583 3.643
R5021 VN.n6582 VN.t2590 3.643
R5022 VN.n12360 VN.n12358 2.799
R5023 VN.n11534 VN.n11532 2.511
R5024 VN.n10714 VN.n10713 2.511
R5025 VN.n9854 VN.n9853 2.511
R5026 VN.n9006 VN.n9005 2.511
R5027 VN.n8173 VN.n8172 2.511
R5028 VN.n7362 VN.n7361 2.511
R5029 VN.n6569 VN.n6568 2.511
R5030 VN.n5793 VN.n5792 2.511
R5031 VN.n5030 VN.n5029 2.511
R5032 VN.n4289 VN.n4288 2.511
R5033 VN.n3561 VN.n3560 2.511
R5034 VN.n2855 VN.n2854 2.511
R5035 VN.n2162 VN.n2161 2.511
R5036 VN.n1488 VN.n1487 2.511
R5037 VN.n838 VN.n837 2.511
R5038 VN.n811 VN.n810 2.511
R5039 VN.n13127 VN.n13126 2.511
R5040 VN.n824 VN.n823 0.21
R5041 VN.n179 VN.n176 0.178
R5042 VN.n11530 VN.n11529 0.172
R5043 VN.n11782 VN.n11779 0.164
R5044 VN VN.n182 0.138
R5045 VN.n252 VN.n251 0.133
R5046 VN.n863 VN.n862 0.133
R5047 VN.n1549 VN.n1548 0.133
R5048 VN.n2254 VN.n2253 0.133
R5049 VN.n2976 VN.n2975 0.133
R5050 VN.n3716 VN.n3715 0.133
R5051 VN.n4473 VN.n4472 0.133
R5052 VN.n5248 VN.n5247 0.133
R5053 VN.n6040 VN.n6039 0.133
R5054 VN.n7283 VN.n7282 0.133
R5055 VN.n7672 VN.n7671 0.133
R5056 VN.n8517 VN.n8516 0.133
R5057 VN.n9379 VN.n9378 0.133
R5058 VN.n10262 VN.n10261 0.133
R5059 VN.n11505 VN.n11504 0.133
R5060 VN.n10711 VN.n10710 0.119
R5061 VN.n9851 VN.n9850 0.119
R5062 VN.n9003 VN.n9002 0.119
R5063 VN.n8170 VN.n8169 0.119
R5064 VN.n7359 VN.n7358 0.119
R5065 VN.n6566 VN.n6565 0.119
R5066 VN.n5790 VN.n5789 0.119
R5067 VN.n5027 VN.n5026 0.119
R5068 VN.n4286 VN.n4285 0.119
R5069 VN.n3558 VN.n3557 0.119
R5070 VN.n2852 VN.n2851 0.119
R5071 VN.n2159 VN.n2158 0.119
R5072 VN.n1485 VN.n1484 0.119
R5073 VN.n835 VN.n834 0.119
R5074 VN.n808 VN.n807 0.119
R5075 VN.n13124 VN.n13123 0.119
R5076 VN.n12201 VN.n11525 0.114
R5077 VN.n12200 VN.n12182 0.111
R5078 VN.n12202 VN.n10707 0.111
R5079 VN.n12203 VN.n9827 0.111
R5080 VN.n12204 VN.n8981 0.111
R5081 VN.n12205 VN.n8148 0.111
R5082 VN.n12206 VN.n7337 0.111
R5083 VN.n12207 VN.n6544 0.111
R5084 VN.n12208 VN.n5768 0.111
R5085 VN.n12209 VN.n5005 0.111
R5086 VN.n12210 VN.n4264 0.111
R5087 VN.n12211 VN.n3536 0.111
R5088 VN.n12212 VN.n2830 0.111
R5089 VN.n12213 VN.n2137 0.111
R5090 VN.n12214 VN.n1463 0.111
R5091 VN.n12215 VN.n821 0.111
R5092 VN.n83 VN.n82 0.11
R5093 VN.n13138 VN.n13137 0.11
R5094 VN.n9777 VN.n9772 0.106
R5095 VN.n8931 VN.n8926 0.106
R5096 VN.n8098 VN.n8093 0.106
R5097 VN.n6923 VN.n6918 0.106
R5098 VN.n6494 VN.n6489 0.106
R5099 VN.n5718 VN.n5713 0.106
R5100 VN.n4955 VN.n4950 0.106
R5101 VN.n4214 VN.n4209 0.106
R5102 VN.n3486 VN.n3481 0.106
R5103 VN.n2780 VN.n2775 0.106
R5104 VN.n2087 VN.n2082 0.106
R5105 VN.n1413 VN.n1408 0.106
R5106 VN.n12735 VN.n12730 0.106
R5107 VN.n10223 VN.n10222 0.097
R5108 VN.n9340 VN.n9339 0.097
R5109 VN.n8478 VN.n8477 0.097
R5110 VN.n7633 VN.n7632 0.097
R5111 VN.n7244 VN.n7243 0.097
R5112 VN.n6001 VN.n6000 0.097
R5113 VN.n5209 VN.n5208 0.097
R5114 VN.n4434 VN.n4433 0.097
R5115 VN.n3677 VN.n3676 0.097
R5116 VN.n2937 VN.n2936 0.097
R5117 VN.n2215 VN.n2214 0.097
R5118 VN.n1507 VN.n1506 0.097
R5119 VN.n913 VN.n912 0.097
R5120 VN.n11410 VN.n11409 0.097
R5121 VN.n11437 VN.n11436 0.097
R5122 VN.n194 VN.n193 0.095
R5123 VN.n76 VN.n75 0.093
R5124 VN.n12354 VN.n12353 0.093
R5125 VN.n12686 VN.n12685 0.093
R5126 VN.n23 VN.n22 0.092
R5127 VN.n89 VN.n88 0.092
R5128 VN.n11056 VN.n11055 0.087
R5129 VN.n74 VN.n73 0.085
R5130 VN.n11542 VN.n11541 0.082
R5131 VN.n10722 VN.n10721 0.082
R5132 VN.n9862 VN.n9861 0.082
R5133 VN.n9014 VN.n9013 0.082
R5134 VN.n8181 VN.n8180 0.082
R5135 VN.n7370 VN.n7369 0.082
R5136 VN.n6577 VN.n6576 0.082
R5137 VN.n5801 VN.n5800 0.082
R5138 VN.n5038 VN.n5037 0.082
R5139 VN.n4297 VN.n4296 0.082
R5140 VN.n3569 VN.n3568 0.082
R5141 VN.n2863 VN.n2862 0.082
R5142 VN.n2170 VN.n2169 0.082
R5143 VN.n1496 VN.n1495 0.082
R5144 VN.n846 VN.n845 0.082
R5145 VN.n819 VN.n818 0.082
R5146 VN.n13135 VN.n13134 0.082
R5147 VN.n908 VN.n907 0.08
R5148 VN.n1502 VN.n1501 0.08
R5149 VN.n2210 VN.n2209 0.08
R5150 VN.n2932 VN.n2931 0.08
R5151 VN.n3672 VN.n3671 0.08
R5152 VN.n4429 VN.n4428 0.08
R5153 VN.n5204 VN.n5203 0.08
R5154 VN.n5996 VN.n5995 0.08
R5155 VN.n7239 VN.n7238 0.08
R5156 VN.n7628 VN.n7627 0.08
R5157 VN.n8473 VN.n8472 0.08
R5158 VN.n9335 VN.n9334 0.08
R5159 VN.n10218 VN.n10217 0.08
R5160 VN.n11439 VN.n11438 0.08
R5161 VN.n11412 VN.n11411 0.08
R5162 VN.n11787 VN.n11786 0.08
R5163 VN.n11787 VN.n11784 0.08
R5164 VN.n181 VN.n180 0.079
R5165 VN.n10577 VN.n10576 0.077
R5166 VN.n9692 VN.n9691 0.077
R5167 VN.n8830 VN.n8829 0.077
R5168 VN.n7981 VN.n7980 0.077
R5169 VN.n6790 VN.n6789 0.077
R5170 VN.n6345 VN.n6344 0.077
R5171 VN.n5553 VN.n5552 0.077
R5172 VN.n4774 VN.n4773 0.077
R5173 VN.n4017 VN.n4016 0.077
R5174 VN.n3273 VN.n3272 0.077
R5175 VN.n2551 VN.n2550 0.077
R5176 VN.n1842 VN.n1841 0.077
R5177 VN.n1152 VN.n1151 0.077
R5178 VN.n11396 VN.n11395 0.077
R5179 VN.n11137 VN.n11136 0.077
R5180 VN.n488 VN.n487 0.076
R5181 VN.n9841 VN.n9840 0.075
R5182 VN.n8995 VN.n8994 0.075
R5183 VN.n8162 VN.n8161 0.075
R5184 VN.n7351 VN.n7350 0.075
R5185 VN.n6558 VN.n6557 0.075
R5186 VN.n5782 VN.n5781 0.075
R5187 VN.n5019 VN.n5018 0.075
R5188 VN.n4278 VN.n4277 0.075
R5189 VN.n3550 VN.n3549 0.075
R5190 VN.n2844 VN.n2843 0.075
R5191 VN.n2151 VN.n2150 0.075
R5192 VN.n1477 VN.n1476 0.075
R5193 VN.n12365 VN.n12364 0.074
R5194 VN.n1140 VN.n1139 0.074
R5195 VN.n12695 VN.n12694 0.074
R5196 VN.n1814 VN.n1813 0.074
R5197 VN.n2505 VN.n2504 0.074
R5198 VN.n3211 VN.n3210 0.074
R5199 VN.n3937 VN.n3936 0.074
R5200 VN.n4678 VN.n4677 0.074
R5201 VN.n5439 VN.n5438 0.074
R5202 VN.n6213 VN.n6212 0.074
R5203 VN.n6642 VN.n6641 0.074
R5204 VN.n7817 VN.n7816 0.074
R5205 VN.n8648 VN.n8647 0.074
R5206 VN.n9494 VN.n9493 0.074
R5207 VN.n10349 VN.n10348 0.074
R5208 VN.n11376 VN.n11375 0.074
R5209 VN.n72 VN.n71 0.073
R5210 VN.n69 VN.n68 0.073
R5211 VN.n66 VN.n65 0.073
R5212 VN.n63 VN.n62 0.073
R5213 VN.n60 VN.n59 0.073
R5214 VN.n57 VN.n56 0.073
R5215 VN.n54 VN.n53 0.073
R5216 VN.n51 VN.n50 0.073
R5217 VN.n48 VN.n47 0.073
R5218 VN.n45 VN.n44 0.073
R5219 VN.n42 VN.n41 0.073
R5220 VN.n39 VN.n38 0.073
R5221 VN.n36 VN.n35 0.073
R5222 VN.n34 VN.n33 0.073
R5223 VN.n2 VN.n1 0.071
R5224 VN.n5 VN.n4 0.071
R5225 VN.n9775 VN.n9774 0.07
R5226 VN.n8929 VN.n8928 0.07
R5227 VN.n8096 VN.n8095 0.07
R5228 VN.n6921 VN.n6920 0.07
R5229 VN.n6492 VN.n6491 0.07
R5230 VN.n5716 VN.n5715 0.07
R5231 VN.n4953 VN.n4952 0.07
R5232 VN.n4212 VN.n4211 0.07
R5233 VN.n3484 VN.n3483 0.07
R5234 VN.n2778 VN.n2777 0.07
R5235 VN.n2085 VN.n2084 0.07
R5236 VN.n1411 VN.n1410 0.07
R5237 VN.n12733 VN.n12732 0.07
R5238 VN.n12067 VN.n12066 0.069
R5239 VN.t51 VN.n77 0.068
R5240 VN.n11672 VN.n11670 0.067
R5241 VN.n11672 VN.n11671 0.067
R5242 VN.n11715 VN.n11713 0.067
R5243 VN.n11715 VN.n11714 0.067
R5244 VN.n11707 VN.n11705 0.067
R5245 VN.n11707 VN.n11706 0.067
R5246 VN.n11692 VN.n11691 0.067
R5247 VN.n11692 VN.n11690 0.067
R5248 VN.n11680 VN.n11678 0.067
R5249 VN.n11680 VN.n11679 0.067
R5250 VN.n11854 VN.n11840 0.067
R5251 VN.n11854 VN.n11839 0.067
R5252 VN.n11726 VN.n11724 0.067
R5253 VN.n11726 VN.n11725 0.067
R5254 VN.n11830 VN.n11829 0.067
R5255 VN.n11830 VN.n11828 0.067
R5256 VN.n11737 VN.n11735 0.067
R5257 VN.n11737 VN.n11736 0.067
R5258 VN.n11819 VN.n11818 0.067
R5259 VN.n11819 VN.n11817 0.067
R5260 VN.n11655 VN.n11654 0.067
R5261 VN.n11748 VN.n11746 0.067
R5262 VN.n11748 VN.n11747 0.067
R5263 VN.n11759 VN.n11757 0.067
R5264 VN.n11759 VN.n11758 0.067
R5265 VN.n11808 VN.n11807 0.067
R5266 VN.n11808 VN.n11806 0.067
R5267 VN.n11797 VN.n11796 0.067
R5268 VN.n11797 VN.n11795 0.067
R5269 VN.n11542 VN.n11528 0.067
R5270 VN.n11542 VN.n11527 0.067
R5271 VN.n9862 VN.n9848 0.067
R5272 VN.n9862 VN.n9846 0.067
R5273 VN.n9014 VN.n9000 0.067
R5274 VN.n9014 VN.n8999 0.067
R5275 VN.n8181 VN.n8167 0.067
R5276 VN.n8181 VN.n8166 0.067
R5277 VN.n7370 VN.n7356 0.067
R5278 VN.n7370 VN.n7355 0.067
R5279 VN.n6577 VN.n6563 0.067
R5280 VN.n6577 VN.n6562 0.067
R5281 VN.n5801 VN.n5787 0.067
R5282 VN.n5801 VN.n5786 0.067
R5283 VN.n5038 VN.n5024 0.067
R5284 VN.n5038 VN.n5023 0.067
R5285 VN.n4297 VN.n4283 0.067
R5286 VN.n4297 VN.n4282 0.067
R5287 VN.n3569 VN.n3555 0.067
R5288 VN.n3569 VN.n3554 0.067
R5289 VN.n2863 VN.n2849 0.067
R5290 VN.n2863 VN.n2848 0.067
R5291 VN.n2170 VN.n2156 0.067
R5292 VN.n2170 VN.n2155 0.067
R5293 VN.n1496 VN.n1482 0.067
R5294 VN.n1496 VN.n1481 0.067
R5295 VN.n846 VN.n832 0.067
R5296 VN.n846 VN.n831 0.067
R5297 VN.n13135 VN.n13119 0.067
R5298 VN.n13135 VN.n13121 0.067
R5299 VN.n11655 VN.n11653 0.067
R5300 VN.n12115 VN.n12114 0.066
R5301 VN.n11543 VN.n11526 0.065
R5302 VN.n820 VN.n819 0.063
R5303 VN.n11681 VN.n11680 0.063
R5304 VN.n12165 VN.n12164 0.063
R5305 VN.n11465 VN.n11464 0.063
R5306 VN.n10297 VN.n10296 0.063
R5307 VN.n9414 VN.n9413 0.063
R5308 VN.n8552 VN.n8551 0.063
R5309 VN.n7707 VN.n7706 0.063
R5310 VN.n7318 VN.n7317 0.063
R5311 VN.n6075 VN.n6074 0.063
R5312 VN.n5283 VN.n5282 0.063
R5313 VN.n4508 VN.n4507 0.063
R5314 VN.n3751 VN.n3750 0.063
R5315 VN.n3011 VN.n3010 0.063
R5316 VN.n2289 VN.n2288 0.063
R5317 VN.n1581 VN.n1580 0.063
R5318 VN.n898 VN.n897 0.063
R5319 VN.n227 VN.n226 0.063
R5320 VN.n11069 VN.n11044 0.063
R5321 VN.n10209 VN.n10208 0.063
R5322 VN.n9326 VN.n9325 0.063
R5323 VN.n8464 VN.n8463 0.063
R5324 VN.n7619 VN.n7618 0.063
R5325 VN.n7230 VN.n7229 0.063
R5326 VN.n5987 VN.n5986 0.063
R5327 VN.n5195 VN.n5194 0.063
R5328 VN.n4420 VN.n4419 0.063
R5329 VN.n3663 VN.n3662 0.063
R5330 VN.n2923 VN.n2922 0.063
R5331 VN.n2201 VN.n2200 0.063
R5332 VN.n11441 VN.n11422 0.063
R5333 VN.n10263 VN.n10250 0.063
R5334 VN.n9380 VN.n9367 0.063
R5335 VN.n8518 VN.n8505 0.063
R5336 VN.n7673 VN.n7660 0.063
R5337 VN.n7284 VN.n7271 0.063
R5338 VN.n6041 VN.n6028 0.063
R5339 VN.n5249 VN.n5236 0.063
R5340 VN.n4474 VN.n4461 0.063
R5341 VN.n3717 VN.n3704 0.063
R5342 VN.n2977 VN.n2964 0.063
R5343 VN.n2255 VN.n2242 0.063
R5344 VN.n1550 VN.n1537 0.063
R5345 VN.n864 VN.n851 0.063
R5346 VN.n12144 VN.n12125 0.063
R5347 VN.n2889 VN.n2868 0.063
R5348 VN.n3629 VN.n3608 0.063
R5349 VN.n4386 VN.n4365 0.063
R5350 VN.n5161 VN.n5140 0.063
R5351 VN.n5953 VN.n5932 0.063
R5352 VN.n7196 VN.n7175 0.063
R5353 VN.n7585 VN.n7564 0.063
R5354 VN.n8430 VN.n8409 0.063
R5355 VN.n9292 VN.n9271 0.063
R5356 VN.n10174 VN.n10153 0.063
R5357 VN.n11036 VN.n11018 0.063
R5358 VN.n12059 VN.n12044 0.063
R5359 VN.n11009 VN.n11008 0.063
R5360 VN.n10145 VN.n10144 0.063
R5361 VN.n9263 VN.n9262 0.063
R5362 VN.n8401 VN.n8400 0.063
R5363 VN.n7556 VN.n7555 0.063
R5364 VN.n7167 VN.n7166 0.063
R5365 VN.n5924 VN.n5923 0.063
R5366 VN.n5132 VN.n5131 0.063
R5367 VN.n4357 VN.n4356 0.063
R5368 VN.n3600 VN.n3599 0.063
R5369 VN.n4323 VN.n4302 0.063
R5370 VN.n5098 VN.n5077 0.063
R5371 VN.n5890 VN.n5869 0.063
R5372 VN.n7133 VN.n7112 0.063
R5373 VN.n7522 VN.n7501 0.063
R5374 VN.n8367 VN.n8346 0.063
R5375 VN.n9229 VN.n9208 0.063
R5376 VN.n10111 VN.n10090 0.063
R5377 VN.n10980 VN.n10960 0.063
R5378 VN.n12014 VN.n11999 0.063
R5379 VN.n10951 VN.n10950 0.063
R5380 VN.n10082 VN.n10081 0.063
R5381 VN.n9200 VN.n9199 0.063
R5382 VN.n8338 VN.n8337 0.063
R5383 VN.n7493 VN.n7492 0.063
R5384 VN.n7104 VN.n7103 0.063
R5385 VN.n5861 VN.n5860 0.063
R5386 VN.n5069 VN.n5068 0.063
R5387 VN.n5827 VN.n5806 0.063
R5388 VN.n7070 VN.n7049 0.063
R5389 VN.n7459 VN.n7438 0.063
R5390 VN.n8304 VN.n8283 0.063
R5391 VN.n9166 VN.n9145 0.063
R5392 VN.n10048 VN.n10027 0.063
R5393 VN.n10922 VN.n10902 0.063
R5394 VN.n11969 VN.n11954 0.063
R5395 VN.n10893 VN.n10892 0.063
R5396 VN.n10019 VN.n10018 0.063
R5397 VN.n9137 VN.n9136 0.063
R5398 VN.n8275 VN.n8274 0.063
R5399 VN.n7430 VN.n7429 0.063
R5400 VN.n7041 VN.n7040 0.063
R5401 VN.n10835 VN.n10834 0.063
R5402 VN.n9956 VN.n9955 0.063
R5403 VN.n9074 VN.n9073 0.063
R5404 VN.n8212 VN.n8211 0.063
R5405 VN.n9040 VN.n9019 0.063
R5406 VN.n9922 VN.n9901 0.063
R5407 VN.n10806 VN.n10786 0.063
R5408 VN.n11876 VN.n11647 0.063
R5409 VN.n10777 VN.n10776 0.063
R5410 VN.n9893 VN.n9892 0.063
R5411 VN.n10748 VN.n10728 0.063
R5412 VN.n11617 VN.n11602 0.063
R5413 VN.n11567 VN.n11566 0.063
R5414 VN.n11924 VN.n11905 0.063
R5415 VN.n10864 VN.n10843 0.063
R5416 VN.n9985 VN.n9964 0.063
R5417 VN.n9103 VN.n9082 0.063
R5418 VN.n8241 VN.n8220 0.063
R5419 VN.n7396 VN.n7375 0.063
R5420 VN.n11673 VN.n11672 0.062
R5421 VN.n11716 VN.n11715 0.062
R5422 VN.n11727 VN.n11726 0.062
R5423 VN.n11738 VN.n11737 0.062
R5424 VN.n11749 VN.n11748 0.062
R5425 VN.n11760 VN.n11759 0.062
R5426 VN.n11769 VN.n11768 0.062
R5427 VN.n11693 VN.n11692 0.061
R5428 VN.n181 VN.n179 0.061
R5429 VN.n11855 VN.n11854 0.06
R5430 VN.n11831 VN.n11830 0.06
R5431 VN.n11820 VN.n11819 0.06
R5432 VN.n11809 VN.n11808 0.06
R5433 VN.n11798 VN.n11797 0.06
R5434 VN.n11660 VN.n11659 0.06
R5435 VN.n12255 VN.n12254 0.059
R5436 VN.n236 VN.n235 0.059
R5437 VN.n10192 VN.n10182 0.059
R5438 VN.n11708 VN.n11707 0.059
R5439 VN.n13136 VN.n13135 0.058
R5440 VN.n9829 VN.n9828 0.058
R5441 VN.n8983 VN.n8982 0.058
R5442 VN.n8150 VN.n8149 0.058
R5443 VN.n7339 VN.n7338 0.058
R5444 VN.n6546 VN.n6545 0.058
R5445 VN.n5770 VN.n5769 0.058
R5446 VN.n5007 VN.n5006 0.058
R5447 VN.n4266 VN.n4265 0.058
R5448 VN.n3538 VN.n3537 0.058
R5449 VN.n2832 VN.n2831 0.058
R5450 VN.n2139 VN.n2138 0.058
R5451 VN.n1465 VN.n1464 0.058
R5452 VN.n11543 VN.n11542 0.058
R5453 VN.n170 VN.n169 0.056
R5454 VN.n11791 VN.n11790 0.055
R5455 VN.n13115 VN.n13114 0.055
R5456 VN.n12174 VN.n12173 0.055
R5457 VN.n11517 VN.n11516 0.055
R5458 VN.n10699 VN.n10698 0.055
R5459 VN.n9819 VN.n9818 0.055
R5460 VN.n8973 VN.n8972 0.055
R5461 VN.n8140 VN.n8139 0.055
R5462 VN.n7329 VN.n7328 0.055
R5463 VN.n6536 VN.n6535 0.055
R5464 VN.n5760 VN.n5759 0.055
R5465 VN.n4997 VN.n4996 0.055
R5466 VN.n4256 VN.n4255 0.055
R5467 VN.n3528 VN.n3527 0.055
R5468 VN.n2822 VN.n2821 0.055
R5469 VN.n2129 VN.n2128 0.055
R5470 VN.n1455 VN.n1454 0.055
R5471 VN.n802 VN.n801 0.055
R5472 VN.n11380 VN.n11366 0.054
R5473 VN.n12367 VN.n12350 0.054
R5474 VN.n2508 VN.n2495 0.054
R5475 VN.n1816 VN.n1802 0.054
R5476 VN.n1143 VN.n1130 0.054
R5477 VN.n490 VN.n473 0.054
R5478 VN.n12698 VN.n12683 0.054
R5479 VN.n3940 VN.n3927 0.054
R5480 VN.n3213 VN.n3199 0.054
R5481 VN.n5442 VN.n5429 0.054
R5482 VN.n4680 VN.n4666 0.054
R5483 VN.n6217 VN.n6203 0.054
R5484 VN.n6645 VN.n6632 0.054
R5485 VN.n8651 VN.n8638 0.054
R5486 VN.n7819 VN.n7805 0.054
R5487 VN.n10352 VN.n10339 0.054
R5488 VN.n9496 VN.n9482 0.054
R5489 VN.n11854 VN.n11853 0.054
R5490 VN.n12168 VN.n12167 0.054
R5491 VN.n12265 VN.n12264 0.054
R5492 VN.n12716 VN.n12715 0.054
R5493 VN.n230 VN.n229 0.054
R5494 VN.n527 VN.n526 0.054
R5495 VN.n901 VN.n900 0.054
R5496 VN.n1202 VN.n1201 0.054
R5497 VN.n1584 VN.n1583 0.054
R5498 VN.n1892 VN.n1891 0.054
R5499 VN.n2292 VN.n2291 0.054
R5500 VN.n2601 VN.n2600 0.054
R5501 VN.n3014 VN.n3013 0.054
R5502 VN.n3323 VN.n3322 0.054
R5503 VN.n3754 VN.n3753 0.054
R5504 VN.n4067 VN.n4066 0.054
R5505 VN.n4511 VN.n4510 0.054
R5506 VN.n4824 VN.n4823 0.054
R5507 VN.n5286 VN.n5285 0.054
R5508 VN.n5603 VN.n5602 0.054
R5509 VN.n6078 VN.n6077 0.054
R5510 VN.n6395 VN.n6394 0.054
R5511 VN.n7321 VN.n7320 0.054
R5512 VN.n6840 VN.n6839 0.054
R5513 VN.n7710 VN.n7709 0.054
R5514 VN.n8031 VN.n8030 0.054
R5515 VN.n8555 VN.n8554 0.054
R5516 VN.n8880 VN.n8879 0.054
R5517 VN.n9417 VN.n9416 0.054
R5518 VN.n9742 VN.n9741 0.054
R5519 VN.n10300 VN.n10299 0.054
R5520 VN.n10630 VN.n10629 0.054
R5521 VN.n11468 VN.n11467 0.054
R5522 VN.n11124 VN.n11123 0.054
R5523 VN.n12039 VN.n12038 0.054
R5524 VN.n3045 VN.n3044 0.054
R5525 VN.n3231 VN.n3230 0.054
R5526 VN.n3603 VN.n3602 0.054
R5527 VN.n3975 VN.n3974 0.054
R5528 VN.n4360 VN.n4359 0.054
R5529 VN.n4732 VN.n4731 0.054
R5530 VN.n5135 VN.n5134 0.054
R5531 VN.n5511 VN.n5510 0.054
R5532 VN.n5927 VN.n5926 0.054
R5533 VN.n6303 VN.n6302 0.054
R5534 VN.n7170 VN.n7169 0.054
R5535 VN.n6748 VN.n6747 0.054
R5536 VN.n7559 VN.n7558 0.054
R5537 VN.n7939 VN.n7938 0.054
R5538 VN.n8404 VN.n8403 0.054
R5539 VN.n8788 VN.n8787 0.054
R5540 VN.n9266 VN.n9265 0.054
R5541 VN.n9650 VN.n9649 0.054
R5542 VN.n10148 VN.n10147 0.054
R5543 VN.n10528 VN.n10527 0.054
R5544 VN.n11012 VN.n11011 0.054
R5545 VN.n11194 VN.n11193 0.054
R5546 VN.n12062 VN.n12061 0.054
R5547 VN.n2326 VN.n2325 0.054
R5548 VN.n2526 VN.n2525 0.054
R5549 VN.n2892 VN.n2891 0.054
R5550 VN.n3248 VN.n3247 0.054
R5551 VN.n3632 VN.n3631 0.054
R5552 VN.n3992 VN.n3991 0.054
R5553 VN.n4389 VN.n4388 0.054
R5554 VN.n4749 VN.n4748 0.054
R5555 VN.n5164 VN.n5163 0.054
R5556 VN.n5528 VN.n5527 0.054
R5557 VN.n5956 VN.n5955 0.054
R5558 VN.n6320 VN.n6319 0.054
R5559 VN.n7199 VN.n7198 0.054
R5560 VN.n6765 VN.n6764 0.054
R5561 VN.n7588 VN.n7587 0.054
R5562 VN.n7956 VN.n7955 0.054
R5563 VN.n8433 VN.n8432 0.054
R5564 VN.n8805 VN.n8804 0.054
R5565 VN.n9295 VN.n9294 0.054
R5566 VN.n9667 VN.n9666 0.054
R5567 VN.n10177 VN.n10176 0.054
R5568 VN.n10548 VN.n10547 0.054
R5569 VN.n10569 VN.n10568 0.054
R5570 VN.n11072 VN.n11071 0.054
R5571 VN.n11160 VN.n11159 0.054
R5572 VN.n12084 VN.n12083 0.054
R5573 VN.n10212 VN.n10211 0.054
R5574 VN.n9329 VN.n9328 0.054
R5575 VN.n8467 VN.n8466 0.054
R5576 VN.n7622 VN.n7621 0.054
R5577 VN.n7233 VN.n7232 0.054
R5578 VN.n5990 VN.n5989 0.054
R5579 VN.n5198 VN.n5197 0.054
R5580 VN.n4423 VN.n4422 0.054
R5581 VN.n3666 VN.n3665 0.054
R5582 VN.n2926 VN.n2925 0.054
R5583 VN.n2204 VN.n2203 0.054
R5584 VN.n1618 VN.n1617 0.054
R5585 VN.n1834 VN.n1833 0.054
R5586 VN.n2543 VN.n2542 0.054
R5587 VN.n3265 VN.n3264 0.054
R5588 VN.n4009 VN.n4008 0.054
R5589 VN.n4766 VN.n4765 0.054
R5590 VN.n5545 VN.n5544 0.054
R5591 VN.n6337 VN.n6336 0.054
R5592 VN.n6782 VN.n6781 0.054
R5593 VN.n7973 VN.n7972 0.054
R5594 VN.n8822 VN.n8821 0.054
R5595 VN.n9684 VN.n9683 0.054
R5596 VN.n11417 VN.n11416 0.054
R5597 VN.n11388 VN.n11387 0.054
R5598 VN.n12118 VN.n12117 0.054
R5599 VN.n931 VN.n930 0.054
R5600 VN.n1166 VN.n1165 0.054
R5601 VN.n1529 VN.n1528 0.054
R5602 VN.n1856 VN.n1855 0.054
R5603 VN.n2237 VN.n2236 0.054
R5604 VN.n2565 VN.n2564 0.054
R5605 VN.n2959 VN.n2958 0.054
R5606 VN.n3287 VN.n3286 0.054
R5607 VN.n3699 VN.n3698 0.054
R5608 VN.n4031 VN.n4030 0.054
R5609 VN.n4456 VN.n4455 0.054
R5610 VN.n4788 VN.n4787 0.054
R5611 VN.n5231 VN.n5230 0.054
R5612 VN.n5567 VN.n5566 0.054
R5613 VN.n6023 VN.n6022 0.054
R5614 VN.n6359 VN.n6358 0.054
R5615 VN.n7266 VN.n7265 0.054
R5616 VN.n6804 VN.n6803 0.054
R5617 VN.n7655 VN.n7654 0.054
R5618 VN.n7995 VN.n7994 0.054
R5619 VN.n8500 VN.n8499 0.054
R5620 VN.n8844 VN.n8843 0.054
R5621 VN.n9362 VN.n9361 0.054
R5622 VN.n9706 VN.n9705 0.054
R5623 VN.n10245 VN.n10244 0.054
R5624 VN.n10591 VN.n10590 0.054
R5625 VN.n11444 VN.n11443 0.054
R5626 VN.n11144 VN.n11143 0.054
R5627 VN.n10612 VN.n10611 0.054
R5628 VN.n10266 VN.n10265 0.054
R5629 VN.n9725 VN.n9724 0.054
R5630 VN.n9383 VN.n9382 0.054
R5631 VN.n8863 VN.n8862 0.054
R5632 VN.n8521 VN.n8520 0.054
R5633 VN.n8014 VN.n8013 0.054
R5634 VN.n7676 VN.n7675 0.054
R5635 VN.n6823 VN.n6822 0.054
R5636 VN.n7287 VN.n7286 0.054
R5637 VN.n6378 VN.n6377 0.054
R5638 VN.n6044 VN.n6043 0.054
R5639 VN.n5586 VN.n5585 0.054
R5640 VN.n5252 VN.n5251 0.054
R5641 VN.n4807 VN.n4806 0.054
R5642 VN.n4477 VN.n4476 0.054
R5643 VN.n4050 VN.n4049 0.054
R5644 VN.n3720 VN.n3719 0.054
R5645 VN.n3306 VN.n3305 0.054
R5646 VN.n2980 VN.n2979 0.054
R5647 VN.n2584 VN.n2583 0.054
R5648 VN.n2258 VN.n2257 0.054
R5649 VN.n1875 VN.n1874 0.054
R5650 VN.n1535 VN.n1534 0.054
R5651 VN.n1185 VN.n1184 0.054
R5652 VN.n867 VN.n866 0.054
R5653 VN.n510 VN.n509 0.054
R5654 VN.n259 VN.n258 0.054
R5655 VN.n12147 VN.n12146 0.054
R5656 VN.n11039 VN.n11038 0.054
R5657 VN.n11178 VN.n11177 0.054
R5658 VN.n11994 VN.n11993 0.054
R5659 VN.n4542 VN.n4541 0.054
R5660 VN.n4698 VN.n4697 0.054
R5661 VN.n5072 VN.n5071 0.054
R5662 VN.n5477 VN.n5476 0.054
R5663 VN.n5864 VN.n5863 0.054
R5664 VN.n6269 VN.n6268 0.054
R5665 VN.n7107 VN.n7106 0.054
R5666 VN.n6714 VN.n6713 0.054
R5667 VN.n7496 VN.n7495 0.054
R5668 VN.n7905 VN.n7904 0.054
R5669 VN.n8341 VN.n8340 0.054
R5670 VN.n8754 VN.n8753 0.054
R5671 VN.n9203 VN.n9202 0.054
R5672 VN.n9616 VN.n9615 0.054
R5673 VN.n10085 VN.n10084 0.054
R5674 VN.n10493 VN.n10492 0.054
R5675 VN.n10954 VN.n10953 0.054
R5676 VN.n11228 VN.n11227 0.054
R5677 VN.n12017 VN.n12016 0.054
R5678 VN.n3788 VN.n3787 0.054
R5679 VN.n3958 VN.n3957 0.054
R5680 VN.n4326 VN.n4325 0.054
R5681 VN.n4715 VN.n4714 0.054
R5682 VN.n5101 VN.n5100 0.054
R5683 VN.n5494 VN.n5493 0.054
R5684 VN.n5893 VN.n5892 0.054
R5685 VN.n6286 VN.n6285 0.054
R5686 VN.n7136 VN.n7135 0.054
R5687 VN.n6731 VN.n6730 0.054
R5688 VN.n7525 VN.n7524 0.054
R5689 VN.n7922 VN.n7921 0.054
R5690 VN.n8370 VN.n8369 0.054
R5691 VN.n8771 VN.n8770 0.054
R5692 VN.n9232 VN.n9231 0.054
R5693 VN.n9633 VN.n9632 0.054
R5694 VN.n10114 VN.n10113 0.054
R5695 VN.n10510 VN.n10509 0.054
R5696 VN.n10983 VN.n10982 0.054
R5697 VN.n11212 VN.n11211 0.054
R5698 VN.n11949 VN.n11948 0.054
R5699 VN.n6109 VN.n6108 0.054
R5700 VN.n6235 VN.n6234 0.054
R5701 VN.n7044 VN.n7043 0.054
R5702 VN.n6680 VN.n6679 0.054
R5703 VN.n7433 VN.n7432 0.054
R5704 VN.n7871 VN.n7870 0.054
R5705 VN.n8278 VN.n8277 0.054
R5706 VN.n8720 VN.n8719 0.054
R5707 VN.n9140 VN.n9139 0.054
R5708 VN.n9582 VN.n9581 0.054
R5709 VN.n10022 VN.n10021 0.054
R5710 VN.n10458 VN.n10457 0.054
R5711 VN.n10896 VN.n10895 0.054
R5712 VN.n11262 VN.n11261 0.054
R5713 VN.n11972 VN.n11971 0.054
R5714 VN.n5320 VN.n5319 0.054
R5715 VN.n5460 VN.n5459 0.054
R5716 VN.n5830 VN.n5829 0.054
R5717 VN.n6252 VN.n6251 0.054
R5718 VN.n7073 VN.n7072 0.054
R5719 VN.n6697 VN.n6696 0.054
R5720 VN.n7462 VN.n7461 0.054
R5721 VN.n7888 VN.n7887 0.054
R5722 VN.n8307 VN.n8306 0.054
R5723 VN.n8737 VN.n8736 0.054
R5724 VN.n9169 VN.n9168 0.054
R5725 VN.n9599 VN.n9598 0.054
R5726 VN.n10051 VN.n10050 0.054
R5727 VN.n10475 VN.n10474 0.054
R5728 VN.n10925 VN.n10924 0.054
R5729 VN.n11246 VN.n11245 0.054
R5730 VN.n6663 VN.n6662 0.054
R5731 VN.n7399 VN.n7398 0.054
R5732 VN.n7854 VN.n7853 0.054
R5733 VN.n8244 VN.n8243 0.054
R5734 VN.n8703 VN.n8702 0.054
R5735 VN.n9106 VN.n9105 0.054
R5736 VN.n9565 VN.n9564 0.054
R5737 VN.n9988 VN.n9987 0.054
R5738 VN.n10440 VN.n10439 0.054
R5739 VN.n10867 VN.n10866 0.054
R5740 VN.n11279 VN.n11278 0.054
R5741 VN.n11927 VN.n11926 0.054
R5742 VN.n11900 VN.n11899 0.054
R5743 VN.n7741 VN.n7740 0.054
R5744 VN.n7837 VN.n7836 0.054
R5745 VN.n8215 VN.n8214 0.054
R5746 VN.n8686 VN.n8685 0.054
R5747 VN.n9077 VN.n9076 0.054
R5748 VN.n9548 VN.n9547 0.054
R5749 VN.n9959 VN.n9958 0.054
R5750 VN.n10423 VN.n10422 0.054
R5751 VN.n10838 VN.n10837 0.054
R5752 VN.n11295 VN.n11294 0.054
R5753 VN.n11642 VN.n11641 0.054
R5754 VN.n9448 VN.n9447 0.054
R5755 VN.n9514 VN.n9513 0.054
R5756 VN.n9896 VN.n9895 0.054
R5757 VN.n10388 VN.n10387 0.054
R5758 VN.n10780 VN.n10779 0.054
R5759 VN.n11329 VN.n11328 0.054
R5760 VN.n11879 VN.n11878 0.054
R5761 VN.n8589 VN.n8588 0.054
R5762 VN.n8669 VN.n8668 0.054
R5763 VN.n9043 VN.n9042 0.054
R5764 VN.n9531 VN.n9530 0.054
R5765 VN.n9925 VN.n9924 0.054
R5766 VN.n10405 VN.n10404 0.054
R5767 VN.n10809 VN.n10808 0.054
R5768 VN.n11313 VN.n11312 0.054
R5769 VN.n11597 VN.n11596 0.054
R5770 VN.n11495 VN.n11494 0.054
R5771 VN.n11363 VN.n11362 0.054
R5772 VN.n11620 VN.n11619 0.054
R5773 VN.n10334 VN.n10333 0.054
R5774 VN.n10370 VN.n10369 0.054
R5775 VN.n10751 VN.n10750 0.054
R5776 VN.n11347 VN.n11346 0.054
R5777 VN.n11103 VN.n11102 0.054
R5778 VN.n11512 VN.n11511 0.054
R5779 VN.n10656 VN.n10655 0.054
R5780 VN.n10682 VN.n10681 0.054
R5781 VN.n9763 VN.n9762 0.054
R5782 VN.n9468 VN.n9467 0.054
R5783 VN.n8901 VN.n8900 0.054
R5784 VN.n8609 VN.n8608 0.054
R5785 VN.n8052 VN.n8051 0.054
R5786 VN.n7761 VN.n7760 0.054
R5787 VN.n6861 VN.n6860 0.054
R5788 VN.n7010 VN.n7009 0.054
R5789 VN.n6416 VN.n6415 0.054
R5790 VN.n6129 VN.n6128 0.054
R5791 VN.n5624 VN.n5623 0.054
R5792 VN.n5340 VN.n5339 0.054
R5793 VN.n4845 VN.n4844 0.054
R5794 VN.n4562 VN.n4561 0.054
R5795 VN.n4088 VN.n4087 0.054
R5796 VN.n3808 VN.n3807 0.054
R5797 VN.n3344 VN.n3343 0.054
R5798 VN.n3065 VN.n3064 0.054
R5799 VN.n2622 VN.n2621 0.054
R5800 VN.n2346 VN.n2345 0.054
R5801 VN.n1913 VN.n1912 0.054
R5802 VN.n1638 VN.n1637 0.054
R5803 VN.n1223 VN.n1222 0.054
R5804 VN.n951 VN.n950 0.054
R5805 VN.n548 VN.n547 0.054
R5806 VN.n279 VN.n278 0.054
R5807 VN.n12293 VN.n12292 0.054
R5808 VN.n12320 VN.n12319 0.054
R5809 VN.n12275 VN.n12274 0.054
R5810 VN.n10650 VN.n10649 0.054
R5811 VN.n10697 VN.n10696 0.054
R5812 VN.n12623 VN.n12622 0.054
R5813 VN.n12638 VN.n12637 0.054
R5814 VN.n12336 VN.n12335 0.054
R5815 VN.n294 VN.n293 0.054
R5816 VN.n564 VN.n563 0.054
R5817 VN.n966 VN.n965 0.054
R5818 VN.n1239 VN.n1238 0.054
R5819 VN.n1653 VN.n1652 0.054
R5820 VN.n1929 VN.n1928 0.054
R5821 VN.n2361 VN.n2360 0.054
R5822 VN.n2638 VN.n2637 0.054
R5823 VN.n3080 VN.n3079 0.054
R5824 VN.n3360 VN.n3359 0.054
R5825 VN.n3823 VN.n3822 0.054
R5826 VN.n4104 VN.n4103 0.054
R5827 VN.n4577 VN.n4576 0.054
R5828 VN.n4861 VN.n4860 0.054
R5829 VN.n5355 VN.n5354 0.054
R5830 VN.n5640 VN.n5639 0.054
R5831 VN.n6144 VN.n6143 0.054
R5832 VN.n6432 VN.n6431 0.054
R5833 VN.n6990 VN.n6989 0.054
R5834 VN.n6877 VN.n6876 0.054
R5835 VN.n7776 VN.n7775 0.054
R5836 VN.n8068 VN.n8067 0.054
R5837 VN.n8624 VN.n8623 0.054
R5838 VN.n8917 VN.n8916 0.054
R5839 VN.n9802 VN.n9801 0.054
R5840 VN.n9788 VN.n9787 0.054
R5841 VN.n9785 VN.n9784 0.054
R5842 VN.n9817 VN.n9816 0.054
R5843 VN.n12428 VN.n12427 0.054
R5844 VN.n12669 VN.n12668 0.054
R5845 VN.n12654 VN.n12653 0.054
R5846 VN.n309 VN.n308 0.054
R5847 VN.n580 VN.n579 0.054
R5848 VN.n981 VN.n980 0.054
R5849 VN.n1255 VN.n1254 0.054
R5850 VN.n1668 VN.n1667 0.054
R5851 VN.n1945 VN.n1944 0.054
R5852 VN.n2376 VN.n2375 0.054
R5853 VN.n2654 VN.n2653 0.054
R5854 VN.n3095 VN.n3094 0.054
R5855 VN.n3376 VN.n3375 0.054
R5856 VN.n3838 VN.n3837 0.054
R5857 VN.n4120 VN.n4119 0.054
R5858 VN.n4592 VN.n4591 0.054
R5859 VN.n4877 VN.n4876 0.054
R5860 VN.n5370 VN.n5369 0.054
R5861 VN.n5656 VN.n5655 0.054
R5862 VN.n6159 VN.n6158 0.054
R5863 VN.n6448 VN.n6447 0.054
R5864 VN.n6975 VN.n6974 0.054
R5865 VN.n6893 VN.n6892 0.054
R5866 VN.n7791 VN.n7790 0.054
R5867 VN.n8084 VN.n8083 0.054
R5868 VN.n8956 VN.n8955 0.054
R5869 VN.n8942 VN.n8941 0.054
R5870 VN.n8939 VN.n8938 0.054
R5871 VN.n8971 VN.n8970 0.054
R5872 VN.n12444 VN.n12443 0.054
R5873 VN.n12780 VN.n12779 0.054
R5874 VN.n12765 VN.n12764 0.054
R5875 VN.n324 VN.n323 0.054
R5876 VN.n596 VN.n595 0.054
R5877 VN.n996 VN.n995 0.054
R5878 VN.n1271 VN.n1270 0.054
R5879 VN.n1683 VN.n1682 0.054
R5880 VN.n1961 VN.n1960 0.054
R5881 VN.n2391 VN.n2390 0.054
R5882 VN.n2670 VN.n2669 0.054
R5883 VN.n3110 VN.n3109 0.054
R5884 VN.n3392 VN.n3391 0.054
R5885 VN.n3853 VN.n3852 0.054
R5886 VN.n4136 VN.n4135 0.054
R5887 VN.n4607 VN.n4606 0.054
R5888 VN.n4893 VN.n4892 0.054
R5889 VN.n5385 VN.n5384 0.054
R5890 VN.n5672 VN.n5671 0.054
R5891 VN.n6174 VN.n6173 0.054
R5892 VN.n6464 VN.n6463 0.054
R5893 VN.n6960 VN.n6959 0.054
R5894 VN.n6909 VN.n6908 0.054
R5895 VN.n8123 VN.n8122 0.054
R5896 VN.n8109 VN.n8108 0.054
R5897 VN.n8106 VN.n8105 0.054
R5898 VN.n8138 VN.n8137 0.054
R5899 VN.n12460 VN.n12459 0.054
R5900 VN.n12788 VN.n12787 0.054
R5901 VN.n12799 VN.n12798 0.054
R5902 VN.n339 VN.n338 0.054
R5903 VN.n612 VN.n611 0.054
R5904 VN.n1011 VN.n1010 0.054
R5905 VN.n1287 VN.n1286 0.054
R5906 VN.n1698 VN.n1697 0.054
R5907 VN.n1977 VN.n1976 0.054
R5908 VN.n2406 VN.n2405 0.054
R5909 VN.n2686 VN.n2685 0.054
R5910 VN.n3125 VN.n3124 0.054
R5911 VN.n3408 VN.n3407 0.054
R5912 VN.n3868 VN.n3867 0.054
R5913 VN.n4152 VN.n4151 0.054
R5914 VN.n4622 VN.n4621 0.054
R5915 VN.n4909 VN.n4908 0.054
R5916 VN.n5400 VN.n5399 0.054
R5917 VN.n5688 VN.n5687 0.054
R5918 VN.n6189 VN.n6188 0.054
R5919 VN.n6480 VN.n6479 0.054
R5920 VN.n6945 VN.n6944 0.054
R5921 VN.n6934 VN.n6933 0.054
R5922 VN.n6931 VN.n6930 0.054
R5923 VN.n6615 VN.n6614 0.054
R5924 VN.n12476 VN.n12475 0.054
R5925 VN.n12819 VN.n12818 0.054
R5926 VN.n12830 VN.n12829 0.054
R5927 VN.n354 VN.n353 0.054
R5928 VN.n628 VN.n627 0.054
R5929 VN.n1026 VN.n1025 0.054
R5930 VN.n1303 VN.n1302 0.054
R5931 VN.n1713 VN.n1712 0.054
R5932 VN.n1993 VN.n1992 0.054
R5933 VN.n2421 VN.n2420 0.054
R5934 VN.n2702 VN.n2701 0.054
R5935 VN.n3140 VN.n3139 0.054
R5936 VN.n3424 VN.n3423 0.054
R5937 VN.n3883 VN.n3882 0.054
R5938 VN.n4168 VN.n4167 0.054
R5939 VN.n4637 VN.n4636 0.054
R5940 VN.n4925 VN.n4924 0.054
R5941 VN.n5415 VN.n5414 0.054
R5942 VN.n5704 VN.n5703 0.054
R5943 VN.n6519 VN.n6518 0.054
R5944 VN.n6505 VN.n6504 0.054
R5945 VN.n6502 VN.n6501 0.054
R5946 VN.n6534 VN.n6533 0.054
R5947 VN.n12492 VN.n12491 0.054
R5948 VN.n12873 VN.n12872 0.054
R5949 VN.n12858 VN.n12857 0.054
R5950 VN.n369 VN.n368 0.054
R5951 VN.n644 VN.n643 0.054
R5952 VN.n1041 VN.n1040 0.054
R5953 VN.n1319 VN.n1318 0.054
R5954 VN.n1728 VN.n1727 0.054
R5955 VN.n2009 VN.n2008 0.054
R5956 VN.n2436 VN.n2435 0.054
R5957 VN.n2718 VN.n2717 0.054
R5958 VN.n3155 VN.n3154 0.054
R5959 VN.n3440 VN.n3439 0.054
R5960 VN.n3898 VN.n3897 0.054
R5961 VN.n4184 VN.n4183 0.054
R5962 VN.n4652 VN.n4651 0.054
R5963 VN.n4941 VN.n4940 0.054
R5964 VN.n5743 VN.n5742 0.054
R5965 VN.n5729 VN.n5728 0.054
R5966 VN.n5726 VN.n5725 0.054
R5967 VN.n5758 VN.n5757 0.054
R5968 VN.n12508 VN.n12507 0.054
R5969 VN.n12904 VN.n12903 0.054
R5970 VN.n12889 VN.n12888 0.054
R5971 VN.n384 VN.n383 0.054
R5972 VN.n660 VN.n659 0.054
R5973 VN.n1056 VN.n1055 0.054
R5974 VN.n1335 VN.n1334 0.054
R5975 VN.n1743 VN.n1742 0.054
R5976 VN.n2025 VN.n2024 0.054
R5977 VN.n2451 VN.n2450 0.054
R5978 VN.n2734 VN.n2733 0.054
R5979 VN.n3170 VN.n3169 0.054
R5980 VN.n3456 VN.n3455 0.054
R5981 VN.n3913 VN.n3912 0.054
R5982 VN.n4200 VN.n4199 0.054
R5983 VN.n4980 VN.n4979 0.054
R5984 VN.n4966 VN.n4965 0.054
R5985 VN.n4963 VN.n4962 0.054
R5986 VN.n4995 VN.n4994 0.054
R5987 VN.n12524 VN.n12523 0.054
R5988 VN.n12935 VN.n12934 0.054
R5989 VN.n12920 VN.n12919 0.054
R5990 VN.n399 VN.n398 0.054
R5991 VN.n676 VN.n675 0.054
R5992 VN.n1071 VN.n1070 0.054
R5993 VN.n1351 VN.n1350 0.054
R5994 VN.n1758 VN.n1757 0.054
R5995 VN.n2041 VN.n2040 0.054
R5996 VN.n2466 VN.n2465 0.054
R5997 VN.n2750 VN.n2749 0.054
R5998 VN.n3185 VN.n3184 0.054
R5999 VN.n3472 VN.n3471 0.054
R6000 VN.n4239 VN.n4238 0.054
R6001 VN.n4225 VN.n4224 0.054
R6002 VN.n4222 VN.n4221 0.054
R6003 VN.n4254 VN.n4253 0.054
R6004 VN.n12540 VN.n12539 0.054
R6005 VN.n12966 VN.n12965 0.054
R6006 VN.n12951 VN.n12950 0.054
R6007 VN.n414 VN.n413 0.054
R6008 VN.n692 VN.n691 0.054
R6009 VN.n1086 VN.n1085 0.054
R6010 VN.n1367 VN.n1366 0.054
R6011 VN.n1773 VN.n1772 0.054
R6012 VN.n2057 VN.n2056 0.054
R6013 VN.n2481 VN.n2480 0.054
R6014 VN.n2766 VN.n2765 0.054
R6015 VN.n3511 VN.n3510 0.054
R6016 VN.n3497 VN.n3496 0.054
R6017 VN.n3494 VN.n3493 0.054
R6018 VN.n3526 VN.n3525 0.054
R6019 VN.n12556 VN.n12555 0.054
R6020 VN.n12997 VN.n12996 0.054
R6021 VN.n12982 VN.n12981 0.054
R6022 VN.n429 VN.n428 0.054
R6023 VN.n708 VN.n707 0.054
R6024 VN.n1101 VN.n1100 0.054
R6025 VN.n1383 VN.n1382 0.054
R6026 VN.n1788 VN.n1787 0.054
R6027 VN.n2073 VN.n2072 0.054
R6028 VN.n2805 VN.n2804 0.054
R6029 VN.n2791 VN.n2790 0.054
R6030 VN.n2788 VN.n2787 0.054
R6031 VN.n2820 VN.n2819 0.054
R6032 VN.n12572 VN.n12571 0.054
R6033 VN.n13028 VN.n13027 0.054
R6034 VN.n13013 VN.n13012 0.054
R6035 VN.n444 VN.n443 0.054
R6036 VN.n724 VN.n723 0.054
R6037 VN.n1116 VN.n1115 0.054
R6038 VN.n1399 VN.n1398 0.054
R6039 VN.n2112 VN.n2111 0.054
R6040 VN.n2098 VN.n2097 0.054
R6041 VN.n2095 VN.n2094 0.054
R6042 VN.n2127 VN.n2126 0.054
R6043 VN.n12588 VN.n12587 0.054
R6044 VN.n13059 VN.n13058 0.054
R6045 VN.n13044 VN.n13043 0.054
R6046 VN.n459 VN.n458 0.054
R6047 VN.n740 VN.n739 0.054
R6048 VN.n1438 VN.n1437 0.054
R6049 VN.n1424 VN.n1423 0.054
R6050 VN.n1421 VN.n1420 0.054
R6051 VN.n1453 VN.n1452 0.054
R6052 VN.n12604 VN.n12603 0.054
R6053 VN.n13090 VN.n13089 0.054
R6054 VN.n13075 VN.n13074 0.054
R6055 VN.n778 VN.n777 0.054
R6056 VN.n764 VN.n763 0.054
R6057 VN.n761 VN.n760 0.054
R6058 VN.n800 VN.n799 0.054
R6059 VN.n12620 VN.n12619 0.054
R6060 VN.n13110 VN.n13109 0.054
R6061 VN.n12762 VN.n12761 0.054
R6062 VN.n12388 VN.n12387 0.054
R6063 VN.n12219 VN.n12218 0.054
R6064 VN.n12740 VN.n12739 0.054
R6065 VN.n11656 VN.n11655 0.053
R6066 VN.n17 VN.n16 0.053
R6067 VN.t76 VN.n6584 0.052
R6068 VN.n11374 VN.n11373 0.052
R6069 VN.n10347 VN.n10346 0.052
R6070 VN.n9492 VN.n9491 0.052
R6071 VN.n8646 VN.n8645 0.052
R6072 VN.n7815 VN.n7814 0.052
R6073 VN.n6640 VN.n6639 0.052
R6074 VN.n6211 VN.n6210 0.052
R6075 VN.n5437 VN.n5436 0.052
R6076 VN.n4676 VN.n4675 0.052
R6077 VN.n3935 VN.n3934 0.052
R6078 VN.n3209 VN.n3208 0.052
R6079 VN.n2503 VN.n2502 0.052
R6080 VN.n1812 VN.n1811 0.052
R6081 VN.n1138 VN.n1137 0.052
R6082 VN.n486 VN.n485 0.052
R6083 VN.n12693 VN.n12692 0.052
R6084 VN.n12363 VN.n12362 0.052
R6085 VN.n10725 VN.n10724 0.052
R6086 VN.n9774 VN.n9773 0.052
R6087 VN.n10705 VN.n10704 0.052
R6088 VN.n8928 VN.n8927 0.052
R6089 VN.n9825 VN.n9824 0.052
R6090 VN.n8095 VN.n8094 0.052
R6091 VN.n8979 VN.n8978 0.052
R6092 VN.n6920 VN.n6919 0.052
R6093 VN.n8146 VN.n8145 0.052
R6094 VN.n6491 VN.n6490 0.052
R6095 VN.n7335 VN.n7334 0.052
R6096 VN.n5715 VN.n5714 0.052
R6097 VN.n6542 VN.n6541 0.052
R6098 VN.n4952 VN.n4951 0.052
R6099 VN.n5766 VN.n5765 0.052
R6100 VN.n4211 VN.n4210 0.052
R6101 VN.n5003 VN.n5002 0.052
R6102 VN.n3483 VN.n3482 0.052
R6103 VN.n4262 VN.n4261 0.052
R6104 VN.n2777 VN.n2776 0.052
R6105 VN.n3534 VN.n3533 0.052
R6106 VN.n2084 VN.n2083 0.052
R6107 VN.n2828 VN.n2827 0.052
R6108 VN.n1410 VN.n1409 0.052
R6109 VN.n2135 VN.n2134 0.052
R6110 VN.n1461 VN.n1460 0.052
R6111 VN.n12732 VN.n12731 0.052
R6112 VN.n197 VN.n196 0.052
R6113 VN.t76 VN.n7327 0.051
R6114 VN.n1610 VN.n1608 0.051
R6115 VN.n2299 VN.n2298 0.051
R6116 VN.n3037 VN.n3035 0.051
R6117 VN.n3761 VN.n3760 0.051
R6118 VN.n4534 VN.n4532 0.051
R6119 VN.n5293 VN.n5292 0.051
R6120 VN.n6101 VN.n6099 0.051
R6121 VN.n6587 VN.n6585 0.051
R6122 VN.n7733 VN.n7731 0.051
R6123 VN.n8562 VN.n8561 0.051
R6124 VN.n9440 VN.n9438 0.051
R6125 VN.n10307 VN.n10306 0.051
R6126 VN.n11487 VN.n11485 0.051
R6127 VN.n11553 VN.n11551 0.051
R6128 VN.n27 VN.n26 0.051
R6129 VN.n29 VN.n28 0.051
R6130 VN.n93 VN.n92 0.051
R6131 VN.n95 VN.n94 0.051
R6132 VN.n11506 VN.n11496 0.051
R6133 VN.n12314 VN.n12300 0.051
R6134 VN.n12632 VN.n12344 0.051
R6135 VN.n12663 VN.n12662 0.051
R6136 VN.n12774 VN.n12773 0.051
R6137 VN.n12808 VN.n12807 0.051
R6138 VN.n12839 VN.n12838 0.051
R6139 VN.n12867 VN.n12866 0.051
R6140 VN.n12898 VN.n12897 0.051
R6141 VN.n12929 VN.n12928 0.051
R6142 VN.n12960 VN.n12959 0.051
R6143 VN.n12991 VN.n12990 0.051
R6144 VN.n13022 VN.n13021 0.051
R6145 VN.n13053 VN.n13052 0.051
R6146 VN.n13084 VN.n13083 0.051
R6147 VN.n12259 VN.n12258 0.05
R6148 VN.n1612 VN.n1611 0.05
R6149 VN.n253 VN.n239 0.05
R6150 VN.n12136 VN.n12135 0.05
R6151 VN.n2315 VN.n2314 0.05
R6152 VN.n2320 VN.n2301 0.05
R6153 VN.n3039 VN.n3038 0.05
R6154 VN.n3779 VN.n3776 0.05
R6155 VN.n3782 VN.n3763 0.05
R6156 VN.n4536 VN.n4535 0.05
R6157 VN.n5311 VN.n5308 0.05
R6158 VN.n5314 VN.n5295 0.05
R6159 VN.n6103 VN.n6102 0.05
R6160 VN.n6599 VN.n6596 0.05
R6161 VN.n7735 VN.n7734 0.05
R6162 VN.n8578 VN.n8577 0.05
R6163 VN.n8583 VN.n8564 0.05
R6164 VN.n9442 VN.n9441 0.05
R6165 VN.n10323 VN.n10322 0.05
R6166 VN.n10328 VN.n10309 0.05
R6167 VN.n11489 VN.n11488 0.05
R6168 VN.n11567 VN.n11554 0.05
R6169 VN.t76 VN.n6589 0.05
R6170 VN.n11414 VN.n11398 0.05
R6171 VN.n12161 VN.n12160 0.05
R6172 VN.n11571 VN.n11570 0.05
R6173 VN.n10580 VN.n10579 0.049
R6174 VN.n9695 VN.n9694 0.049
R6175 VN.n8833 VN.n8832 0.049
R6176 VN.n7984 VN.n7983 0.049
R6177 VN.n6793 VN.n6792 0.049
R6178 VN.n6348 VN.n6347 0.049
R6179 VN.n5556 VN.n5555 0.049
R6180 VN.n4777 VN.n4776 0.049
R6181 VN.n4020 VN.n4019 0.049
R6182 VN.n3276 VN.n3275 0.049
R6183 VN.n2554 VN.n2553 0.049
R6184 VN.n1845 VN.n1844 0.049
R6185 VN.n1155 VN.n1154 0.049
R6186 VN.n11394 VN.n11393 0.049
R6187 VN.n11135 VN.n11134 0.049
R6188 VN.n824 VN.n822 0.049
R6189 VN.n754 VN.n753 0.048
R6190 VN.n10723 VN.n10722 0.048
R6191 VN.n9863 VN.n9862 0.048
R6192 VN.n9015 VN.n9014 0.048
R6193 VN.n8182 VN.n8181 0.048
R6194 VN.n7371 VN.n7370 0.048
R6195 VN.n6578 VN.n6577 0.048
R6196 VN.n5802 VN.n5801 0.048
R6197 VN.n5039 VN.n5038 0.048
R6198 VN.n4298 VN.n4297 0.048
R6199 VN.n3570 VN.n3569 0.048
R6200 VN.n2864 VN.n2863 0.048
R6201 VN.n2171 VN.n2170 0.048
R6202 VN.n1497 VN.n1496 0.048
R6203 VN.n847 VN.n846 0.048
R6204 VN.n13137 VN.n13117 0.047
R6205 VN.n12165 VN.n12155 0.047
R6206 VN.n12259 VN.n12242 0.047
R6207 VN.n12713 VN.n12707 0.047
R6208 VN.n227 VN.n213 0.047
R6209 VN.n524 VN.n518 0.047
R6210 VN.n898 VN.n884 0.047
R6211 VN.n1199 VN.n1193 0.047
R6212 VN.n1581 VN.n1567 0.047
R6213 VN.n1889 VN.n1883 0.047
R6214 VN.n2289 VN.n2275 0.047
R6215 VN.n2598 VN.n2592 0.047
R6216 VN.n3011 VN.n2997 0.047
R6217 VN.n3320 VN.n3314 0.047
R6218 VN.n3751 VN.n3737 0.047
R6219 VN.n4064 VN.n4058 0.047
R6220 VN.n4508 VN.n4494 0.047
R6221 VN.n4821 VN.n4815 0.047
R6222 VN.n5283 VN.n5269 0.047
R6223 VN.n5600 VN.n5594 0.047
R6224 VN.n6075 VN.n6061 0.047
R6225 VN.n6392 VN.n6386 0.047
R6226 VN.n7318 VN.n7304 0.047
R6227 VN.n6837 VN.n6831 0.047
R6228 VN.n7707 VN.n7693 0.047
R6229 VN.n8028 VN.n8022 0.047
R6230 VN.n8552 VN.n8538 0.047
R6231 VN.n8877 VN.n8871 0.047
R6232 VN.n9414 VN.n9400 0.047
R6233 VN.n9739 VN.n9733 0.047
R6234 VN.n10297 VN.n10283 0.047
R6235 VN.n10627 VN.n10620 0.047
R6236 VN.n11465 VN.n11452 0.047
R6237 VN.n11118 VN.n11112 0.047
R6238 VN.n12036 VN.n12034 0.047
R6239 VN.n3039 VN.n3023 0.047
R6240 VN.n3228 VN.n3222 0.047
R6241 VN.n3600 VN.n3586 0.047
R6242 VN.n3972 VN.n3966 0.047
R6243 VN.n4357 VN.n4343 0.047
R6244 VN.n4729 VN.n4723 0.047
R6245 VN.n5132 VN.n5118 0.047
R6246 VN.n5508 VN.n5502 0.047
R6247 VN.n5924 VN.n5910 0.047
R6248 VN.n6300 VN.n6294 0.047
R6249 VN.n7167 VN.n7153 0.047
R6250 VN.n6745 VN.n6739 0.047
R6251 VN.n7556 VN.n7542 0.047
R6252 VN.n7936 VN.n7930 0.047
R6253 VN.n8401 VN.n8387 0.047
R6254 VN.n8785 VN.n8779 0.047
R6255 VN.n9263 VN.n9249 0.047
R6256 VN.n9647 VN.n9641 0.047
R6257 VN.n10145 VN.n10131 0.047
R6258 VN.n10525 VN.n10518 0.047
R6259 VN.n11009 VN.n11000 0.047
R6260 VN.n11188 VN.n11182 0.047
R6261 VN.n12059 VN.n12057 0.047
R6262 VN.n2320 VN.n2311 0.047
R6263 VN.n2523 VN.n2521 0.047
R6264 VN.n2889 VN.n2878 0.047
R6265 VN.n3245 VN.n3243 0.047
R6266 VN.n3629 VN.n3618 0.047
R6267 VN.n3989 VN.n3987 0.047
R6268 VN.n4386 VN.n4375 0.047
R6269 VN.n4746 VN.n4744 0.047
R6270 VN.n5161 VN.n5150 0.047
R6271 VN.n5525 VN.n5523 0.047
R6272 VN.n5953 VN.n5942 0.047
R6273 VN.n6317 VN.n6315 0.047
R6274 VN.n7196 VN.n7185 0.047
R6275 VN.n6762 VN.n6760 0.047
R6276 VN.n7585 VN.n7574 0.047
R6277 VN.n7953 VN.n7951 0.047
R6278 VN.n8430 VN.n8419 0.047
R6279 VN.n8802 VN.n8800 0.047
R6280 VN.n9292 VN.n9281 0.047
R6281 VN.n9664 VN.n9662 0.047
R6282 VN.n10174 VN.n10163 0.047
R6283 VN.n10545 VN.n10540 0.047
R6284 VN.n10566 VN.n10561 0.047
R6285 VN.n11069 VN.n11054 0.047
R6286 VN.n11154 VN.n11152 0.047
R6287 VN.n12081 VN.n12074 0.047
R6288 VN.n10209 VN.n10195 0.047
R6289 VN.n9326 VN.n9312 0.047
R6290 VN.n8464 VN.n8450 0.047
R6291 VN.n7619 VN.n7605 0.047
R6292 VN.n7230 VN.n7216 0.047
R6293 VN.n5987 VN.n5973 0.047
R6294 VN.n5195 VN.n5181 0.047
R6295 VN.n4420 VN.n4406 0.047
R6296 VN.n3663 VN.n3649 0.047
R6297 VN.n2923 VN.n2909 0.047
R6298 VN.n2201 VN.n2187 0.047
R6299 VN.n1612 VN.n1596 0.047
R6300 VN.n1831 VN.n1825 0.047
R6301 VN.n2540 VN.n2534 0.047
R6302 VN.n3262 VN.n3256 0.047
R6303 VN.n4006 VN.n4000 0.047
R6304 VN.n4763 VN.n4757 0.047
R6305 VN.n5542 VN.n5536 0.047
R6306 VN.n6334 VN.n6328 0.047
R6307 VN.n6779 VN.n6773 0.047
R6308 VN.n7970 VN.n7964 0.047
R6309 VN.n8819 VN.n8813 0.047
R6310 VN.n9681 VN.n9675 0.047
R6311 VN.n11414 VN.n11405 0.047
R6312 VN.n11397 VN.n11391 0.047
R6313 VN.n12115 VN.n12108 0.047
R6314 VN.n925 VN.n917 0.047
R6315 VN.n1163 VN.n1158 0.047
R6316 VN.n1526 VN.n1511 0.047
R6317 VN.n1853 VN.n1848 0.047
R6318 VN.n2234 VN.n2219 0.047
R6319 VN.n2562 VN.n2557 0.047
R6320 VN.n2956 VN.n2941 0.047
R6321 VN.n3284 VN.n3279 0.047
R6322 VN.n3696 VN.n3681 0.047
R6323 VN.n4028 VN.n4023 0.047
R6324 VN.n4453 VN.n4438 0.047
R6325 VN.n4785 VN.n4780 0.047
R6326 VN.n5228 VN.n5213 0.047
R6327 VN.n5564 VN.n5559 0.047
R6328 VN.n6020 VN.n6005 0.047
R6329 VN.n6356 VN.n6351 0.047
R6330 VN.n7263 VN.n7248 0.047
R6331 VN.n6801 VN.n6796 0.047
R6332 VN.n7652 VN.n7637 0.047
R6333 VN.n7992 VN.n7987 0.047
R6334 VN.n8497 VN.n8482 0.047
R6335 VN.n8841 VN.n8836 0.047
R6336 VN.n9359 VN.n9344 0.047
R6337 VN.n9703 VN.n9698 0.047
R6338 VN.n10242 VN.n10227 0.047
R6339 VN.n10588 VN.n10583 0.047
R6340 VN.n11441 VN.n11432 0.047
R6341 VN.n11138 VN.n11133 0.047
R6342 VN.n10609 VN.n10603 0.047
R6343 VN.n10263 VN.n10260 0.047
R6344 VN.n9722 VN.n9718 0.047
R6345 VN.n9380 VN.n9377 0.047
R6346 VN.n8860 VN.n8856 0.047
R6347 VN.n8518 VN.n8515 0.047
R6348 VN.n8011 VN.n8007 0.047
R6349 VN.n7673 VN.n7670 0.047
R6350 VN.n6820 VN.n6816 0.047
R6351 VN.n7284 VN.n7281 0.047
R6352 VN.n6375 VN.n6371 0.047
R6353 VN.n6041 VN.n6038 0.047
R6354 VN.n5583 VN.n5579 0.047
R6355 VN.n5249 VN.n5246 0.047
R6356 VN.n4804 VN.n4800 0.047
R6357 VN.n4474 VN.n4471 0.047
R6358 VN.n4047 VN.n4043 0.047
R6359 VN.n3717 VN.n3714 0.047
R6360 VN.n3303 VN.n3299 0.047
R6361 VN.n2977 VN.n2974 0.047
R6362 VN.n2581 VN.n2577 0.047
R6363 VN.n2255 VN.n2252 0.047
R6364 VN.n1872 VN.n1868 0.047
R6365 VN.n1550 VN.n1547 0.047
R6366 VN.n1182 VN.n1178 0.047
R6367 VN.n864 VN.n861 0.047
R6368 VN.n507 VN.n503 0.047
R6369 VN.n253 VN.n250 0.047
R6370 VN.n12144 VN.n12134 0.047
R6371 VN.n11036 VN.n11027 0.047
R6372 VN.n11172 VN.n11170 0.047
R6373 VN.n11991 VN.n11989 0.047
R6374 VN.n4536 VN.n4520 0.047
R6375 VN.n4695 VN.n4689 0.047
R6376 VN.n5069 VN.n5055 0.047
R6377 VN.n5474 VN.n5468 0.047
R6378 VN.n5861 VN.n5847 0.047
R6379 VN.n6266 VN.n6260 0.047
R6380 VN.n7104 VN.n7090 0.047
R6381 VN.n6711 VN.n6705 0.047
R6382 VN.n7493 VN.n7479 0.047
R6383 VN.n7902 VN.n7896 0.047
R6384 VN.n8338 VN.n8324 0.047
R6385 VN.n8751 VN.n8745 0.047
R6386 VN.n9200 VN.n9186 0.047
R6387 VN.n9613 VN.n9607 0.047
R6388 VN.n10082 VN.n10068 0.047
R6389 VN.n10490 VN.n10483 0.047
R6390 VN.n10951 VN.n10942 0.047
R6391 VN.n11222 VN.n11216 0.047
R6392 VN.n12014 VN.n12012 0.047
R6393 VN.n3782 VN.n3773 0.047
R6394 VN.n3955 VN.n3953 0.047
R6395 VN.n4323 VN.n4312 0.047
R6396 VN.n4712 VN.n4710 0.047
R6397 VN.n5098 VN.n5087 0.047
R6398 VN.n5491 VN.n5489 0.047
R6399 VN.n5890 VN.n5879 0.047
R6400 VN.n6283 VN.n6281 0.047
R6401 VN.n7133 VN.n7122 0.047
R6402 VN.n6728 VN.n6726 0.047
R6403 VN.n7522 VN.n7511 0.047
R6404 VN.n7919 VN.n7917 0.047
R6405 VN.n8367 VN.n8356 0.047
R6406 VN.n8768 VN.n8766 0.047
R6407 VN.n9229 VN.n9218 0.047
R6408 VN.n9630 VN.n9628 0.047
R6409 VN.n10111 VN.n10100 0.047
R6410 VN.n10507 VN.n10505 0.047
R6411 VN.n10980 VN.n10969 0.047
R6412 VN.n11206 VN.n11204 0.047
R6413 VN.n11946 VN.n11944 0.047
R6414 VN.n6103 VN.n6087 0.047
R6415 VN.n6232 VN.n6226 0.047
R6416 VN.n7041 VN.n7027 0.047
R6417 VN.n6677 VN.n6671 0.047
R6418 VN.n7430 VN.n7416 0.047
R6419 VN.n7868 VN.n7862 0.047
R6420 VN.n8275 VN.n8261 0.047
R6421 VN.n8717 VN.n8711 0.047
R6422 VN.n9137 VN.n9123 0.047
R6423 VN.n9579 VN.n9573 0.047
R6424 VN.n10019 VN.n10005 0.047
R6425 VN.n10455 VN.n10448 0.047
R6426 VN.n10893 VN.n10884 0.047
R6427 VN.n11256 VN.n11250 0.047
R6428 VN.n11969 VN.n11967 0.047
R6429 VN.n5314 VN.n5305 0.047
R6430 VN.n5457 VN.n5455 0.047
R6431 VN.n5827 VN.n5816 0.047
R6432 VN.n6249 VN.n6247 0.047
R6433 VN.n7070 VN.n7059 0.047
R6434 VN.n6694 VN.n6692 0.047
R6435 VN.n7459 VN.n7448 0.047
R6436 VN.n7885 VN.n7883 0.047
R6437 VN.n8304 VN.n8293 0.047
R6438 VN.n8734 VN.n8732 0.047
R6439 VN.n9166 VN.n9155 0.047
R6440 VN.n9596 VN.n9594 0.047
R6441 VN.n10048 VN.n10037 0.047
R6442 VN.n10472 VN.n10470 0.047
R6443 VN.n10922 VN.n10911 0.047
R6444 VN.n11240 VN.n11238 0.047
R6445 VN.n6660 VN.n6658 0.047
R6446 VN.n7396 VN.n7385 0.047
R6447 VN.n7851 VN.n7849 0.047
R6448 VN.n8241 VN.n8230 0.047
R6449 VN.n8700 VN.n8698 0.047
R6450 VN.n9103 VN.n9092 0.047
R6451 VN.n9562 VN.n9560 0.047
R6452 VN.n9985 VN.n9974 0.047
R6453 VN.n10437 VN.n10435 0.047
R6454 VN.n10864 VN.n10853 0.047
R6455 VN.n11273 VN.n11271 0.047
R6456 VN.n11924 VN.n11918 0.047
R6457 VN.n11897 VN.n11895 0.047
R6458 VN.n7735 VN.n7719 0.047
R6459 VN.n7834 VN.n7828 0.047
R6460 VN.n8212 VN.n8198 0.047
R6461 VN.n8683 VN.n8677 0.047
R6462 VN.n9074 VN.n9060 0.047
R6463 VN.n9545 VN.n9539 0.047
R6464 VN.n9956 VN.n9942 0.047
R6465 VN.n10420 VN.n10413 0.047
R6466 VN.n10835 VN.n10826 0.047
R6467 VN.n11289 VN.n11284 0.047
R6468 VN.n11639 VN.n11637 0.047
R6469 VN.n9442 VN.n9426 0.047
R6470 VN.n9511 VN.n9505 0.047
R6471 VN.n9893 VN.n9879 0.047
R6472 VN.n10385 VN.n10378 0.047
R6473 VN.n10777 VN.n10768 0.047
R6474 VN.n11323 VN.n11317 0.047
R6475 VN.n11876 VN.n11874 0.047
R6476 VN.n8583 VN.n8574 0.047
R6477 VN.n8666 VN.n8664 0.047
R6478 VN.n9040 VN.n9029 0.047
R6479 VN.n9528 VN.n9526 0.047
R6480 VN.n9922 VN.n9911 0.047
R6481 VN.n10402 VN.n10400 0.047
R6482 VN.n10806 VN.n10795 0.047
R6483 VN.n11307 VN.n11305 0.047
R6484 VN.n11594 VN.n11592 0.047
R6485 VN.n11489 VN.n11477 0.047
R6486 VN.n11357 VN.n11351 0.047
R6487 VN.n11617 VN.n11615 0.047
R6488 VN.n10328 VN.n10319 0.047
R6489 VN.n10367 VN.n10365 0.047
R6490 VN.n10748 VN.n10737 0.047
R6491 VN.n11341 VN.n11339 0.047
R6492 VN.n12182 VN.n11545 0.047
R6493 VN.n11100 VN.n11097 0.047
R6494 VN.n11506 VN.n11503 0.047
R6495 VN.n10662 VN.n10659 0.047
R6496 VN.n10676 VN.n10669 0.047
R6497 VN.n9757 VN.n9754 0.047
R6498 VN.n9462 VN.n9455 0.047
R6499 VN.n8895 VN.n8892 0.047
R6500 VN.n8603 VN.n8596 0.047
R6501 VN.n8046 VN.n8043 0.047
R6502 VN.n7755 VN.n7748 0.047
R6503 VN.n6855 VN.n6852 0.047
R6504 VN.n7007 VN.n7000 0.047
R6505 VN.n6410 VN.n6407 0.047
R6506 VN.n6123 VN.n6116 0.047
R6507 VN.n5618 VN.n5615 0.047
R6508 VN.n5334 VN.n5327 0.047
R6509 VN.n4839 VN.n4836 0.047
R6510 VN.n4556 VN.n4549 0.047
R6511 VN.n4082 VN.n4079 0.047
R6512 VN.n3802 VN.n3795 0.047
R6513 VN.n3338 VN.n3335 0.047
R6514 VN.n3059 VN.n3052 0.047
R6515 VN.n2616 VN.n2613 0.047
R6516 VN.n2340 VN.n2333 0.047
R6517 VN.n1907 VN.n1904 0.047
R6518 VN.n1632 VN.n1625 0.047
R6519 VN.n1217 VN.n1214 0.047
R6520 VN.n945 VN.n938 0.047
R6521 VN.n542 VN.n539 0.047
R6522 VN.n273 VN.n266 0.047
R6523 VN.n12299 VN.n12296 0.047
R6524 VN.n12314 VN.n12307 0.047
R6525 VN.n12282 VN.n12278 0.047
R6526 VN.n11524 VN.n11519 0.047
R6527 VN.n10644 VN.n10642 0.047
R6528 VN.n10691 VN.n10687 0.047
R6529 VN.n12630 VN.n12349 0.047
R6530 VN.n12632 VN.n12325 0.047
R6531 VN.n12343 VN.n12333 0.047
R6532 VN.n288 VN.n284 0.047
R6533 VN.n558 VN.n553 0.047
R6534 VN.n960 VN.n956 0.047
R6535 VN.n1233 VN.n1228 0.047
R6536 VN.n1647 VN.n1643 0.047
R6537 VN.n1923 VN.n1918 0.047
R6538 VN.n2355 VN.n2351 0.047
R6539 VN.n2632 VN.n2627 0.047
R6540 VN.n3074 VN.n3070 0.047
R6541 VN.n3354 VN.n3349 0.047
R6542 VN.n3817 VN.n3813 0.047
R6543 VN.n4098 VN.n4093 0.047
R6544 VN.n4571 VN.n4567 0.047
R6545 VN.n4855 VN.n4850 0.047
R6546 VN.n5349 VN.n5345 0.047
R6547 VN.n5634 VN.n5629 0.047
R6548 VN.n6138 VN.n6134 0.047
R6549 VN.n6426 VN.n6421 0.047
R6550 VN.n6987 VN.n6983 0.047
R6551 VN.n6871 VN.n6866 0.047
R6552 VN.n7770 VN.n7766 0.047
R6553 VN.n8062 VN.n8057 0.047
R6554 VN.n8618 VN.n8614 0.047
R6555 VN.n8911 VN.n8906 0.047
R6556 VN.n9796 VN.n9473 0.047
R6557 VN.n9795 VN.n9481 0.047
R6558 VN.n10707 VN.n9865 0.047
R6559 VN.n9779 VN.n9771 0.047
R6560 VN.n9811 VN.n9807 0.047
R6561 VN.n12422 VN.n12417 0.047
R6562 VN.n12663 VN.n12643 0.047
R6563 VN.n12661 VN.n12651 0.047
R6564 VN.n303 VN.n299 0.047
R6565 VN.n574 VN.n569 0.047
R6566 VN.n975 VN.n971 0.047
R6567 VN.n1249 VN.n1244 0.047
R6568 VN.n1662 VN.n1658 0.047
R6569 VN.n1939 VN.n1934 0.047
R6570 VN.n2370 VN.n2366 0.047
R6571 VN.n2648 VN.n2643 0.047
R6572 VN.n3089 VN.n3085 0.047
R6573 VN.n3370 VN.n3365 0.047
R6574 VN.n3832 VN.n3828 0.047
R6575 VN.n4114 VN.n4109 0.047
R6576 VN.n4586 VN.n4582 0.047
R6577 VN.n4871 VN.n4866 0.047
R6578 VN.n5364 VN.n5360 0.047
R6579 VN.n5650 VN.n5645 0.047
R6580 VN.n6153 VN.n6149 0.047
R6581 VN.n6442 VN.n6437 0.047
R6582 VN.n6972 VN.n6968 0.047
R6583 VN.n6887 VN.n6882 0.047
R6584 VN.n7785 VN.n7781 0.047
R6585 VN.n8078 VN.n8073 0.047
R6586 VN.n8950 VN.n8629 0.047
R6587 VN.n8949 VN.n8637 0.047
R6588 VN.n9827 VN.n9017 0.047
R6589 VN.n8933 VN.n8925 0.047
R6590 VN.n8965 VN.n8961 0.047
R6591 VN.n12438 VN.n12433 0.047
R6592 VN.n12774 VN.n12674 0.047
R6593 VN.n12772 VN.n12682 0.047
R6594 VN.n318 VN.n314 0.047
R6595 VN.n590 VN.n585 0.047
R6596 VN.n990 VN.n986 0.047
R6597 VN.n1265 VN.n1260 0.047
R6598 VN.n1677 VN.n1673 0.047
R6599 VN.n1955 VN.n1950 0.047
R6600 VN.n2385 VN.n2381 0.047
R6601 VN.n2664 VN.n2659 0.047
R6602 VN.n3104 VN.n3100 0.047
R6603 VN.n3386 VN.n3381 0.047
R6604 VN.n3847 VN.n3843 0.047
R6605 VN.n4130 VN.n4125 0.047
R6606 VN.n4601 VN.n4597 0.047
R6607 VN.n4887 VN.n4882 0.047
R6608 VN.n5379 VN.n5375 0.047
R6609 VN.n5666 VN.n5661 0.047
R6610 VN.n6168 VN.n6164 0.047
R6611 VN.n6458 VN.n6453 0.047
R6612 VN.n6957 VN.n6953 0.047
R6613 VN.n6903 VN.n6898 0.047
R6614 VN.n8117 VN.n7796 0.047
R6615 VN.n8116 VN.n7804 0.047
R6616 VN.n8981 VN.n8184 0.047
R6617 VN.n8100 VN.n8092 0.047
R6618 VN.n8132 VN.n8128 0.047
R6619 VN.n12454 VN.n12449 0.047
R6620 VN.n12808 VN.n12785 0.047
R6621 VN.n12806 VN.n12796 0.047
R6622 VN.n333 VN.n329 0.047
R6623 VN.n606 VN.n601 0.047
R6624 VN.n1005 VN.n1001 0.047
R6625 VN.n1281 VN.n1276 0.047
R6626 VN.n1692 VN.n1688 0.047
R6627 VN.n1971 VN.n1966 0.047
R6628 VN.n2400 VN.n2396 0.047
R6629 VN.n2680 VN.n2675 0.047
R6630 VN.n3119 VN.n3115 0.047
R6631 VN.n3402 VN.n3397 0.047
R6632 VN.n3862 VN.n3858 0.047
R6633 VN.n4146 VN.n4141 0.047
R6634 VN.n4616 VN.n4612 0.047
R6635 VN.n4903 VN.n4898 0.047
R6636 VN.n5394 VN.n5390 0.047
R6637 VN.n5682 VN.n5677 0.047
R6638 VN.n6183 VN.n6179 0.047
R6639 VN.n6474 VN.n6469 0.047
R6640 VN.n6942 VN.n6623 0.047
R6641 VN.n6941 VN.n6631 0.047
R6642 VN.n8148 VN.n7373 0.047
R6643 VN.n6925 VN.n6917 0.047
R6644 VN.n6612 VN.n6608 0.047
R6645 VN.n12470 VN.n12465 0.047
R6646 VN.n12839 VN.n12816 0.047
R6647 VN.n12837 VN.n12827 0.047
R6648 VN.n348 VN.n344 0.047
R6649 VN.n622 VN.n617 0.047
R6650 VN.n1020 VN.n1016 0.047
R6651 VN.n1297 VN.n1292 0.047
R6652 VN.n1707 VN.n1703 0.047
R6653 VN.n1987 VN.n1982 0.047
R6654 VN.n2415 VN.n2411 0.047
R6655 VN.n2696 VN.n2691 0.047
R6656 VN.n3134 VN.n3130 0.047
R6657 VN.n3418 VN.n3413 0.047
R6658 VN.n3877 VN.n3873 0.047
R6659 VN.n4162 VN.n4157 0.047
R6660 VN.n4631 VN.n4627 0.047
R6661 VN.n4919 VN.n4914 0.047
R6662 VN.n5409 VN.n5405 0.047
R6663 VN.n5698 VN.n5693 0.047
R6664 VN.n6513 VN.n6194 0.047
R6665 VN.n6512 VN.n6202 0.047
R6666 VN.n7337 VN.n6580 0.047
R6667 VN.n6496 VN.n6488 0.047
R6668 VN.n6528 VN.n6524 0.047
R6669 VN.n12486 VN.n12481 0.047
R6670 VN.n12867 VN.n12847 0.047
R6671 VN.n12865 VN.n12855 0.047
R6672 VN.n363 VN.n359 0.047
R6673 VN.n638 VN.n633 0.047
R6674 VN.n1035 VN.n1031 0.047
R6675 VN.n1313 VN.n1308 0.047
R6676 VN.n1722 VN.n1718 0.047
R6677 VN.n2003 VN.n1998 0.047
R6678 VN.n2430 VN.n2426 0.047
R6679 VN.n2712 VN.n2707 0.047
R6680 VN.n3149 VN.n3145 0.047
R6681 VN.n3434 VN.n3429 0.047
R6682 VN.n3892 VN.n3888 0.047
R6683 VN.n4178 VN.n4173 0.047
R6684 VN.n4646 VN.n4642 0.047
R6685 VN.n4935 VN.n4930 0.047
R6686 VN.n5737 VN.n5420 0.047
R6687 VN.n5736 VN.n5428 0.047
R6688 VN.n6544 VN.n5804 0.047
R6689 VN.n5720 VN.n5712 0.047
R6690 VN.n5752 VN.n5748 0.047
R6691 VN.n12502 VN.n12497 0.047
R6692 VN.n12898 VN.n12878 0.047
R6693 VN.n12896 VN.n12886 0.047
R6694 VN.n378 VN.n374 0.047
R6695 VN.n654 VN.n649 0.047
R6696 VN.n1050 VN.n1046 0.047
R6697 VN.n1329 VN.n1324 0.047
R6698 VN.n1737 VN.n1733 0.047
R6699 VN.n2019 VN.n2014 0.047
R6700 VN.n2445 VN.n2441 0.047
R6701 VN.n2728 VN.n2723 0.047
R6702 VN.n3164 VN.n3160 0.047
R6703 VN.n3450 VN.n3445 0.047
R6704 VN.n3907 VN.n3903 0.047
R6705 VN.n4194 VN.n4189 0.047
R6706 VN.n4974 VN.n4657 0.047
R6707 VN.n4973 VN.n4665 0.047
R6708 VN.n5768 VN.n5041 0.047
R6709 VN.n4957 VN.n4949 0.047
R6710 VN.n4989 VN.n4985 0.047
R6711 VN.n12518 VN.n12513 0.047
R6712 VN.n12929 VN.n12909 0.047
R6713 VN.n12927 VN.n12917 0.047
R6714 VN.n393 VN.n389 0.047
R6715 VN.n670 VN.n665 0.047
R6716 VN.n1065 VN.n1061 0.047
R6717 VN.n1345 VN.n1340 0.047
R6718 VN.n1752 VN.n1748 0.047
R6719 VN.n2035 VN.n2030 0.047
R6720 VN.n2460 VN.n2456 0.047
R6721 VN.n2744 VN.n2739 0.047
R6722 VN.n3179 VN.n3175 0.047
R6723 VN.n3466 VN.n3461 0.047
R6724 VN.n4233 VN.n3918 0.047
R6725 VN.n4232 VN.n3926 0.047
R6726 VN.n5005 VN.n4300 0.047
R6727 VN.n4216 VN.n4208 0.047
R6728 VN.n4248 VN.n4244 0.047
R6729 VN.n12534 VN.n12529 0.047
R6730 VN.n12960 VN.n12940 0.047
R6731 VN.n12958 VN.n12948 0.047
R6732 VN.n408 VN.n404 0.047
R6733 VN.n686 VN.n681 0.047
R6734 VN.n1080 VN.n1076 0.047
R6735 VN.n1361 VN.n1356 0.047
R6736 VN.n1767 VN.n1763 0.047
R6737 VN.n2051 VN.n2046 0.047
R6738 VN.n2475 VN.n2471 0.047
R6739 VN.n2760 VN.n2755 0.047
R6740 VN.n3505 VN.n3190 0.047
R6741 VN.n3504 VN.n3198 0.047
R6742 VN.n4264 VN.n3572 0.047
R6743 VN.n3488 VN.n3480 0.047
R6744 VN.n3520 VN.n3516 0.047
R6745 VN.n12550 VN.n12545 0.047
R6746 VN.n12991 VN.n12971 0.047
R6747 VN.n12989 VN.n12979 0.047
R6748 VN.n423 VN.n419 0.047
R6749 VN.n702 VN.n697 0.047
R6750 VN.n1095 VN.n1091 0.047
R6751 VN.n1377 VN.n1372 0.047
R6752 VN.n1782 VN.n1778 0.047
R6753 VN.n2067 VN.n2062 0.047
R6754 VN.n2799 VN.n2486 0.047
R6755 VN.n2798 VN.n2494 0.047
R6756 VN.n3536 VN.n2866 0.047
R6757 VN.n2782 VN.n2774 0.047
R6758 VN.n2814 VN.n2810 0.047
R6759 VN.n12566 VN.n12561 0.047
R6760 VN.n13022 VN.n13002 0.047
R6761 VN.n13020 VN.n13010 0.047
R6762 VN.n438 VN.n434 0.047
R6763 VN.n718 VN.n713 0.047
R6764 VN.n1110 VN.n1106 0.047
R6765 VN.n1393 VN.n1388 0.047
R6766 VN.n2106 VN.n1793 0.047
R6767 VN.n2105 VN.n1801 0.047
R6768 VN.n2830 VN.n2173 0.047
R6769 VN.n2089 VN.n2081 0.047
R6770 VN.n2121 VN.n2117 0.047
R6771 VN.n12582 VN.n12577 0.047
R6772 VN.n13053 VN.n13033 0.047
R6773 VN.n13051 VN.n13041 0.047
R6774 VN.n453 VN.n449 0.047
R6775 VN.n734 VN.n729 0.047
R6776 VN.n1432 VN.n1121 0.047
R6777 VN.n1431 VN.n1129 0.047
R6778 VN.n2137 VN.n1499 0.047
R6779 VN.n1415 VN.n1407 0.047
R6780 VN.n1447 VN.n1443 0.047
R6781 VN.n12598 VN.n12593 0.047
R6782 VN.n13084 VN.n13064 0.047
R6783 VN.n13082 VN.n13072 0.047
R6784 VN.n772 VN.n464 0.047
R6785 VN.n771 VN.n472 0.047
R6786 VN.n1463 VN.n849 0.047
R6787 VN.n755 VN.n746 0.047
R6788 VN.n794 VN.n791 0.047
R6789 VN.n12614 VN.n12612 0.047
R6790 VN.n13104 VN.n13102 0.047
R6791 VN.n12756 VN.n12754 0.047
R6792 VN.n821 VN.n199 0.047
R6793 VN.n12385 VN.n12383 0.047
R6794 VN.n12233 VN.n12231 0.047
R6795 VN.n12737 VN.n12728 0.047
R6796 VN.n12405 VN.n12401 0.047
R6797 VN.n11067 VN.n11062 0.047
R6798 VN.n2183 VN.n2182 0.047
R6799 VN.n2905 VN.n2904 0.047
R6800 VN.n3645 VN.n3644 0.047
R6801 VN.n4402 VN.n4401 0.047
R6802 VN.n5177 VN.n5176 0.047
R6803 VN.n5969 VN.n5968 0.047
R6804 VN.n7212 VN.n7211 0.047
R6805 VN.n7601 VN.n7600 0.047
R6806 VN.n8446 VN.n8445 0.047
R6807 VN.n9308 VN.n9307 0.047
R6808 VN.n10191 VN.n10190 0.047
R6809 VN.n10676 VN.n10662 0.046
R6810 VN.n9796 VN.n9795 0.046
R6811 VN.n8950 VN.n8949 0.045
R6812 VN.n8117 VN.n8116 0.045
R6813 VN.n6942 VN.n6941 0.045
R6814 VN.n6513 VN.n6512 0.045
R6815 VN.n5737 VN.n5736 0.045
R6816 VN.n4974 VN.n4973 0.045
R6817 VN.n4233 VN.n4232 0.045
R6818 VN.n3505 VN.n3504 0.045
R6819 VN.n2799 VN.n2798 0.045
R6820 VN.n2106 VN.n2105 0.045
R6821 VN.n1432 VN.n1431 0.045
R6822 VN.n772 VN.n771 0.045
R6823 VN.n11701 VN.n11700 0.045
R6824 VN.n793 VN.n792 0.045
R6825 VN.n12099 VN.n12098 0.045
R6826 VN.n11084 VN.n11076 0.045
R6827 VN.n10239 VN.n10231 0.045
R6828 VN.n9356 VN.n9348 0.045
R6829 VN.n8494 VN.n8486 0.045
R6830 VN.n7649 VN.n7641 0.045
R6831 VN.n7260 VN.n7252 0.045
R6832 VN.n6017 VN.n6009 0.045
R6833 VN.n5225 VN.n5217 0.045
R6834 VN.n4450 VN.n4442 0.045
R6835 VN.n3693 VN.n3685 0.045
R6836 VN.n2953 VN.n2945 0.045
R6837 VN.n2231 VN.n2223 0.045
R6838 VN.n1523 VN.n1515 0.045
R6839 VN.n9831 VN.n9830 0.045
R6840 VN.n8985 VN.n8984 0.045
R6841 VN.n8152 VN.n8151 0.045
R6842 VN.n7341 VN.n7340 0.045
R6843 VN.n6548 VN.n6547 0.045
R6844 VN.n5772 VN.n5771 0.045
R6845 VN.n5009 VN.n5008 0.045
R6846 VN.n4268 VN.n4267 0.045
R6847 VN.n3540 VN.n3539 0.045
R6848 VN.n2834 VN.n2833 0.045
R6849 VN.n2141 VN.n2140 0.045
R6850 VN.n1467 VN.n1466 0.045
R6851 VN.n20 VN.n19 0.045
R6852 VN.n87 VN.n86 0.045
R6853 VN.n12314 VN.n12283 0.044
R6854 VN.n12632 VN.n12631 0.044
R6855 VN.n18 VN.n17 0.044
R6856 VN.n83 VN.n81 0.044
R6857 VN.n11909 VN.n11908 0.044
R6858 VN.n12048 VN.n12047 0.044
R6859 VN.n12003 VN.n12002 0.044
R6860 VN.n11958 VN.n11957 0.044
R6861 VN.n11651 VN.n11650 0.044
R6862 VN.n11606 VN.n11605 0.044
R6863 VN.n12023 VN.n12022 0.044
R6864 VN.n11978 VN.n11977 0.044
R6865 VN.n11933 VN.n11932 0.044
R6866 VN.n11885 VN.n11884 0.044
R6867 VN.n11626 VN.n11625 0.044
R6868 VN.n11581 VN.n11580 0.044
R6869 VN.n100 VN.n99 0.043
R6870 VN.n12258 VN.n12257 0.043
R6871 VN.n12078 VN.n12077 0.043
R6872 VN.n239 VN.n238 0.043
R6873 VN.n11561 VN.n11560 0.043
R6874 VN.n11046 VN.n11045 0.043
R6875 VN.n11912 VN.n11911 0.043
R6876 VN.n12123 VN.n12122 0.043
R6877 VN.n11020 VN.n11019 0.042
R6878 VN.n10155 VN.n10154 0.042
R6879 VN.n9273 VN.n9272 0.042
R6880 VN.n8411 VN.n8410 0.042
R6881 VN.n7566 VN.n7565 0.042
R6882 VN.n7177 VN.n7176 0.042
R6883 VN.n5934 VN.n5933 0.042
R6884 VN.n5142 VN.n5141 0.042
R6885 VN.n4367 VN.n4366 0.042
R6886 VN.n3610 VN.n3609 0.042
R6887 VN.n2870 VN.n2869 0.042
R6888 VN.n10962 VN.n10961 0.042
R6889 VN.n10092 VN.n10091 0.042
R6890 VN.n9210 VN.n9209 0.042
R6891 VN.n8348 VN.n8347 0.042
R6892 VN.n7503 VN.n7502 0.042
R6893 VN.n7114 VN.n7113 0.042
R6894 VN.n5871 VN.n5870 0.042
R6895 VN.n5079 VN.n5078 0.042
R6896 VN.n4304 VN.n4303 0.042
R6897 VN.n10904 VN.n10903 0.042
R6898 VN.n10029 VN.n10028 0.042
R6899 VN.n9147 VN.n9146 0.042
R6900 VN.n8285 VN.n8284 0.042
R6901 VN.n7440 VN.n7439 0.042
R6902 VN.n7051 VN.n7050 0.042
R6903 VN.n5808 VN.n5807 0.042
R6904 VN.n10788 VN.n10787 0.042
R6905 VN.n9903 VN.n9902 0.042
R6906 VN.n9021 VN.n9020 0.042
R6907 VN.n10730 VN.n10729 0.042
R6908 VN.n11005 VN.n11004 0.042
R6909 VN.n10947 VN.n10946 0.042
R6910 VN.n10889 VN.n10888 0.042
R6911 VN.n10831 VN.n10830 0.042
R6912 VN.n10773 VN.n10772 0.042
R6913 VN.n11563 VN.n11562 0.042
R6914 VN.n223 VN.n218 0.042
R6915 VN.n894 VN.n889 0.042
R6916 VN.n1577 VN.n1572 0.042
R6917 VN.n2285 VN.n2280 0.042
R6918 VN.n3007 VN.n3002 0.042
R6919 VN.n3747 VN.n3742 0.042
R6920 VN.n4504 VN.n4499 0.042
R6921 VN.n5279 VN.n5274 0.042
R6922 VN.n6071 VN.n6066 0.042
R6923 VN.n7314 VN.n7309 0.042
R6924 VN.n7703 VN.n7698 0.042
R6925 VN.n8548 VN.n8543 0.042
R6926 VN.n9410 VN.n9405 0.042
R6927 VN.n10293 VN.n10288 0.042
R6928 VN.n11461 VN.n11456 0.042
R6929 VN.n3596 VN.n3591 0.042
R6930 VN.n4353 VN.n4348 0.042
R6931 VN.n5128 VN.n5123 0.042
R6932 VN.n5920 VN.n5915 0.042
R6933 VN.n7163 VN.n7158 0.042
R6934 VN.n7552 VN.n7547 0.042
R6935 VN.n8397 VN.n8392 0.042
R6936 VN.n9259 VN.n9254 0.042
R6937 VN.n10141 VN.n10136 0.042
R6938 VN.n2197 VN.n2192 0.042
R6939 VN.n2919 VN.n2914 0.042
R6940 VN.n3659 VN.n3654 0.042
R6941 VN.n4416 VN.n4411 0.042
R6942 VN.n5191 VN.n5186 0.042
R6943 VN.n5983 VN.n5978 0.042
R6944 VN.n7226 VN.n7221 0.042
R6945 VN.n7615 VN.n7610 0.042
R6946 VN.n8460 VN.n8455 0.042
R6947 VN.n9322 VN.n9317 0.042
R6948 VN.n10205 VN.n10200 0.042
R6949 VN.n5065 VN.n5060 0.042
R6950 VN.n5857 VN.n5852 0.042
R6951 VN.n7100 VN.n7095 0.042
R6952 VN.n7489 VN.n7484 0.042
R6953 VN.n8334 VN.n8329 0.042
R6954 VN.n9196 VN.n9191 0.042
R6955 VN.n10078 VN.n10073 0.042
R6956 VN.n7037 VN.n7032 0.042
R6957 VN.n7426 VN.n7421 0.042
R6958 VN.n8271 VN.n8266 0.042
R6959 VN.n9133 VN.n9128 0.042
R6960 VN.n10015 VN.n10010 0.042
R6961 VN.n8208 VN.n8203 0.042
R6962 VN.n9070 VN.n9065 0.042
R6963 VN.n9952 VN.n9947 0.042
R6964 VN.n9889 VN.n9884 0.042
R6965 VN.n12051 VN.n12050 0.042
R6966 VN.n12102 VN.n12101 0.042
R6967 VN.n12006 VN.n12005 0.042
R6968 VN.n11961 VN.n11960 0.042
R6969 VN.n11868 VN.n11867 0.042
R6970 VN.n11609 VN.n11608 0.042
R6971 VN.n7377 VN.n7376 0.042
R6972 VN.n8222 VN.n8221 0.042
R6973 VN.n9084 VN.n9083 0.042
R6974 VN.n9966 VN.n9965 0.042
R6975 VN.n10845 VN.n10844 0.042
R6976 VN.n853 VN.n852 0.042
R6977 VN.n1539 VN.n1538 0.042
R6978 VN.n2244 VN.n2243 0.042
R6979 VN.n2966 VN.n2965 0.042
R6980 VN.n3706 VN.n3705 0.042
R6981 VN.n4463 VN.n4462 0.042
R6982 VN.n5238 VN.n5237 0.042
R6983 VN.n6030 VN.n6029 0.042
R6984 VN.n7273 VN.n7272 0.042
R6985 VN.n7662 VN.n7661 0.042
R6986 VN.n8507 VN.n8506 0.042
R6987 VN.n9369 VN.n9368 0.042
R6988 VN.n10252 VN.n10251 0.042
R6989 VN.n11424 VN.n11423 0.042
R6990 VN.n12127 VN.n12126 0.041
R6991 VN.n1593 VN.n1592 0.041
R6992 VN.n11788 VN.n11782 0.041
R6993 VN.n12179 VN.n12178 0.041
R6994 VN.n11374 VN.n11368 0.04
R6995 VN.n10347 VN.n10341 0.04
R6996 VN.n9492 VN.n9486 0.04
R6997 VN.n8646 VN.n8640 0.04
R6998 VN.n7815 VN.n7809 0.04
R6999 VN.n6640 VN.n6634 0.04
R7000 VN.n6211 VN.n6205 0.04
R7001 VN.n5437 VN.n5431 0.04
R7002 VN.n4676 VN.n4670 0.04
R7003 VN.n3935 VN.n3929 0.04
R7004 VN.n3209 VN.n3203 0.04
R7005 VN.n2503 VN.n2497 0.04
R7006 VN.n1812 VN.n1806 0.04
R7007 VN.n1138 VN.n1132 0.04
R7008 VN.n486 VN.n480 0.04
R7009 VN.n12693 VN.n12687 0.04
R7010 VN.n11781 VN.n11780 0.039
R7011 VN.n9832 VN.n9831 0.039
R7012 VN.n9837 VN.n9836 0.039
R7013 VN.n8986 VN.n8985 0.039
R7014 VN.n8991 VN.n8990 0.039
R7015 VN.n8153 VN.n8152 0.039
R7016 VN.n8158 VN.n8157 0.039
R7017 VN.n7342 VN.n7341 0.039
R7018 VN.n7347 VN.n7346 0.039
R7019 VN.n6549 VN.n6548 0.039
R7020 VN.n6554 VN.n6553 0.039
R7021 VN.n5773 VN.n5772 0.039
R7022 VN.n5778 VN.n5777 0.039
R7023 VN.n5010 VN.n5009 0.039
R7024 VN.n5015 VN.n5014 0.039
R7025 VN.n4269 VN.n4268 0.039
R7026 VN.n4274 VN.n4273 0.039
R7027 VN.n3541 VN.n3540 0.039
R7028 VN.n3546 VN.n3545 0.039
R7029 VN.n2835 VN.n2834 0.039
R7030 VN.n2840 VN.n2839 0.039
R7031 VN.n2142 VN.n2141 0.039
R7032 VN.n2147 VN.n2146 0.039
R7033 VN.n1468 VN.n1467 0.039
R7034 VN.n1473 VN.n1472 0.039
R7035 VN.n190 VN.n189 0.039
R7036 VN.n16 VN.n2 0.039
R7037 VN.n6 VN.n5 0.039
R7038 VN.n11373 VN.n11369 0.039
R7039 VN.n10346 VN.n10342 0.039
R7040 VN.n9491 VN.n9487 0.039
R7041 VN.n8645 VN.n8641 0.039
R7042 VN.n7814 VN.n7810 0.039
R7043 VN.n6639 VN.n6635 0.039
R7044 VN.n6210 VN.n6206 0.039
R7045 VN.n5436 VN.n5432 0.039
R7046 VN.n4675 VN.n4671 0.039
R7047 VN.n3934 VN.n3930 0.039
R7048 VN.n3208 VN.n3204 0.039
R7049 VN.n2502 VN.n2498 0.039
R7050 VN.n1811 VN.n1807 0.039
R7051 VN.n1137 VN.n1133 0.039
R7052 VN.n485 VN.n481 0.039
R7053 VN.n12692 VN.n12688 0.039
R7054 VN.n12362 VN.n12355 0.039
R7055 VN.n12354 VN.n12352 0.038
R7056 VN.n12686 VN.n12684 0.038
R7057 VN.n209 VN.n208 0.038
R7058 VN.n880 VN.n879 0.038
R7059 VN.n1563 VN.n1562 0.038
R7060 VN.n2271 VN.n2270 0.038
R7061 VN.n2993 VN.n2992 0.038
R7062 VN.n3733 VN.n3732 0.038
R7063 VN.n4490 VN.n4489 0.038
R7064 VN.n5265 VN.n5264 0.038
R7065 VN.n6057 VN.n6056 0.038
R7066 VN.n7300 VN.n7299 0.038
R7067 VN.n7689 VN.n7688 0.038
R7068 VN.n8534 VN.n8533 0.038
R7069 VN.n9396 VN.n9395 0.038
R7070 VN.n10279 VN.n10278 0.038
R7071 VN.n3582 VN.n3581 0.038
R7072 VN.n4339 VN.n4338 0.038
R7073 VN.n5114 VN.n5113 0.038
R7074 VN.n5906 VN.n5905 0.038
R7075 VN.n7149 VN.n7148 0.038
R7076 VN.n7538 VN.n7537 0.038
R7077 VN.n8383 VN.n8382 0.038
R7078 VN.n9245 VN.n9244 0.038
R7079 VN.n10127 VN.n10126 0.038
R7080 VN.n10996 VN.n10995 0.038
R7081 VN.n2887 VN.n2882 0.038
R7082 VN.n3627 VN.n3622 0.038
R7083 VN.n4384 VN.n4379 0.038
R7084 VN.n5159 VN.n5154 0.038
R7085 VN.n5951 VN.n5946 0.038
R7086 VN.n7194 VN.n7189 0.038
R7087 VN.n7583 VN.n7578 0.038
R7088 VN.n8428 VN.n8423 0.038
R7089 VN.n9290 VN.n9285 0.038
R7090 VN.n10172 VN.n10167 0.038
R7091 VN.n11034 VN.n11031 0.038
R7092 VN.n5051 VN.n5050 0.038
R7093 VN.n5843 VN.n5842 0.038
R7094 VN.n7086 VN.n7085 0.038
R7095 VN.n7475 VN.n7474 0.038
R7096 VN.n8320 VN.n8319 0.038
R7097 VN.n9182 VN.n9181 0.038
R7098 VN.n10064 VN.n10063 0.038
R7099 VN.n10938 VN.n10937 0.038
R7100 VN.n4321 VN.n4316 0.038
R7101 VN.n5096 VN.n5091 0.038
R7102 VN.n5888 VN.n5883 0.038
R7103 VN.n7131 VN.n7126 0.038
R7104 VN.n7520 VN.n7515 0.038
R7105 VN.n8365 VN.n8360 0.038
R7106 VN.n9227 VN.n9222 0.038
R7107 VN.n10109 VN.n10104 0.038
R7108 VN.n10978 VN.n10973 0.038
R7109 VN.n7023 VN.n7022 0.038
R7110 VN.n7412 VN.n7411 0.038
R7111 VN.n8257 VN.n8256 0.038
R7112 VN.n9119 VN.n9118 0.038
R7113 VN.n10001 VN.n10000 0.038
R7114 VN.n10880 VN.n10879 0.038
R7115 VN.n5825 VN.n5820 0.038
R7116 VN.n7068 VN.n7063 0.038
R7117 VN.n7457 VN.n7452 0.038
R7118 VN.n8302 VN.n8297 0.038
R7119 VN.n9164 VN.n9159 0.038
R7120 VN.n10046 VN.n10041 0.038
R7121 VN.n10920 VN.n10915 0.038
R7122 VN.n7394 VN.n7389 0.038
R7123 VN.n8239 VN.n8234 0.038
R7124 VN.n9101 VN.n9096 0.038
R7125 VN.n9983 VN.n9978 0.038
R7126 VN.n10862 VN.n10857 0.038
R7127 VN.n8194 VN.n8193 0.038
R7128 VN.n9056 VN.n9055 0.038
R7129 VN.n9938 VN.n9937 0.038
R7130 VN.n10822 VN.n10821 0.038
R7131 VN.n9875 VN.n9874 0.038
R7132 VN.n10764 VN.n10763 0.038
R7133 VN.n9038 VN.n9033 0.038
R7134 VN.n9920 VN.n9915 0.038
R7135 VN.n10804 VN.n10799 0.038
R7136 VN.n10746 VN.n10741 0.038
R7137 VN.n12200 VN.n12199 0.038
R7138 VN.n12076 VN.n12075 0.038
R7139 VN.n924 VN.n922 0.037
R7140 VN.n10242 VN.n10224 0.037
R7141 VN.n9359 VN.n9341 0.037
R7142 VN.n8497 VN.n8479 0.037
R7143 VN.n7652 VN.n7634 0.037
R7144 VN.n7263 VN.n7245 0.037
R7145 VN.n6020 VN.n6002 0.037
R7146 VN.n5228 VN.n5210 0.037
R7147 VN.n4453 VN.n4435 0.037
R7148 VN.n3696 VN.n3678 0.037
R7149 VN.n2956 VN.n2938 0.037
R7150 VN.n2234 VN.n2216 0.037
R7151 VN.n1526 VN.n1508 0.037
R7152 VN.n925 VN.n914 0.037
R7153 VN.n11441 VN.n11433 0.037
R7154 VN.n11414 VN.n11406 0.037
R7155 VN.n9837 VN.n9834 0.037
R7156 VN.n9836 VN.n9835 0.037
R7157 VN.n8991 VN.n8988 0.037
R7158 VN.n8990 VN.n8989 0.037
R7159 VN.n8158 VN.n8155 0.037
R7160 VN.n8157 VN.n8156 0.037
R7161 VN.n7347 VN.n7344 0.037
R7162 VN.n7346 VN.n7345 0.037
R7163 VN.n6554 VN.n6551 0.037
R7164 VN.n6553 VN.n6552 0.037
R7165 VN.n5778 VN.n5775 0.037
R7166 VN.n5777 VN.n5776 0.037
R7167 VN.n5015 VN.n5012 0.037
R7168 VN.n5014 VN.n5013 0.037
R7169 VN.n4274 VN.n4271 0.037
R7170 VN.n4273 VN.n4272 0.037
R7171 VN.n3546 VN.n3543 0.037
R7172 VN.n3545 VN.n3544 0.037
R7173 VN.n2840 VN.n2837 0.037
R7174 VN.n2839 VN.n2838 0.037
R7175 VN.n2147 VN.n2144 0.037
R7176 VN.n2146 VN.n2145 0.037
R7177 VN.n1473 VN.n1470 0.037
R7178 VN.n1472 VN.n1471 0.037
R7179 VN.n190 VN.n187 0.037
R7180 VN.n189 VN.n188 0.037
R7181 VN.n13095 VN.n13094 0.037
R7182 VN.n784 VN.n783 0.037
R7183 VN.n11378 VN.n11377 0.036
R7184 VN.n12182 VN.n12179 0.036
R7185 VN.n11126 VN.n11125 0.036
R7186 VN.n10608 VN.n10607 0.036
R7187 VN.n9711 VN.n9710 0.036
R7188 VN.n8849 VN.n8848 0.036
R7189 VN.n8000 VN.n7999 0.036
R7190 VN.n6809 VN.n6808 0.036
R7191 VN.n6364 VN.n6363 0.036
R7192 VN.n5572 VN.n5571 0.036
R7193 VN.n4793 VN.n4792 0.036
R7194 VN.n4036 VN.n4035 0.036
R7195 VN.n3292 VN.n3291 0.036
R7196 VN.n2570 VN.n2569 0.036
R7197 VN.n1861 VN.n1860 0.036
R7198 VN.n1171 VN.n1170 0.036
R7199 VN.n496 VN.n495 0.036
R7200 VN.n11163 VN.n11161 0.036
R7201 VN.n11197 VN.n11195 0.036
R7202 VN.n11231 VN.n11229 0.036
R7203 VN.n11298 VN.n11296 0.036
R7204 VN.n11332 VN.n11330 0.036
R7205 VN.n11264 VN.n11263 0.036
R7206 VN.n10428 VN.n10427 0.036
R7207 VN.n9553 VN.n9552 0.036
R7208 VN.n8691 VN.n8690 0.036
R7209 VN.n7842 VN.n7841 0.036
R7210 VN.n6651 VN.n6650 0.036
R7211 VN.n2514 VN.n2513 0.035
R7212 VN.n3236 VN.n3235 0.035
R7213 VN.n3980 VN.n3979 0.035
R7214 VN.n4737 VN.n4736 0.035
R7215 VN.n5516 VN.n5515 0.035
R7216 VN.n6308 VN.n6307 0.035
R7217 VN.n6753 VN.n6752 0.035
R7218 VN.n7944 VN.n7943 0.035
R7219 VN.n8793 VN.n8792 0.035
R7220 VN.n9655 VN.n9654 0.035
R7221 VN.n10533 VN.n10532 0.035
R7222 VN.n3946 VN.n3945 0.035
R7223 VN.n4703 VN.n4702 0.035
R7224 VN.n5482 VN.n5481 0.035
R7225 VN.n6274 VN.n6273 0.035
R7226 VN.n6719 VN.n6718 0.035
R7227 VN.n7910 VN.n7909 0.035
R7228 VN.n8759 VN.n8758 0.035
R7229 VN.n9621 VN.n9620 0.035
R7230 VN.n10498 VN.n10497 0.035
R7231 VN.n5448 VN.n5447 0.035
R7232 VN.n6240 VN.n6239 0.035
R7233 VN.n6685 VN.n6684 0.035
R7234 VN.n7876 VN.n7875 0.035
R7235 VN.n8725 VN.n8724 0.035
R7236 VN.n9587 VN.n9586 0.035
R7237 VN.n10463 VN.n10462 0.035
R7238 VN.n8657 VN.n8656 0.035
R7239 VN.n9519 VN.n9518 0.035
R7240 VN.n10393 VN.n10392 0.035
R7241 VN.n10358 VN.n10357 0.035
R7242 VN.n12224 VN.n12223 0.035
R7243 VN.n11365 VN.n11364 0.035
R7244 VN.n12371 VN.n12370 0.035
R7245 VN.n2512 VN.n2511 0.035
R7246 VN.n1820 VN.n1819 0.035
R7247 VN.n1147 VN.n1146 0.035
R7248 VN.n494 VN.n493 0.035
R7249 VN.n12702 VN.n12701 0.035
R7250 VN.n3944 VN.n3943 0.035
R7251 VN.n3217 VN.n3216 0.035
R7252 VN.n5446 VN.n5445 0.035
R7253 VN.n4684 VN.n4683 0.035
R7254 VN.n6221 VN.n6220 0.035
R7255 VN.n6649 VN.n6648 0.035
R7256 VN.n8655 VN.n8654 0.035
R7257 VN.n7823 VN.n7822 0.035
R7258 VN.n10356 VN.n10355 0.035
R7259 VN.n9500 VN.n9499 0.035
R7260 VN.n209 VN.n204 0.035
R7261 VN.n880 VN.n875 0.035
R7262 VN.n1563 VN.n1558 0.035
R7263 VN.n2271 VN.n2266 0.035
R7264 VN.n2993 VN.n2988 0.035
R7265 VN.n3733 VN.n3728 0.035
R7266 VN.n4490 VN.n4485 0.035
R7267 VN.n5265 VN.n5260 0.035
R7268 VN.n6057 VN.n6052 0.035
R7269 VN.n7300 VN.n7295 0.035
R7270 VN.n7689 VN.n7684 0.035
R7271 VN.n8534 VN.n8529 0.035
R7272 VN.n9396 VN.n9391 0.035
R7273 VN.n10279 VN.n10274 0.035
R7274 VN.n3582 VN.n3577 0.035
R7275 VN.n4339 VN.n4334 0.035
R7276 VN.n5114 VN.n5109 0.035
R7277 VN.n5906 VN.n5901 0.035
R7278 VN.n7149 VN.n7144 0.035
R7279 VN.n7538 VN.n7533 0.035
R7280 VN.n8383 VN.n8378 0.035
R7281 VN.n9245 VN.n9240 0.035
R7282 VN.n10127 VN.n10122 0.035
R7283 VN.n10996 VN.n10991 0.035
R7284 VN.n1612 VN.n1593 0.035
R7285 VN.n11034 VN.n11033 0.035
R7286 VN.n10172 VN.n10171 0.035
R7287 VN.n9290 VN.n9289 0.035
R7288 VN.n8428 VN.n8427 0.035
R7289 VN.n7583 VN.n7582 0.035
R7290 VN.n7194 VN.n7193 0.035
R7291 VN.n5951 VN.n5950 0.035
R7292 VN.n5159 VN.n5158 0.035
R7293 VN.n4384 VN.n4383 0.035
R7294 VN.n3627 VN.n3626 0.035
R7295 VN.n2887 VN.n2886 0.035
R7296 VN.n5051 VN.n5046 0.035
R7297 VN.n5843 VN.n5838 0.035
R7298 VN.n7086 VN.n7081 0.035
R7299 VN.n7475 VN.n7470 0.035
R7300 VN.n8320 VN.n8315 0.035
R7301 VN.n9182 VN.n9177 0.035
R7302 VN.n10064 VN.n10059 0.035
R7303 VN.n10938 VN.n10933 0.035
R7304 VN.n10978 VN.n10977 0.035
R7305 VN.n10109 VN.n10108 0.035
R7306 VN.n9227 VN.n9226 0.035
R7307 VN.n8365 VN.n8364 0.035
R7308 VN.n7520 VN.n7519 0.035
R7309 VN.n7131 VN.n7130 0.035
R7310 VN.n5888 VN.n5887 0.035
R7311 VN.n5096 VN.n5095 0.035
R7312 VN.n4321 VN.n4320 0.035
R7313 VN.n7023 VN.n7018 0.035
R7314 VN.n7412 VN.n7407 0.035
R7315 VN.n8257 VN.n8252 0.035
R7316 VN.n9119 VN.n9114 0.035
R7317 VN.n10001 VN.n9996 0.035
R7318 VN.n10880 VN.n10875 0.035
R7319 VN.n10920 VN.n10919 0.035
R7320 VN.n10046 VN.n10045 0.035
R7321 VN.n9164 VN.n9163 0.035
R7322 VN.n8302 VN.n8301 0.035
R7323 VN.n7457 VN.n7456 0.035
R7324 VN.n7068 VN.n7067 0.035
R7325 VN.n5825 VN.n5824 0.035
R7326 VN.n10862 VN.n10861 0.035
R7327 VN.n9983 VN.n9982 0.035
R7328 VN.n9101 VN.n9100 0.035
R7329 VN.n8239 VN.n8238 0.035
R7330 VN.n7394 VN.n7393 0.035
R7331 VN.n8194 VN.n8189 0.035
R7332 VN.n9056 VN.n9051 0.035
R7333 VN.n9938 VN.n9933 0.035
R7334 VN.n10822 VN.n10817 0.035
R7335 VN.n9875 VN.n9870 0.035
R7336 VN.n10764 VN.n10759 0.035
R7337 VN.n10804 VN.n10803 0.035
R7338 VN.n9920 VN.n9919 0.035
R7339 VN.n9038 VN.n9037 0.035
R7340 VN.n10746 VN.n10745 0.035
R7341 VN.n9830 VN.n9829 0.035
R7342 VN.n9838 VN.n9837 0.035
R7343 VN.n8984 VN.n8983 0.035
R7344 VN.n8992 VN.n8991 0.035
R7345 VN.n8151 VN.n8150 0.035
R7346 VN.n8159 VN.n8158 0.035
R7347 VN.n7340 VN.n7339 0.035
R7348 VN.n7348 VN.n7347 0.035
R7349 VN.n6547 VN.n6546 0.035
R7350 VN.n6555 VN.n6554 0.035
R7351 VN.n5771 VN.n5770 0.035
R7352 VN.n5779 VN.n5778 0.035
R7353 VN.n5008 VN.n5007 0.035
R7354 VN.n5016 VN.n5015 0.035
R7355 VN.n4267 VN.n4266 0.035
R7356 VN.n4275 VN.n4274 0.035
R7357 VN.n3539 VN.n3538 0.035
R7358 VN.n3547 VN.n3546 0.035
R7359 VN.n2833 VN.n2832 0.035
R7360 VN.n2841 VN.n2840 0.035
R7361 VN.n2140 VN.n2139 0.035
R7362 VN.n2148 VN.n2147 0.035
R7363 VN.n1466 VN.n1465 0.035
R7364 VN.n1474 VN.n1473 0.035
R7365 VN.n191 VN.n190 0.035
R7366 VN.t8 VN.n11664 0.035
R7367 VN.t51 VN.n85 0.035
R7368 VN.t8 VN.n11674 0.035
R7369 VN.t8 VN.n11720 0.035
R7370 VN.t8 VN.n11856 0.035
R7371 VN.t8 VN.n11709 0.035
R7372 VN.t8 VN.n11696 0.035
R7373 VN.t8 VN.n11683 0.035
R7374 VN.t8 VN.n11731 0.035
R7375 VN.t8 VN.n11832 0.035
R7376 VN.t8 VN.n11742 0.035
R7377 VN.t8 VN.n11821 0.035
R7378 VN.t8 VN.n11862 0.035
R7379 VN.t8 VN.n11753 0.035
R7380 VN.t8 VN.n11764 0.035
R7381 VN.t8 VN.n11810 0.035
R7382 VN.t8 VN.n11773 0.035
R7383 VN.t8 VN.n11799 0.035
R7384 VN.t51 VN.n104 0.035
R7385 VN.t51 VN.n108 0.035
R7386 VN.t51 VN.n112 0.035
R7387 VN.t51 VN.n116 0.035
R7388 VN.t51 VN.n120 0.035
R7389 VN.t51 VN.n124 0.035
R7390 VN.t51 VN.n128 0.035
R7391 VN.t51 VN.n132 0.035
R7392 VN.t51 VN.n136 0.035
R7393 VN.t51 VN.n140 0.035
R7394 VN.t51 VN.n144 0.035
R7395 VN.t51 VN.n148 0.035
R7396 VN.t51 VN.n152 0.035
R7397 VN.t51 VN.n156 0.035
R7398 VN.t51 VN.n160 0.035
R7399 VN.t51 VN.n164 0.035
R7400 VN.n80 VN.n79 0.035
R7401 VN.n829 VN.n828 0.034
R7402 VN.n11558 VN.n11557 0.034
R7403 VN.n11719 VN.n11718 0.034
R7404 VN.n11708 VN.n11704 0.034
R7405 VN.n11730 VN.n11729 0.034
R7406 VN.n11741 VN.n11740 0.034
R7407 VN.n11752 VN.n11751 0.034
R7408 VN.n11763 VN.n11762 0.034
R7409 VN.n11772 VN.n11771 0.034
R7410 VN.n12282 VN.n12279 0.034
R7411 VN.n12314 VN.n12309 0.034
R7412 VN.n273 VN.n268 0.034
R7413 VN.n945 VN.n940 0.034
R7414 VN.n1632 VN.n1627 0.034
R7415 VN.n2340 VN.n2335 0.034
R7416 VN.n3059 VN.n3054 0.034
R7417 VN.n3802 VN.n3797 0.034
R7418 VN.n4556 VN.n4551 0.034
R7419 VN.n5334 VN.n5329 0.034
R7420 VN.n6123 VN.n6118 0.034
R7421 VN.n7007 VN.n7002 0.034
R7422 VN.n7755 VN.n7750 0.034
R7423 VN.n8603 VN.n8598 0.034
R7424 VN.n9462 VN.n9457 0.034
R7425 VN.n10676 VN.n10671 0.034
R7426 VN.n11524 VN.n10708 0.034
R7427 VN.n10707 VN.n10706 0.034
R7428 VN.n9827 VN.n9826 0.034
R7429 VN.n8981 VN.n8980 0.034
R7430 VN.n8148 VN.n8147 0.034
R7431 VN.n7337 VN.n7336 0.034
R7432 VN.n6544 VN.n6543 0.034
R7433 VN.n5768 VN.n5767 0.034
R7434 VN.n5005 VN.n5004 0.034
R7435 VN.n4264 VN.n4263 0.034
R7436 VN.n3536 VN.n3535 0.034
R7437 VN.n2830 VN.n2829 0.034
R7438 VN.n2137 VN.n2136 0.034
R7439 VN.n1463 VN.n1462 0.034
R7440 VN.n821 VN.n184 0.034
R7441 VN.n11372 VN.n11370 0.034
R7442 VN.n10345 VN.n10343 0.034
R7443 VN.n9490 VN.n9488 0.034
R7444 VN.n8644 VN.n8642 0.034
R7445 VN.n7813 VN.n7811 0.034
R7446 VN.n6638 VN.n6636 0.034
R7447 VN.n6209 VN.n6207 0.034
R7448 VN.n5435 VN.n5433 0.034
R7449 VN.n4674 VN.n4672 0.034
R7450 VN.n3933 VN.n3931 0.034
R7451 VN.n3207 VN.n3205 0.034
R7452 VN.n2501 VN.n2499 0.034
R7453 VN.n1810 VN.n1808 0.034
R7454 VN.n1136 VN.n1134 0.034
R7455 VN.n484 VN.n482 0.034
R7456 VN.n12691 VN.n12689 0.034
R7457 VN.n12361 VN.n12356 0.034
R7458 VN.n175 VN.n171 0.034
R7459 VN.n1140 VN.n1131 0.034
R7460 VN.n1814 VN.n1805 0.034
R7461 VN.n2505 VN.n2496 0.034
R7462 VN.n3211 VN.n3202 0.034
R7463 VN.n3937 VN.n3928 0.034
R7464 VN.n4678 VN.n4669 0.034
R7465 VN.n5439 VN.n5430 0.034
R7466 VN.n6213 VN.n6204 0.034
R7467 VN.n6642 VN.n6633 0.034
R7468 VN.n7817 VN.n7808 0.034
R7469 VN.n8648 VN.n8639 0.034
R7470 VN.n9494 VN.n9485 0.034
R7471 VN.n10349 VN.n10340 0.034
R7472 VN.n11376 VN.n11367 0.034
R7473 VN.n25 VN.n24 0.034
R7474 VN.n91 VN.n90 0.034
R7475 VN.t8 VN.n11667 0.034
R7476 VN.t51 VN.n84 0.034
R7477 VN.t8 VN.n11677 0.034
R7478 VN.t8 VN.n11723 0.034
R7479 VN.t8 VN.n11859 0.034
R7480 VN.t8 VN.n11712 0.034
R7481 VN.t8 VN.n11699 0.034
R7482 VN.t8 VN.n11686 0.034
R7483 VN.t8 VN.n11734 0.034
R7484 VN.t8 VN.n11835 0.034
R7485 VN.t8 VN.n11745 0.034
R7486 VN.t8 VN.n11824 0.034
R7487 VN.t8 VN.n11863 0.034
R7488 VN.t8 VN.n11756 0.034
R7489 VN.t8 VN.n11767 0.034
R7490 VN.t8 VN.n11813 0.034
R7491 VN.t8 VN.n11776 0.034
R7492 VN.t8 VN.n11802 0.034
R7493 VN.t51 VN.n107 0.034
R7494 VN.t51 VN.n111 0.034
R7495 VN.t51 VN.n115 0.034
R7496 VN.t51 VN.n119 0.034
R7497 VN.t51 VN.n123 0.034
R7498 VN.t51 VN.n127 0.034
R7499 VN.t51 VN.n131 0.034
R7500 VN.t51 VN.n135 0.034
R7501 VN.t51 VN.n139 0.034
R7502 VN.t51 VN.n143 0.034
R7503 VN.t51 VN.n147 0.034
R7504 VN.t51 VN.n151 0.034
R7505 VN.t51 VN.n155 0.034
R7506 VN.t51 VN.n159 0.034
R7507 VN.t51 VN.n163 0.034
R7508 VN.t51 VN.n167 0.034
R7509 VN.n11538 VN.n11534 0.034
R7510 VN.n10718 VN.n10714 0.034
R7511 VN.n9858 VN.n9854 0.034
R7512 VN.n9010 VN.n9006 0.034
R7513 VN.n8177 VN.n8173 0.034
R7514 VN.n7366 VN.n7362 0.034
R7515 VN.n6573 VN.n6569 0.034
R7516 VN.n5797 VN.n5793 0.034
R7517 VN.n5034 VN.n5030 0.034
R7518 VN.n4293 VN.n4289 0.034
R7519 VN.n3565 VN.n3561 0.034
R7520 VN.n2859 VN.n2855 0.034
R7521 VN.n2166 VN.n2162 0.034
R7522 VN.n1492 VN.n1488 0.034
R7523 VN.n842 VN.n838 0.034
R7524 VN.n815 VN.n811 0.034
R7525 VN.n13131 VN.n13127 0.034
R7526 VN.n10565 VN.n10564 0.033
R7527 VN.n12404 VN.n12403 0.033
R7528 VN.n11788 VN.n11787 0.032
R7529 VN.n12365 VN.n12354 0.032
R7530 VN.n12695 VN.n12686 0.032
R7531 VN.n10575 VN.n10574 0.032
R7532 VN.n9690 VN.n9689 0.032
R7533 VN.n8828 VN.n8827 0.032
R7534 VN.n7979 VN.n7978 0.032
R7535 VN.n6788 VN.n6787 0.032
R7536 VN.n6343 VN.n6342 0.032
R7537 VN.n5551 VN.n5550 0.032
R7538 VN.n4772 VN.n4771 0.032
R7539 VN.n4015 VN.n4014 0.032
R7540 VN.n3271 VN.n3270 0.032
R7541 VN.n2549 VN.n2548 0.032
R7542 VN.n1840 VN.n1839 0.032
R7543 VN.n1150 VN.n1149 0.032
R7544 VN.n475 VN.n474 0.032
R7545 VN.n10597 VN.n10596 0.032
R7546 VN.t35 VN.n11365 0.031
R7547 VN.t82 VN.n12371 0.031
R7548 VN.t57 VN.n2512 0.031
R7549 VN.t108 VN.n1820 0.031
R7550 VN.t94 VN.n1147 0.031
R7551 VN.t41 VN.n494 0.031
R7552 VN.t101 VN.n12702 0.031
R7553 VN.t28 VN.n3944 0.031
R7554 VN.t183 VN.n3217 0.031
R7555 VN.t176 VN.n5446 0.031
R7556 VN.t32 VN.n4684 0.031
R7557 VN.t146 VN.n6221 0.031
R7558 VN.t253 VN.n6649 0.031
R7559 VN.t39 VN.n8655 0.031
R7560 VN.t73 VN.n7823 0.031
R7561 VN.t241 VN.n10356 0.031
R7562 VN.t0 VN.n9500 0.031
R7563 VN.n11572 VN.n11549 0.031
R7564 VN.n204 VN.n203 0.031
R7565 VN.n875 VN.n874 0.031
R7566 VN.n1558 VN.n1557 0.031
R7567 VN.n2266 VN.n2265 0.031
R7568 VN.n2988 VN.n2987 0.031
R7569 VN.n3728 VN.n3727 0.031
R7570 VN.n4485 VN.n4484 0.031
R7571 VN.n5260 VN.n5259 0.031
R7572 VN.n6052 VN.n6051 0.031
R7573 VN.n7295 VN.n7294 0.031
R7574 VN.n7684 VN.n7683 0.031
R7575 VN.n8529 VN.n8528 0.031
R7576 VN.n9391 VN.n9390 0.031
R7577 VN.n10274 VN.n10273 0.031
R7578 VN.n3577 VN.n3576 0.031
R7579 VN.n4334 VN.n4333 0.031
R7580 VN.n5109 VN.n5108 0.031
R7581 VN.n5901 VN.n5900 0.031
R7582 VN.n7144 VN.n7143 0.031
R7583 VN.n7533 VN.n7532 0.031
R7584 VN.n8378 VN.n8377 0.031
R7585 VN.n9240 VN.n9239 0.031
R7586 VN.n10122 VN.n10121 0.031
R7587 VN.n10991 VN.n10990 0.031
R7588 VN.n11033 VN.n11032 0.031
R7589 VN.n10171 VN.n10170 0.031
R7590 VN.n9289 VN.n9288 0.031
R7591 VN.n8427 VN.n8426 0.031
R7592 VN.n7582 VN.n7581 0.031
R7593 VN.n7193 VN.n7192 0.031
R7594 VN.n5950 VN.n5949 0.031
R7595 VN.n5158 VN.n5157 0.031
R7596 VN.n4383 VN.n4382 0.031
R7597 VN.n3626 VN.n3625 0.031
R7598 VN.n2886 VN.n2885 0.031
R7599 VN.n5046 VN.n5045 0.031
R7600 VN.n5838 VN.n5837 0.031
R7601 VN.n7081 VN.n7080 0.031
R7602 VN.n7470 VN.n7469 0.031
R7603 VN.n8315 VN.n8314 0.031
R7604 VN.n9177 VN.n9176 0.031
R7605 VN.n10059 VN.n10058 0.031
R7606 VN.n10933 VN.n10932 0.031
R7607 VN.n10977 VN.n10976 0.031
R7608 VN.n10108 VN.n10107 0.031
R7609 VN.n9226 VN.n9225 0.031
R7610 VN.n8364 VN.n8363 0.031
R7611 VN.n7519 VN.n7518 0.031
R7612 VN.n7130 VN.n7129 0.031
R7613 VN.n5887 VN.n5886 0.031
R7614 VN.n5095 VN.n5094 0.031
R7615 VN.n4320 VN.n4319 0.031
R7616 VN.n7018 VN.n7017 0.031
R7617 VN.n7407 VN.n7406 0.031
R7618 VN.n8252 VN.n8251 0.031
R7619 VN.n9114 VN.n9113 0.031
R7620 VN.n9996 VN.n9995 0.031
R7621 VN.n10875 VN.n10874 0.031
R7622 VN.n10919 VN.n10918 0.031
R7623 VN.n10045 VN.n10044 0.031
R7624 VN.n9163 VN.n9162 0.031
R7625 VN.n8301 VN.n8300 0.031
R7626 VN.n7456 VN.n7455 0.031
R7627 VN.n7067 VN.n7066 0.031
R7628 VN.n5824 VN.n5823 0.031
R7629 VN.n10861 VN.n10860 0.031
R7630 VN.n9982 VN.n9981 0.031
R7631 VN.n9100 VN.n9099 0.031
R7632 VN.n8238 VN.n8237 0.031
R7633 VN.n7393 VN.n7392 0.031
R7634 VN.n8189 VN.n8188 0.031
R7635 VN.n9051 VN.n9050 0.031
R7636 VN.n9933 VN.n9932 0.031
R7637 VN.n10817 VN.n10816 0.031
R7638 VN.n9870 VN.n9869 0.031
R7639 VN.n10759 VN.n10758 0.031
R7640 VN.n10803 VN.n10802 0.031
R7641 VN.n9919 VN.n9918 0.031
R7642 VN.n9037 VN.n9036 0.031
R7643 VN.n10745 VN.n10744 0.031
R7644 VN.n12181 VN.n12180 0.031
R7645 VN.n12312 VN.n12311 0.031
R7646 VN.n271 VN.n270 0.031
R7647 VN.n943 VN.n942 0.031
R7648 VN.n1630 VN.n1629 0.031
R7649 VN.n2338 VN.n2337 0.031
R7650 VN.n3057 VN.n3056 0.031
R7651 VN.n3800 VN.n3799 0.031
R7652 VN.n4554 VN.n4553 0.031
R7653 VN.n5332 VN.n5331 0.031
R7654 VN.n6121 VN.n6120 0.031
R7655 VN.n7005 VN.n7004 0.031
R7656 VN.n7753 VN.n7752 0.031
R7657 VN.n8601 VN.n8600 0.031
R7658 VN.n9460 VN.n9459 0.031
R7659 VN.n10674 VN.n10673 0.031
R7660 VN.n11482 VN.n11481 0.031
R7661 VN.n11549 VN.n11548 0.031
R7662 VN.n2318 VN.n2317 0.031
R7663 VN.n8581 VN.n8580 0.031
R7664 VN.n10326 VN.n10325 0.031
R7665 VN.n2303 VN.n2302 0.03
R7666 VN.n3765 VN.n3764 0.03
R7667 VN.n5297 VN.n5296 0.03
R7668 VN.n8566 VN.n8565 0.03
R7669 VN.n10311 VN.n10310 0.03
R7670 VN.n1520 VN.n1519 0.03
R7671 VN.n2228 VN.n2227 0.03
R7672 VN.n2950 VN.n2949 0.03
R7673 VN.n3690 VN.n3689 0.03
R7674 VN.n4447 VN.n4446 0.03
R7675 VN.n5222 VN.n5221 0.03
R7676 VN.n6014 VN.n6013 0.03
R7677 VN.n7257 VN.n7256 0.03
R7678 VN.n7646 VN.n7645 0.03
R7679 VN.n8491 VN.n8490 0.03
R7680 VN.n9353 VN.n9352 0.03
R7681 VN.n10236 VN.n10235 0.03
R7682 VN.n11081 VN.n11080 0.03
R7683 VN.n12092 VN.n12091 0.03
R7684 VN.n6591 VN.n6590 0.03
R7685 VN.n3032 VN.n3027 0.029
R7686 VN.n1605 VN.n1600 0.029
R7687 VN.n4529 VN.n4524 0.029
R7688 VN.n6096 VN.n6091 0.029
R7689 VN.n7728 VN.n7723 0.029
R7690 VN.n9435 VN.n9430 0.029
R7691 VN.n11461 VN.n11460 0.029
R7692 VN.n10625 VN.n10624 0.029
R7693 VN.n10293 VN.n10292 0.029
R7694 VN.n9410 VN.n9409 0.029
R7695 VN.n8548 VN.n8547 0.029
R7696 VN.n7703 VN.n7702 0.029
R7697 VN.n7314 VN.n7313 0.029
R7698 VN.n6071 VN.n6070 0.029
R7699 VN.n5279 VN.n5278 0.029
R7700 VN.n4504 VN.n4503 0.029
R7701 VN.n3747 VN.n3746 0.029
R7702 VN.n3007 VN.n3006 0.029
R7703 VN.n2285 VN.n2284 0.029
R7704 VN.n1577 VN.n1576 0.029
R7705 VN.n894 VN.n893 0.029
R7706 VN.n223 VN.n222 0.029
R7707 VN.n10553 VN.n10552 0.029
R7708 VN.n10205 VN.n10204 0.029
R7709 VN.n9322 VN.n9321 0.029
R7710 VN.n8460 VN.n8459 0.029
R7711 VN.n7615 VN.n7614 0.029
R7712 VN.n7226 VN.n7225 0.029
R7713 VN.n5983 VN.n5982 0.029
R7714 VN.n5191 VN.n5190 0.029
R7715 VN.n4416 VN.n4415 0.029
R7716 VN.n3659 VN.n3658 0.029
R7717 VN.n2919 VN.n2918 0.029
R7718 VN.n2197 VN.n2196 0.029
R7719 VN.n10523 VN.n10522 0.029
R7720 VN.n10141 VN.n10140 0.029
R7721 VN.n9259 VN.n9258 0.029
R7722 VN.n8397 VN.n8396 0.029
R7723 VN.n7552 VN.n7551 0.029
R7724 VN.n7163 VN.n7162 0.029
R7725 VN.n5920 VN.n5919 0.029
R7726 VN.n5128 VN.n5127 0.029
R7727 VN.n4353 VN.n4352 0.029
R7728 VN.n3596 VN.n3595 0.029
R7729 VN.n10488 VN.n10487 0.029
R7730 VN.n10078 VN.n10077 0.029
R7731 VN.n9196 VN.n9195 0.029
R7732 VN.n8334 VN.n8333 0.029
R7733 VN.n7489 VN.n7488 0.029
R7734 VN.n7100 VN.n7099 0.029
R7735 VN.n5857 VN.n5856 0.029
R7736 VN.n5065 VN.n5064 0.029
R7737 VN.n10453 VN.n10452 0.029
R7738 VN.n10015 VN.n10014 0.029
R7739 VN.n9133 VN.n9132 0.029
R7740 VN.n8271 VN.n8270 0.029
R7741 VN.n7426 VN.n7425 0.029
R7742 VN.n7037 VN.n7036 0.029
R7743 VN.n10418 VN.n10417 0.029
R7744 VN.n9952 VN.n9951 0.029
R7745 VN.n9070 VN.n9069 0.029
R7746 VN.n8208 VN.n8207 0.029
R7747 VN.n10383 VN.n10382 0.029
R7748 VN.n9889 VN.n9888 0.029
R7749 VN.n9309 VN.n9308 0.029
R7750 VN.n8447 VN.n8446 0.029
R7751 VN.n7602 VN.n7601 0.029
R7752 VN.n7213 VN.n7212 0.029
R7753 VN.n5970 VN.n5969 0.029
R7754 VN.n5178 VN.n5177 0.029
R7755 VN.n4403 VN.n4402 0.029
R7756 VN.n3646 VN.n3645 0.029
R7757 VN.n2906 VN.n2905 0.029
R7758 VN.n2184 VN.n2183 0.029
R7759 VN.n1519 VN.n1518 0.029
R7760 VN.n2227 VN.n2226 0.029
R7761 VN.n2949 VN.n2948 0.029
R7762 VN.n3689 VN.n3688 0.029
R7763 VN.n4446 VN.n4445 0.029
R7764 VN.n5221 VN.n5220 0.029
R7765 VN.n6013 VN.n6012 0.029
R7766 VN.n7256 VN.n7255 0.029
R7767 VN.n7645 VN.n7644 0.029
R7768 VN.n8490 VN.n8489 0.029
R7769 VN.n9352 VN.n9351 0.029
R7770 VN.n10235 VN.n10234 0.029
R7771 VN.n11080 VN.n11079 0.029
R7772 VN.n12091 VN.n12090 0.029
R7773 VN.n195 VN.n194 0.028
R7774 VN.n204 VN.n201 0.028
R7775 VN.n875 VN.n872 0.028
R7776 VN.n1558 VN.n1555 0.028
R7777 VN.n2266 VN.n2263 0.028
R7778 VN.n2988 VN.n2985 0.028
R7779 VN.n3728 VN.n3725 0.028
R7780 VN.n4485 VN.n4482 0.028
R7781 VN.n5260 VN.n5257 0.028
R7782 VN.n6052 VN.n6049 0.028
R7783 VN.n7295 VN.n7292 0.028
R7784 VN.n7684 VN.n7681 0.028
R7785 VN.n8529 VN.n8526 0.028
R7786 VN.n9391 VN.n9388 0.028
R7787 VN.n10274 VN.n10271 0.028
R7788 VN.n3577 VN.n3574 0.028
R7789 VN.n4334 VN.n4331 0.028
R7790 VN.n5109 VN.n5106 0.028
R7791 VN.n5901 VN.n5898 0.028
R7792 VN.n7144 VN.n7141 0.028
R7793 VN.n7533 VN.n7530 0.028
R7794 VN.n8378 VN.n8375 0.028
R7795 VN.n9240 VN.n9237 0.028
R7796 VN.n10122 VN.n10119 0.028
R7797 VN.n10991 VN.n10988 0.028
R7798 VN.n10171 VN.n10168 0.028
R7799 VN.n9289 VN.n9286 0.028
R7800 VN.n8427 VN.n8424 0.028
R7801 VN.n7582 VN.n7579 0.028
R7802 VN.n7193 VN.n7190 0.028
R7803 VN.n5950 VN.n5947 0.028
R7804 VN.n5158 VN.n5155 0.028
R7805 VN.n4383 VN.n4380 0.028
R7806 VN.n3626 VN.n3623 0.028
R7807 VN.n2886 VN.n2883 0.028
R7808 VN.n5046 VN.n5043 0.028
R7809 VN.n5838 VN.n5835 0.028
R7810 VN.n7081 VN.n7078 0.028
R7811 VN.n7470 VN.n7467 0.028
R7812 VN.n8315 VN.n8312 0.028
R7813 VN.n9177 VN.n9174 0.028
R7814 VN.n10059 VN.n10056 0.028
R7815 VN.n10933 VN.n10930 0.028
R7816 VN.n10977 VN.n10974 0.028
R7817 VN.n10108 VN.n10105 0.028
R7818 VN.n9226 VN.n9223 0.028
R7819 VN.n8364 VN.n8361 0.028
R7820 VN.n7519 VN.n7516 0.028
R7821 VN.n7130 VN.n7127 0.028
R7822 VN.n5887 VN.n5884 0.028
R7823 VN.n5095 VN.n5092 0.028
R7824 VN.n4320 VN.n4317 0.028
R7825 VN.n7018 VN.n7015 0.028
R7826 VN.n7407 VN.n7404 0.028
R7827 VN.n8252 VN.n8249 0.028
R7828 VN.n9114 VN.n9111 0.028
R7829 VN.n9996 VN.n9993 0.028
R7830 VN.n10875 VN.n10872 0.028
R7831 VN.n10919 VN.n10916 0.028
R7832 VN.n10045 VN.n10042 0.028
R7833 VN.n9163 VN.n9160 0.028
R7834 VN.n8301 VN.n8298 0.028
R7835 VN.n7456 VN.n7453 0.028
R7836 VN.n7067 VN.n7064 0.028
R7837 VN.n5824 VN.n5821 0.028
R7838 VN.n10861 VN.n10858 0.028
R7839 VN.n9982 VN.n9979 0.028
R7840 VN.n9100 VN.n9097 0.028
R7841 VN.n8238 VN.n8235 0.028
R7842 VN.n7393 VN.n7390 0.028
R7843 VN.n8189 VN.n8186 0.028
R7844 VN.n9051 VN.n9048 0.028
R7845 VN.n9933 VN.n9930 0.028
R7846 VN.n10817 VN.n10814 0.028
R7847 VN.n9870 VN.n9867 0.028
R7848 VN.n10759 VN.n10756 0.028
R7849 VN.n10803 VN.n10800 0.028
R7850 VN.n9919 VN.n9916 0.028
R7851 VN.n9037 VN.n9034 0.028
R7852 VN.n10745 VN.n10742 0.028
R7853 VN.n10221 VN.n10220 0.028
R7854 VN.n10223 VN.n10221 0.028
R7855 VN.n9338 VN.n9337 0.028
R7856 VN.n9340 VN.n9338 0.028
R7857 VN.n8476 VN.n8475 0.028
R7858 VN.n8478 VN.n8476 0.028
R7859 VN.n7631 VN.n7630 0.028
R7860 VN.n7633 VN.n7631 0.028
R7861 VN.n7242 VN.n7241 0.028
R7862 VN.n7244 VN.n7242 0.028
R7863 VN.n5999 VN.n5998 0.028
R7864 VN.n6001 VN.n5999 0.028
R7865 VN.n5207 VN.n5206 0.028
R7866 VN.n5209 VN.n5207 0.028
R7867 VN.n4432 VN.n4431 0.028
R7868 VN.n4434 VN.n4432 0.028
R7869 VN.n3675 VN.n3674 0.028
R7870 VN.n3677 VN.n3675 0.028
R7871 VN.n2935 VN.n2934 0.028
R7872 VN.n2937 VN.n2935 0.028
R7873 VN.n2213 VN.n2212 0.028
R7874 VN.n2215 VN.n2213 0.028
R7875 VN.n1505 VN.n1504 0.028
R7876 VN.n1507 VN.n1505 0.028
R7877 VN.n911 VN.n910 0.028
R7878 VN.n913 VN.n911 0.028
R7879 VN.n11408 VN.n11407 0.028
R7880 VN.n11410 VN.n11408 0.028
R7881 VN.n11435 VN.n11434 0.028
R7882 VN.n11437 VN.n11435 0.028
R7883 VN.n11537 VN.n11536 0.028
R7884 VN.n10717 VN.n10716 0.028
R7885 VN.n9857 VN.n9856 0.028
R7886 VN.n9009 VN.n9008 0.028
R7887 VN.n8176 VN.n8175 0.028
R7888 VN.n7365 VN.n7364 0.028
R7889 VN.n6572 VN.n6571 0.028
R7890 VN.n5796 VN.n5795 0.028
R7891 VN.n5033 VN.n5032 0.028
R7892 VN.n4292 VN.n4291 0.028
R7893 VN.n3564 VN.n3563 0.028
R7894 VN.n2858 VN.n2857 0.028
R7895 VN.n2165 VN.n2164 0.028
R7896 VN.n1491 VN.n1490 0.028
R7897 VN.n841 VN.n840 0.028
R7898 VN.n814 VN.n813 0.028
R7899 VN.n13130 VN.n13129 0.028
R7900 VN.n12252 VN.n12251 0.028
R7901 VN.n1605 VN.n1604 0.028
R7902 VN.n3032 VN.n3031 0.028
R7903 VN.n4529 VN.n4528 0.028
R7904 VN.n6096 VN.n6095 0.028
R7905 VN.n7728 VN.n7727 0.028
R7906 VN.n9435 VN.n9434 0.028
R7907 VN.n10192 VN.n10191 0.028
R7908 VN.n13095 VN.n13093 0.027
R7909 VN.n784 VN.n782 0.027
R7910 VN.n12115 VN.n12110 0.027
R7911 VN.n12138 VN.n12137 0.027
R7912 VN.n2317 VN.n2316 0.027
R7913 VN.n3778 VN.n3777 0.027
R7914 VN.n5310 VN.n5309 0.027
R7915 VN.n6598 VN.n6597 0.027
R7916 VN.n8580 VN.n8579 0.027
R7917 VN.n10325 VN.n10324 0.027
R7918 VN.n11524 VN.n11523 0.027
R7919 VN.n10673 VN.n10672 0.027
R7920 VN.n10671 VN.n10670 0.027
R7921 VN.n9459 VN.n9458 0.027
R7922 VN.n9457 VN.n9456 0.027
R7923 VN.n8600 VN.n8599 0.027
R7924 VN.n8598 VN.n8597 0.027
R7925 VN.n7752 VN.n7751 0.027
R7926 VN.n7750 VN.n7749 0.027
R7927 VN.n7004 VN.n7003 0.027
R7928 VN.n7002 VN.n7001 0.027
R7929 VN.n6120 VN.n6119 0.027
R7930 VN.n6118 VN.n6117 0.027
R7931 VN.n5331 VN.n5330 0.027
R7932 VN.n5329 VN.n5328 0.027
R7933 VN.n4553 VN.n4552 0.027
R7934 VN.n4551 VN.n4550 0.027
R7935 VN.n3799 VN.n3798 0.027
R7936 VN.n3797 VN.n3796 0.027
R7937 VN.n3056 VN.n3055 0.027
R7938 VN.n3054 VN.n3053 0.027
R7939 VN.n2337 VN.n2336 0.027
R7940 VN.n2335 VN.n2334 0.027
R7941 VN.n1629 VN.n1628 0.027
R7942 VN.n1627 VN.n1626 0.027
R7943 VN.n942 VN.n941 0.027
R7944 VN.n940 VN.n939 0.027
R7945 VN.n270 VN.n269 0.027
R7946 VN.n268 VN.n267 0.027
R7947 VN.n12311 VN.n12310 0.027
R7948 VN.n12309 VN.n12308 0.027
R7949 VN.n10543 VN.n10542 0.027
R7950 VN.n11118 VN.n11117 0.026
R7951 VN.n11465 VN.n11462 0.026
R7952 VN.n10627 VN.n10626 0.026
R7953 VN.n10297 VN.n10294 0.026
R7954 VN.n9739 VN.n9738 0.026
R7955 VN.n9414 VN.n9411 0.026
R7956 VN.n8877 VN.n8876 0.026
R7957 VN.n8552 VN.n8549 0.026
R7958 VN.n8028 VN.n8027 0.026
R7959 VN.n7707 VN.n7704 0.026
R7960 VN.n6837 VN.n6836 0.026
R7961 VN.n7318 VN.n7315 0.026
R7962 VN.n6392 VN.n6391 0.026
R7963 VN.n6075 VN.n6072 0.026
R7964 VN.n5600 VN.n5599 0.026
R7965 VN.n5283 VN.n5280 0.026
R7966 VN.n4821 VN.n4820 0.026
R7967 VN.n4508 VN.n4505 0.026
R7968 VN.n4064 VN.n4063 0.026
R7969 VN.n3751 VN.n3748 0.026
R7970 VN.n3320 VN.n3319 0.026
R7971 VN.n3011 VN.n3008 0.026
R7972 VN.n2598 VN.n2597 0.026
R7973 VN.n2289 VN.n2286 0.026
R7974 VN.n1889 VN.n1888 0.026
R7975 VN.n1581 VN.n1578 0.026
R7976 VN.n1199 VN.n1198 0.026
R7977 VN.n898 VN.n895 0.026
R7978 VN.n524 VN.n523 0.026
R7979 VN.n227 VN.n224 0.026
R7980 VN.n12713 VN.n12712 0.026
R7981 VN.n12259 VN.n12253 0.026
R7982 VN.n11069 VN.n11047 0.026
R7983 VN.n10566 VN.n10554 0.026
R7984 VN.n10209 VN.n10206 0.026
R7985 VN.n9681 VN.n9680 0.026
R7986 VN.n9326 VN.n9323 0.026
R7987 VN.n8819 VN.n8818 0.026
R7988 VN.n8464 VN.n8461 0.026
R7989 VN.n7970 VN.n7969 0.026
R7990 VN.n7619 VN.n7616 0.026
R7991 VN.n6779 VN.n6778 0.026
R7992 VN.n7230 VN.n7227 0.026
R7993 VN.n6334 VN.n6333 0.026
R7994 VN.n5987 VN.n5984 0.026
R7995 VN.n5542 VN.n5541 0.026
R7996 VN.n5195 VN.n5192 0.026
R7997 VN.n4763 VN.n4762 0.026
R7998 VN.n4420 VN.n4417 0.026
R7999 VN.n4006 VN.n4005 0.026
R8000 VN.n3663 VN.n3660 0.026
R8001 VN.n3262 VN.n3261 0.026
R8002 VN.n2923 VN.n2920 0.026
R8003 VN.n2540 VN.n2539 0.026
R8004 VN.n2201 VN.n2198 0.026
R8005 VN.n1831 VN.n1830 0.026
R8006 VN.n1612 VN.n1606 0.026
R8007 VN.n10577 VN.n10575 0.026
R8008 VN.n9692 VN.n9690 0.026
R8009 VN.n8830 VN.n8828 0.026
R8010 VN.n7981 VN.n7979 0.026
R8011 VN.n6790 VN.n6788 0.026
R8012 VN.n6345 VN.n6343 0.026
R8013 VN.n5553 VN.n5551 0.026
R8014 VN.n4774 VN.n4772 0.026
R8015 VN.n4017 VN.n4015 0.026
R8016 VN.n3273 VN.n3271 0.026
R8017 VN.n2551 VN.n2549 0.026
R8018 VN.n1842 VN.n1840 0.026
R8019 VN.n1152 VN.n1150 0.026
R8020 VN.n506 VN.n505 0.026
R8021 VN.n1181 VN.n1180 0.026
R8022 VN.n1871 VN.n1870 0.026
R8023 VN.n2580 VN.n2579 0.026
R8024 VN.n3302 VN.n3301 0.026
R8025 VN.n4046 VN.n4045 0.026
R8026 VN.n4803 VN.n4802 0.026
R8027 VN.n5582 VN.n5581 0.026
R8028 VN.n6374 VN.n6373 0.026
R8029 VN.n6819 VN.n6818 0.026
R8030 VN.n8010 VN.n8009 0.026
R8031 VN.n8859 VN.n8858 0.026
R8032 VN.n9721 VN.n9720 0.026
R8033 VN.n10598 VN.n10597 0.026
R8034 VN.n11441 VN.n11425 0.026
R8035 VN.n10263 VN.n10253 0.026
R8036 VN.n9380 VN.n9370 0.026
R8037 VN.n8518 VN.n8508 0.026
R8038 VN.n7673 VN.n7663 0.026
R8039 VN.n7284 VN.n7274 0.026
R8040 VN.n6041 VN.n6031 0.026
R8041 VN.n5249 VN.n5239 0.026
R8042 VN.n4474 VN.n4464 0.026
R8043 VN.n3717 VN.n3707 0.026
R8044 VN.n2977 VN.n2967 0.026
R8045 VN.n2255 VN.n2245 0.026
R8046 VN.n1550 VN.n1540 0.026
R8047 VN.n864 VN.n854 0.026
R8048 VN.n253 VN.n243 0.026
R8049 VN.n12144 VN.n12128 0.026
R8050 VN.n2320 VN.n2304 0.026
R8051 VN.n2889 VN.n2871 0.026
R8052 VN.n3629 VN.n3611 0.026
R8053 VN.n4386 VN.n4368 0.026
R8054 VN.n5161 VN.n5143 0.026
R8055 VN.n5953 VN.n5935 0.026
R8056 VN.n7196 VN.n7178 0.026
R8057 VN.n7585 VN.n7567 0.026
R8058 VN.n8430 VN.n8412 0.026
R8059 VN.n9292 VN.n9274 0.026
R8060 VN.n10174 VN.n10156 0.026
R8061 VN.n11036 VN.n11021 0.026
R8062 VN.n11009 VN.n11006 0.026
R8063 VN.n10525 VN.n10524 0.026
R8064 VN.n10145 VN.n10142 0.026
R8065 VN.n9647 VN.n9646 0.026
R8066 VN.n9263 VN.n9260 0.026
R8067 VN.n8785 VN.n8784 0.026
R8068 VN.n8401 VN.n8398 0.026
R8069 VN.n7936 VN.n7935 0.026
R8070 VN.n7556 VN.n7553 0.026
R8071 VN.n6745 VN.n6744 0.026
R8072 VN.n7167 VN.n7164 0.026
R8073 VN.n6300 VN.n6299 0.026
R8074 VN.n5924 VN.n5921 0.026
R8075 VN.n5508 VN.n5507 0.026
R8076 VN.n5132 VN.n5129 0.026
R8077 VN.n4729 VN.n4728 0.026
R8078 VN.n4357 VN.n4354 0.026
R8079 VN.n3972 VN.n3971 0.026
R8080 VN.n3600 VN.n3597 0.026
R8081 VN.n3228 VN.n3227 0.026
R8082 VN.n3039 VN.n3033 0.026
R8083 VN.n3782 VN.n3766 0.026
R8084 VN.n4323 VN.n4305 0.026
R8085 VN.n5098 VN.n5080 0.026
R8086 VN.n5890 VN.n5872 0.026
R8087 VN.n7133 VN.n7115 0.026
R8088 VN.n7522 VN.n7504 0.026
R8089 VN.n8367 VN.n8349 0.026
R8090 VN.n9229 VN.n9211 0.026
R8091 VN.n10111 VN.n10093 0.026
R8092 VN.n10980 VN.n10963 0.026
R8093 VN.n10951 VN.n10948 0.026
R8094 VN.n10490 VN.n10489 0.026
R8095 VN.n10082 VN.n10079 0.026
R8096 VN.n9613 VN.n9612 0.026
R8097 VN.n9200 VN.n9197 0.026
R8098 VN.n8751 VN.n8750 0.026
R8099 VN.n8338 VN.n8335 0.026
R8100 VN.n7902 VN.n7901 0.026
R8101 VN.n7493 VN.n7490 0.026
R8102 VN.n6711 VN.n6710 0.026
R8103 VN.n7104 VN.n7101 0.026
R8104 VN.n6266 VN.n6265 0.026
R8105 VN.n5861 VN.n5858 0.026
R8106 VN.n5474 VN.n5473 0.026
R8107 VN.n5069 VN.n5066 0.026
R8108 VN.n4695 VN.n4694 0.026
R8109 VN.n4536 VN.n4530 0.026
R8110 VN.n5314 VN.n5298 0.026
R8111 VN.n5827 VN.n5809 0.026
R8112 VN.n7070 VN.n7052 0.026
R8113 VN.n7459 VN.n7441 0.026
R8114 VN.n8304 VN.n8286 0.026
R8115 VN.n9166 VN.n9148 0.026
R8116 VN.n10048 VN.n10030 0.026
R8117 VN.n10922 VN.n10905 0.026
R8118 VN.n10893 VN.n10890 0.026
R8119 VN.n10455 VN.n10454 0.026
R8120 VN.n10019 VN.n10016 0.026
R8121 VN.n9579 VN.n9578 0.026
R8122 VN.n9137 VN.n9134 0.026
R8123 VN.n8717 VN.n8716 0.026
R8124 VN.n8275 VN.n8272 0.026
R8125 VN.n7868 VN.n7867 0.026
R8126 VN.n7430 VN.n7427 0.026
R8127 VN.n6677 VN.n6676 0.026
R8128 VN.n7041 VN.n7038 0.026
R8129 VN.n6232 VN.n6231 0.026
R8130 VN.n6103 VN.n6097 0.026
R8131 VN.n10835 VN.n10832 0.026
R8132 VN.n10420 VN.n10419 0.026
R8133 VN.n9956 VN.n9953 0.026
R8134 VN.n9545 VN.n9544 0.026
R8135 VN.n9074 VN.n9071 0.026
R8136 VN.n8683 VN.n8682 0.026
R8137 VN.n8212 VN.n8209 0.026
R8138 VN.n7834 VN.n7833 0.026
R8139 VN.n7735 VN.n7729 0.026
R8140 VN.n8583 VN.n8567 0.026
R8141 VN.n9040 VN.n9022 0.026
R8142 VN.n9922 VN.n9904 0.026
R8143 VN.n10806 VN.n10789 0.026
R8144 VN.n10777 VN.n10774 0.026
R8145 VN.n10385 VN.n10384 0.026
R8146 VN.n9893 VN.n9890 0.026
R8147 VN.n9511 VN.n9510 0.026
R8148 VN.n9442 VN.n9436 0.026
R8149 VN.n10328 VN.n10312 0.026
R8150 VN.n10748 VN.n10731 0.026
R8151 VN.n11489 VN.n11483 0.026
R8152 VN.n11567 VN.n11559 0.026
R8153 VN.n12737 VN.n12722 0.026
R8154 VN.n184 VN.n183 0.026
R8155 VN.n11567 VN.n11564 0.026
R8156 VN.n10864 VN.n10846 0.026
R8157 VN.n9985 VN.n9967 0.026
R8158 VN.n9103 VN.n9085 0.026
R8159 VN.n8241 VN.n8223 0.026
R8160 VN.n7396 VN.n7378 0.026
R8161 VN.t76 VN.n6592 0.026
R8162 VN.n11558 VN.n11556 0.026
R8163 VN.n12081 VN.n12080 0.026
R8164 VN.n11924 VN.n11923 0.026
R8165 VN.n12376 VN.n12375 0.026
R8166 VN.n12396 VN.n12395 0.025
R8167 VN.n10542 VN.n10541 0.025
R8168 VN.t8 VN.n11658 0.025
R8169 VN.t8 VN.n11838 0.025
R8170 VN.t8 VN.n11827 0.025
R8171 VN.t8 VN.n11816 0.025
R8172 VN.t8 VN.n11865 0.025
R8173 VN.t8 VN.n11805 0.025
R8174 VN.t8 VN.n11794 0.025
R8175 VN.t8 VN.n11662 0.025
R8176 VN.n11689 VN.n11688 0.024
R8177 VN.n178 VN.n177 0.024
R8178 VN.n2183 VN.n2178 0.024
R8179 VN.n2905 VN.n2900 0.024
R8180 VN.n3645 VN.n3640 0.024
R8181 VN.n4402 VN.n4397 0.024
R8182 VN.n5177 VN.n5172 0.024
R8183 VN.n5969 VN.n5964 0.024
R8184 VN.n7212 VN.n7207 0.024
R8185 VN.n7601 VN.n7596 0.024
R8186 VN.n8446 VN.n8441 0.024
R8187 VN.n9308 VN.n9303 0.024
R8188 VN.n10191 VN.n10186 0.024
R8189 VN.n10242 VN.n10219 0.024
R8190 VN.n9359 VN.n9336 0.024
R8191 VN.n8497 VN.n8474 0.024
R8192 VN.n7652 VN.n7629 0.024
R8193 VN.n7263 VN.n7240 0.024
R8194 VN.n6020 VN.n5997 0.024
R8195 VN.n5228 VN.n5205 0.024
R8196 VN.n4453 VN.n4430 0.024
R8197 VN.n3696 VN.n3673 0.024
R8198 VN.n2956 VN.n2933 0.024
R8199 VN.n2234 VN.n2211 0.024
R8200 VN.n1526 VN.n1503 0.024
R8201 VN.n925 VN.n909 0.024
R8202 VN.n11441 VN.n11440 0.024
R8203 VN.n11414 VN.n11413 0.024
R8204 VN.n11067 VN.n11066 0.024
R8205 VN.n11523 VN.n11522 0.024
R8206 VN.n11688 VN.n11687 0.024
R8207 VN.n11910 VN.n11907 0.023
R8208 VN.n12026 VN.n12025 0.023
R8209 VN.n12027 VN.n12023 0.023
R8210 VN.n12049 VN.n12046 0.023
R8211 VN.n12079 VN.n12076 0.023
R8212 VN.n11413 VN.n11412 0.023
R8213 VN.t8 VN.n11689 0.023
R8214 VN.n476 VN.n475 0.023
R8215 VN.n909 VN.n908 0.023
R8216 VN.n1503 VN.n1502 0.023
R8217 VN.n2211 VN.n2210 0.023
R8218 VN.n2933 VN.n2932 0.023
R8219 VN.n3673 VN.n3672 0.023
R8220 VN.n4430 VN.n4429 0.023
R8221 VN.n5205 VN.n5204 0.023
R8222 VN.n5997 VN.n5996 0.023
R8223 VN.n7240 VN.n7239 0.023
R8224 VN.n7629 VN.n7628 0.023
R8225 VN.n8474 VN.n8473 0.023
R8226 VN.n9336 VN.n9335 0.023
R8227 VN.n10219 VN.n10218 0.023
R8228 VN.n10242 VN.n10223 0.023
R8229 VN.n9359 VN.n9340 0.023
R8230 VN.n8497 VN.n8478 0.023
R8231 VN.n7652 VN.n7633 0.023
R8232 VN.n7263 VN.n7244 0.023
R8233 VN.n6020 VN.n6001 0.023
R8234 VN.n5228 VN.n5209 0.023
R8235 VN.n4453 VN.n4434 0.023
R8236 VN.n3696 VN.n3677 0.023
R8237 VN.n2956 VN.n2937 0.023
R8238 VN.n2234 VN.n2215 0.023
R8239 VN.n1526 VN.n1507 0.023
R8240 VN.n925 VN.n913 0.023
R8241 VN.n11394 VN.n11392 0.023
R8242 VN.n11440 VN.n11439 0.023
R8243 VN.n12139 VN.n12138 0.023
R8244 VN.n11441 VN.n11437 0.023
R8245 VN.n11414 VN.n11410 0.023
R8246 VN.n11981 VN.n11980 0.023
R8247 VN.n11982 VN.n11978 0.023
R8248 VN.n12004 VN.n12001 0.023
R8249 VN.n3779 VN.n3778 0.023
R8250 VN.n11936 VN.n11935 0.023
R8251 VN.n11937 VN.n11933 0.023
R8252 VN.n11959 VN.n11956 0.023
R8253 VN.n5311 VN.n5310 0.023
R8254 VN.n11920 VN.n11919 0.023
R8255 VN.n11922 VN.n11920 0.023
R8256 VN.n6599 VN.n6598 0.023
R8257 VN.n11887 VN.n11886 0.023
R8258 VN.n11888 VN.n11885 0.023
R8259 VN.n11629 VN.n11628 0.023
R8260 VN.n11630 VN.n11626 0.023
R8261 VN.n11652 VN.n11649 0.023
R8262 VN.n11584 VN.n11583 0.023
R8263 VN.n11585 VN.n11581 0.023
R8264 VN.n11607 VN.n11604 0.023
R8265 VN.n11559 VN.n11555 0.023
R8266 VN.n80 VN.n78 0.023
R8267 VN.n10725 VN.n10723 0.023
R8268 VN.n11521 VN.n11520 0.023
R8269 VN.n10705 VN.n10703 0.023
R8270 VN.n9834 VN.n9833 0.023
R8271 VN.n9825 VN.n9823 0.023
R8272 VN.n8988 VN.n8987 0.023
R8273 VN.n8979 VN.n8977 0.023
R8274 VN.n8155 VN.n8154 0.023
R8275 VN.n8146 VN.n8144 0.023
R8276 VN.n7344 VN.n7343 0.023
R8277 VN.n7335 VN.n7333 0.023
R8278 VN.n6551 VN.n6550 0.023
R8279 VN.n6542 VN.n6540 0.023
R8280 VN.n5775 VN.n5774 0.023
R8281 VN.n5766 VN.n5764 0.023
R8282 VN.n5012 VN.n5011 0.023
R8283 VN.n5003 VN.n5001 0.023
R8284 VN.n4271 VN.n4270 0.023
R8285 VN.n4262 VN.n4260 0.023
R8286 VN.n3543 VN.n3542 0.023
R8287 VN.n3534 VN.n3532 0.023
R8288 VN.n2837 VN.n2836 0.023
R8289 VN.n2828 VN.n2826 0.023
R8290 VN.n2144 VN.n2143 0.023
R8291 VN.n2135 VN.n2133 0.023
R8292 VN.n1470 VN.n1469 0.023
R8293 VN.n1461 VN.n1459 0.023
R8294 VN.n31 VN.n20 0.023
R8295 VN.n12730 VN.n12729 0.023
R8296 VN.n197 VN.n185 0.023
R8297 VN.n98 VN.n87 0.023
R8298 VN.n2178 VN.n2175 0.023
R8299 VN.n2900 VN.n2897 0.023
R8300 VN.n3640 VN.n3637 0.023
R8301 VN.n4397 VN.n4395 0.023
R8302 VN.n5172 VN.n5169 0.023
R8303 VN.n5964 VN.n5962 0.023
R8304 VN.n7207 VN.n7204 0.023
R8305 VN.n7596 VN.n7593 0.023
R8306 VN.n8441 VN.n8438 0.023
R8307 VN.n9303 VN.n9300 0.023
R8308 VN.n10186 VN.n10184 0.023
R8309 VN.n11066 VN.n11064 0.023
R8310 VN.n11058 VN.n11057 0.023
R8311 VN.n12257 VN.n12256 0.022
R8312 VN.n11057 VN.n11056 0.022
R8313 VN.n1521 VN.n1517 0.022
R8314 VN.n2229 VN.n2225 0.022
R8315 VN.n2951 VN.n2947 0.022
R8316 VN.n3691 VN.n3687 0.022
R8317 VN.n4448 VN.n4444 0.022
R8318 VN.n5223 VN.n5219 0.022
R8319 VN.n6015 VN.n6011 0.022
R8320 VN.n7258 VN.n7254 0.022
R8321 VN.n7647 VN.n7643 0.022
R8322 VN.n8492 VN.n8488 0.022
R8323 VN.n9354 VN.n9350 0.022
R8324 VN.n10237 VN.n10233 0.022
R8325 VN.n11082 VN.n11078 0.022
R8326 VN.n12093 VN.n12089 0.022
R8327 VN.n238 VN.n237 0.022
R8328 VN.n9841 VN.n9839 0.022
R8329 VN.n8995 VN.n8993 0.022
R8330 VN.n8162 VN.n8160 0.022
R8331 VN.n7351 VN.n7349 0.022
R8332 VN.n6558 VN.n6556 0.022
R8333 VN.n5782 VN.n5780 0.022
R8334 VN.n5019 VN.n5017 0.022
R8335 VN.n4278 VN.n4276 0.022
R8336 VN.n3550 VN.n3548 0.022
R8337 VN.n2844 VN.n2842 0.022
R8338 VN.n2151 VN.n2149 0.022
R8339 VN.n1477 VN.n1475 0.022
R8340 VN.n1610 VN.n1609 0.022
R8341 VN.n2299 VN.n2297 0.022
R8342 VN.n3037 VN.n3036 0.022
R8343 VN.n3761 VN.n3759 0.022
R8344 VN.n4534 VN.n4533 0.022
R8345 VN.n5293 VN.n5291 0.022
R8346 VN.n6101 VN.n6100 0.022
R8347 VN.n6587 VN.n6586 0.022
R8348 VN.n7733 VN.n7732 0.022
R8349 VN.n8562 VN.n8560 0.022
R8350 VN.n9440 VN.n9439 0.022
R8351 VN.n10307 VN.n10305 0.022
R8352 VN.n11487 VN.n11486 0.022
R8353 VN.n11553 VN.n11552 0.022
R8354 VN.n242 VN.n241 0.022
R8355 VN.n12252 VN.n12247 0.021
R8356 VN.n12405 VN.n12404 0.021
R8357 VN.n12160 VN.n12159 0.021
R8358 VN.n11460 VN.n11459 0.021
R8359 VN.n10292 VN.n10291 0.021
R8360 VN.n10288 VN.n10287 0.021
R8361 VN.n9409 VN.n9408 0.021
R8362 VN.n9405 VN.n9404 0.021
R8363 VN.n8547 VN.n8546 0.021
R8364 VN.n8543 VN.n8542 0.021
R8365 VN.n7702 VN.n7701 0.021
R8366 VN.n7698 VN.n7697 0.021
R8367 VN.n7313 VN.n7312 0.021
R8368 VN.n7309 VN.n7308 0.021
R8369 VN.n6070 VN.n6069 0.021
R8370 VN.n6066 VN.n6065 0.021
R8371 VN.n5278 VN.n5277 0.021
R8372 VN.n5274 VN.n5273 0.021
R8373 VN.n4503 VN.n4502 0.021
R8374 VN.n4499 VN.n4498 0.021
R8375 VN.n3746 VN.n3745 0.021
R8376 VN.n3742 VN.n3741 0.021
R8377 VN.n3006 VN.n3005 0.021
R8378 VN.n3002 VN.n3001 0.021
R8379 VN.n2284 VN.n2283 0.021
R8380 VN.n2280 VN.n2279 0.021
R8381 VN.n1576 VN.n1575 0.021
R8382 VN.n1572 VN.n1571 0.021
R8383 VN.n893 VN.n892 0.021
R8384 VN.n889 VN.n888 0.021
R8385 VN.n222 VN.n221 0.021
R8386 VN.n218 VN.n217 0.021
R8387 VN.n12251 VN.n12250 0.021
R8388 VN.n10204 VN.n10203 0.021
R8389 VN.n10200 VN.n10199 0.021
R8390 VN.n9321 VN.n9320 0.021
R8391 VN.n9317 VN.n9316 0.021
R8392 VN.n8459 VN.n8458 0.021
R8393 VN.n8455 VN.n8454 0.021
R8394 VN.n7614 VN.n7613 0.021
R8395 VN.n7610 VN.n7609 0.021
R8396 VN.n7225 VN.n7224 0.021
R8397 VN.n7221 VN.n7220 0.021
R8398 VN.n5982 VN.n5981 0.021
R8399 VN.n5978 VN.n5977 0.021
R8400 VN.n5190 VN.n5189 0.021
R8401 VN.n5186 VN.n5185 0.021
R8402 VN.n4415 VN.n4414 0.021
R8403 VN.n4411 VN.n4410 0.021
R8404 VN.n3658 VN.n3657 0.021
R8405 VN.n3654 VN.n3653 0.021
R8406 VN.n2918 VN.n2917 0.021
R8407 VN.n2914 VN.n2913 0.021
R8408 VN.n2196 VN.n2195 0.021
R8409 VN.n2192 VN.n2191 0.021
R8410 VN.n1604 VN.n1603 0.021
R8411 VN.n10140 VN.n10139 0.021
R8412 VN.n10136 VN.n10135 0.021
R8413 VN.n9258 VN.n9257 0.021
R8414 VN.n9254 VN.n9253 0.021
R8415 VN.n8396 VN.n8395 0.021
R8416 VN.n8392 VN.n8391 0.021
R8417 VN.n7551 VN.n7550 0.021
R8418 VN.n7547 VN.n7546 0.021
R8419 VN.n7162 VN.n7161 0.021
R8420 VN.n7158 VN.n7157 0.021
R8421 VN.n5919 VN.n5918 0.021
R8422 VN.n5915 VN.n5914 0.021
R8423 VN.n5127 VN.n5126 0.021
R8424 VN.n5123 VN.n5122 0.021
R8425 VN.n4352 VN.n4351 0.021
R8426 VN.n4348 VN.n4347 0.021
R8427 VN.n3595 VN.n3594 0.021
R8428 VN.n3591 VN.n3590 0.021
R8429 VN.n3031 VN.n3030 0.021
R8430 VN.n10077 VN.n10076 0.021
R8431 VN.n10073 VN.n10072 0.021
R8432 VN.n9195 VN.n9194 0.021
R8433 VN.n9191 VN.n9190 0.021
R8434 VN.n8333 VN.n8332 0.021
R8435 VN.n8329 VN.n8328 0.021
R8436 VN.n7488 VN.n7487 0.021
R8437 VN.n7484 VN.n7483 0.021
R8438 VN.n7099 VN.n7098 0.021
R8439 VN.n7095 VN.n7094 0.021
R8440 VN.n5856 VN.n5855 0.021
R8441 VN.n5852 VN.n5851 0.021
R8442 VN.n5064 VN.n5063 0.021
R8443 VN.n5060 VN.n5059 0.021
R8444 VN.n4528 VN.n4527 0.021
R8445 VN.n10014 VN.n10013 0.021
R8446 VN.n10010 VN.n10009 0.021
R8447 VN.n9132 VN.n9131 0.021
R8448 VN.n9128 VN.n9127 0.021
R8449 VN.n8270 VN.n8269 0.021
R8450 VN.n8266 VN.n8265 0.021
R8451 VN.n7425 VN.n7424 0.021
R8452 VN.n7421 VN.n7420 0.021
R8453 VN.n7036 VN.n7035 0.021
R8454 VN.n7032 VN.n7031 0.021
R8455 VN.n6095 VN.n6094 0.021
R8456 VN.n9951 VN.n9950 0.021
R8457 VN.n9947 VN.n9946 0.021
R8458 VN.n9069 VN.n9068 0.021
R8459 VN.n9065 VN.n9064 0.021
R8460 VN.n8207 VN.n8206 0.021
R8461 VN.n8203 VN.n8202 0.021
R8462 VN.n7727 VN.n7726 0.021
R8463 VN.n9888 VN.n9887 0.021
R8464 VN.n9884 VN.n9883 0.021
R8465 VN.n9434 VN.n9433 0.021
R8466 VN.n479 VN.n478 0.021
R8467 VN.n203 VN.n202 0.021
R8468 VN.n874 VN.n873 0.021
R8469 VN.n1557 VN.n1556 0.021
R8470 VN.n2265 VN.n2264 0.021
R8471 VN.n2987 VN.n2986 0.021
R8472 VN.n3727 VN.n3726 0.021
R8473 VN.n4484 VN.n4483 0.021
R8474 VN.n5259 VN.n5258 0.021
R8475 VN.n6051 VN.n6050 0.021
R8476 VN.n7294 VN.n7293 0.021
R8477 VN.n7683 VN.n7682 0.021
R8478 VN.n8528 VN.n8527 0.021
R8479 VN.n9390 VN.n9389 0.021
R8480 VN.n10273 VN.n10272 0.021
R8481 VN.n12164 VN.n12163 0.021
R8482 VN.n3576 VN.n3575 0.021
R8483 VN.n4333 VN.n4332 0.021
R8484 VN.n5108 VN.n5107 0.021
R8485 VN.n5900 VN.n5899 0.021
R8486 VN.n7143 VN.n7142 0.021
R8487 VN.n7532 VN.n7531 0.021
R8488 VN.n8377 VN.n8376 0.021
R8489 VN.n9239 VN.n9238 0.021
R8490 VN.n10121 VN.n10120 0.021
R8491 VN.n10990 VN.n10989 0.021
R8492 VN.n1611 VN.n1610 0.021
R8493 VN.n924 VN.n923 0.021
R8494 VN.n10170 VN.n10169 0.021
R8495 VN.n9288 VN.n9287 0.021
R8496 VN.n8426 VN.n8425 0.021
R8497 VN.n7581 VN.n7580 0.021
R8498 VN.n7192 VN.n7191 0.021
R8499 VN.n5949 VN.n5948 0.021
R8500 VN.n5157 VN.n5156 0.021
R8501 VN.n4382 VN.n4381 0.021
R8502 VN.n3625 VN.n3624 0.021
R8503 VN.n2885 VN.n2884 0.021
R8504 VN.n2301 VN.n2299 0.021
R8505 VN.n12044 VN.n12043 0.021
R8506 VN.n3038 VN.n3037 0.021
R8507 VN.n5045 VN.n5044 0.021
R8508 VN.n5837 VN.n5836 0.021
R8509 VN.n7080 VN.n7079 0.021
R8510 VN.n7469 VN.n7468 0.021
R8511 VN.n8314 VN.n8313 0.021
R8512 VN.n9176 VN.n9175 0.021
R8513 VN.n10058 VN.n10057 0.021
R8514 VN.n10932 VN.n10931 0.021
R8515 VN.n10976 VN.n10975 0.021
R8516 VN.n10107 VN.n10106 0.021
R8517 VN.n9225 VN.n9224 0.021
R8518 VN.n8363 VN.n8362 0.021
R8519 VN.n7518 VN.n7517 0.021
R8520 VN.n7129 VN.n7128 0.021
R8521 VN.n5886 VN.n5885 0.021
R8522 VN.n5094 VN.n5093 0.021
R8523 VN.n4319 VN.n4318 0.021
R8524 VN.n3763 VN.n3761 0.021
R8525 VN.n11999 VN.n11998 0.021
R8526 VN.n4535 VN.n4534 0.021
R8527 VN.n7017 VN.n7016 0.021
R8528 VN.n7406 VN.n7405 0.021
R8529 VN.n8251 VN.n8250 0.021
R8530 VN.n9113 VN.n9112 0.021
R8531 VN.n9995 VN.n9994 0.021
R8532 VN.n10874 VN.n10873 0.021
R8533 VN.n10918 VN.n10917 0.021
R8534 VN.n10044 VN.n10043 0.021
R8535 VN.n9162 VN.n9161 0.021
R8536 VN.n8300 VN.n8299 0.021
R8537 VN.n7455 VN.n7454 0.021
R8538 VN.n7066 VN.n7065 0.021
R8539 VN.n5823 VN.n5822 0.021
R8540 VN.n5295 VN.n5293 0.021
R8541 VN.n11954 VN.n11953 0.021
R8542 VN.n6102 VN.n6101 0.021
R8543 VN.n10860 VN.n10859 0.021
R8544 VN.n9981 VN.n9980 0.021
R8545 VN.n9099 VN.n9098 0.021
R8546 VN.n8237 VN.n8236 0.021
R8547 VN.n7392 VN.n7391 0.021
R8548 VN.n6589 VN.n6587 0.021
R8549 VN.n8188 VN.n8187 0.021
R8550 VN.n9050 VN.n9049 0.021
R8551 VN.n9932 VN.n9931 0.021
R8552 VN.n10816 VN.n10815 0.021
R8553 VN.n7734 VN.n7733 0.021
R8554 VN.n9869 VN.n9868 0.021
R8555 VN.n10758 VN.n10757 0.021
R8556 VN.n10802 VN.n10801 0.021
R8557 VN.n9918 VN.n9917 0.021
R8558 VN.n9036 VN.n9035 0.021
R8559 VN.n8564 VN.n8562 0.021
R8560 VN.n11647 VN.n11646 0.021
R8561 VN.n9441 VN.n9440 0.021
R8562 VN.n10744 VN.n10743 0.021
R8563 VN.n10309 VN.n10307 0.021
R8564 VN.n11602 VN.n11601 0.021
R8565 VN.n11488 VN.n11487 0.021
R8566 VN.n11554 VN.n11553 0.021
R8567 VN.n76 VN.n74 0.021
R8568 VN.n11905 VN.n11904 0.021
R8569 VN.n825 VN.n824 0.021
R8570 VN.n30 VN.n21 0.02
R8571 VN.n97 VN.n96 0.02
R8572 VN.n12223 VN.n12222 0.02
R8573 VN.n12258 VN.n12255 0.02
R8574 VN.n2178 VN.n2177 0.02
R8575 VN.n2900 VN.n2899 0.02
R8576 VN.n3640 VN.n3639 0.02
R8577 VN.n4397 VN.n4396 0.02
R8578 VN.n5172 VN.n5171 0.02
R8579 VN.n5964 VN.n5963 0.02
R8580 VN.n7207 VN.n7206 0.02
R8581 VN.n7596 VN.n7595 0.02
R8582 VN.n8441 VN.n8440 0.02
R8583 VN.n9303 VN.n9302 0.02
R8584 VN.n10186 VN.n10185 0.02
R8585 VN.n1611 VN.n1607 0.02
R8586 VN.n239 VN.n236 0.02
R8587 VN.n11066 VN.n11065 0.02
R8588 VN.n2301 VN.n2300 0.02
R8589 VN.n3038 VN.n3034 0.02
R8590 VN.n3763 VN.n3762 0.02
R8591 VN.n4535 VN.n4531 0.02
R8592 VN.n5295 VN.n5294 0.02
R8593 VN.n6102 VN.n6098 0.02
R8594 VN.n7734 VN.n7730 0.02
R8595 VN.n8564 VN.n8563 0.02
R8596 VN.n9441 VN.n9437 0.02
R8597 VN.n10309 VN.n10308 0.02
R8598 VN.n11488 VN.n11484 0.02
R8599 VN.n11554 VN.n11550 0.02
R8600 VN.n6589 VN.n6588 0.02
R8601 VN.n12143 VN.n12142 0.02
R8602 VN.t8 VN.n11701 0.019
R8603 VN.n10580 VN.n10578 0.019
R8604 VN.n9695 VN.n9693 0.019
R8605 VN.n8833 VN.n8831 0.019
R8606 VN.n7984 VN.n7982 0.019
R8607 VN.n6793 VN.n6791 0.019
R8608 VN.n6348 VN.n6346 0.019
R8609 VN.n5556 VN.n5554 0.019
R8610 VN.n4777 VN.n4775 0.019
R8611 VN.n4020 VN.n4018 0.019
R8612 VN.n3276 VN.n3274 0.019
R8613 VN.n2554 VN.n2552 0.019
R8614 VN.n1845 VN.n1843 0.019
R8615 VN.n1155 VN.n1153 0.019
R8616 VN.n12100 VN.n12099 0.019
R8617 VN.n10600 VN.n10599 0.019
R8618 VN.n1525 VN.n1524 0.019
R8619 VN.n2233 VN.n2232 0.019
R8620 VN.n2955 VN.n2954 0.019
R8621 VN.n3695 VN.n3694 0.019
R8622 VN.n4452 VN.n4451 0.019
R8623 VN.n5227 VN.n5226 0.019
R8624 VN.n6019 VN.n6018 0.019
R8625 VN.n7262 VN.n7261 0.019
R8626 VN.n7651 VN.n7650 0.019
R8627 VN.n8496 VN.n8495 0.019
R8628 VN.n9358 VN.n9357 0.019
R8629 VN.n10241 VN.n10240 0.019
R8630 VN.n11086 VN.n11085 0.019
R8631 VN.n12747 VN.n12746 0.019
R8632 VN.n12112 VN.n12111 0.018
R8633 VN.n12023 VN.n12021 0.018
R8634 VN.n12046 VN.n12045 0.018
R8635 VN.n11978 VN.n11976 0.018
R8636 VN.n12001 VN.n12000 0.018
R8637 VN.n11933 VN.n11931 0.018
R8638 VN.n11956 VN.n11955 0.018
R8639 VN.n11885 VN.n11883 0.018
R8640 VN.n11626 VN.n11624 0.018
R8641 VN.n11649 VN.n11648 0.018
R8642 VN.n11581 VN.n11579 0.018
R8643 VN.n11604 VN.n11603 0.018
R8644 VN.n751 VN.n750 0.018
R8645 VN.n11907 VN.n11906 0.018
R8646 VN.n11695 VN.n11694 0.018
R8647 VN.n2177 VN.n2176 0.018
R8648 VN.n2899 VN.n2898 0.018
R8649 VN.n3639 VN.n3638 0.018
R8650 VN.n5171 VN.n5170 0.018
R8651 VN.n7206 VN.n7205 0.018
R8652 VN.n7595 VN.n7594 0.018
R8653 VN.n8440 VN.n8439 0.018
R8654 VN.n9302 VN.n9301 0.018
R8655 VN.n749 VN.n748 0.017
R8656 VN.n12373 VN.n12372 0.017
R8657 VN.n12398 VN.n12397 0.017
R8658 VN.n755 VN.n752 0.017
R8659 VN.n9844 VN.n9843 0.017
R8660 VN.n8998 VN.n8997 0.017
R8661 VN.n8165 VN.n8164 0.017
R8662 VN.n7354 VN.n7353 0.017
R8663 VN.n6561 VN.n6560 0.017
R8664 VN.n5785 VN.n5784 0.017
R8665 VN.n5022 VN.n5021 0.017
R8666 VN.n4281 VN.n4280 0.017
R8667 VN.n3553 VN.n3552 0.017
R8668 VN.n2847 VN.n2846 0.017
R8669 VN.n2154 VN.n2153 0.017
R8670 VN.n1480 VN.n1479 0.017
R8671 VN.n11069 VN.n11058 0.016
R8672 VN.n10566 VN.n10562 0.016
R8673 VN.n2320 VN.n2312 0.016
R8674 VN.n3782 VN.n3774 0.016
R8675 VN.n5314 VN.n5306 0.016
R8676 VN.t76 VN.n6594 0.016
R8677 VN.n8583 VN.n8575 0.016
R8678 VN.n10328 VN.n10320 0.016
R8679 VN.n9842 VN.n9841 0.016
R8680 VN.n8996 VN.n8995 0.016
R8681 VN.n8163 VN.n8162 0.016
R8682 VN.n7352 VN.n7351 0.016
R8683 VN.n6559 VN.n6558 0.016
R8684 VN.n5783 VN.n5782 0.016
R8685 VN.n5020 VN.n5019 0.016
R8686 VN.n4279 VN.n4278 0.016
R8687 VN.n3551 VN.n3550 0.016
R8688 VN.n2845 VN.n2844 0.016
R8689 VN.n2152 VN.n2151 0.016
R8690 VN.n1478 VN.n1477 0.016
R8691 VN.n4395 VN.n4394 0.015
R8692 VN.n5962 VN.n5961 0.015
R8693 VN.n10184 VN.n10183 0.015
R8694 VN.n11064 VN.n11063 0.015
R8695 VN.n13093 VN.n13092 0.015
R8696 VN.n782 VN.n781 0.015
R8697 VN.n11069 VN.n11068 0.015
R8698 VN.n12247 VN.n12246 0.015
R8699 VN.n1523 VN.n1522 0.015
R8700 VN.n1522 VN.n1521 0.015
R8701 VN.n1521 VN.n1520 0.015
R8702 VN.n2231 VN.n2230 0.015
R8703 VN.n2230 VN.n2229 0.015
R8704 VN.n2229 VN.n2228 0.015
R8705 VN.n2953 VN.n2952 0.015
R8706 VN.n2952 VN.n2951 0.015
R8707 VN.n2951 VN.n2950 0.015
R8708 VN.n3693 VN.n3692 0.015
R8709 VN.n3692 VN.n3691 0.015
R8710 VN.n3691 VN.n3690 0.015
R8711 VN.n4450 VN.n4449 0.015
R8712 VN.n4449 VN.n4448 0.015
R8713 VN.n4448 VN.n4447 0.015
R8714 VN.n5225 VN.n5224 0.015
R8715 VN.n5224 VN.n5223 0.015
R8716 VN.n5223 VN.n5222 0.015
R8717 VN.n6017 VN.n6016 0.015
R8718 VN.n6016 VN.n6015 0.015
R8719 VN.n6015 VN.n6014 0.015
R8720 VN.n7260 VN.n7259 0.015
R8721 VN.n7259 VN.n7258 0.015
R8722 VN.n7258 VN.n7257 0.015
R8723 VN.n7649 VN.n7648 0.015
R8724 VN.n7648 VN.n7647 0.015
R8725 VN.n7647 VN.n7646 0.015
R8726 VN.n8494 VN.n8493 0.015
R8727 VN.n8493 VN.n8492 0.015
R8728 VN.n8492 VN.n8491 0.015
R8729 VN.n9356 VN.n9355 0.015
R8730 VN.n9355 VN.n9354 0.015
R8731 VN.n9354 VN.n9353 0.015
R8732 VN.n10239 VN.n10238 0.015
R8733 VN.n10238 VN.n10237 0.015
R8734 VN.n10237 VN.n10236 0.015
R8735 VN.n11084 VN.n11083 0.015
R8736 VN.n11083 VN.n11082 0.015
R8737 VN.n11082 VN.n11081 0.015
R8738 VN.n12094 VN.n12093 0.015
R8739 VN.n12093 VN.n12092 0.015
R8740 VN.n241 VN.n240 0.015
R8741 VN.n12141 VN.n12140 0.015
R8742 VN.t51 VN.n80 0.015
R8743 VN.n10707 VN.n9863 0.015
R8744 VN.n9827 VN.n9015 0.015
R8745 VN.n8981 VN.n8182 0.015
R8746 VN.n8148 VN.n7371 0.015
R8747 VN.n7337 VN.n6578 0.015
R8748 VN.n6544 VN.n5802 0.015
R8749 VN.n5768 VN.n5039 0.015
R8750 VN.n5005 VN.n4298 0.015
R8751 VN.n4264 VN.n3570 0.015
R8752 VN.n3536 VN.n2864 0.015
R8753 VN.n2830 VN.n2171 0.015
R8754 VN.n2137 VN.n1497 0.015
R8755 VN.n13092 VN.n13091 0.015
R8756 VN.n781 VN.n780 0.015
R8757 VN.n1463 VN.n847 0.015
R8758 VN.n9848 VN.n9847 0.015
R8759 VN.n13119 VN.n13118 0.015
R8760 VN.n9846 VN.n9845 0.015
R8761 VN.n13121 VN.n13120 0.015
R8762 VN.n206 VN.n205 0.015
R8763 VN.n877 VN.n876 0.015
R8764 VN.n1560 VN.n1559 0.015
R8765 VN.n2268 VN.n2267 0.015
R8766 VN.n2990 VN.n2989 0.015
R8767 VN.n3730 VN.n3729 0.015
R8768 VN.n4487 VN.n4486 0.015
R8769 VN.n5262 VN.n5261 0.015
R8770 VN.n6054 VN.n6053 0.015
R8771 VN.n7297 VN.n7296 0.015
R8772 VN.n7686 VN.n7685 0.015
R8773 VN.n8531 VN.n8530 0.015
R8774 VN.n9393 VN.n9392 0.015
R8775 VN.n10276 VN.n10275 0.015
R8776 VN.n3579 VN.n3578 0.015
R8777 VN.n4336 VN.n4335 0.015
R8778 VN.n5111 VN.n5110 0.015
R8779 VN.n5903 VN.n5902 0.015
R8780 VN.n7146 VN.n7145 0.015
R8781 VN.n7535 VN.n7534 0.015
R8782 VN.n8380 VN.n8379 0.015
R8783 VN.n9242 VN.n9241 0.015
R8784 VN.n10124 VN.n10123 0.015
R8785 VN.n10993 VN.n10992 0.015
R8786 VN.n2880 VN.n2879 0.015
R8787 VN.n3620 VN.n3619 0.015
R8788 VN.n4377 VN.n4376 0.015
R8789 VN.n5152 VN.n5151 0.015
R8790 VN.n5944 VN.n5943 0.015
R8791 VN.n7187 VN.n7186 0.015
R8792 VN.n7576 VN.n7575 0.015
R8793 VN.n8421 VN.n8420 0.015
R8794 VN.n9283 VN.n9282 0.015
R8795 VN.n10165 VN.n10164 0.015
R8796 VN.n11029 VN.n11028 0.015
R8797 VN.n5048 VN.n5047 0.015
R8798 VN.n5840 VN.n5839 0.015
R8799 VN.n7083 VN.n7082 0.015
R8800 VN.n7472 VN.n7471 0.015
R8801 VN.n8317 VN.n8316 0.015
R8802 VN.n9179 VN.n9178 0.015
R8803 VN.n10061 VN.n10060 0.015
R8804 VN.n10935 VN.n10934 0.015
R8805 VN.n4314 VN.n4313 0.015
R8806 VN.n5089 VN.n5088 0.015
R8807 VN.n5881 VN.n5880 0.015
R8808 VN.n7124 VN.n7123 0.015
R8809 VN.n7513 VN.n7512 0.015
R8810 VN.n8358 VN.n8357 0.015
R8811 VN.n9220 VN.n9219 0.015
R8812 VN.n10102 VN.n10101 0.015
R8813 VN.n10971 VN.n10970 0.015
R8814 VN.n7020 VN.n7019 0.015
R8815 VN.n7409 VN.n7408 0.015
R8816 VN.n8254 VN.n8253 0.015
R8817 VN.n9116 VN.n9115 0.015
R8818 VN.n9998 VN.n9997 0.015
R8819 VN.n10877 VN.n10876 0.015
R8820 VN.n5818 VN.n5817 0.015
R8821 VN.n7061 VN.n7060 0.015
R8822 VN.n7450 VN.n7449 0.015
R8823 VN.n8295 VN.n8294 0.015
R8824 VN.n9157 VN.n9156 0.015
R8825 VN.n10039 VN.n10038 0.015
R8826 VN.n10913 VN.n10912 0.015
R8827 VN.n7387 VN.n7386 0.015
R8828 VN.n8232 VN.n8231 0.015
R8829 VN.n9094 VN.n9093 0.015
R8830 VN.n9976 VN.n9975 0.015
R8831 VN.n10855 VN.n10854 0.015
R8832 VN.n8191 VN.n8190 0.015
R8833 VN.n9053 VN.n9052 0.015
R8834 VN.n9935 VN.n9934 0.015
R8835 VN.n10819 VN.n10818 0.015
R8836 VN.n9872 VN.n9871 0.015
R8837 VN.n10761 VN.n10760 0.015
R8838 VN.n9031 VN.n9030 0.015
R8839 VN.n9913 VN.n9912 0.015
R8840 VN.n10797 VN.n10796 0.015
R8841 VN.n10739 VN.n10738 0.015
R8842 VN.n12097 VN.n12096 0.014
R8843 VN.n828 VN.n826 0.014
R8844 VN.n10173 VN.n10172 0.014
R8845 VN.n9291 VN.n9290 0.014
R8846 VN.n8429 VN.n8428 0.014
R8847 VN.n7584 VN.n7583 0.014
R8848 VN.n7195 VN.n7194 0.014
R8849 VN.n5952 VN.n5951 0.014
R8850 VN.n5160 VN.n5159 0.014
R8851 VN.n4385 VN.n4384 0.014
R8852 VN.n3628 VN.n3627 0.014
R8853 VN.n2888 VN.n2887 0.014
R8854 VN.n10110 VN.n10109 0.014
R8855 VN.n9228 VN.n9227 0.014
R8856 VN.n8366 VN.n8365 0.014
R8857 VN.n7521 VN.n7520 0.014
R8858 VN.n7132 VN.n7131 0.014
R8859 VN.n5889 VN.n5888 0.014
R8860 VN.n5097 VN.n5096 0.014
R8861 VN.n4322 VN.n4321 0.014
R8862 VN.n10047 VN.n10046 0.014
R8863 VN.n9165 VN.n9164 0.014
R8864 VN.n8303 VN.n8302 0.014
R8865 VN.n7458 VN.n7457 0.014
R8866 VN.n7069 VN.n7068 0.014
R8867 VN.n5826 VN.n5825 0.014
R8868 VN.n10863 VN.n10862 0.014
R8869 VN.n9984 VN.n9983 0.014
R8870 VN.n9102 VN.n9101 0.014
R8871 VN.n8240 VN.n8239 0.014
R8872 VN.n7395 VN.n7394 0.014
R8873 VN.n9921 VN.n9920 0.014
R8874 VN.n9039 VN.n9038 0.014
R8875 VN.n13104 VN.n13095 0.014
R8876 VN.n794 VN.n784 0.014
R8877 VN.n11068 VN.n11067 0.014
R8878 VN.n10544 VN.n10543 0.014
R8879 VN.n9778 VN.n9777 0.014
R8880 VN.n8932 VN.n8931 0.014
R8881 VN.n8099 VN.n8098 0.014
R8882 VN.n6924 VN.n6923 0.014
R8883 VN.n6495 VN.n6494 0.014
R8884 VN.n5719 VN.n5718 0.014
R8885 VN.n4956 VN.n4955 0.014
R8886 VN.n4215 VN.n4214 0.014
R8887 VN.n3487 VN.n3486 0.014
R8888 VN.n2781 VN.n2780 0.014
R8889 VN.n2088 VN.n2087 0.014
R8890 VN.n1414 VN.n1413 0.014
R8891 VN.n12736 VN.n12735 0.014
R8892 VN.n210 VN.n209 0.013
R8893 VN.n881 VN.n880 0.013
R8894 VN.n1564 VN.n1563 0.013
R8895 VN.n2272 VN.n2271 0.013
R8896 VN.n2994 VN.n2993 0.013
R8897 VN.n3734 VN.n3733 0.013
R8898 VN.n4491 VN.n4490 0.013
R8899 VN.n5266 VN.n5265 0.013
R8900 VN.n6058 VN.n6057 0.013
R8901 VN.n7301 VN.n7300 0.013
R8902 VN.n7690 VN.n7689 0.013
R8903 VN.n8535 VN.n8534 0.013
R8904 VN.n9397 VN.n9396 0.013
R8905 VN.n10280 VN.n10279 0.013
R8906 VN.n3583 VN.n3582 0.013
R8907 VN.n4340 VN.n4339 0.013
R8908 VN.n5115 VN.n5114 0.013
R8909 VN.n5907 VN.n5906 0.013
R8910 VN.n7150 VN.n7149 0.013
R8911 VN.n7539 VN.n7538 0.013
R8912 VN.n8384 VN.n8383 0.013
R8913 VN.n9246 VN.n9245 0.013
R8914 VN.n10128 VN.n10127 0.013
R8915 VN.n10997 VN.n10996 0.013
R8916 VN.n11035 VN.n11034 0.013
R8917 VN.n5052 VN.n5051 0.013
R8918 VN.n5844 VN.n5843 0.013
R8919 VN.n7087 VN.n7086 0.013
R8920 VN.n7476 VN.n7475 0.013
R8921 VN.n8321 VN.n8320 0.013
R8922 VN.n9183 VN.n9182 0.013
R8923 VN.n10065 VN.n10064 0.013
R8924 VN.n10939 VN.n10938 0.013
R8925 VN.n10979 VN.n10978 0.013
R8926 VN.n7024 VN.n7023 0.013
R8927 VN.n7413 VN.n7412 0.013
R8928 VN.n8258 VN.n8257 0.013
R8929 VN.n9120 VN.n9119 0.013
R8930 VN.n10002 VN.n10001 0.013
R8931 VN.n10881 VN.n10880 0.013
R8932 VN.n10921 VN.n10920 0.013
R8933 VN.n8195 VN.n8194 0.013
R8934 VN.n9057 VN.n9056 0.013
R8935 VN.n9939 VN.n9938 0.013
R8936 VN.n10823 VN.n10822 0.013
R8937 VN.n9876 VN.n9875 0.013
R8938 VN.n10765 VN.n10764 0.013
R8939 VN.n10805 VN.n10804 0.013
R8940 VN.n10747 VN.n10746 0.013
R8941 VN.n922 VN.n921 0.013
R8942 VN.n11786 VN.n11785 0.013
R8943 VN.n11784 VN.n11783 0.013
R8944 VN.n9777 VN.n9776 0.013
R8945 VN.n8931 VN.n8930 0.013
R8946 VN.n8098 VN.n8097 0.013
R8947 VN.n6923 VN.n6922 0.013
R8948 VN.n6494 VN.n6493 0.013
R8949 VN.n5718 VN.n5717 0.013
R8950 VN.n4955 VN.n4954 0.013
R8951 VN.n4214 VN.n4213 0.013
R8952 VN.n3486 VN.n3485 0.013
R8953 VN.n2780 VN.n2779 0.013
R8954 VN.n2087 VN.n2086 0.013
R8955 VN.n1413 VN.n1412 0.013
R8956 VN.n12735 VN.n12734 0.013
R8957 VN.t8 VN.n11836 0.012
R8958 VN.t8 VN.n11825 0.012
R8959 VN.t8 VN.n11814 0.012
R8960 VN.t8 VN.n11866 0.012
R8961 VN.t8 VN.n11803 0.012
R8962 VN.t8 VN.n11792 0.012
R8963 VN.t8 VN.n11663 0.012
R8964 VN.t8 VN.n11656 0.012
R8965 VN.n847 VN.n830 0.012
R8966 VN.n207 VN.n206 0.012
R8967 VN.n878 VN.n877 0.012
R8968 VN.n1561 VN.n1560 0.012
R8969 VN.n2269 VN.n2268 0.012
R8970 VN.n2991 VN.n2990 0.012
R8971 VN.n3731 VN.n3730 0.012
R8972 VN.n4488 VN.n4487 0.012
R8973 VN.n5263 VN.n5262 0.012
R8974 VN.n6055 VN.n6054 0.012
R8975 VN.n7298 VN.n7297 0.012
R8976 VN.n7687 VN.n7686 0.012
R8977 VN.n8532 VN.n8531 0.012
R8978 VN.n9394 VN.n9393 0.012
R8979 VN.n10277 VN.n10276 0.012
R8980 VN.n12165 VN.n12162 0.012
R8981 VN.n3580 VN.n3579 0.012
R8982 VN.n4337 VN.n4336 0.012
R8983 VN.n5112 VN.n5111 0.012
R8984 VN.n5904 VN.n5903 0.012
R8985 VN.n7147 VN.n7146 0.012
R8986 VN.n7536 VN.n7535 0.012
R8987 VN.n8381 VN.n8380 0.012
R8988 VN.n9243 VN.n9242 0.012
R8989 VN.n10125 VN.n10124 0.012
R8990 VN.n10994 VN.n10993 0.012
R8991 VN.n2881 VN.n2880 0.012
R8992 VN.n3621 VN.n3620 0.012
R8993 VN.n4378 VN.n4377 0.012
R8994 VN.n5153 VN.n5152 0.012
R8995 VN.n5945 VN.n5944 0.012
R8996 VN.n7188 VN.n7187 0.012
R8997 VN.n7577 VN.n7576 0.012
R8998 VN.n8422 VN.n8421 0.012
R8999 VN.n9284 VN.n9283 0.012
R9000 VN.n10166 VN.n10165 0.012
R9001 VN.n11061 VN.n11060 0.012
R9002 VN.n2181 VN.n2180 0.012
R9003 VN.n2903 VN.n2902 0.012
R9004 VN.n3643 VN.n3642 0.012
R9005 VN.n4400 VN.n4399 0.012
R9006 VN.n5175 VN.n5174 0.012
R9007 VN.n5967 VN.n5966 0.012
R9008 VN.n7210 VN.n7209 0.012
R9009 VN.n7599 VN.n7598 0.012
R9010 VN.n8444 VN.n8443 0.012
R9011 VN.n9306 VN.n9305 0.012
R9012 VN.n10189 VN.n10188 0.012
R9013 VN.n11030 VN.n11029 0.012
R9014 VN.n12059 VN.n12049 0.012
R9015 VN.n5049 VN.n5048 0.012
R9016 VN.n5841 VN.n5840 0.012
R9017 VN.n7084 VN.n7083 0.012
R9018 VN.n7473 VN.n7472 0.012
R9019 VN.n8318 VN.n8317 0.012
R9020 VN.n9180 VN.n9179 0.012
R9021 VN.n10062 VN.n10061 0.012
R9022 VN.n10936 VN.n10935 0.012
R9023 VN.n4315 VN.n4314 0.012
R9024 VN.n5090 VN.n5089 0.012
R9025 VN.n5882 VN.n5881 0.012
R9026 VN.n7125 VN.n7124 0.012
R9027 VN.n7514 VN.n7513 0.012
R9028 VN.n8359 VN.n8358 0.012
R9029 VN.n9221 VN.n9220 0.012
R9030 VN.n10103 VN.n10102 0.012
R9031 VN.n10972 VN.n10971 0.012
R9032 VN.n12014 VN.n12004 0.012
R9033 VN.n7021 VN.n7020 0.012
R9034 VN.n7410 VN.n7409 0.012
R9035 VN.n8255 VN.n8254 0.012
R9036 VN.n9117 VN.n9116 0.012
R9037 VN.n9999 VN.n9998 0.012
R9038 VN.n10878 VN.n10877 0.012
R9039 VN.n5819 VN.n5818 0.012
R9040 VN.n7062 VN.n7061 0.012
R9041 VN.n7451 VN.n7450 0.012
R9042 VN.n8296 VN.n8295 0.012
R9043 VN.n9158 VN.n9157 0.012
R9044 VN.n10040 VN.n10039 0.012
R9045 VN.n10914 VN.n10913 0.012
R9046 VN.n11969 VN.n11959 0.012
R9047 VN.n7388 VN.n7387 0.012
R9048 VN.n8233 VN.n8232 0.012
R9049 VN.n9095 VN.n9094 0.012
R9050 VN.n9977 VN.n9976 0.012
R9051 VN.n10856 VN.n10855 0.012
R9052 VN.n8192 VN.n8191 0.012
R9053 VN.n9054 VN.n9053 0.012
R9054 VN.n9936 VN.n9935 0.012
R9055 VN.n10820 VN.n10819 0.012
R9056 VN.n9873 VN.n9872 0.012
R9057 VN.n10762 VN.n10761 0.012
R9058 VN.n9032 VN.n9031 0.012
R9059 VN.n9914 VN.n9913 0.012
R9060 VN.n10798 VN.n10797 0.012
R9061 VN.n11876 VN.n11652 0.012
R9062 VN.n10740 VN.n10739 0.012
R9063 VN.n11617 VN.n11607 0.012
R9064 VN.n9776 VN.n9775 0.012
R9065 VN.n9839 VN.n9838 0.012
R9066 VN.n8930 VN.n8929 0.012
R9067 VN.n8993 VN.n8992 0.012
R9068 VN.n8097 VN.n8096 0.012
R9069 VN.n8160 VN.n8159 0.012
R9070 VN.n6922 VN.n6921 0.012
R9071 VN.n7349 VN.n7348 0.012
R9072 VN.n6493 VN.n6492 0.012
R9073 VN.n6556 VN.n6555 0.012
R9074 VN.n5717 VN.n5716 0.012
R9075 VN.n5780 VN.n5779 0.012
R9076 VN.n4954 VN.n4953 0.012
R9077 VN.n5017 VN.n5016 0.012
R9078 VN.n4213 VN.n4212 0.012
R9079 VN.n4276 VN.n4275 0.012
R9080 VN.n3485 VN.n3484 0.012
R9081 VN.n3548 VN.n3547 0.012
R9082 VN.n2779 VN.n2778 0.012
R9083 VN.n2842 VN.n2841 0.012
R9084 VN.n2086 VN.n2085 0.012
R9085 VN.n2149 VN.n2148 0.012
R9086 VN.n1412 VN.n1411 0.012
R9087 VN.n1475 VN.n1474 0.012
R9088 VN.n28 VN.n27 0.012
R9089 VN.n12734 VN.n12733 0.012
R9090 VN.n192 VN.n191 0.012
R9091 VN.n94 VN.n93 0.012
R9092 VN.n11924 VN.n11910 0.012
R9093 VN.n12405 VN.n12396 0.012
R9094 VN.n12385 VN.n12376 0.011
R9095 VN.n755 VN.n749 0.01
R9096 VN.n11163 VN.n11162 0.01
R9097 VN.n11197 VN.n11196 0.01
R9098 VN.n11231 VN.n11230 0.01
R9099 VN.n11298 VN.n11297 0.01
R9100 VN.n11332 VN.n11331 0.01
R9101 VN.n1591 VN.n1590 0.01
R9102 VN.n12027 VN.n12026 0.01
R9103 VN.n12081 VN.n12079 0.01
R9104 VN.n10588 VN.n10580 0.01
R9105 VN.n9703 VN.n9695 0.01
R9106 VN.n8841 VN.n8833 0.01
R9107 VN.n7992 VN.n7984 0.01
R9108 VN.n6801 VN.n6793 0.01
R9109 VN.n6356 VN.n6348 0.01
R9110 VN.n5564 VN.n5556 0.01
R9111 VN.n4785 VN.n4777 0.01
R9112 VN.n4028 VN.n4020 0.01
R9113 VN.n3284 VN.n3276 0.01
R9114 VN.n2562 VN.n2554 0.01
R9115 VN.n1853 VN.n1845 0.01
R9116 VN.n1163 VN.n1155 0.01
R9117 VN.n11397 VN.n11394 0.01
R9118 VN.n507 VN.n504 0.01
R9119 VN.n1182 VN.n1179 0.01
R9120 VN.n1872 VN.n1869 0.01
R9121 VN.n2581 VN.n2578 0.01
R9122 VN.n3303 VN.n3300 0.01
R9123 VN.n4047 VN.n4044 0.01
R9124 VN.n4804 VN.n4801 0.01
R9125 VN.n5583 VN.n5580 0.01
R9126 VN.n6375 VN.n6372 0.01
R9127 VN.n6820 VN.n6817 0.01
R9128 VN.n8011 VN.n8008 0.01
R9129 VN.n8860 VN.n8857 0.01
R9130 VN.n9722 VN.n9719 0.01
R9131 VN.n10609 VN.n10600 0.01
R9132 VN.n12144 VN.n12143 0.01
R9133 VN.n11138 VN.n11135 0.01
R9134 VN.n11982 VN.n11981 0.01
R9135 VN.n11937 VN.n11936 0.01
R9136 VN.n11924 VN.n11922 0.01
R9137 VN.n11888 VN.n11887 0.01
R9138 VN.n11630 VN.n11629 0.01
R9139 VN.n11585 VN.n11584 0.01
R9140 VN.n11100 VN.n11098 0.01
R9141 VN.n11524 VN.n11521 0.01
R9142 VN.n11524 VN.n10725 0.01
R9143 VN.n10707 VN.n10705 0.01
R9144 VN.n9827 VN.n9825 0.01
R9145 VN.n8981 VN.n8979 0.01
R9146 VN.n8148 VN.n8146 0.01
R9147 VN.n7337 VN.n7335 0.01
R9148 VN.n6544 VN.n6542 0.01
R9149 VN.n5768 VN.n5766 0.01
R9150 VN.n5005 VN.n5003 0.01
R9151 VN.n4264 VN.n4262 0.01
R9152 VN.n3536 VN.n3534 0.01
R9153 VN.n2830 VN.n2828 0.01
R9154 VN.n2137 VN.n2135 0.01
R9155 VN.n1463 VN.n1461 0.01
R9156 VN.n12385 VN.n12373 0.01
R9157 VN.n821 VN.n197 0.01
R9158 VN.n12405 VN.n12398 0.01
R9159 VN.n12115 VN.n12097 0.01
R9160 VN.n12049 VN.n12048 0.01
R9161 VN.n12004 VN.n12003 0.01
R9162 VN.n11959 VN.n11958 0.01
R9163 VN.n11652 VN.n11651 0.01
R9164 VN.n11607 VN.n11606 0.01
R9165 VN.n11910 VN.n11909 0.01
R9166 VN.n194 VN.n192 0.01
R9167 VN.n10565 VN.n10563 0.01
R9168 VN.n12025 VN.n12024 0.01
R9169 VN.n11980 VN.n11979 0.01
R9170 VN.n11935 VN.n11934 0.01
R9171 VN.n11628 VN.n11627 0.01
R9172 VN.n11583 VN.n11582 0.01
R9173 VN.n489 VN.n479 0.01
R9174 VN.n1815 VN.n1804 0.01
R9175 VN.n3212 VN.n3201 0.01
R9176 VN.n4679 VN.n4668 0.01
R9177 VN.n6216 VN.n6214 0.01
R9178 VN.n7818 VN.n7807 0.01
R9179 VN.n9495 VN.n9484 0.01
R9180 VN.n13137 VN.n12216 0.009
R9181 VN.n925 VN.n924 0.009
R9182 VN.t51 VN.n76 0.009
R9183 VN.n12201 VN.n12200 0.009
R9184 VN.n12202 VN.n12201 0.009
R9185 VN.n12203 VN.n12202 0.009
R9186 VN.n12204 VN.n12203 0.009
R9187 VN.n12205 VN.n12204 0.009
R9188 VN.n12206 VN.n12205 0.009
R9189 VN.n12207 VN.n12206 0.009
R9190 VN.n12208 VN.n12207 0.009
R9191 VN.n12209 VN.n12208 0.009
R9192 VN.n12210 VN.n12209 0.009
R9193 VN.n12211 VN.n12210 0.009
R9194 VN.n12212 VN.n12211 0.009
R9195 VN.n12213 VN.n12212 0.009
R9196 VN.n12214 VN.n12213 0.009
R9197 VN.n12215 VN.n12214 0.009
R9198 VN.n13138 VN.n12215 0.009
R9199 VN.n821 VN.n820 0.009
R9200 VN.n30 VN.n29 0.008
R9201 VN.n97 VN.n95 0.008
R9202 VN.n208 VN.n207 0.008
R9203 VN.n879 VN.n878 0.008
R9204 VN.n1562 VN.n1561 0.008
R9205 VN.n2270 VN.n2269 0.008
R9206 VN.n2992 VN.n2991 0.008
R9207 VN.n3732 VN.n3731 0.008
R9208 VN.n4489 VN.n4488 0.008
R9209 VN.n5264 VN.n5263 0.008
R9210 VN.n6056 VN.n6055 0.008
R9211 VN.n7299 VN.n7298 0.008
R9212 VN.n7688 VN.n7687 0.008
R9213 VN.n8533 VN.n8532 0.008
R9214 VN.n9395 VN.n9394 0.008
R9215 VN.n10278 VN.n10277 0.008
R9216 VN.n3581 VN.n3580 0.008
R9217 VN.n4338 VN.n4337 0.008
R9218 VN.n5113 VN.n5112 0.008
R9219 VN.n5905 VN.n5904 0.008
R9220 VN.n7148 VN.n7147 0.008
R9221 VN.n7537 VN.n7536 0.008
R9222 VN.n8382 VN.n8381 0.008
R9223 VN.n9244 VN.n9243 0.008
R9224 VN.n10126 VN.n10125 0.008
R9225 VN.n10995 VN.n10994 0.008
R9226 VN.n2882 VN.n2881 0.008
R9227 VN.n3622 VN.n3621 0.008
R9228 VN.n4379 VN.n4378 0.008
R9229 VN.n5154 VN.n5153 0.008
R9230 VN.n5946 VN.n5945 0.008
R9231 VN.n7189 VN.n7188 0.008
R9232 VN.n7578 VN.n7577 0.008
R9233 VN.n8423 VN.n8422 0.008
R9234 VN.n9285 VN.n9284 0.008
R9235 VN.n10167 VN.n10166 0.008
R9236 VN.n11031 VN.n11030 0.008
R9237 VN.n5050 VN.n5049 0.008
R9238 VN.n5842 VN.n5841 0.008
R9239 VN.n7085 VN.n7084 0.008
R9240 VN.n7474 VN.n7473 0.008
R9241 VN.n8319 VN.n8318 0.008
R9242 VN.n9181 VN.n9180 0.008
R9243 VN.n10063 VN.n10062 0.008
R9244 VN.n10937 VN.n10936 0.008
R9245 VN.n4316 VN.n4315 0.008
R9246 VN.n5091 VN.n5090 0.008
R9247 VN.n5883 VN.n5882 0.008
R9248 VN.n7126 VN.n7125 0.008
R9249 VN.n7515 VN.n7514 0.008
R9250 VN.n8360 VN.n8359 0.008
R9251 VN.n9222 VN.n9221 0.008
R9252 VN.n10104 VN.n10103 0.008
R9253 VN.n10973 VN.n10972 0.008
R9254 VN.n7022 VN.n7021 0.008
R9255 VN.n7411 VN.n7410 0.008
R9256 VN.n8256 VN.n8255 0.008
R9257 VN.n9118 VN.n9117 0.008
R9258 VN.n10000 VN.n9999 0.008
R9259 VN.n10879 VN.n10878 0.008
R9260 VN.n5820 VN.n5819 0.008
R9261 VN.n7063 VN.n7062 0.008
R9262 VN.n7452 VN.n7451 0.008
R9263 VN.n8297 VN.n8296 0.008
R9264 VN.n9159 VN.n9158 0.008
R9265 VN.n10041 VN.n10040 0.008
R9266 VN.n10915 VN.n10914 0.008
R9267 VN.n7389 VN.n7388 0.008
R9268 VN.n8234 VN.n8233 0.008
R9269 VN.n9096 VN.n9095 0.008
R9270 VN.n9978 VN.n9977 0.008
R9271 VN.n10857 VN.n10856 0.008
R9272 VN.n8193 VN.n8192 0.008
R9273 VN.n9055 VN.n9054 0.008
R9274 VN.n9937 VN.n9936 0.008
R9275 VN.n10821 VN.n10820 0.008
R9276 VN.n9874 VN.n9873 0.008
R9277 VN.n10763 VN.n10762 0.008
R9278 VN.n9033 VN.n9032 0.008
R9279 VN.n9915 VN.n9914 0.008
R9280 VN.n10799 VN.n10798 0.008
R9281 VN.n10741 VN.n10740 0.008
R9282 VN.n11458 VN.n11457 0.008
R9283 VN.n11464 VN.n11463 0.008
R9284 VN.n10290 VN.n10289 0.008
R9285 VN.n10296 VN.n10295 0.008
R9286 VN.n9407 VN.n9406 0.008
R9287 VN.n9413 VN.n9412 0.008
R9288 VN.n8545 VN.n8544 0.008
R9289 VN.n8551 VN.n8550 0.008
R9290 VN.n7700 VN.n7699 0.008
R9291 VN.n7706 VN.n7705 0.008
R9292 VN.n7311 VN.n7310 0.008
R9293 VN.n7317 VN.n7316 0.008
R9294 VN.n6068 VN.n6067 0.008
R9295 VN.n6074 VN.n6073 0.008
R9296 VN.n5276 VN.n5275 0.008
R9297 VN.n5282 VN.n5281 0.008
R9298 VN.n4501 VN.n4500 0.008
R9299 VN.n4507 VN.n4506 0.008
R9300 VN.n3744 VN.n3743 0.008
R9301 VN.n3750 VN.n3749 0.008
R9302 VN.n3004 VN.n3003 0.008
R9303 VN.n3010 VN.n3009 0.008
R9304 VN.n2282 VN.n2281 0.008
R9305 VN.n2288 VN.n2287 0.008
R9306 VN.n1574 VN.n1573 0.008
R9307 VN.n1580 VN.n1579 0.008
R9308 VN.n891 VN.n890 0.008
R9309 VN.n897 VN.n896 0.008
R9310 VN.n220 VN.n219 0.008
R9311 VN.n226 VN.n225 0.008
R9312 VN.n12249 VN.n12248 0.008
R9313 VN.n11044 VN.n11043 0.008
R9314 VN.n10202 VN.n10201 0.008
R9315 VN.n10208 VN.n10207 0.008
R9316 VN.n9319 VN.n9318 0.008
R9317 VN.n9325 VN.n9324 0.008
R9318 VN.n8457 VN.n8456 0.008
R9319 VN.n8463 VN.n8462 0.008
R9320 VN.n7612 VN.n7611 0.008
R9321 VN.n7618 VN.n7617 0.008
R9322 VN.n7223 VN.n7222 0.008
R9323 VN.n7229 VN.n7228 0.008
R9324 VN.n5980 VN.n5979 0.008
R9325 VN.n5986 VN.n5985 0.008
R9326 VN.n5188 VN.n5187 0.008
R9327 VN.n5194 VN.n5193 0.008
R9328 VN.n4413 VN.n4412 0.008
R9329 VN.n4419 VN.n4418 0.008
R9330 VN.n3656 VN.n3655 0.008
R9331 VN.n3662 VN.n3661 0.008
R9332 VN.n2916 VN.n2915 0.008
R9333 VN.n2922 VN.n2921 0.008
R9334 VN.n2194 VN.n2193 0.008
R9335 VN.n2200 VN.n2199 0.008
R9336 VN.n1602 VN.n1601 0.008
R9337 VN.n10588 VN.n10577 0.008
R9338 VN.n9703 VN.n9692 0.008
R9339 VN.n8841 VN.n8830 0.008
R9340 VN.n7992 VN.n7981 0.008
R9341 VN.n6801 VN.n6790 0.008
R9342 VN.n6356 VN.n6345 0.008
R9343 VN.n5564 VN.n5553 0.008
R9344 VN.n4785 VN.n4774 0.008
R9345 VN.n4028 VN.n4017 0.008
R9346 VN.n3284 VN.n3273 0.008
R9347 VN.n2562 VN.n2551 0.008
R9348 VN.n1853 VN.n1842 0.008
R9349 VN.n1163 VN.n1152 0.008
R9350 VN.n11397 VN.n11396 0.008
R9351 VN.n507 VN.n506 0.008
R9352 VN.n1182 VN.n1181 0.008
R9353 VN.n1872 VN.n1871 0.008
R9354 VN.n2581 VN.n2580 0.008
R9355 VN.n3303 VN.n3302 0.008
R9356 VN.n4047 VN.n4046 0.008
R9357 VN.n4804 VN.n4803 0.008
R9358 VN.n5583 VN.n5582 0.008
R9359 VN.n6375 VN.n6374 0.008
R9360 VN.n6820 VN.n6819 0.008
R9361 VN.n8011 VN.n8010 0.008
R9362 VN.n8860 VN.n8859 0.008
R9363 VN.n9722 VN.n9721 0.008
R9364 VN.n10609 VN.n10598 0.008
R9365 VN.n11422 VN.n11421 0.008
R9366 VN.n10250 VN.n10249 0.008
R9367 VN.n9367 VN.n9366 0.008
R9368 VN.n8505 VN.n8504 0.008
R9369 VN.n7660 VN.n7659 0.008
R9370 VN.n7271 VN.n7270 0.008
R9371 VN.n6028 VN.n6027 0.008
R9372 VN.n5236 VN.n5235 0.008
R9373 VN.n4461 VN.n4460 0.008
R9374 VN.n3704 VN.n3703 0.008
R9375 VN.n2964 VN.n2963 0.008
R9376 VN.n2242 VN.n2241 0.008
R9377 VN.n1537 VN.n1536 0.008
R9378 VN.n851 VN.n850 0.008
R9379 VN.n12125 VN.n12124 0.008
R9380 VN.n12140 VN.n12136 0.008
R9381 VN.n12140 VN.n12139 0.008
R9382 VN.n11138 VN.n11137 0.008
R9383 VN.n2319 VN.n2315 0.008
R9384 VN.n2868 VN.n2867 0.008
R9385 VN.n3608 VN.n3607 0.008
R9386 VN.n4365 VN.n4364 0.008
R9387 VN.n5140 VN.n5139 0.008
R9388 VN.n5932 VN.n5931 0.008
R9389 VN.n7175 VN.n7174 0.008
R9390 VN.n7564 VN.n7563 0.008
R9391 VN.n8409 VN.n8408 0.008
R9392 VN.n9271 VN.n9270 0.008
R9393 VN.n10153 VN.n10152 0.008
R9394 VN.n11018 VN.n11017 0.008
R9395 VN.n11008 VN.n11007 0.008
R9396 VN.n10138 VN.n10137 0.008
R9397 VN.n10144 VN.n10143 0.008
R9398 VN.n9256 VN.n9255 0.008
R9399 VN.n9262 VN.n9261 0.008
R9400 VN.n8394 VN.n8393 0.008
R9401 VN.n8400 VN.n8399 0.008
R9402 VN.n7549 VN.n7548 0.008
R9403 VN.n7555 VN.n7554 0.008
R9404 VN.n7160 VN.n7159 0.008
R9405 VN.n7166 VN.n7165 0.008
R9406 VN.n5917 VN.n5916 0.008
R9407 VN.n5923 VN.n5922 0.008
R9408 VN.n5125 VN.n5124 0.008
R9409 VN.n5131 VN.n5130 0.008
R9410 VN.n4350 VN.n4349 0.008
R9411 VN.n4356 VN.n4355 0.008
R9412 VN.n3593 VN.n3592 0.008
R9413 VN.n3599 VN.n3598 0.008
R9414 VN.n3029 VN.n3028 0.008
R9415 VN.n3781 VN.n3779 0.008
R9416 VN.n4302 VN.n4301 0.008
R9417 VN.n5077 VN.n5076 0.008
R9418 VN.n5869 VN.n5868 0.008
R9419 VN.n7112 VN.n7111 0.008
R9420 VN.n7501 VN.n7500 0.008
R9421 VN.n8346 VN.n8345 0.008
R9422 VN.n9208 VN.n9207 0.008
R9423 VN.n10090 VN.n10089 0.008
R9424 VN.n10960 VN.n10959 0.008
R9425 VN.n10950 VN.n10949 0.008
R9426 VN.n10075 VN.n10074 0.008
R9427 VN.n10081 VN.n10080 0.008
R9428 VN.n9193 VN.n9192 0.008
R9429 VN.n9199 VN.n9198 0.008
R9430 VN.n8331 VN.n8330 0.008
R9431 VN.n8337 VN.n8336 0.008
R9432 VN.n7486 VN.n7485 0.008
R9433 VN.n7492 VN.n7491 0.008
R9434 VN.n7097 VN.n7096 0.008
R9435 VN.n7103 VN.n7102 0.008
R9436 VN.n5854 VN.n5853 0.008
R9437 VN.n5860 VN.n5859 0.008
R9438 VN.n5062 VN.n5061 0.008
R9439 VN.n5068 VN.n5067 0.008
R9440 VN.n4526 VN.n4525 0.008
R9441 VN.n5313 VN.n5311 0.008
R9442 VN.n5806 VN.n5805 0.008
R9443 VN.n7049 VN.n7048 0.008
R9444 VN.n7438 VN.n7437 0.008
R9445 VN.n8283 VN.n8282 0.008
R9446 VN.n9145 VN.n9144 0.008
R9447 VN.n10027 VN.n10026 0.008
R9448 VN.n10902 VN.n10901 0.008
R9449 VN.n10892 VN.n10891 0.008
R9450 VN.n10012 VN.n10011 0.008
R9451 VN.n10018 VN.n10017 0.008
R9452 VN.n9130 VN.n9129 0.008
R9453 VN.n9136 VN.n9135 0.008
R9454 VN.n8268 VN.n8267 0.008
R9455 VN.n8274 VN.n8273 0.008
R9456 VN.n7423 VN.n7422 0.008
R9457 VN.n7429 VN.n7428 0.008
R9458 VN.n7034 VN.n7033 0.008
R9459 VN.n7040 VN.n7039 0.008
R9460 VN.n6093 VN.n6092 0.008
R9461 VN.n6601 VN.n6599 0.008
R9462 VN.n10834 VN.n10833 0.008
R9463 VN.n9949 VN.n9948 0.008
R9464 VN.n9955 VN.n9954 0.008
R9465 VN.n9067 VN.n9066 0.008
R9466 VN.n9073 VN.n9072 0.008
R9467 VN.n8205 VN.n8204 0.008
R9468 VN.n8211 VN.n8210 0.008
R9469 VN.n7725 VN.n7724 0.008
R9470 VN.n8582 VN.n8578 0.008
R9471 VN.n9019 VN.n9018 0.008
R9472 VN.n9901 VN.n9900 0.008
R9473 VN.n10786 VN.n10785 0.008
R9474 VN.n10776 VN.n10775 0.008
R9475 VN.n9886 VN.n9885 0.008
R9476 VN.n9892 VN.n9891 0.008
R9477 VN.n9432 VN.n9431 0.008
R9478 VN.n10327 VN.n10323 0.008
R9479 VN.n10728 VN.n10727 0.008
R9480 VN.n12184 VN.n12183 0.008
R9481 VN.n12185 VN.n12184 0.008
R9482 VN.n12186 VN.n12185 0.008
R9483 VN.n12187 VN.n12186 0.008
R9484 VN.n12188 VN.n12187 0.008
R9485 VN.n12189 VN.n12188 0.008
R9486 VN.n12190 VN.n12189 0.008
R9487 VN.n12191 VN.n12190 0.008
R9488 VN.n12192 VN.n12191 0.008
R9489 VN.n12193 VN.n12192 0.008
R9490 VN.n12194 VN.n12193 0.008
R9491 VN.n12195 VN.n12194 0.008
R9492 VN.n12196 VN.n12195 0.008
R9493 VN.n12197 VN.n12196 0.008
R9494 VN.n12198 VN.n12197 0.008
R9495 VN.n12199 VN.n12198 0.008
R9496 VN.n11100 VN.n11099 0.008
R9497 VN.n12182 VN.n12181 0.008
R9498 VN.n755 VN.n754 0.008
R9499 VN.n12221 VN.n12220 0.008
R9500 VN VN.n13138 0.008
R9501 VN.n11566 VN.n11565 0.008
R9502 VN.n10843 VN.n10842 0.008
R9503 VN.n9964 VN.n9963 0.008
R9504 VN.n9082 VN.n9081 0.008
R9505 VN.n8220 VN.n8219 0.008
R9506 VN.n7375 VN.n7374 0.008
R9507 VN.n12114 VN.n12113 0.008
R9508 VN.n12114 VN.n12112 0.007
R9509 VN.t8 VN.n11719 0.007
R9510 VN.t8 VN.n11708 0.007
R9511 VN.t8 VN.n11730 0.007
R9512 VN.t8 VN.n11741 0.007
R9513 VN.t8 VN.n11752 0.007
R9514 VN.t8 VN.n11763 0.007
R9515 VN.t8 VN.n11772 0.007
R9516 VN.n196 VN.n195 0.007
R9517 VN.n12096 VN.n12095 0.007
R9518 VN.n11559 VN.n11558 0.007
R9519 VN.t51 VN.n70 0.006
R9520 VN.t51 VN.n67 0.006
R9521 VN.t51 VN.n64 0.006
R9522 VN.t51 VN.n61 0.006
R9523 VN.t51 VN.n58 0.006
R9524 VN.t51 VN.n55 0.006
R9525 VN.t51 VN.n52 0.006
R9526 VN.t51 VN.n49 0.006
R9527 VN.t51 VN.n46 0.006
R9528 VN.t51 VN.n43 0.006
R9529 VN.t51 VN.n40 0.006
R9530 VN.t51 VN.n37 0.006
R9531 VN.t51 VN.n32 0.006
R9532 VN.n11459 VN.n11458 0.006
R9533 VN.n10291 VN.n10290 0.006
R9534 VN.n9408 VN.n9407 0.006
R9535 VN.n8546 VN.n8545 0.006
R9536 VN.n7701 VN.n7700 0.006
R9537 VN.n7312 VN.n7311 0.006
R9538 VN.n6069 VN.n6068 0.006
R9539 VN.n5277 VN.n5276 0.006
R9540 VN.n4502 VN.n4501 0.006
R9541 VN.n3745 VN.n3744 0.006
R9542 VN.n3005 VN.n3004 0.006
R9543 VN.n2283 VN.n2282 0.006
R9544 VN.n1575 VN.n1574 0.006
R9545 VN.n892 VN.n891 0.006
R9546 VN.n221 VN.n220 0.006
R9547 VN.n12250 VN.n12249 0.006
R9548 VN.n10203 VN.n10202 0.006
R9549 VN.n9320 VN.n9319 0.006
R9550 VN.n8458 VN.n8457 0.006
R9551 VN.n7613 VN.n7612 0.006
R9552 VN.n7224 VN.n7223 0.006
R9553 VN.n5981 VN.n5980 0.006
R9554 VN.n5189 VN.n5188 0.006
R9555 VN.n4414 VN.n4413 0.006
R9556 VN.n3657 VN.n3656 0.006
R9557 VN.n2917 VN.n2916 0.006
R9558 VN.n2195 VN.n2194 0.006
R9559 VN.n1603 VN.n1602 0.006
R9560 VN.n10139 VN.n10138 0.006
R9561 VN.n9257 VN.n9256 0.006
R9562 VN.n8395 VN.n8394 0.006
R9563 VN.n7550 VN.n7549 0.006
R9564 VN.n7161 VN.n7160 0.006
R9565 VN.n5918 VN.n5917 0.006
R9566 VN.n5126 VN.n5125 0.006
R9567 VN.n4351 VN.n4350 0.006
R9568 VN.n3594 VN.n3593 0.006
R9569 VN.n3030 VN.n3029 0.006
R9570 VN.n10076 VN.n10075 0.006
R9571 VN.n9194 VN.n9193 0.006
R9572 VN.n8332 VN.n8331 0.006
R9573 VN.n7487 VN.n7486 0.006
R9574 VN.n7098 VN.n7097 0.006
R9575 VN.n5855 VN.n5854 0.006
R9576 VN.n5063 VN.n5062 0.006
R9577 VN.n4527 VN.n4526 0.006
R9578 VN.n10013 VN.n10012 0.006
R9579 VN.n9131 VN.n9130 0.006
R9580 VN.n8269 VN.n8268 0.006
R9581 VN.n7424 VN.n7423 0.006
R9582 VN.n7035 VN.n7034 0.006
R9583 VN.n6094 VN.n6093 0.006
R9584 VN.n9950 VN.n9949 0.006
R9585 VN.n9068 VN.n9067 0.006
R9586 VN.n8206 VN.n8205 0.006
R9587 VN.n7726 VN.n7725 0.006
R9588 VN.n9887 VN.n9886 0.006
R9589 VN.n9433 VN.n9432 0.006
R9590 VN.n12222 VN.n12221 0.006
R9591 VN.n31 VN.n30 0.006
R9592 VN.n98 VN.n97 0.006
R9593 VN.n12036 VN.n12027 0.006
R9594 VN.n11991 VN.n11982 0.006
R9595 VN.n11946 VN.n11937 0.006
R9596 VN.n11897 VN.n11888 0.006
R9597 VN.n11639 VN.n11630 0.006
R9598 VN.n11594 VN.n11585 0.006
R9599 VN.n12081 VN.n12067 0.005
R9600 VN.n11062 VN.n11061 0.005
R9601 VN.n2182 VN.n2181 0.005
R9602 VN.n2904 VN.n2903 0.005
R9603 VN.n3644 VN.n3643 0.005
R9604 VN.n4401 VN.n4400 0.005
R9605 VN.n5176 VN.n5175 0.005
R9606 VN.n5968 VN.n5967 0.005
R9607 VN.n7211 VN.n7210 0.005
R9608 VN.n7600 VN.n7599 0.005
R9609 VN.n8445 VN.n8444 0.005
R9610 VN.n9307 VN.n9306 0.005
R9611 VN.n10190 VN.n10189 0.005
R9612 VN.t8 VN.n11702 0.005
R9613 VN.n2314 VN.n2313 0.005
R9614 VN.n3776 VN.n3775 0.005
R9615 VN.n5308 VN.n5307 0.005
R9616 VN.n6596 VN.n6595 0.005
R9617 VN.n8577 VN.n8576 0.005
R9618 VN.n10322 VN.n10321 0.005
R9619 VN.n29 VN.n25 0.005
R9620 VN.n95 VN.n91 0.005
R9621 VN.t8 VN.n11693 0.005
R9622 VN.n11570 VN.n11569 0.004
R9623 VN.n13117 VN.n13116 0.004
R9624 VN.n12155 VN.n12154 0.004
R9625 VN.n12242 VN.n12241 0.004
R9626 VN.n12707 VN.n12706 0.004
R9627 VN.n213 VN.n212 0.004
R9628 VN.n518 VN.n517 0.004
R9629 VN.n884 VN.n883 0.004
R9630 VN.n1193 VN.n1192 0.004
R9631 VN.n1567 VN.n1566 0.004
R9632 VN.n1883 VN.n1882 0.004
R9633 VN.n2275 VN.n2274 0.004
R9634 VN.n2592 VN.n2591 0.004
R9635 VN.n2997 VN.n2996 0.004
R9636 VN.n3314 VN.n3313 0.004
R9637 VN.n3737 VN.n3736 0.004
R9638 VN.n4058 VN.n4057 0.004
R9639 VN.n4494 VN.n4493 0.004
R9640 VN.n4815 VN.n4814 0.004
R9641 VN.n5269 VN.n5268 0.004
R9642 VN.n5594 VN.n5593 0.004
R9643 VN.n6061 VN.n6060 0.004
R9644 VN.n6386 VN.n6385 0.004
R9645 VN.n7304 VN.n7303 0.004
R9646 VN.n6831 VN.n6830 0.004
R9647 VN.n7693 VN.n7692 0.004
R9648 VN.n8022 VN.n8021 0.004
R9649 VN.n8538 VN.n8537 0.004
R9650 VN.n8871 VN.n8870 0.004
R9651 VN.n9400 VN.n9399 0.004
R9652 VN.n9733 VN.n9732 0.004
R9653 VN.n10283 VN.n10282 0.004
R9654 VN.n10620 VN.n10619 0.004
R9655 VN.n11452 VN.n11451 0.004
R9656 VN.n11112 VN.n11111 0.004
R9657 VN.n12034 VN.n12033 0.004
R9658 VN.n3023 VN.n3022 0.004
R9659 VN.n3222 VN.n3221 0.004
R9660 VN.n3586 VN.n3585 0.004
R9661 VN.n3966 VN.n3965 0.004
R9662 VN.n4343 VN.n4342 0.004
R9663 VN.n4723 VN.n4722 0.004
R9664 VN.n5118 VN.n5117 0.004
R9665 VN.n5502 VN.n5501 0.004
R9666 VN.n5910 VN.n5909 0.004
R9667 VN.n6294 VN.n6293 0.004
R9668 VN.n7153 VN.n7152 0.004
R9669 VN.n6739 VN.n6738 0.004
R9670 VN.n7542 VN.n7541 0.004
R9671 VN.n7930 VN.n7929 0.004
R9672 VN.n8387 VN.n8386 0.004
R9673 VN.n8779 VN.n8778 0.004
R9674 VN.n9249 VN.n9248 0.004
R9675 VN.n9641 VN.n9640 0.004
R9676 VN.n10131 VN.n10130 0.004
R9677 VN.n10518 VN.n10517 0.004
R9678 VN.n11000 VN.n10999 0.004
R9679 VN.n11182 VN.n11181 0.004
R9680 VN.n12057 VN.n12056 0.004
R9681 VN.n2311 VN.n2310 0.004
R9682 VN.n2521 VN.n2520 0.004
R9683 VN.n2878 VN.n2877 0.004
R9684 VN.n3243 VN.n3242 0.004
R9685 VN.n3618 VN.n3617 0.004
R9686 VN.n3987 VN.n3986 0.004
R9687 VN.n4375 VN.n4374 0.004
R9688 VN.n4744 VN.n4743 0.004
R9689 VN.n5150 VN.n5149 0.004
R9690 VN.n5523 VN.n5522 0.004
R9691 VN.n5942 VN.n5941 0.004
R9692 VN.n6315 VN.n6314 0.004
R9693 VN.n7185 VN.n7184 0.004
R9694 VN.n6760 VN.n6759 0.004
R9695 VN.n7574 VN.n7573 0.004
R9696 VN.n7951 VN.n7950 0.004
R9697 VN.n8419 VN.n8418 0.004
R9698 VN.n8800 VN.n8799 0.004
R9699 VN.n9281 VN.n9280 0.004
R9700 VN.n9662 VN.n9661 0.004
R9701 VN.n10163 VN.n10162 0.004
R9702 VN.n10540 VN.n10539 0.004
R9703 VN.n10561 VN.n10560 0.004
R9704 VN.n11054 VN.n11053 0.004
R9705 VN.n11152 VN.n11151 0.004
R9706 VN.n12074 VN.n12073 0.004
R9707 VN.n10195 VN.n10194 0.004
R9708 VN.n9312 VN.n9311 0.004
R9709 VN.n8450 VN.n8449 0.004
R9710 VN.n7605 VN.n7604 0.004
R9711 VN.n7216 VN.n7215 0.004
R9712 VN.n5973 VN.n5972 0.004
R9713 VN.n5181 VN.n5180 0.004
R9714 VN.n4406 VN.n4405 0.004
R9715 VN.n3649 VN.n3648 0.004
R9716 VN.n2909 VN.n2908 0.004
R9717 VN.n2187 VN.n2186 0.004
R9718 VN.n1596 VN.n1595 0.004
R9719 VN.n1825 VN.n1824 0.004
R9720 VN.n2534 VN.n2533 0.004
R9721 VN.n3256 VN.n3255 0.004
R9722 VN.n4000 VN.n3999 0.004
R9723 VN.n4757 VN.n4756 0.004
R9724 VN.n5536 VN.n5535 0.004
R9725 VN.n6328 VN.n6327 0.004
R9726 VN.n6773 VN.n6772 0.004
R9727 VN.n7964 VN.n7963 0.004
R9728 VN.n8813 VN.n8812 0.004
R9729 VN.n9675 VN.n9674 0.004
R9730 VN.n11405 VN.n11404 0.004
R9731 VN.n11391 VN.n11390 0.004
R9732 VN.n12108 VN.n12107 0.004
R9733 VN.n917 VN.n916 0.004
R9734 VN.n1158 VN.n1157 0.004
R9735 VN.n1511 VN.n1510 0.004
R9736 VN.n1848 VN.n1847 0.004
R9737 VN.n2219 VN.n2218 0.004
R9738 VN.n2557 VN.n2556 0.004
R9739 VN.n2941 VN.n2940 0.004
R9740 VN.n3279 VN.n3278 0.004
R9741 VN.n3681 VN.n3680 0.004
R9742 VN.n4023 VN.n4022 0.004
R9743 VN.n4438 VN.n4437 0.004
R9744 VN.n4780 VN.n4779 0.004
R9745 VN.n5213 VN.n5212 0.004
R9746 VN.n5559 VN.n5558 0.004
R9747 VN.n6005 VN.n6004 0.004
R9748 VN.n6351 VN.n6350 0.004
R9749 VN.n7248 VN.n7247 0.004
R9750 VN.n6796 VN.n6795 0.004
R9751 VN.n7637 VN.n7636 0.004
R9752 VN.n7987 VN.n7986 0.004
R9753 VN.n8482 VN.n8481 0.004
R9754 VN.n8836 VN.n8835 0.004
R9755 VN.n9344 VN.n9343 0.004
R9756 VN.n9698 VN.n9697 0.004
R9757 VN.n10227 VN.n10226 0.004
R9758 VN.n10583 VN.n10582 0.004
R9759 VN.n11432 VN.n11431 0.004
R9760 VN.n11133 VN.n11132 0.004
R9761 VN.n10603 VN.n10602 0.004
R9762 VN.n10260 VN.n10259 0.004
R9763 VN.n9718 VN.n9717 0.004
R9764 VN.n9377 VN.n9376 0.004
R9765 VN.n8856 VN.n8855 0.004
R9766 VN.n8515 VN.n8514 0.004
R9767 VN.n8007 VN.n8006 0.004
R9768 VN.n7670 VN.n7669 0.004
R9769 VN.n6816 VN.n6815 0.004
R9770 VN.n7281 VN.n7280 0.004
R9771 VN.n6371 VN.n6370 0.004
R9772 VN.n6038 VN.n6037 0.004
R9773 VN.n5579 VN.n5578 0.004
R9774 VN.n5246 VN.n5245 0.004
R9775 VN.n4800 VN.n4799 0.004
R9776 VN.n4471 VN.n4470 0.004
R9777 VN.n4043 VN.n4042 0.004
R9778 VN.n3714 VN.n3713 0.004
R9779 VN.n3299 VN.n3298 0.004
R9780 VN.n2974 VN.n2973 0.004
R9781 VN.n2577 VN.n2576 0.004
R9782 VN.n2252 VN.n2251 0.004
R9783 VN.n1868 VN.n1867 0.004
R9784 VN.n1547 VN.n1546 0.004
R9785 VN.n1178 VN.n1177 0.004
R9786 VN.n861 VN.n860 0.004
R9787 VN.n503 VN.n502 0.004
R9788 VN.n250 VN.n249 0.004
R9789 VN.n12134 VN.n12133 0.004
R9790 VN.n11027 VN.n11026 0.004
R9791 VN.n11170 VN.n11169 0.004
R9792 VN.n11989 VN.n11988 0.004
R9793 VN.n4520 VN.n4519 0.004
R9794 VN.n4689 VN.n4688 0.004
R9795 VN.n5055 VN.n5054 0.004
R9796 VN.n5468 VN.n5467 0.004
R9797 VN.n5847 VN.n5846 0.004
R9798 VN.n6260 VN.n6259 0.004
R9799 VN.n7090 VN.n7089 0.004
R9800 VN.n6705 VN.n6704 0.004
R9801 VN.n7479 VN.n7478 0.004
R9802 VN.n7896 VN.n7895 0.004
R9803 VN.n8324 VN.n8323 0.004
R9804 VN.n8745 VN.n8744 0.004
R9805 VN.n9186 VN.n9185 0.004
R9806 VN.n9607 VN.n9606 0.004
R9807 VN.n10068 VN.n10067 0.004
R9808 VN.n10483 VN.n10482 0.004
R9809 VN.n10942 VN.n10941 0.004
R9810 VN.n11216 VN.n11215 0.004
R9811 VN.n12012 VN.n12011 0.004
R9812 VN.n3773 VN.n3772 0.004
R9813 VN.n3953 VN.n3952 0.004
R9814 VN.n4312 VN.n4311 0.004
R9815 VN.n4710 VN.n4709 0.004
R9816 VN.n5087 VN.n5086 0.004
R9817 VN.n5489 VN.n5488 0.004
R9818 VN.n5879 VN.n5878 0.004
R9819 VN.n6281 VN.n6280 0.004
R9820 VN.n7122 VN.n7121 0.004
R9821 VN.n6726 VN.n6725 0.004
R9822 VN.n7511 VN.n7510 0.004
R9823 VN.n7917 VN.n7916 0.004
R9824 VN.n8356 VN.n8355 0.004
R9825 VN.n8766 VN.n8765 0.004
R9826 VN.n9218 VN.n9217 0.004
R9827 VN.n9628 VN.n9627 0.004
R9828 VN.n10100 VN.n10099 0.004
R9829 VN.n10505 VN.n10504 0.004
R9830 VN.n10969 VN.n10968 0.004
R9831 VN.n11204 VN.n11203 0.004
R9832 VN.n11944 VN.n11943 0.004
R9833 VN.n6087 VN.n6086 0.004
R9834 VN.n6226 VN.n6225 0.004
R9835 VN.n7027 VN.n7026 0.004
R9836 VN.n6671 VN.n6670 0.004
R9837 VN.n7416 VN.n7415 0.004
R9838 VN.n7862 VN.n7861 0.004
R9839 VN.n8261 VN.n8260 0.004
R9840 VN.n8711 VN.n8710 0.004
R9841 VN.n9123 VN.n9122 0.004
R9842 VN.n9573 VN.n9572 0.004
R9843 VN.n10005 VN.n10004 0.004
R9844 VN.n10448 VN.n10447 0.004
R9845 VN.n10884 VN.n10883 0.004
R9846 VN.n11250 VN.n11249 0.004
R9847 VN.n11967 VN.n11966 0.004
R9848 VN.n5305 VN.n5304 0.004
R9849 VN.n5455 VN.n5454 0.004
R9850 VN.n5816 VN.n5815 0.004
R9851 VN.n6247 VN.n6246 0.004
R9852 VN.n7059 VN.n7058 0.004
R9853 VN.n6692 VN.n6691 0.004
R9854 VN.n7448 VN.n7447 0.004
R9855 VN.n7883 VN.n7882 0.004
R9856 VN.n8293 VN.n8292 0.004
R9857 VN.n8732 VN.n8731 0.004
R9858 VN.n9155 VN.n9154 0.004
R9859 VN.n9594 VN.n9593 0.004
R9860 VN.n10037 VN.n10036 0.004
R9861 VN.n10470 VN.n10469 0.004
R9862 VN.n10911 VN.n10910 0.004
R9863 VN.n11238 VN.n11237 0.004
R9864 VN.n6658 VN.n6657 0.004
R9865 VN.n7385 VN.n7384 0.004
R9866 VN.n7849 VN.n7848 0.004
R9867 VN.n8230 VN.n8229 0.004
R9868 VN.n8698 VN.n8697 0.004
R9869 VN.n9092 VN.n9091 0.004
R9870 VN.n9560 VN.n9559 0.004
R9871 VN.n9974 VN.n9973 0.004
R9872 VN.n10435 VN.n10434 0.004
R9873 VN.n10853 VN.n10852 0.004
R9874 VN.n11271 VN.n11270 0.004
R9875 VN.n11918 VN.n11917 0.004
R9876 VN.n11895 VN.n11894 0.004
R9877 VN.n7719 VN.n7718 0.004
R9878 VN.n7828 VN.n7827 0.004
R9879 VN.n8198 VN.n8197 0.004
R9880 VN.n8677 VN.n8676 0.004
R9881 VN.n9060 VN.n9059 0.004
R9882 VN.n9539 VN.n9538 0.004
R9883 VN.n9942 VN.n9941 0.004
R9884 VN.n10413 VN.n10412 0.004
R9885 VN.n10826 VN.n10825 0.004
R9886 VN.n11284 VN.n11283 0.004
R9887 VN.n11637 VN.n11636 0.004
R9888 VN.n9426 VN.n9425 0.004
R9889 VN.n9505 VN.n9504 0.004
R9890 VN.n9879 VN.n9878 0.004
R9891 VN.n10378 VN.n10377 0.004
R9892 VN.n10768 VN.n10767 0.004
R9893 VN.n11317 VN.n11316 0.004
R9894 VN.n11874 VN.n11873 0.004
R9895 VN.n8574 VN.n8573 0.004
R9896 VN.n8664 VN.n8663 0.004
R9897 VN.n9029 VN.n9028 0.004
R9898 VN.n9526 VN.n9525 0.004
R9899 VN.n9911 VN.n9910 0.004
R9900 VN.n10400 VN.n10399 0.004
R9901 VN.n10795 VN.n10794 0.004
R9902 VN.n11305 VN.n11304 0.004
R9903 VN.n11592 VN.n11591 0.004
R9904 VN.n11477 VN.n11476 0.004
R9905 VN.n11351 VN.n11350 0.004
R9906 VN.n11615 VN.n11614 0.004
R9907 VN.n10319 VN.n10318 0.004
R9908 VN.n10365 VN.n10364 0.004
R9909 VN.n10737 VN.n10736 0.004
R9910 VN.n11339 VN.n11338 0.004
R9911 VN.n11545 VN.n11544 0.004
R9912 VN.n11097 VN.n11096 0.004
R9913 VN.n11503 VN.n11502 0.004
R9914 VN.n10659 VN.n10658 0.004
R9915 VN.n10669 VN.n10668 0.004
R9916 VN.n9754 VN.n9753 0.004
R9917 VN.n9455 VN.n9454 0.004
R9918 VN.n8892 VN.n8891 0.004
R9919 VN.n8596 VN.n8595 0.004
R9920 VN.n8043 VN.n8042 0.004
R9921 VN.n7748 VN.n7747 0.004
R9922 VN.n6852 VN.n6851 0.004
R9923 VN.n7000 VN.n6999 0.004
R9924 VN.n6407 VN.n6406 0.004
R9925 VN.n6116 VN.n6115 0.004
R9926 VN.n5615 VN.n5614 0.004
R9927 VN.n5327 VN.n5326 0.004
R9928 VN.n4836 VN.n4835 0.004
R9929 VN.n4549 VN.n4548 0.004
R9930 VN.n4079 VN.n4078 0.004
R9931 VN.n3795 VN.n3794 0.004
R9932 VN.n3335 VN.n3334 0.004
R9933 VN.n3052 VN.n3051 0.004
R9934 VN.n2613 VN.n2612 0.004
R9935 VN.n2333 VN.n2332 0.004
R9936 VN.n1904 VN.n1903 0.004
R9937 VN.n1625 VN.n1624 0.004
R9938 VN.n1214 VN.n1213 0.004
R9939 VN.n938 VN.n937 0.004
R9940 VN.n539 VN.n538 0.004
R9941 VN.n266 VN.n265 0.004
R9942 VN.n12296 VN.n12295 0.004
R9943 VN.n12307 VN.n12306 0.004
R9944 VN.n12278 VN.n12277 0.004
R9945 VN.n11519 VN.n11518 0.004
R9946 VN.n10642 VN.n10641 0.004
R9947 VN.n10687 VN.n10686 0.004
R9948 VN.n12349 VN.n12348 0.004
R9949 VN.n12325 VN.n12324 0.004
R9950 VN.n12333 VN.n12332 0.004
R9951 VN.n284 VN.n283 0.004
R9952 VN.n553 VN.n552 0.004
R9953 VN.n956 VN.n955 0.004
R9954 VN.n1228 VN.n1227 0.004
R9955 VN.n1643 VN.n1642 0.004
R9956 VN.n1918 VN.n1917 0.004
R9957 VN.n2351 VN.n2350 0.004
R9958 VN.n2627 VN.n2626 0.004
R9959 VN.n3070 VN.n3069 0.004
R9960 VN.n3349 VN.n3348 0.004
R9961 VN.n3813 VN.n3812 0.004
R9962 VN.n4093 VN.n4092 0.004
R9963 VN.n4567 VN.n4566 0.004
R9964 VN.n4850 VN.n4849 0.004
R9965 VN.n5345 VN.n5344 0.004
R9966 VN.n5629 VN.n5628 0.004
R9967 VN.n6134 VN.n6133 0.004
R9968 VN.n6421 VN.n6420 0.004
R9969 VN.n6983 VN.n6982 0.004
R9970 VN.n6866 VN.n6865 0.004
R9971 VN.n7766 VN.n7765 0.004
R9972 VN.n8057 VN.n8056 0.004
R9973 VN.n8614 VN.n8613 0.004
R9974 VN.n8906 VN.n8905 0.004
R9975 VN.n9473 VN.n9472 0.004
R9976 VN.n9481 VN.n9480 0.004
R9977 VN.n9865 VN.n9864 0.004
R9978 VN.n9771 VN.n9770 0.004
R9979 VN.n9807 VN.n9806 0.004
R9980 VN.n12417 VN.n12416 0.004
R9981 VN.n12643 VN.n12642 0.004
R9982 VN.n12651 VN.n12650 0.004
R9983 VN.n299 VN.n298 0.004
R9984 VN.n569 VN.n568 0.004
R9985 VN.n971 VN.n970 0.004
R9986 VN.n1244 VN.n1243 0.004
R9987 VN.n1658 VN.n1657 0.004
R9988 VN.n1934 VN.n1933 0.004
R9989 VN.n2366 VN.n2365 0.004
R9990 VN.n2643 VN.n2642 0.004
R9991 VN.n3085 VN.n3084 0.004
R9992 VN.n3365 VN.n3364 0.004
R9993 VN.n3828 VN.n3827 0.004
R9994 VN.n4109 VN.n4108 0.004
R9995 VN.n4582 VN.n4581 0.004
R9996 VN.n4866 VN.n4865 0.004
R9997 VN.n5360 VN.n5359 0.004
R9998 VN.n5645 VN.n5644 0.004
R9999 VN.n6149 VN.n6148 0.004
R10000 VN.n6437 VN.n6436 0.004
R10001 VN.n6968 VN.n6967 0.004
R10002 VN.n6882 VN.n6881 0.004
R10003 VN.n7781 VN.n7780 0.004
R10004 VN.n8073 VN.n8072 0.004
R10005 VN.n8629 VN.n8628 0.004
R10006 VN.n8637 VN.n8636 0.004
R10007 VN.n9017 VN.n9016 0.004
R10008 VN.n8925 VN.n8924 0.004
R10009 VN.n8961 VN.n8960 0.004
R10010 VN.n12433 VN.n12432 0.004
R10011 VN.n12674 VN.n12673 0.004
R10012 VN.n12682 VN.n12681 0.004
R10013 VN.n314 VN.n313 0.004
R10014 VN.n585 VN.n584 0.004
R10015 VN.n986 VN.n985 0.004
R10016 VN.n1260 VN.n1259 0.004
R10017 VN.n1673 VN.n1672 0.004
R10018 VN.n1950 VN.n1949 0.004
R10019 VN.n2381 VN.n2380 0.004
R10020 VN.n2659 VN.n2658 0.004
R10021 VN.n3100 VN.n3099 0.004
R10022 VN.n3381 VN.n3380 0.004
R10023 VN.n3843 VN.n3842 0.004
R10024 VN.n4125 VN.n4124 0.004
R10025 VN.n4597 VN.n4596 0.004
R10026 VN.n4882 VN.n4881 0.004
R10027 VN.n5375 VN.n5374 0.004
R10028 VN.n5661 VN.n5660 0.004
R10029 VN.n6164 VN.n6163 0.004
R10030 VN.n6453 VN.n6452 0.004
R10031 VN.n6953 VN.n6952 0.004
R10032 VN.n6898 VN.n6897 0.004
R10033 VN.n7796 VN.n7795 0.004
R10034 VN.n7804 VN.n7803 0.004
R10035 VN.n8184 VN.n8183 0.004
R10036 VN.n8092 VN.n8091 0.004
R10037 VN.n8128 VN.n8127 0.004
R10038 VN.n12449 VN.n12448 0.004
R10039 VN.n12785 VN.n12784 0.004
R10040 VN.n12796 VN.n12795 0.004
R10041 VN.n329 VN.n328 0.004
R10042 VN.n601 VN.n600 0.004
R10043 VN.n1001 VN.n1000 0.004
R10044 VN.n1276 VN.n1275 0.004
R10045 VN.n1688 VN.n1687 0.004
R10046 VN.n1966 VN.n1965 0.004
R10047 VN.n2396 VN.n2395 0.004
R10048 VN.n2675 VN.n2674 0.004
R10049 VN.n3115 VN.n3114 0.004
R10050 VN.n3397 VN.n3396 0.004
R10051 VN.n3858 VN.n3857 0.004
R10052 VN.n4141 VN.n4140 0.004
R10053 VN.n4612 VN.n4611 0.004
R10054 VN.n4898 VN.n4897 0.004
R10055 VN.n5390 VN.n5389 0.004
R10056 VN.n5677 VN.n5676 0.004
R10057 VN.n6179 VN.n6178 0.004
R10058 VN.n6469 VN.n6468 0.004
R10059 VN.n6623 VN.n6622 0.004
R10060 VN.n6631 VN.n6630 0.004
R10061 VN.n7373 VN.n7372 0.004
R10062 VN.n6917 VN.n6916 0.004
R10063 VN.n6608 VN.n6607 0.004
R10064 VN.n12465 VN.n12464 0.004
R10065 VN.n12816 VN.n12815 0.004
R10066 VN.n12827 VN.n12826 0.004
R10067 VN.n344 VN.n343 0.004
R10068 VN.n617 VN.n616 0.004
R10069 VN.n1016 VN.n1015 0.004
R10070 VN.n1292 VN.n1291 0.004
R10071 VN.n1703 VN.n1702 0.004
R10072 VN.n1982 VN.n1981 0.004
R10073 VN.n2411 VN.n2410 0.004
R10074 VN.n2691 VN.n2690 0.004
R10075 VN.n3130 VN.n3129 0.004
R10076 VN.n3413 VN.n3412 0.004
R10077 VN.n3873 VN.n3872 0.004
R10078 VN.n4157 VN.n4156 0.004
R10079 VN.n4627 VN.n4626 0.004
R10080 VN.n4914 VN.n4913 0.004
R10081 VN.n5405 VN.n5404 0.004
R10082 VN.n5693 VN.n5692 0.004
R10083 VN.n6194 VN.n6193 0.004
R10084 VN.n6202 VN.n6201 0.004
R10085 VN.n6580 VN.n6579 0.004
R10086 VN.n6488 VN.n6487 0.004
R10087 VN.n6524 VN.n6523 0.004
R10088 VN.n12481 VN.n12480 0.004
R10089 VN.n12847 VN.n12846 0.004
R10090 VN.n12855 VN.n12854 0.004
R10091 VN.n359 VN.n358 0.004
R10092 VN.n633 VN.n632 0.004
R10093 VN.n1031 VN.n1030 0.004
R10094 VN.n1308 VN.n1307 0.004
R10095 VN.n1718 VN.n1717 0.004
R10096 VN.n1998 VN.n1997 0.004
R10097 VN.n2426 VN.n2425 0.004
R10098 VN.n2707 VN.n2706 0.004
R10099 VN.n3145 VN.n3144 0.004
R10100 VN.n3429 VN.n3428 0.004
R10101 VN.n3888 VN.n3887 0.004
R10102 VN.n4173 VN.n4172 0.004
R10103 VN.n4642 VN.n4641 0.004
R10104 VN.n4930 VN.n4929 0.004
R10105 VN.n5420 VN.n5419 0.004
R10106 VN.n5428 VN.n5427 0.004
R10107 VN.n5804 VN.n5803 0.004
R10108 VN.n5712 VN.n5711 0.004
R10109 VN.n5748 VN.n5747 0.004
R10110 VN.n12497 VN.n12496 0.004
R10111 VN.n12878 VN.n12877 0.004
R10112 VN.n12886 VN.n12885 0.004
R10113 VN.n374 VN.n373 0.004
R10114 VN.n649 VN.n648 0.004
R10115 VN.n1046 VN.n1045 0.004
R10116 VN.n1324 VN.n1323 0.004
R10117 VN.n1733 VN.n1732 0.004
R10118 VN.n2014 VN.n2013 0.004
R10119 VN.n2441 VN.n2440 0.004
R10120 VN.n2723 VN.n2722 0.004
R10121 VN.n3160 VN.n3159 0.004
R10122 VN.n3445 VN.n3444 0.004
R10123 VN.n3903 VN.n3902 0.004
R10124 VN.n4189 VN.n4188 0.004
R10125 VN.n4657 VN.n4656 0.004
R10126 VN.n4665 VN.n4664 0.004
R10127 VN.n5041 VN.n5040 0.004
R10128 VN.n4949 VN.n4948 0.004
R10129 VN.n4985 VN.n4984 0.004
R10130 VN.n12513 VN.n12512 0.004
R10131 VN.n12909 VN.n12908 0.004
R10132 VN.n12917 VN.n12916 0.004
R10133 VN.n389 VN.n388 0.004
R10134 VN.n665 VN.n664 0.004
R10135 VN.n1061 VN.n1060 0.004
R10136 VN.n1340 VN.n1339 0.004
R10137 VN.n1748 VN.n1747 0.004
R10138 VN.n2030 VN.n2029 0.004
R10139 VN.n2456 VN.n2455 0.004
R10140 VN.n2739 VN.n2738 0.004
R10141 VN.n3175 VN.n3174 0.004
R10142 VN.n3461 VN.n3460 0.004
R10143 VN.n3918 VN.n3917 0.004
R10144 VN.n3926 VN.n3925 0.004
R10145 VN.n4300 VN.n4299 0.004
R10146 VN.n4208 VN.n4207 0.004
R10147 VN.n4244 VN.n4243 0.004
R10148 VN.n12529 VN.n12528 0.004
R10149 VN.n12940 VN.n12939 0.004
R10150 VN.n12948 VN.n12947 0.004
R10151 VN.n404 VN.n403 0.004
R10152 VN.n681 VN.n680 0.004
R10153 VN.n1076 VN.n1075 0.004
R10154 VN.n1356 VN.n1355 0.004
R10155 VN.n1763 VN.n1762 0.004
R10156 VN.n2046 VN.n2045 0.004
R10157 VN.n2471 VN.n2470 0.004
R10158 VN.n2755 VN.n2754 0.004
R10159 VN.n3190 VN.n3189 0.004
R10160 VN.n3198 VN.n3197 0.004
R10161 VN.n3572 VN.n3571 0.004
R10162 VN.n3480 VN.n3479 0.004
R10163 VN.n3516 VN.n3515 0.004
R10164 VN.n12545 VN.n12544 0.004
R10165 VN.n12971 VN.n12970 0.004
R10166 VN.n12979 VN.n12978 0.004
R10167 VN.n419 VN.n418 0.004
R10168 VN.n697 VN.n696 0.004
R10169 VN.n1091 VN.n1090 0.004
R10170 VN.n1372 VN.n1371 0.004
R10171 VN.n1778 VN.n1777 0.004
R10172 VN.n2062 VN.n2061 0.004
R10173 VN.n2486 VN.n2485 0.004
R10174 VN.n2494 VN.n2493 0.004
R10175 VN.n2866 VN.n2865 0.004
R10176 VN.n2774 VN.n2773 0.004
R10177 VN.n2810 VN.n2809 0.004
R10178 VN.n12561 VN.n12560 0.004
R10179 VN.n13002 VN.n13001 0.004
R10180 VN.n13010 VN.n13009 0.004
R10181 VN.n434 VN.n433 0.004
R10182 VN.n713 VN.n712 0.004
R10183 VN.n1106 VN.n1105 0.004
R10184 VN.n1388 VN.n1387 0.004
R10185 VN.n1793 VN.n1792 0.004
R10186 VN.n1801 VN.n1800 0.004
R10187 VN.n2173 VN.n2172 0.004
R10188 VN.n2081 VN.n2080 0.004
R10189 VN.n2117 VN.n2116 0.004
R10190 VN.n12577 VN.n12576 0.004
R10191 VN.n13033 VN.n13032 0.004
R10192 VN.n13041 VN.n13040 0.004
R10193 VN.n449 VN.n448 0.004
R10194 VN.n729 VN.n728 0.004
R10195 VN.n1121 VN.n1120 0.004
R10196 VN.n1129 VN.n1128 0.004
R10197 VN.n1499 VN.n1498 0.004
R10198 VN.n1407 VN.n1406 0.004
R10199 VN.n1443 VN.n1442 0.004
R10200 VN.n12593 VN.n12592 0.004
R10201 VN.n13064 VN.n13063 0.004
R10202 VN.n13072 VN.n13071 0.004
R10203 VN.n464 VN.n463 0.004
R10204 VN.n472 VN.n471 0.004
R10205 VN.n849 VN.n848 0.004
R10206 VN.n746 VN.n745 0.004
R10207 VN.n791 VN.n790 0.004
R10208 VN.n12612 VN.n12611 0.004
R10209 VN.n13102 VN.n13101 0.004
R10210 VN.n12754 VN.n12753 0.004
R10211 VN.n199 VN.n198 0.004
R10212 VN.n12383 VN.n12382 0.004
R10213 VN.n12231 VN.n12230 0.004
R10214 VN.n12728 VN.n12727 0.004
R10215 VN.n12401 VN.n12400 0.004
R10216 VN.n11548 VN.n11547 0.004
R10217 VN.t8 VN.n11695 0.004
R10218 VN.n12165 VN.n12152 0.004
R10219 VN.n12036 VN.n12035 0.004
R10220 VN.n12059 VN.n12058 0.004
R10221 VN.n11991 VN.n11990 0.004
R10222 VN.n12014 VN.n12013 0.004
R10223 VN.n11946 VN.n11945 0.004
R10224 VN.n11969 VN.n11968 0.004
R10225 VN.n11897 VN.n11896 0.004
R10226 VN.n11639 VN.n11638 0.004
R10227 VN.n11876 VN.n11875 0.004
R10228 VN.n11594 VN.n11593 0.004
R10229 VN.n11617 VN.n11616 0.004
R10230 VN.t8 VN.n11682 0.004
R10231 VN.n1142 VN.n1141 0.004
R10232 VN.n11379 VN.n11378 0.004
R10233 VN.n1517 VN.n1516 0.004
R10234 VN.n2225 VN.n2224 0.004
R10235 VN.n2947 VN.n2946 0.004
R10236 VN.n3687 VN.n3686 0.004
R10237 VN.n4444 VN.n4443 0.004
R10238 VN.n5219 VN.n5218 0.004
R10239 VN.n6011 VN.n6010 0.004
R10240 VN.n7254 VN.n7253 0.004
R10241 VN.n7643 VN.n7642 0.004
R10242 VN.n8488 VN.n8487 0.004
R10243 VN.n9350 VN.n9349 0.004
R10244 VN.n10233 VN.n10232 0.004
R10245 VN.n11078 VN.n11077 0.004
R10246 VN.n12089 VN.n12088 0.004
R10247 VN.n12366 VN.n12365 0.004
R10248 VN.n1142 VN.n1140 0.004
R10249 VN.n11138 VN.n11126 0.004
R10250 VN.n10609 VN.n10608 0.004
R10251 VN.n9722 VN.n9711 0.004
R10252 VN.n8860 VN.n8849 0.004
R10253 VN.n8011 VN.n8000 0.004
R10254 VN.n6820 VN.n6809 0.004
R10255 VN.n6375 VN.n6364 0.004
R10256 VN.n5583 VN.n5572 0.004
R10257 VN.n4804 VN.n4793 0.004
R10258 VN.n4047 VN.n4036 0.004
R10259 VN.n3303 VN.n3292 0.004
R10260 VN.n2581 VN.n2570 0.004
R10261 VN.n1872 VN.n1861 0.004
R10262 VN.n1182 VN.n1171 0.004
R10263 VN.n507 VN.n496 0.004
R10264 VN.n12697 VN.n12695 0.004
R10265 VN.n1815 VN.n1814 0.004
R10266 VN.n11172 VN.n11163 0.004
R10267 VN.n2507 VN.n2505 0.004
R10268 VN.n3212 VN.n3211 0.004
R10269 VN.n11206 VN.n11197 0.004
R10270 VN.n3939 VN.n3937 0.004
R10271 VN.n4679 VN.n4678 0.004
R10272 VN.n11240 VN.n11231 0.004
R10273 VN.n5441 VN.n5439 0.004
R10274 VN.n6216 VN.n6213 0.004
R10275 VN.n6644 VN.n6642 0.004
R10276 VN.n7818 VN.n7817 0.004
R10277 VN.n11307 VN.n11298 0.004
R10278 VN.n8650 VN.n8648 0.004
R10279 VN.n9495 VN.n9494 0.004
R10280 VN.n11341 VN.n11332 0.004
R10281 VN.n10351 VN.n10349 0.004
R10282 VN.n11379 VN.n11376 0.004
R10283 VN.n11273 VN.n11264 0.004
R10284 VN.n10437 VN.n10428 0.004
R10285 VN.n9562 VN.n9553 0.004
R10286 VN.n8700 VN.n8691 0.004
R10287 VN.n7851 VN.n7842 0.004
R10288 VN.n6660 VN.n6651 0.004
R10289 VN.n11060 VN.n11059 0.004
R10290 VN.n2180 VN.n2179 0.004
R10291 VN.n2902 VN.n2901 0.004
R10292 VN.n3642 VN.n3641 0.004
R10293 VN.n4399 VN.n4398 0.004
R10294 VN.n5174 VN.n5173 0.004
R10295 VN.n5966 VN.n5965 0.004
R10296 VN.n7209 VN.n7208 0.004
R10297 VN.n7598 VN.n7597 0.004
R10298 VN.n8443 VN.n8442 0.004
R10299 VN.n9305 VN.n9304 0.004
R10300 VN.n10188 VN.n10187 0.004
R10301 VN.n489 VN.n476 0.004
R10302 VN.n1525 VN.n1523 0.004
R10303 VN.n2233 VN.n2231 0.004
R10304 VN.n2955 VN.n2953 0.004
R10305 VN.n3695 VN.n3693 0.004
R10306 VN.n4452 VN.n4450 0.004
R10307 VN.n5227 VN.n5225 0.004
R10308 VN.n6019 VN.n6017 0.004
R10309 VN.n7262 VN.n7260 0.004
R10310 VN.n7651 VN.n7649 0.004
R10311 VN.n8496 VN.n8494 0.004
R10312 VN.n9358 VN.n9356 0.004
R10313 VN.n10241 VN.n10239 0.004
R10314 VN.n11086 VN.n11084 0.004
R10315 VN.n10566 VN.n10565 0.004
R10316 VN.n2320 VN.n2319 0.004
R10317 VN.n1815 VN.n1803 0.004
R10318 VN.n3782 VN.n3781 0.004
R10319 VN.n3212 VN.n3200 0.004
R10320 VN.n5314 VN.n5313 0.004
R10321 VN.n4679 VN.n4667 0.004
R10322 VN.t76 VN.n6601 0.004
R10323 VN.n6216 VN.n6215 0.004
R10324 VN.n8583 VN.n8582 0.004
R10325 VN.n7818 VN.n7806 0.004
R10326 VN.n10328 VN.n10327 0.004
R10327 VN.n9495 VN.n9483 0.004
R10328 VN.n9844 VN.n9832 0.004
R10329 VN.n10707 VN.n9844 0.004
R10330 VN.n8998 VN.n8986 0.004
R10331 VN.n9827 VN.n8998 0.004
R10332 VN.n8165 VN.n8153 0.004
R10333 VN.n8981 VN.n8165 0.004
R10334 VN.n7354 VN.n7342 0.004
R10335 VN.n8148 VN.n7354 0.004
R10336 VN.n6561 VN.n6549 0.004
R10337 VN.n7337 VN.n6561 0.004
R10338 VN.n5785 VN.n5773 0.004
R10339 VN.n6544 VN.n5785 0.004
R10340 VN.n5022 VN.n5010 0.004
R10341 VN.n5768 VN.n5022 0.004
R10342 VN.n4281 VN.n4269 0.004
R10343 VN.n5005 VN.n4281 0.004
R10344 VN.n3553 VN.n3541 0.004
R10345 VN.n4264 VN.n3553 0.004
R10346 VN.n2847 VN.n2835 0.004
R10347 VN.n3536 VN.n2847 0.004
R10348 VN.n2154 VN.n2142 0.004
R10349 VN.n2830 VN.n2154 0.004
R10350 VN.n1480 VN.n1468 0.004
R10351 VN.n2137 VN.n1480 0.004
R10352 VN.n12747 VN.n12745 0.004
R10353 VN.n830 VN.n829 0.004
R10354 VN.n1463 VN.n825 0.004
R10355 VN.t51 VN.n72 0.004
R10356 VN.t51 VN.n69 0.004
R10357 VN.t51 VN.n66 0.004
R10358 VN.t51 VN.n63 0.004
R10359 VN.t51 VN.n60 0.004
R10360 VN.t51 VN.n57 0.004
R10361 VN.t51 VN.n54 0.004
R10362 VN.t51 VN.n51 0.004
R10363 VN.t51 VN.n48 0.004
R10364 VN.t51 VN.n45 0.004
R10365 VN.t51 VN.n42 0.004
R10366 VN.t51 VN.n39 0.004
R10367 VN.t51 VN.n36 0.004
R10368 VN.t51 VN.n34 0.004
R10369 VN.n11575 VN.n11574 0.004
R10370 VN.t8 VN.n11676 0.004
R10371 VN.t82 VN.n12369 0.004
R10372 VN.t8 VN.n11722 0.004
R10373 VN.t57 VN.n2510 0.004
R10374 VN.t8 VN.n11858 0.004
R10375 VN.t108 VN.n1818 0.004
R10376 VN.t8 VN.n11711 0.004
R10377 VN.t94 VN.n1145 0.004
R10378 VN.t8 VN.n11698 0.004
R10379 VN.t41 VN.n492 0.004
R10380 VN.t101 VN.n12700 0.004
R10381 VN.t8 VN.n11685 0.004
R10382 VN.t8 VN.n11733 0.004
R10383 VN.t28 VN.n3942 0.004
R10384 VN.t8 VN.n11834 0.004
R10385 VN.t183 VN.n3215 0.004
R10386 VN.t8 VN.n11744 0.004
R10387 VN.t176 VN.n5444 0.004
R10388 VN.t8 VN.n11823 0.004
R10389 VN.t32 VN.n4682 0.004
R10390 VN.t146 VN.n6219 0.004
R10391 VN.t8 VN.n11861 0.004
R10392 VN.t8 VN.n11755 0.004
R10393 VN.t253 VN.n6647 0.004
R10394 VN.t8 VN.n11766 0.004
R10395 VN.t39 VN.n8653 0.004
R10396 VN.t8 VN.n11812 0.004
R10397 VN.t73 VN.n7821 0.004
R10398 VN.t8 VN.n11775 0.004
R10399 VN.t241 VN.n10354 0.004
R10400 VN.t8 VN.n11801 0.004
R10401 VN.t0 VN.n9498 0.004
R10402 VN.t51 VN.n168 0.004
R10403 VN.t51 VN.n102 0.004
R10404 VN.t51 VN.n106 0.004
R10405 VN.t51 VN.n110 0.004
R10406 VN.t51 VN.n114 0.004
R10407 VN.t51 VN.n118 0.004
R10408 VN.t51 VN.n122 0.004
R10409 VN.t51 VN.n126 0.004
R10410 VN.t51 VN.n130 0.004
R10411 VN.t51 VN.n134 0.004
R10412 VN.t51 VN.n138 0.004
R10413 VN.t51 VN.n142 0.004
R10414 VN.t51 VN.n146 0.004
R10415 VN.t51 VN.n150 0.004
R10416 VN.t51 VN.n154 0.004
R10417 VN.t51 VN.n158 0.004
R10418 VN.t51 VN.n162 0.004
R10419 VN.t51 VN.n166 0.004
R10420 VN.t8 VN.n11668 0.004
R10421 VN.t51 VN.n83 0.004
R10422 VN.t76 VN.n6582 0.004
R10423 VN.t35 VN.n11382 0.004
R10424 VN.t8 VN.n11666 0.004
R10425 VN.t8 VN.n11855 0.004
R10426 VN.t8 VN.n11831 0.004
R10427 VN.t8 VN.n11820 0.004
R10428 VN.t8 VN.n11809 0.004
R10429 VN.t8 VN.n11798 0.004
R10430 VN.t8 VN.n11660 0.004
R10431 VN.n11154 VN.n11153 0.004
R10432 VN.t8 VN.n11673 0.004
R10433 VN.t8 VN.n11716 0.004
R10434 VN.t8 VN.n11727 0.004
R10435 VN.t8 VN.n11738 0.004
R10436 VN.t8 VN.n11749 0.004
R10437 VN.t8 VN.n11760 0.004
R10438 VN.t8 VN.n11769 0.004
R10439 VN.n12697 VN.n12696 0.004
R10440 VN.n1831 VN.n1822 0.004
R10441 VN.n2540 VN.n2531 0.004
R10442 VN.n3262 VN.n3253 0.004
R10443 VN.n4006 VN.n3997 0.004
R10444 VN.n4763 VN.n4754 0.004
R10445 VN.n5542 VN.n5533 0.004
R10446 VN.n6334 VN.n6325 0.004
R10447 VN.n6779 VN.n6770 0.004
R10448 VN.n7970 VN.n7961 0.004
R10449 VN.n8819 VN.n8810 0.004
R10450 VN.n9681 VN.n9672 0.004
R10451 VN.n12408 VN.n12407 0.003
R10452 VN.n11578 VN.n11577 0.003
R10453 VN.n12411 VN.n12410 0.003
R10454 VN.n13113 VN.n13112 0.003
R10455 VN.n12171 VN.n12170 0.003
R10456 VN.n12262 VN.n12261 0.003
R10457 VN.n12719 VN.n12718 0.003
R10458 VN.n233 VN.n232 0.003
R10459 VN.n530 VN.n529 0.003
R10460 VN.n904 VN.n903 0.003
R10461 VN.n1205 VN.n1204 0.003
R10462 VN.n1587 VN.n1586 0.003
R10463 VN.n1895 VN.n1894 0.003
R10464 VN.n2295 VN.n2294 0.003
R10465 VN.n2604 VN.n2603 0.003
R10466 VN.n3017 VN.n3016 0.003
R10467 VN.n3326 VN.n3325 0.003
R10468 VN.n3757 VN.n3756 0.003
R10469 VN.n4070 VN.n4069 0.003
R10470 VN.n4514 VN.n4513 0.003
R10471 VN.n4827 VN.n4826 0.003
R10472 VN.n5289 VN.n5288 0.003
R10473 VN.n5606 VN.n5605 0.003
R10474 VN.n6081 VN.n6080 0.003
R10475 VN.n6398 VN.n6397 0.003
R10476 VN.n7324 VN.n7323 0.003
R10477 VN.n6843 VN.n6842 0.003
R10478 VN.n7713 VN.n7712 0.003
R10479 VN.n8034 VN.n8033 0.003
R10480 VN.n8558 VN.n8557 0.003
R10481 VN.n8883 VN.n8882 0.003
R10482 VN.n9420 VN.n9419 0.003
R10483 VN.n9745 VN.n9744 0.003
R10484 VN.n10303 VN.n10302 0.003
R10485 VN.n10633 VN.n10632 0.003
R10486 VN.n11471 VN.n11470 0.003
R10487 VN.n11121 VN.n11120 0.003
R10488 VN.n12042 VN.n12041 0.003
R10489 VN.n3042 VN.n3041 0.003
R10490 VN.n3234 VN.n3233 0.003
R10491 VN.n3606 VN.n3605 0.003
R10492 VN.n3978 VN.n3977 0.003
R10493 VN.n4363 VN.n4362 0.003
R10494 VN.n4735 VN.n4734 0.003
R10495 VN.n5138 VN.n5137 0.003
R10496 VN.n5514 VN.n5513 0.003
R10497 VN.n5930 VN.n5929 0.003
R10498 VN.n6306 VN.n6305 0.003
R10499 VN.n7173 VN.n7172 0.003
R10500 VN.n6751 VN.n6750 0.003
R10501 VN.n7562 VN.n7561 0.003
R10502 VN.n7942 VN.n7941 0.003
R10503 VN.n8407 VN.n8406 0.003
R10504 VN.n8791 VN.n8790 0.003
R10505 VN.n9269 VN.n9268 0.003
R10506 VN.n9653 VN.n9652 0.003
R10507 VN.n10151 VN.n10150 0.003
R10508 VN.n10531 VN.n10530 0.003
R10509 VN.n11015 VN.n11014 0.003
R10510 VN.n11191 VN.n11190 0.003
R10511 VN.n12065 VN.n12064 0.003
R10512 VN.n2323 VN.n2322 0.003
R10513 VN.n2529 VN.n2528 0.003
R10514 VN.n2895 VN.n2894 0.003
R10515 VN.n3251 VN.n3250 0.003
R10516 VN.n3635 VN.n3634 0.003
R10517 VN.n3995 VN.n3994 0.003
R10518 VN.n4392 VN.n4391 0.003
R10519 VN.n4752 VN.n4751 0.003
R10520 VN.n5167 VN.n5166 0.003
R10521 VN.n5531 VN.n5530 0.003
R10522 VN.n5959 VN.n5958 0.003
R10523 VN.n6323 VN.n6322 0.003
R10524 VN.n7202 VN.n7201 0.003
R10525 VN.n6768 VN.n6767 0.003
R10526 VN.n7591 VN.n7590 0.003
R10527 VN.n7959 VN.n7958 0.003
R10528 VN.n8436 VN.n8435 0.003
R10529 VN.n8808 VN.n8807 0.003
R10530 VN.n9298 VN.n9297 0.003
R10531 VN.n9670 VN.n9669 0.003
R10532 VN.n10180 VN.n10179 0.003
R10533 VN.n10551 VN.n10550 0.003
R10534 VN.n10572 VN.n10571 0.003
R10535 VN.n11075 VN.n11074 0.003
R10536 VN.n11157 VN.n11156 0.003
R10537 VN.n12087 VN.n12086 0.003
R10538 VN.n10215 VN.n10214 0.003
R10539 VN.n9332 VN.n9331 0.003
R10540 VN.n8470 VN.n8469 0.003
R10541 VN.n7625 VN.n7624 0.003
R10542 VN.n7236 VN.n7235 0.003
R10543 VN.n5993 VN.n5992 0.003
R10544 VN.n5201 VN.n5200 0.003
R10545 VN.n4426 VN.n4425 0.003
R10546 VN.n3669 VN.n3668 0.003
R10547 VN.n2929 VN.n2928 0.003
R10548 VN.n2207 VN.n2206 0.003
R10549 VN.n1615 VN.n1614 0.003
R10550 VN.n1837 VN.n1836 0.003
R10551 VN.n2546 VN.n2545 0.003
R10552 VN.n3268 VN.n3267 0.003
R10553 VN.n4012 VN.n4011 0.003
R10554 VN.n4769 VN.n4768 0.003
R10555 VN.n5548 VN.n5547 0.003
R10556 VN.n6340 VN.n6339 0.003
R10557 VN.n6785 VN.n6784 0.003
R10558 VN.n7976 VN.n7975 0.003
R10559 VN.n8825 VN.n8824 0.003
R10560 VN.n9687 VN.n9686 0.003
R10561 VN.n11420 VN.n11419 0.003
R10562 VN.n11385 VN.n11384 0.003
R10563 VN.n12121 VN.n12120 0.003
R10564 VN.n928 VN.n927 0.003
R10565 VN.n1169 VN.n1168 0.003
R10566 VN.n1532 VN.n1531 0.003
R10567 VN.n1859 VN.n1858 0.003
R10568 VN.n2240 VN.n2239 0.003
R10569 VN.n2568 VN.n2567 0.003
R10570 VN.n2962 VN.n2961 0.003
R10571 VN.n3290 VN.n3289 0.003
R10572 VN.n3702 VN.n3701 0.003
R10573 VN.n4034 VN.n4033 0.003
R10574 VN.n4459 VN.n4458 0.003
R10575 VN.n4791 VN.n4790 0.003
R10576 VN.n5234 VN.n5233 0.003
R10577 VN.n5570 VN.n5569 0.003
R10578 VN.n6026 VN.n6025 0.003
R10579 VN.n6362 VN.n6361 0.003
R10580 VN.n7269 VN.n7268 0.003
R10581 VN.n6807 VN.n6806 0.003
R10582 VN.n7658 VN.n7657 0.003
R10583 VN.n7998 VN.n7997 0.003
R10584 VN.n8503 VN.n8502 0.003
R10585 VN.n8847 VN.n8846 0.003
R10586 VN.n9365 VN.n9364 0.003
R10587 VN.n9709 VN.n9708 0.003
R10588 VN.n10248 VN.n10247 0.003
R10589 VN.n10594 VN.n10593 0.003
R10590 VN.n11447 VN.n11446 0.003
R10591 VN.n11141 VN.n11140 0.003
R10592 VN.n10615 VN.n10614 0.003
R10593 VN.n10269 VN.n10268 0.003
R10594 VN.n9728 VN.n9727 0.003
R10595 VN.n9386 VN.n9385 0.003
R10596 VN.n8866 VN.n8865 0.003
R10597 VN.n8524 VN.n8523 0.003
R10598 VN.n8017 VN.n8016 0.003
R10599 VN.n7679 VN.n7678 0.003
R10600 VN.n6826 VN.n6825 0.003
R10601 VN.n7290 VN.n7289 0.003
R10602 VN.n6381 VN.n6380 0.003
R10603 VN.n6047 VN.n6046 0.003
R10604 VN.n5589 VN.n5588 0.003
R10605 VN.n5255 VN.n5254 0.003
R10606 VN.n4810 VN.n4809 0.003
R10607 VN.n4480 VN.n4479 0.003
R10608 VN.n4053 VN.n4052 0.003
R10609 VN.n3723 VN.n3722 0.003
R10610 VN.n3309 VN.n3308 0.003
R10611 VN.n2983 VN.n2982 0.003
R10612 VN.n2587 VN.n2586 0.003
R10613 VN.n2261 VN.n2260 0.003
R10614 VN.n1878 VN.n1877 0.003
R10615 VN.n1553 VN.n1552 0.003
R10616 VN.n1188 VN.n1187 0.003
R10617 VN.n870 VN.n869 0.003
R10618 VN.n513 VN.n512 0.003
R10619 VN.n256 VN.n255 0.003
R10620 VN.n12150 VN.n12149 0.003
R10621 VN.n11042 VN.n11041 0.003
R10622 VN.n11175 VN.n11174 0.003
R10623 VN.n11997 VN.n11996 0.003
R10624 VN.n4539 VN.n4538 0.003
R10625 VN.n4701 VN.n4700 0.003
R10626 VN.n5075 VN.n5074 0.003
R10627 VN.n5480 VN.n5479 0.003
R10628 VN.n5867 VN.n5866 0.003
R10629 VN.n6272 VN.n6271 0.003
R10630 VN.n7110 VN.n7109 0.003
R10631 VN.n6717 VN.n6716 0.003
R10632 VN.n7499 VN.n7498 0.003
R10633 VN.n7908 VN.n7907 0.003
R10634 VN.n8344 VN.n8343 0.003
R10635 VN.n8757 VN.n8756 0.003
R10636 VN.n9206 VN.n9205 0.003
R10637 VN.n9619 VN.n9618 0.003
R10638 VN.n10088 VN.n10087 0.003
R10639 VN.n10496 VN.n10495 0.003
R10640 VN.n10957 VN.n10956 0.003
R10641 VN.n11225 VN.n11224 0.003
R10642 VN.n12020 VN.n12019 0.003
R10643 VN.n3785 VN.n3784 0.003
R10644 VN.n3961 VN.n3960 0.003
R10645 VN.n4329 VN.n4328 0.003
R10646 VN.n4718 VN.n4717 0.003
R10647 VN.n5104 VN.n5103 0.003
R10648 VN.n5497 VN.n5496 0.003
R10649 VN.n5896 VN.n5895 0.003
R10650 VN.n6289 VN.n6288 0.003
R10651 VN.n7139 VN.n7138 0.003
R10652 VN.n6734 VN.n6733 0.003
R10653 VN.n7528 VN.n7527 0.003
R10654 VN.n7925 VN.n7924 0.003
R10655 VN.n8373 VN.n8372 0.003
R10656 VN.n8774 VN.n8773 0.003
R10657 VN.n9235 VN.n9234 0.003
R10658 VN.n9636 VN.n9635 0.003
R10659 VN.n10117 VN.n10116 0.003
R10660 VN.n10513 VN.n10512 0.003
R10661 VN.n10986 VN.n10985 0.003
R10662 VN.n11209 VN.n11208 0.003
R10663 VN.n11952 VN.n11951 0.003
R10664 VN.n6106 VN.n6105 0.003
R10665 VN.n6238 VN.n6237 0.003
R10666 VN.n7047 VN.n7046 0.003
R10667 VN.n6683 VN.n6682 0.003
R10668 VN.n7436 VN.n7435 0.003
R10669 VN.n7874 VN.n7873 0.003
R10670 VN.n8281 VN.n8280 0.003
R10671 VN.n8723 VN.n8722 0.003
R10672 VN.n9143 VN.n9142 0.003
R10673 VN.n9585 VN.n9584 0.003
R10674 VN.n10025 VN.n10024 0.003
R10675 VN.n10461 VN.n10460 0.003
R10676 VN.n10899 VN.n10898 0.003
R10677 VN.n11259 VN.n11258 0.003
R10678 VN.n11975 VN.n11974 0.003
R10679 VN.n5317 VN.n5316 0.003
R10680 VN.n5463 VN.n5462 0.003
R10681 VN.n5833 VN.n5832 0.003
R10682 VN.n6255 VN.n6254 0.003
R10683 VN.n7076 VN.n7075 0.003
R10684 VN.n6700 VN.n6699 0.003
R10685 VN.n7465 VN.n7464 0.003
R10686 VN.n7891 VN.n7890 0.003
R10687 VN.n8310 VN.n8309 0.003
R10688 VN.n8740 VN.n8739 0.003
R10689 VN.n9172 VN.n9171 0.003
R10690 VN.n9602 VN.n9601 0.003
R10691 VN.n10054 VN.n10053 0.003
R10692 VN.n10478 VN.n10477 0.003
R10693 VN.n10928 VN.n10927 0.003
R10694 VN.n11243 VN.n11242 0.003
R10695 VN.n6666 VN.n6665 0.003
R10696 VN.n7402 VN.n7401 0.003
R10697 VN.n7857 VN.n7856 0.003
R10698 VN.n8247 VN.n8246 0.003
R10699 VN.n8706 VN.n8705 0.003
R10700 VN.n9109 VN.n9108 0.003
R10701 VN.n9568 VN.n9567 0.003
R10702 VN.n9991 VN.n9990 0.003
R10703 VN.n10443 VN.n10442 0.003
R10704 VN.n10870 VN.n10869 0.003
R10705 VN.n11276 VN.n11275 0.003
R10706 VN.n11930 VN.n11929 0.003
R10707 VN.n11903 VN.n11902 0.003
R10708 VN.n7738 VN.n7737 0.003
R10709 VN.n7840 VN.n7839 0.003
R10710 VN.n8218 VN.n8217 0.003
R10711 VN.n8689 VN.n8688 0.003
R10712 VN.n9080 VN.n9079 0.003
R10713 VN.n9551 VN.n9550 0.003
R10714 VN.n9962 VN.n9961 0.003
R10715 VN.n10426 VN.n10425 0.003
R10716 VN.n10841 VN.n10840 0.003
R10717 VN.n11292 VN.n11291 0.003
R10718 VN.n11645 VN.n11644 0.003
R10719 VN.n9445 VN.n9444 0.003
R10720 VN.n9517 VN.n9516 0.003
R10721 VN.n9899 VN.n9898 0.003
R10722 VN.n10391 VN.n10390 0.003
R10723 VN.n10783 VN.n10782 0.003
R10724 VN.n11326 VN.n11325 0.003
R10725 VN.n11882 VN.n11881 0.003
R10726 VN.n8586 VN.n8585 0.003
R10727 VN.n8672 VN.n8671 0.003
R10728 VN.n9046 VN.n9045 0.003
R10729 VN.n9534 VN.n9533 0.003
R10730 VN.n9928 VN.n9927 0.003
R10731 VN.n10408 VN.n10407 0.003
R10732 VN.n10812 VN.n10811 0.003
R10733 VN.n11310 VN.n11309 0.003
R10734 VN.n11600 VN.n11599 0.003
R10735 VN.n11492 VN.n11491 0.003
R10736 VN.n11360 VN.n11359 0.003
R10737 VN.n11623 VN.n11622 0.003
R10738 VN.n10331 VN.n10330 0.003
R10739 VN.n10373 VN.n10372 0.003
R10740 VN.n10754 VN.n10753 0.003
R10741 VN.n11344 VN.n11343 0.003
R10742 VN.n12177 VN.n12176 0.003
R10743 VN.n11106 VN.n11105 0.003
R10744 VN.n11509 VN.n11508 0.003
R10745 VN.n10653 VN.n10652 0.003
R10746 VN.n10679 VN.n10678 0.003
R10747 VN.n9760 VN.n9759 0.003
R10748 VN.n9465 VN.n9464 0.003
R10749 VN.n8898 VN.n8897 0.003
R10750 VN.n8606 VN.n8605 0.003
R10751 VN.n8049 VN.n8048 0.003
R10752 VN.n7758 VN.n7757 0.003
R10753 VN.n6858 VN.n6857 0.003
R10754 VN.n7013 VN.n7012 0.003
R10755 VN.n6413 VN.n6412 0.003
R10756 VN.n6126 VN.n6125 0.003
R10757 VN.n5621 VN.n5620 0.003
R10758 VN.n5337 VN.n5336 0.003
R10759 VN.n4842 VN.n4841 0.003
R10760 VN.n4559 VN.n4558 0.003
R10761 VN.n4085 VN.n4084 0.003
R10762 VN.n3805 VN.n3804 0.003
R10763 VN.n3341 VN.n3340 0.003
R10764 VN.n3062 VN.n3061 0.003
R10765 VN.n2619 VN.n2618 0.003
R10766 VN.n2343 VN.n2342 0.003
R10767 VN.n1910 VN.n1909 0.003
R10768 VN.n1635 VN.n1634 0.003
R10769 VN.n1220 VN.n1219 0.003
R10770 VN.n948 VN.n947 0.003
R10771 VN.n545 VN.n544 0.003
R10772 VN.n276 VN.n275 0.003
R10773 VN.n12290 VN.n12289 0.003
R10774 VN.n12317 VN.n12316 0.003
R10775 VN.n12272 VN.n12271 0.003
R10776 VN.n11515 VN.n11514 0.003
R10777 VN.n10647 VN.n10646 0.003
R10778 VN.n10694 VN.n10693 0.003
R10779 VN.n12626 VN.n12625 0.003
R10780 VN.n12635 VN.n12634 0.003
R10781 VN.n12339 VN.n12338 0.003
R10782 VN.n291 VN.n290 0.003
R10783 VN.n561 VN.n560 0.003
R10784 VN.n963 VN.n962 0.003
R10785 VN.n1236 VN.n1235 0.003
R10786 VN.n1650 VN.n1649 0.003
R10787 VN.n1926 VN.n1925 0.003
R10788 VN.n2358 VN.n2357 0.003
R10789 VN.n2635 VN.n2634 0.003
R10790 VN.n3077 VN.n3076 0.003
R10791 VN.n3357 VN.n3356 0.003
R10792 VN.n3820 VN.n3819 0.003
R10793 VN.n4101 VN.n4100 0.003
R10794 VN.n4574 VN.n4573 0.003
R10795 VN.n4858 VN.n4857 0.003
R10796 VN.n5352 VN.n5351 0.003
R10797 VN.n5637 VN.n5636 0.003
R10798 VN.n6141 VN.n6140 0.003
R10799 VN.n6429 VN.n6428 0.003
R10800 VN.n6993 VN.n6992 0.003
R10801 VN.n6874 VN.n6873 0.003
R10802 VN.n7773 VN.n7772 0.003
R10803 VN.n8065 VN.n8064 0.003
R10804 VN.n8621 VN.n8620 0.003
R10805 VN.n8914 VN.n8913 0.003
R10806 VN.n9799 VN.n9798 0.003
R10807 VN.n9791 VN.n9790 0.003
R10808 VN.n10702 VN.n10701 0.003
R10809 VN.n9782 VN.n9781 0.003
R10810 VN.n9814 VN.n9813 0.003
R10811 VN.n12425 VN.n12424 0.003
R10812 VN.n12666 VN.n12665 0.003
R10813 VN.n12657 VN.n12656 0.003
R10814 VN.n306 VN.n305 0.003
R10815 VN.n577 VN.n576 0.003
R10816 VN.n978 VN.n977 0.003
R10817 VN.n1252 VN.n1251 0.003
R10818 VN.n1665 VN.n1664 0.003
R10819 VN.n1942 VN.n1941 0.003
R10820 VN.n2373 VN.n2372 0.003
R10821 VN.n2651 VN.n2650 0.003
R10822 VN.n3092 VN.n3091 0.003
R10823 VN.n3373 VN.n3372 0.003
R10824 VN.n3835 VN.n3834 0.003
R10825 VN.n4117 VN.n4116 0.003
R10826 VN.n4589 VN.n4588 0.003
R10827 VN.n4874 VN.n4873 0.003
R10828 VN.n5367 VN.n5366 0.003
R10829 VN.n5653 VN.n5652 0.003
R10830 VN.n6156 VN.n6155 0.003
R10831 VN.n6445 VN.n6444 0.003
R10832 VN.n6978 VN.n6977 0.003
R10833 VN.n6890 VN.n6889 0.003
R10834 VN.n7788 VN.n7787 0.003
R10835 VN.n8081 VN.n8080 0.003
R10836 VN.n8953 VN.n8952 0.003
R10837 VN.n8945 VN.n8944 0.003
R10838 VN.n9822 VN.n9821 0.003
R10839 VN.n8936 VN.n8935 0.003
R10840 VN.n8968 VN.n8967 0.003
R10841 VN.n12441 VN.n12440 0.003
R10842 VN.n12777 VN.n12776 0.003
R10843 VN.n12768 VN.n12767 0.003
R10844 VN.n321 VN.n320 0.003
R10845 VN.n593 VN.n592 0.003
R10846 VN.n993 VN.n992 0.003
R10847 VN.n1268 VN.n1267 0.003
R10848 VN.n1680 VN.n1679 0.003
R10849 VN.n1958 VN.n1957 0.003
R10850 VN.n2388 VN.n2387 0.003
R10851 VN.n2667 VN.n2666 0.003
R10852 VN.n3107 VN.n3106 0.003
R10853 VN.n3389 VN.n3388 0.003
R10854 VN.n3850 VN.n3849 0.003
R10855 VN.n4133 VN.n4132 0.003
R10856 VN.n4604 VN.n4603 0.003
R10857 VN.n4890 VN.n4889 0.003
R10858 VN.n5382 VN.n5381 0.003
R10859 VN.n5669 VN.n5668 0.003
R10860 VN.n6171 VN.n6170 0.003
R10861 VN.n6461 VN.n6460 0.003
R10862 VN.n6963 VN.n6962 0.003
R10863 VN.n6906 VN.n6905 0.003
R10864 VN.n8120 VN.n8119 0.003
R10865 VN.n8112 VN.n8111 0.003
R10866 VN.n8976 VN.n8975 0.003
R10867 VN.n8103 VN.n8102 0.003
R10868 VN.n8135 VN.n8134 0.003
R10869 VN.n12457 VN.n12456 0.003
R10870 VN.n12811 VN.n12810 0.003
R10871 VN.n12802 VN.n12801 0.003
R10872 VN.n336 VN.n335 0.003
R10873 VN.n609 VN.n608 0.003
R10874 VN.n1008 VN.n1007 0.003
R10875 VN.n1284 VN.n1283 0.003
R10876 VN.n1695 VN.n1694 0.003
R10877 VN.n1974 VN.n1973 0.003
R10878 VN.n2403 VN.n2402 0.003
R10879 VN.n2683 VN.n2682 0.003
R10880 VN.n3122 VN.n3121 0.003
R10881 VN.n3405 VN.n3404 0.003
R10882 VN.n3865 VN.n3864 0.003
R10883 VN.n4149 VN.n4148 0.003
R10884 VN.n4619 VN.n4618 0.003
R10885 VN.n4906 VN.n4905 0.003
R10886 VN.n5397 VN.n5396 0.003
R10887 VN.n5685 VN.n5684 0.003
R10888 VN.n6186 VN.n6185 0.003
R10889 VN.n6477 VN.n6476 0.003
R10890 VN.n6948 VN.n6947 0.003
R10891 VN.n6937 VN.n6936 0.003
R10892 VN.n8143 VN.n8142 0.003
R10893 VN.n6928 VN.n6927 0.003
R10894 VN.n6618 VN.n6617 0.003
R10895 VN.n12473 VN.n12472 0.003
R10896 VN.n12842 VN.n12841 0.003
R10897 VN.n12833 VN.n12832 0.003
R10898 VN.n351 VN.n350 0.003
R10899 VN.n625 VN.n624 0.003
R10900 VN.n1023 VN.n1022 0.003
R10901 VN.n1300 VN.n1299 0.003
R10902 VN.n1710 VN.n1709 0.003
R10903 VN.n1990 VN.n1989 0.003
R10904 VN.n2418 VN.n2417 0.003
R10905 VN.n2699 VN.n2698 0.003
R10906 VN.n3137 VN.n3136 0.003
R10907 VN.n3421 VN.n3420 0.003
R10908 VN.n3880 VN.n3879 0.003
R10909 VN.n4165 VN.n4164 0.003
R10910 VN.n4634 VN.n4633 0.003
R10911 VN.n4922 VN.n4921 0.003
R10912 VN.n5412 VN.n5411 0.003
R10913 VN.n5701 VN.n5700 0.003
R10914 VN.n6516 VN.n6515 0.003
R10915 VN.n6508 VN.n6507 0.003
R10916 VN.n7332 VN.n7331 0.003
R10917 VN.n6499 VN.n6498 0.003
R10918 VN.n6531 VN.n6530 0.003
R10919 VN.n12489 VN.n12488 0.003
R10920 VN.n12870 VN.n12869 0.003
R10921 VN.n12861 VN.n12860 0.003
R10922 VN.n366 VN.n365 0.003
R10923 VN.n641 VN.n640 0.003
R10924 VN.n1038 VN.n1037 0.003
R10925 VN.n1316 VN.n1315 0.003
R10926 VN.n1725 VN.n1724 0.003
R10927 VN.n2006 VN.n2005 0.003
R10928 VN.n2433 VN.n2432 0.003
R10929 VN.n2715 VN.n2714 0.003
R10930 VN.n3152 VN.n3151 0.003
R10931 VN.n3437 VN.n3436 0.003
R10932 VN.n3895 VN.n3894 0.003
R10933 VN.n4181 VN.n4180 0.003
R10934 VN.n4649 VN.n4648 0.003
R10935 VN.n4938 VN.n4937 0.003
R10936 VN.n5740 VN.n5739 0.003
R10937 VN.n5732 VN.n5731 0.003
R10938 VN.n6539 VN.n6538 0.003
R10939 VN.n5723 VN.n5722 0.003
R10940 VN.n5755 VN.n5754 0.003
R10941 VN.n12505 VN.n12504 0.003
R10942 VN.n12901 VN.n12900 0.003
R10943 VN.n12892 VN.n12891 0.003
R10944 VN.n381 VN.n380 0.003
R10945 VN.n657 VN.n656 0.003
R10946 VN.n1053 VN.n1052 0.003
R10947 VN.n1332 VN.n1331 0.003
R10948 VN.n1740 VN.n1739 0.003
R10949 VN.n2022 VN.n2021 0.003
R10950 VN.n2448 VN.n2447 0.003
R10951 VN.n2731 VN.n2730 0.003
R10952 VN.n3167 VN.n3166 0.003
R10953 VN.n3453 VN.n3452 0.003
R10954 VN.n3910 VN.n3909 0.003
R10955 VN.n4197 VN.n4196 0.003
R10956 VN.n4977 VN.n4976 0.003
R10957 VN.n4969 VN.n4968 0.003
R10958 VN.n5763 VN.n5762 0.003
R10959 VN.n4960 VN.n4959 0.003
R10960 VN.n4992 VN.n4991 0.003
R10961 VN.n12521 VN.n12520 0.003
R10962 VN.n12932 VN.n12931 0.003
R10963 VN.n12923 VN.n12922 0.003
R10964 VN.n396 VN.n395 0.003
R10965 VN.n673 VN.n672 0.003
R10966 VN.n1068 VN.n1067 0.003
R10967 VN.n1348 VN.n1347 0.003
R10968 VN.n1755 VN.n1754 0.003
R10969 VN.n2038 VN.n2037 0.003
R10970 VN.n2463 VN.n2462 0.003
R10971 VN.n2747 VN.n2746 0.003
R10972 VN.n3182 VN.n3181 0.003
R10973 VN.n3469 VN.n3468 0.003
R10974 VN.n4236 VN.n4235 0.003
R10975 VN.n4228 VN.n4227 0.003
R10976 VN.n5000 VN.n4999 0.003
R10977 VN.n4219 VN.n4218 0.003
R10978 VN.n4251 VN.n4250 0.003
R10979 VN.n12537 VN.n12536 0.003
R10980 VN.n12963 VN.n12962 0.003
R10981 VN.n12954 VN.n12953 0.003
R10982 VN.n411 VN.n410 0.003
R10983 VN.n689 VN.n688 0.003
R10984 VN.n1083 VN.n1082 0.003
R10985 VN.n1364 VN.n1363 0.003
R10986 VN.n1770 VN.n1769 0.003
R10987 VN.n2054 VN.n2053 0.003
R10988 VN.n2478 VN.n2477 0.003
R10989 VN.n2763 VN.n2762 0.003
R10990 VN.n3508 VN.n3507 0.003
R10991 VN.n3500 VN.n3499 0.003
R10992 VN.n4259 VN.n4258 0.003
R10993 VN.n3491 VN.n3490 0.003
R10994 VN.n3523 VN.n3522 0.003
R10995 VN.n12553 VN.n12552 0.003
R10996 VN.n12994 VN.n12993 0.003
R10997 VN.n12985 VN.n12984 0.003
R10998 VN.n426 VN.n425 0.003
R10999 VN.n705 VN.n704 0.003
R11000 VN.n1098 VN.n1097 0.003
R11001 VN.n1380 VN.n1379 0.003
R11002 VN.n1785 VN.n1784 0.003
R11003 VN.n2070 VN.n2069 0.003
R11004 VN.n2802 VN.n2801 0.003
R11005 VN.n2794 VN.n2793 0.003
R11006 VN.n3531 VN.n3530 0.003
R11007 VN.n2785 VN.n2784 0.003
R11008 VN.n2817 VN.n2816 0.003
R11009 VN.n12569 VN.n12568 0.003
R11010 VN.n13025 VN.n13024 0.003
R11011 VN.n13016 VN.n13015 0.003
R11012 VN.n441 VN.n440 0.003
R11013 VN.n721 VN.n720 0.003
R11014 VN.n1113 VN.n1112 0.003
R11015 VN.n1396 VN.n1395 0.003
R11016 VN.n2109 VN.n2108 0.003
R11017 VN.n2101 VN.n2100 0.003
R11018 VN.n2825 VN.n2824 0.003
R11019 VN.n2092 VN.n2091 0.003
R11020 VN.n2124 VN.n2123 0.003
R11021 VN.n12585 VN.n12584 0.003
R11022 VN.n13056 VN.n13055 0.003
R11023 VN.n13047 VN.n13046 0.003
R11024 VN.n456 VN.n455 0.003
R11025 VN.n737 VN.n736 0.003
R11026 VN.n1435 VN.n1434 0.003
R11027 VN.n1427 VN.n1426 0.003
R11028 VN.n2132 VN.n2131 0.003
R11029 VN.n1418 VN.n1417 0.003
R11030 VN.n1450 VN.n1449 0.003
R11031 VN.n12601 VN.n12600 0.003
R11032 VN.n13087 VN.n13086 0.003
R11033 VN.n13078 VN.n13077 0.003
R11034 VN.n775 VN.n774 0.003
R11035 VN.n767 VN.n766 0.003
R11036 VN.n1458 VN.n1457 0.003
R11037 VN.n758 VN.n757 0.003
R11038 VN.n797 VN.n796 0.003
R11039 VN.n12617 VN.n12616 0.003
R11040 VN.n13107 VN.n13106 0.003
R11041 VN.n12759 VN.n12758 0.003
R11042 VN.n805 VN.n804 0.003
R11043 VN.n12391 VN.n12390 0.003
R11044 VN.n12236 VN.n12235 0.003
R11045 VN.n12743 VN.n12742 0.003
R11046 VN.n10545 VN.n10544 0.003
R11047 VN.n12165 VN.n12158 0.003
R11048 VN.n12259 VN.n12245 0.003
R11049 VN.n12713 VN.n12710 0.003
R11050 VN.n227 VN.n216 0.003
R11051 VN.n524 VN.n521 0.003
R11052 VN.n898 VN.n887 0.003
R11053 VN.n1199 VN.n1196 0.003
R11054 VN.n1581 VN.n1570 0.003
R11055 VN.n1889 VN.n1886 0.003
R11056 VN.n2289 VN.n2278 0.003
R11057 VN.n2598 VN.n2595 0.003
R11058 VN.n3011 VN.n3000 0.003
R11059 VN.n3320 VN.n3317 0.003
R11060 VN.n3751 VN.n3740 0.003
R11061 VN.n4064 VN.n4061 0.003
R11062 VN.n4508 VN.n4497 0.003
R11063 VN.n4821 VN.n4818 0.003
R11064 VN.n5283 VN.n5272 0.003
R11065 VN.n5600 VN.n5597 0.003
R11066 VN.n6075 VN.n6064 0.003
R11067 VN.n6392 VN.n6389 0.003
R11068 VN.n7318 VN.n7307 0.003
R11069 VN.n6837 VN.n6834 0.003
R11070 VN.n7707 VN.n7696 0.003
R11071 VN.n8028 VN.n8025 0.003
R11072 VN.n8552 VN.n8541 0.003
R11073 VN.n8877 VN.n8874 0.003
R11074 VN.n9414 VN.n9403 0.003
R11075 VN.n9739 VN.n9736 0.003
R11076 VN.n10297 VN.n10286 0.003
R11077 VN.n10627 VN.n10623 0.003
R11078 VN.n11465 VN.n11455 0.003
R11079 VN.n11118 VN.n11115 0.003
R11080 VN.n12036 VN.n12031 0.003
R11081 VN.n3039 VN.n3026 0.003
R11082 VN.n3228 VN.n3225 0.003
R11083 VN.n3600 VN.n3589 0.003
R11084 VN.n3972 VN.n3969 0.003
R11085 VN.n4357 VN.n4346 0.003
R11086 VN.n4729 VN.n4726 0.003
R11087 VN.n5132 VN.n5121 0.003
R11088 VN.n5508 VN.n5505 0.003
R11089 VN.n5924 VN.n5913 0.003
R11090 VN.n6300 VN.n6297 0.003
R11091 VN.n7167 VN.n7156 0.003
R11092 VN.n6745 VN.n6742 0.003
R11093 VN.n7556 VN.n7545 0.003
R11094 VN.n7936 VN.n7933 0.003
R11095 VN.n8401 VN.n8390 0.003
R11096 VN.n8785 VN.n8782 0.003
R11097 VN.n9263 VN.n9252 0.003
R11098 VN.n9647 VN.n9644 0.003
R11099 VN.n10145 VN.n10134 0.003
R11100 VN.n10525 VN.n10521 0.003
R11101 VN.n11009 VN.n11003 0.003
R11102 VN.n11188 VN.n11185 0.003
R11103 VN.n12059 VN.n12054 0.003
R11104 VN.n2320 VN.n2308 0.003
R11105 VN.n2523 VN.n2518 0.003
R11106 VN.n2889 VN.n2875 0.003
R11107 VN.n3245 VN.n3240 0.003
R11108 VN.n3629 VN.n3615 0.003
R11109 VN.n3989 VN.n3984 0.003
R11110 VN.n4386 VN.n4372 0.003
R11111 VN.n4746 VN.n4741 0.003
R11112 VN.n5161 VN.n5147 0.003
R11113 VN.n5525 VN.n5520 0.003
R11114 VN.n5953 VN.n5939 0.003
R11115 VN.n6317 VN.n6312 0.003
R11116 VN.n7196 VN.n7182 0.003
R11117 VN.n6762 VN.n6757 0.003
R11118 VN.n7585 VN.n7571 0.003
R11119 VN.n7953 VN.n7948 0.003
R11120 VN.n8430 VN.n8416 0.003
R11121 VN.n8802 VN.n8797 0.003
R11122 VN.n9292 VN.n9278 0.003
R11123 VN.n9664 VN.n9659 0.003
R11124 VN.n10174 VN.n10160 0.003
R11125 VN.n10545 VN.n10537 0.003
R11126 VN.n10566 VN.n10558 0.003
R11127 VN.n11069 VN.n11051 0.003
R11128 VN.n11154 VN.n11149 0.003
R11129 VN.n12081 VN.n12071 0.003
R11130 VN.n10209 VN.n10198 0.003
R11131 VN.n9326 VN.n9315 0.003
R11132 VN.n8464 VN.n8453 0.003
R11133 VN.n7619 VN.n7608 0.003
R11134 VN.n7230 VN.n7219 0.003
R11135 VN.n5987 VN.n5976 0.003
R11136 VN.n5195 VN.n5184 0.003
R11137 VN.n4420 VN.n4409 0.003
R11138 VN.n3663 VN.n3652 0.003
R11139 VN.n2923 VN.n2912 0.003
R11140 VN.n2201 VN.n2190 0.003
R11141 VN.n1612 VN.n1599 0.003
R11142 VN.n1831 VN.n1828 0.003
R11143 VN.n2540 VN.n2537 0.003
R11144 VN.n3262 VN.n3259 0.003
R11145 VN.n4006 VN.n4003 0.003
R11146 VN.n4763 VN.n4760 0.003
R11147 VN.n5542 VN.n5539 0.003
R11148 VN.n6334 VN.n6331 0.003
R11149 VN.n6779 VN.n6776 0.003
R11150 VN.n7970 VN.n7967 0.003
R11151 VN.n8819 VN.n8816 0.003
R11152 VN.n9681 VN.n9678 0.003
R11153 VN.n11414 VN.n11402 0.003
R11154 VN.n11397 VN.n11090 0.003
R11155 VN.n12115 VN.n12105 0.003
R11156 VN.n925 VN.n920 0.003
R11157 VN.n1163 VN.n1161 0.003
R11158 VN.n1526 VN.n1514 0.003
R11159 VN.n1853 VN.n1851 0.003
R11160 VN.n2234 VN.n2222 0.003
R11161 VN.n2562 VN.n2560 0.003
R11162 VN.n2956 VN.n2944 0.003
R11163 VN.n3284 VN.n3282 0.003
R11164 VN.n3696 VN.n3684 0.003
R11165 VN.n4028 VN.n4026 0.003
R11166 VN.n4453 VN.n4441 0.003
R11167 VN.n4785 VN.n4783 0.003
R11168 VN.n5228 VN.n5216 0.003
R11169 VN.n5564 VN.n5562 0.003
R11170 VN.n6020 VN.n6008 0.003
R11171 VN.n6356 VN.n6354 0.003
R11172 VN.n7263 VN.n7251 0.003
R11173 VN.n6801 VN.n6799 0.003
R11174 VN.n7652 VN.n7640 0.003
R11175 VN.n7992 VN.n7990 0.003
R11176 VN.n8497 VN.n8485 0.003
R11177 VN.n8841 VN.n8839 0.003
R11178 VN.n9359 VN.n9347 0.003
R11179 VN.n9703 VN.n9701 0.003
R11180 VN.n10242 VN.n10230 0.003
R11181 VN.n10588 VN.n10586 0.003
R11182 VN.n11441 VN.n11429 0.003
R11183 VN.n11138 VN.n11130 0.003
R11184 VN.n10609 VN.n10606 0.003
R11185 VN.n10263 VN.n10257 0.003
R11186 VN.n9722 VN.n9715 0.003
R11187 VN.n9380 VN.n9374 0.003
R11188 VN.n8860 VN.n8853 0.003
R11189 VN.n8518 VN.n8512 0.003
R11190 VN.n8011 VN.n8004 0.003
R11191 VN.n7673 VN.n7667 0.003
R11192 VN.n6820 VN.n6813 0.003
R11193 VN.n7284 VN.n7278 0.003
R11194 VN.n6375 VN.n6368 0.003
R11195 VN.n6041 VN.n6035 0.003
R11196 VN.n5583 VN.n5576 0.003
R11197 VN.n5249 VN.n5243 0.003
R11198 VN.n4804 VN.n4797 0.003
R11199 VN.n4474 VN.n4468 0.003
R11200 VN.n4047 VN.n4040 0.003
R11201 VN.n3717 VN.n3711 0.003
R11202 VN.n3303 VN.n3296 0.003
R11203 VN.n2977 VN.n2971 0.003
R11204 VN.n2581 VN.n2574 0.003
R11205 VN.n2255 VN.n2249 0.003
R11206 VN.n1872 VN.n1865 0.003
R11207 VN.n1550 VN.n1544 0.003
R11208 VN.n1182 VN.n1175 0.003
R11209 VN.n864 VN.n858 0.003
R11210 VN.n507 VN.n500 0.003
R11211 VN.n253 VN.n247 0.003
R11212 VN.n12144 VN.n12131 0.003
R11213 VN.n11036 VN.n11024 0.003
R11214 VN.n11172 VN.n11167 0.003
R11215 VN.n11991 VN.n11986 0.003
R11216 VN.n4536 VN.n4523 0.003
R11217 VN.n4695 VN.n4692 0.003
R11218 VN.n5069 VN.n5058 0.003
R11219 VN.n5474 VN.n5471 0.003
R11220 VN.n5861 VN.n5850 0.003
R11221 VN.n6266 VN.n6263 0.003
R11222 VN.n7104 VN.n7093 0.003
R11223 VN.n6711 VN.n6708 0.003
R11224 VN.n7493 VN.n7482 0.003
R11225 VN.n7902 VN.n7899 0.003
R11226 VN.n8338 VN.n8327 0.003
R11227 VN.n8751 VN.n8748 0.003
R11228 VN.n9200 VN.n9189 0.003
R11229 VN.n9613 VN.n9610 0.003
R11230 VN.n10082 VN.n10071 0.003
R11231 VN.n10490 VN.n10486 0.003
R11232 VN.n10951 VN.n10945 0.003
R11233 VN.n11222 VN.n11219 0.003
R11234 VN.n12014 VN.n12009 0.003
R11235 VN.n3782 VN.n3770 0.003
R11236 VN.n3955 VN.n3950 0.003
R11237 VN.n4323 VN.n4309 0.003
R11238 VN.n4712 VN.n4707 0.003
R11239 VN.n5098 VN.n5084 0.003
R11240 VN.n5491 VN.n5486 0.003
R11241 VN.n5890 VN.n5876 0.003
R11242 VN.n6283 VN.n6278 0.003
R11243 VN.n7133 VN.n7119 0.003
R11244 VN.n6728 VN.n6723 0.003
R11245 VN.n7522 VN.n7508 0.003
R11246 VN.n7919 VN.n7914 0.003
R11247 VN.n8367 VN.n8353 0.003
R11248 VN.n8768 VN.n8763 0.003
R11249 VN.n9229 VN.n9215 0.003
R11250 VN.n9630 VN.n9625 0.003
R11251 VN.n10111 VN.n10097 0.003
R11252 VN.n10507 VN.n10502 0.003
R11253 VN.n10980 VN.n10966 0.003
R11254 VN.n11206 VN.n11201 0.003
R11255 VN.n11946 VN.n11941 0.003
R11256 VN.n6103 VN.n6090 0.003
R11257 VN.n6232 VN.n6229 0.003
R11258 VN.n7041 VN.n7030 0.003
R11259 VN.n6677 VN.n6674 0.003
R11260 VN.n7430 VN.n7419 0.003
R11261 VN.n7868 VN.n7865 0.003
R11262 VN.n8275 VN.n8264 0.003
R11263 VN.n8717 VN.n8714 0.003
R11264 VN.n9137 VN.n9126 0.003
R11265 VN.n9579 VN.n9576 0.003
R11266 VN.n10019 VN.n10008 0.003
R11267 VN.n10455 VN.n10451 0.003
R11268 VN.n10893 VN.n10887 0.003
R11269 VN.n11256 VN.n11253 0.003
R11270 VN.n11969 VN.n11964 0.003
R11271 VN.n5314 VN.n5302 0.003
R11272 VN.n5457 VN.n5452 0.003
R11273 VN.n5827 VN.n5813 0.003
R11274 VN.n6249 VN.n6244 0.003
R11275 VN.n7070 VN.n7056 0.003
R11276 VN.n6694 VN.n6689 0.003
R11277 VN.n7459 VN.n7445 0.003
R11278 VN.n7885 VN.n7880 0.003
R11279 VN.n8304 VN.n8290 0.003
R11280 VN.n8734 VN.n8729 0.003
R11281 VN.n9166 VN.n9152 0.003
R11282 VN.n9596 VN.n9591 0.003
R11283 VN.n10048 VN.n10034 0.003
R11284 VN.n10472 VN.n10467 0.003
R11285 VN.n10922 VN.n10908 0.003
R11286 VN.n11240 VN.n11235 0.003
R11287 VN.n6660 VN.n6655 0.003
R11288 VN.n7396 VN.n7382 0.003
R11289 VN.n7851 VN.n7846 0.003
R11290 VN.n8241 VN.n8227 0.003
R11291 VN.n8700 VN.n8695 0.003
R11292 VN.n9103 VN.n9089 0.003
R11293 VN.n9562 VN.n9557 0.003
R11294 VN.n9985 VN.n9971 0.003
R11295 VN.n10437 VN.n10432 0.003
R11296 VN.n10864 VN.n10850 0.003
R11297 VN.n11273 VN.n11268 0.003
R11298 VN.n11924 VN.n11915 0.003
R11299 VN.n11897 VN.n11892 0.003
R11300 VN.n7735 VN.n7722 0.003
R11301 VN.n7834 VN.n7831 0.003
R11302 VN.n8212 VN.n8201 0.003
R11303 VN.n8683 VN.n8680 0.003
R11304 VN.n9074 VN.n9063 0.003
R11305 VN.n9545 VN.n9542 0.003
R11306 VN.n9956 VN.n9945 0.003
R11307 VN.n10420 VN.n10416 0.003
R11308 VN.n10835 VN.n10829 0.003
R11309 VN.n11289 VN.n11287 0.003
R11310 VN.n11639 VN.n11634 0.003
R11311 VN.n9442 VN.n9429 0.003
R11312 VN.n9511 VN.n9508 0.003
R11313 VN.n9893 VN.n9882 0.003
R11314 VN.n10385 VN.n10381 0.003
R11315 VN.n10777 VN.n10771 0.003
R11316 VN.n11323 VN.n11320 0.003
R11317 VN.n11876 VN.n11871 0.003
R11318 VN.n8583 VN.n8571 0.003
R11319 VN.n8666 VN.n8661 0.003
R11320 VN.n9040 VN.n9026 0.003
R11321 VN.n9528 VN.n9523 0.003
R11322 VN.n9922 VN.n9908 0.003
R11323 VN.n10402 VN.n10397 0.003
R11324 VN.n10806 VN.n10792 0.003
R11325 VN.n11307 VN.n11302 0.003
R11326 VN.n11594 VN.n11589 0.003
R11327 VN.n11489 VN.n11480 0.003
R11328 VN.n11357 VN.n11354 0.003
R11329 VN.n11617 VN.n11612 0.003
R11330 VN.n10328 VN.n10316 0.003
R11331 VN.n10367 VN.n10362 0.003
R11332 VN.n10748 VN.n10734 0.003
R11333 VN.n11341 VN.n11336 0.003
R11334 VN.n11100 VN.n11094 0.003
R11335 VN.n11506 VN.n11500 0.003
R11336 VN.n10662 VN.n10338 0.003
R11337 VN.n10676 VN.n10666 0.003
R11338 VN.n9757 VN.n9751 0.003
R11339 VN.n9462 VN.n9452 0.003
R11340 VN.n8895 VN.n8889 0.003
R11341 VN.n8603 VN.n8593 0.003
R11342 VN.n8046 VN.n8040 0.003
R11343 VN.n7755 VN.n7745 0.003
R11344 VN.n6855 VN.n6849 0.003
R11345 VN.n7007 VN.n6997 0.003
R11346 VN.n6410 VN.n6404 0.003
R11347 VN.n6123 VN.n6113 0.003
R11348 VN.n5618 VN.n5612 0.003
R11349 VN.n5334 VN.n5324 0.003
R11350 VN.n4839 VN.n4833 0.003
R11351 VN.n4556 VN.n4546 0.003
R11352 VN.n4082 VN.n4076 0.003
R11353 VN.n3802 VN.n3792 0.003
R11354 VN.n3338 VN.n3332 0.003
R11355 VN.n3059 VN.n3049 0.003
R11356 VN.n2616 VN.n2610 0.003
R11357 VN.n2340 VN.n2330 0.003
R11358 VN.n1907 VN.n1901 0.003
R11359 VN.n1632 VN.n1622 0.003
R11360 VN.n1217 VN.n1211 0.003
R11361 VN.n945 VN.n935 0.003
R11362 VN.n542 VN.n536 0.003
R11363 VN.n273 VN.n263 0.003
R11364 VN.n12299 VN.n12287 0.003
R11365 VN.n12314 VN.n12304 0.003
R11366 VN.n12282 VN.n12269 0.003
R11367 VN.n10644 VN.n10639 0.003
R11368 VN.n10691 VN.n10690 0.003
R11369 VN.n12630 VN.n12629 0.003
R11370 VN.n12632 VN.n12328 0.003
R11371 VN.n12343 VN.n12342 0.003
R11372 VN.n288 VN.n287 0.003
R11373 VN.n558 VN.n556 0.003
R11374 VN.n960 VN.n959 0.003
R11375 VN.n1233 VN.n1231 0.003
R11376 VN.n1647 VN.n1646 0.003
R11377 VN.n1923 VN.n1921 0.003
R11378 VN.n2355 VN.n2354 0.003
R11379 VN.n2632 VN.n2630 0.003
R11380 VN.n3074 VN.n3073 0.003
R11381 VN.n3354 VN.n3352 0.003
R11382 VN.n3817 VN.n3816 0.003
R11383 VN.n4098 VN.n4096 0.003
R11384 VN.n4571 VN.n4570 0.003
R11385 VN.n4855 VN.n4853 0.003
R11386 VN.n5349 VN.n5348 0.003
R11387 VN.n5634 VN.n5632 0.003
R11388 VN.n6138 VN.n6137 0.003
R11389 VN.n6426 VN.n6424 0.003
R11390 VN.n6987 VN.n6986 0.003
R11391 VN.n6871 VN.n6869 0.003
R11392 VN.n7770 VN.n7769 0.003
R11393 VN.n8062 VN.n8060 0.003
R11394 VN.n8618 VN.n8617 0.003
R11395 VN.n8911 VN.n8909 0.003
R11396 VN.n9796 VN.n9476 0.003
R11397 VN.n9795 VN.n9794 0.003
R11398 VN.n9779 VN.n9768 0.003
R11399 VN.n9811 VN.n9810 0.003
R11400 VN.n12422 VN.n12420 0.003
R11401 VN.n12663 VN.n12646 0.003
R11402 VN.n12661 VN.n12660 0.003
R11403 VN.n303 VN.n302 0.003
R11404 VN.n574 VN.n572 0.003
R11405 VN.n975 VN.n974 0.003
R11406 VN.n1249 VN.n1247 0.003
R11407 VN.n1662 VN.n1661 0.003
R11408 VN.n1939 VN.n1937 0.003
R11409 VN.n2370 VN.n2369 0.003
R11410 VN.n2648 VN.n2646 0.003
R11411 VN.n3089 VN.n3088 0.003
R11412 VN.n3370 VN.n3368 0.003
R11413 VN.n3832 VN.n3831 0.003
R11414 VN.n4114 VN.n4112 0.003
R11415 VN.n4586 VN.n4585 0.003
R11416 VN.n4871 VN.n4869 0.003
R11417 VN.n5364 VN.n5363 0.003
R11418 VN.n5650 VN.n5648 0.003
R11419 VN.n6153 VN.n6152 0.003
R11420 VN.n6442 VN.n6440 0.003
R11421 VN.n6972 VN.n6971 0.003
R11422 VN.n6887 VN.n6885 0.003
R11423 VN.n7785 VN.n7784 0.003
R11424 VN.n8078 VN.n8076 0.003
R11425 VN.n8950 VN.n8632 0.003
R11426 VN.n8949 VN.n8948 0.003
R11427 VN.n8933 VN.n8922 0.003
R11428 VN.n8965 VN.n8964 0.003
R11429 VN.n12438 VN.n12436 0.003
R11430 VN.n12774 VN.n12677 0.003
R11431 VN.n12772 VN.n12771 0.003
R11432 VN.n318 VN.n317 0.003
R11433 VN.n590 VN.n588 0.003
R11434 VN.n990 VN.n989 0.003
R11435 VN.n1265 VN.n1263 0.003
R11436 VN.n1677 VN.n1676 0.003
R11437 VN.n1955 VN.n1953 0.003
R11438 VN.n2385 VN.n2384 0.003
R11439 VN.n2664 VN.n2662 0.003
R11440 VN.n3104 VN.n3103 0.003
R11441 VN.n3386 VN.n3384 0.003
R11442 VN.n3847 VN.n3846 0.003
R11443 VN.n4130 VN.n4128 0.003
R11444 VN.n4601 VN.n4600 0.003
R11445 VN.n4887 VN.n4885 0.003
R11446 VN.n5379 VN.n5378 0.003
R11447 VN.n5666 VN.n5664 0.003
R11448 VN.n6168 VN.n6167 0.003
R11449 VN.n6458 VN.n6456 0.003
R11450 VN.n6957 VN.n6956 0.003
R11451 VN.n6903 VN.n6901 0.003
R11452 VN.n8117 VN.n7799 0.003
R11453 VN.n8116 VN.n8115 0.003
R11454 VN.n8100 VN.n8089 0.003
R11455 VN.n8132 VN.n8131 0.003
R11456 VN.n12454 VN.n12452 0.003
R11457 VN.n12808 VN.n12791 0.003
R11458 VN.n12806 VN.n12805 0.003
R11459 VN.n333 VN.n332 0.003
R11460 VN.n606 VN.n604 0.003
R11461 VN.n1005 VN.n1004 0.003
R11462 VN.n1281 VN.n1279 0.003
R11463 VN.n1692 VN.n1691 0.003
R11464 VN.n1971 VN.n1969 0.003
R11465 VN.n2400 VN.n2399 0.003
R11466 VN.n2680 VN.n2678 0.003
R11467 VN.n3119 VN.n3118 0.003
R11468 VN.n3402 VN.n3400 0.003
R11469 VN.n3862 VN.n3861 0.003
R11470 VN.n4146 VN.n4144 0.003
R11471 VN.n4616 VN.n4615 0.003
R11472 VN.n4903 VN.n4901 0.003
R11473 VN.n5394 VN.n5393 0.003
R11474 VN.n5682 VN.n5680 0.003
R11475 VN.n6183 VN.n6182 0.003
R11476 VN.n6474 VN.n6472 0.003
R11477 VN.n6942 VN.n6626 0.003
R11478 VN.n6941 VN.n6940 0.003
R11479 VN.n6925 VN.n6914 0.003
R11480 VN.n6612 VN.n6611 0.003
R11481 VN.n12470 VN.n12468 0.003
R11482 VN.n12839 VN.n12822 0.003
R11483 VN.n12837 VN.n12836 0.003
R11484 VN.n348 VN.n347 0.003
R11485 VN.n622 VN.n620 0.003
R11486 VN.n1020 VN.n1019 0.003
R11487 VN.n1297 VN.n1295 0.003
R11488 VN.n1707 VN.n1706 0.003
R11489 VN.n1987 VN.n1985 0.003
R11490 VN.n2415 VN.n2414 0.003
R11491 VN.n2696 VN.n2694 0.003
R11492 VN.n3134 VN.n3133 0.003
R11493 VN.n3418 VN.n3416 0.003
R11494 VN.n3877 VN.n3876 0.003
R11495 VN.n4162 VN.n4160 0.003
R11496 VN.n4631 VN.n4630 0.003
R11497 VN.n4919 VN.n4917 0.003
R11498 VN.n5409 VN.n5408 0.003
R11499 VN.n5698 VN.n5696 0.003
R11500 VN.n6513 VN.n6197 0.003
R11501 VN.n6512 VN.n6511 0.003
R11502 VN.n6496 VN.n6485 0.003
R11503 VN.n6528 VN.n6527 0.003
R11504 VN.n12486 VN.n12484 0.003
R11505 VN.n12867 VN.n12850 0.003
R11506 VN.n12865 VN.n12864 0.003
R11507 VN.n363 VN.n362 0.003
R11508 VN.n638 VN.n636 0.003
R11509 VN.n1035 VN.n1034 0.003
R11510 VN.n1313 VN.n1311 0.003
R11511 VN.n1722 VN.n1721 0.003
R11512 VN.n2003 VN.n2001 0.003
R11513 VN.n2430 VN.n2429 0.003
R11514 VN.n2712 VN.n2710 0.003
R11515 VN.n3149 VN.n3148 0.003
R11516 VN.n3434 VN.n3432 0.003
R11517 VN.n3892 VN.n3891 0.003
R11518 VN.n4178 VN.n4176 0.003
R11519 VN.n4646 VN.n4645 0.003
R11520 VN.n4935 VN.n4933 0.003
R11521 VN.n5737 VN.n5423 0.003
R11522 VN.n5736 VN.n5735 0.003
R11523 VN.n5720 VN.n5709 0.003
R11524 VN.n5752 VN.n5751 0.003
R11525 VN.n12502 VN.n12500 0.003
R11526 VN.n12898 VN.n12881 0.003
R11527 VN.n12896 VN.n12895 0.003
R11528 VN.n378 VN.n377 0.003
R11529 VN.n654 VN.n652 0.003
R11530 VN.n1050 VN.n1049 0.003
R11531 VN.n1329 VN.n1327 0.003
R11532 VN.n1737 VN.n1736 0.003
R11533 VN.n2019 VN.n2017 0.003
R11534 VN.n2445 VN.n2444 0.003
R11535 VN.n2728 VN.n2726 0.003
R11536 VN.n3164 VN.n3163 0.003
R11537 VN.n3450 VN.n3448 0.003
R11538 VN.n3907 VN.n3906 0.003
R11539 VN.n4194 VN.n4192 0.003
R11540 VN.n4974 VN.n4660 0.003
R11541 VN.n4973 VN.n4972 0.003
R11542 VN.n4957 VN.n4946 0.003
R11543 VN.n4989 VN.n4988 0.003
R11544 VN.n12518 VN.n12516 0.003
R11545 VN.n12929 VN.n12912 0.003
R11546 VN.n12927 VN.n12926 0.003
R11547 VN.n393 VN.n392 0.003
R11548 VN.n670 VN.n668 0.003
R11549 VN.n1065 VN.n1064 0.003
R11550 VN.n1345 VN.n1343 0.003
R11551 VN.n1752 VN.n1751 0.003
R11552 VN.n2035 VN.n2033 0.003
R11553 VN.n2460 VN.n2459 0.003
R11554 VN.n2744 VN.n2742 0.003
R11555 VN.n3179 VN.n3178 0.003
R11556 VN.n3466 VN.n3464 0.003
R11557 VN.n4233 VN.n3921 0.003
R11558 VN.n4232 VN.n4231 0.003
R11559 VN.n4216 VN.n4205 0.003
R11560 VN.n4248 VN.n4247 0.003
R11561 VN.n12534 VN.n12532 0.003
R11562 VN.n12960 VN.n12943 0.003
R11563 VN.n12958 VN.n12957 0.003
R11564 VN.n408 VN.n407 0.003
R11565 VN.n686 VN.n684 0.003
R11566 VN.n1080 VN.n1079 0.003
R11567 VN.n1361 VN.n1359 0.003
R11568 VN.n1767 VN.n1766 0.003
R11569 VN.n2051 VN.n2049 0.003
R11570 VN.n2475 VN.n2474 0.003
R11571 VN.n2760 VN.n2758 0.003
R11572 VN.n3505 VN.n3193 0.003
R11573 VN.n3504 VN.n3503 0.003
R11574 VN.n3488 VN.n3477 0.003
R11575 VN.n3520 VN.n3519 0.003
R11576 VN.n12550 VN.n12548 0.003
R11577 VN.n12991 VN.n12974 0.003
R11578 VN.n12989 VN.n12988 0.003
R11579 VN.n423 VN.n422 0.003
R11580 VN.n702 VN.n700 0.003
R11581 VN.n1095 VN.n1094 0.003
R11582 VN.n1377 VN.n1375 0.003
R11583 VN.n1782 VN.n1781 0.003
R11584 VN.n2067 VN.n2065 0.003
R11585 VN.n2799 VN.n2489 0.003
R11586 VN.n2798 VN.n2797 0.003
R11587 VN.n2782 VN.n2771 0.003
R11588 VN.n2814 VN.n2813 0.003
R11589 VN.n12566 VN.n12564 0.003
R11590 VN.n13022 VN.n13005 0.003
R11591 VN.n13020 VN.n13019 0.003
R11592 VN.n438 VN.n437 0.003
R11593 VN.n718 VN.n716 0.003
R11594 VN.n1110 VN.n1109 0.003
R11595 VN.n1393 VN.n1391 0.003
R11596 VN.n2106 VN.n1796 0.003
R11597 VN.n2105 VN.n2104 0.003
R11598 VN.n2089 VN.n2078 0.003
R11599 VN.n2121 VN.n2120 0.003
R11600 VN.n12582 VN.n12580 0.003
R11601 VN.n13053 VN.n13036 0.003
R11602 VN.n13051 VN.n13050 0.003
R11603 VN.n453 VN.n452 0.003
R11604 VN.n734 VN.n732 0.003
R11605 VN.n1432 VN.n1124 0.003
R11606 VN.n1431 VN.n1430 0.003
R11607 VN.n1415 VN.n1404 0.003
R11608 VN.n1447 VN.n1446 0.003
R11609 VN.n12598 VN.n12596 0.003
R11610 VN.n13084 VN.n13067 0.003
R11611 VN.n13082 VN.n13081 0.003
R11612 VN.n772 VN.n467 0.003
R11613 VN.n771 VN.n770 0.003
R11614 VN.n755 VN.n743 0.003
R11615 VN.n794 VN.n788 0.003
R11616 VN.n12614 VN.n12609 0.003
R11617 VN.n13104 VN.n13099 0.003
R11618 VN.n12756 VN.n12751 0.003
R11619 VN.n12385 VN.n12380 0.003
R11620 VN.n12233 VN.n12228 0.003
R11621 VN.n12737 VN.n12725 0.003
R11622 VN.n12182 VN.n11543 0.003
R11623 VN.n11838 VN.n11837 0.003
R11624 VN.n11827 VN.n11826 0.003
R11625 VN.n11816 VN.n11815 0.003
R11626 VN.n11865 VN.n11864 0.003
R11627 VN.n11805 VN.n11804 0.003
R11628 VN.n11794 VN.n11793 0.003
R11629 VN.n11662 VN.n11661 0.003
R11630 VN.n11658 VN.n11657 0.003
R11631 VN.n182 VN.n0 0.003
R11632 VN.n182 VN.n181 0.003
R11633 VN.n489 VN.n488 0.003
R11634 VN.n12079 VN.n12078 0.003
R11635 VN.n478 VN.n477 0.003
R11636 VN.n1526 VN.n1525 0.003
R11637 VN.n2234 VN.n2233 0.003
R11638 VN.n2956 VN.n2955 0.003
R11639 VN.n3696 VN.n3695 0.003
R11640 VN.n4453 VN.n4452 0.003
R11641 VN.n5228 VN.n5227 0.003
R11642 VN.n6020 VN.n6019 0.003
R11643 VN.n7263 VN.n7262 0.003
R11644 VN.n7652 VN.n7651 0.003
R11645 VN.n8497 VN.n8496 0.003
R11646 VN.n9359 VN.n9358 0.003
R11647 VN.n10242 VN.n10241 0.003
R11648 VN.n11414 VN.n11086 0.003
R11649 VN.n11922 VN.n11921 0.003
R11650 VN.n12756 VN.n12747 0.003
R11651 VN.n13137 VN.n13136 0.003
R11652 VN.t8 VN.n11777 0.003
R11653 VN.t76 VN.n6603 0.003
R11654 VN.n12366 VN.n12351 0.003
R11655 VN.n2507 VN.n2506 0.003
R11656 VN.n3939 VN.n3938 0.003
R11657 VN.n5441 VN.n5440 0.003
R11658 VN.n6644 VN.n6643 0.003
R11659 VN.n8650 VN.n8649 0.003
R11660 VN.n10351 VN.n10350 0.003
R11661 VN.t51 VN.n18 0.003
R11662 VN.t51 VN.n100 0.003
R11663 VN.n6592 VN.n6591 0.003
R11664 VN.n243 VN.n242 0.003
R11665 VN.n2523 VN.n2514 0.003
R11666 VN.n3245 VN.n3236 0.003
R11667 VN.n3989 VN.n3980 0.003
R11668 VN.n4746 VN.n4737 0.003
R11669 VN.n5525 VN.n5516 0.003
R11670 VN.n6317 VN.n6308 0.003
R11671 VN.n6762 VN.n6753 0.003
R11672 VN.n7953 VN.n7944 0.003
R11673 VN.n8802 VN.n8793 0.003
R11674 VN.n9664 VN.n9655 0.003
R11675 VN.n10545 VN.n10533 0.003
R11676 VN.n3955 VN.n3946 0.003
R11677 VN.n4712 VN.n4703 0.003
R11678 VN.n5491 VN.n5482 0.003
R11679 VN.n6283 VN.n6274 0.003
R11680 VN.n6728 VN.n6719 0.003
R11681 VN.n7919 VN.n7910 0.003
R11682 VN.n8768 VN.n8759 0.003
R11683 VN.n9630 VN.n9621 0.003
R11684 VN.n10507 VN.n10498 0.003
R11685 VN.n5457 VN.n5448 0.003
R11686 VN.n6249 VN.n6240 0.003
R11687 VN.n6694 VN.n6685 0.003
R11688 VN.n7885 VN.n7876 0.003
R11689 VN.n8734 VN.n8725 0.003
R11690 VN.n9596 VN.n9587 0.003
R11691 VN.n10472 VN.n10463 0.003
R11692 VN.n8666 VN.n8657 0.003
R11693 VN.n9528 VN.n9519 0.003
R11694 VN.n10402 VN.n10393 0.003
R11695 VN.n10367 VN.n10358 0.003
R11696 VN.n12233 VN.n12224 0.003
R11697 VN.n195 VN.n186 0.003
R11698 VN.n12162 VN.n12161 0.003
R11699 VN.n11483 VN.n11482 0.003
R11700 VN.n12095 VN.n12094 0.003
R11701 VN.n780 VN.n779 0.003
R11702 VN.n12059 VN.n12051 0.002
R11703 VN.n11172 VN.n11164 0.002
R11704 VN.n11036 VN.n11016 0.002
R11705 VN.n10545 VN.n10534 0.002
R11706 VN.n10174 VN.n10157 0.002
R11707 VN.n9664 VN.n9656 0.002
R11708 VN.n9292 VN.n9275 0.002
R11709 VN.n8802 VN.n8794 0.002
R11710 VN.n8430 VN.n8413 0.002
R11711 VN.n7953 VN.n7945 0.002
R11712 VN.n7585 VN.n7568 0.002
R11713 VN.n6762 VN.n6754 0.002
R11714 VN.n7196 VN.n7179 0.002
R11715 VN.n6317 VN.n6309 0.002
R11716 VN.n5953 VN.n5936 0.002
R11717 VN.n5525 VN.n5517 0.002
R11718 VN.n5161 VN.n5144 0.002
R11719 VN.n4746 VN.n4738 0.002
R11720 VN.n4386 VN.n4369 0.002
R11721 VN.n3989 VN.n3981 0.002
R11722 VN.n3629 VN.n3612 0.002
R11723 VN.n3245 VN.n3237 0.002
R11724 VN.n2889 VN.n2872 0.002
R11725 VN.n2523 VN.n2515 0.002
R11726 VN.n12115 VN.n12102 0.002
R11727 VN.n11397 VN.n11087 0.002
R11728 VN.n11414 VN.n11399 0.002
R11729 VN.n10588 VN.n10573 0.002
R11730 VN.n10242 VN.n10216 0.002
R11731 VN.n9703 VN.n9688 0.002
R11732 VN.n9359 VN.n9333 0.002
R11733 VN.n8841 VN.n8826 0.002
R11734 VN.n8497 VN.n8471 0.002
R11735 VN.n7992 VN.n7977 0.002
R11736 VN.n7652 VN.n7626 0.002
R11737 VN.n6801 VN.n6786 0.002
R11738 VN.n7263 VN.n7237 0.002
R11739 VN.n6356 VN.n6341 0.002
R11740 VN.n6020 VN.n5994 0.002
R11741 VN.n5564 VN.n5549 0.002
R11742 VN.n5228 VN.n5202 0.002
R11743 VN.n4785 VN.n4770 0.002
R11744 VN.n4453 VN.n4427 0.002
R11745 VN.n4028 VN.n4013 0.002
R11746 VN.n3696 VN.n3670 0.002
R11747 VN.n3284 VN.n3269 0.002
R11748 VN.n2956 VN.n2930 0.002
R11749 VN.n2562 VN.n2547 0.002
R11750 VN.n2234 VN.n2208 0.002
R11751 VN.n1853 VN.n1838 0.002
R11752 VN.n1526 VN.n1500 0.002
R11753 VN.n1163 VN.n1148 0.002
R11754 VN.n507 VN.n497 0.002
R11755 VN.n864 VN.n855 0.002
R11756 VN.n1182 VN.n1172 0.002
R11757 VN.n1550 VN.n1541 0.002
R11758 VN.n1872 VN.n1862 0.002
R11759 VN.n2255 VN.n2246 0.002
R11760 VN.n2581 VN.n2571 0.002
R11761 VN.n2977 VN.n2968 0.002
R11762 VN.n3303 VN.n3293 0.002
R11763 VN.n3717 VN.n3708 0.002
R11764 VN.n4047 VN.n4037 0.002
R11765 VN.n4474 VN.n4465 0.002
R11766 VN.n4804 VN.n4794 0.002
R11767 VN.n5249 VN.n5240 0.002
R11768 VN.n5583 VN.n5573 0.002
R11769 VN.n6041 VN.n6032 0.002
R11770 VN.n6375 VN.n6365 0.002
R11771 VN.n7284 VN.n7275 0.002
R11772 VN.n6820 VN.n6810 0.002
R11773 VN.n7673 VN.n7664 0.002
R11774 VN.n8011 VN.n8001 0.002
R11775 VN.n8518 VN.n8509 0.002
R11776 VN.n8860 VN.n8850 0.002
R11777 VN.n9380 VN.n9371 0.002
R11778 VN.n9722 VN.n9712 0.002
R11779 VN.n10263 VN.n10254 0.002
R11780 VN.n10609 VN.n10595 0.002
R11781 VN.n11441 VN.n11426 0.002
R11782 VN.n11138 VN.n11127 0.002
R11783 VN.n12144 VN.n12123 0.002
R11784 VN.n12014 VN.n12006 0.002
R11785 VN.n11206 VN.n11198 0.002
R11786 VN.n10980 VN.n10958 0.002
R11787 VN.n10507 VN.n10499 0.002
R11788 VN.n10111 VN.n10094 0.002
R11789 VN.n9630 VN.n9622 0.002
R11790 VN.n9229 VN.n9212 0.002
R11791 VN.n8768 VN.n8760 0.002
R11792 VN.n8367 VN.n8350 0.002
R11793 VN.n7919 VN.n7911 0.002
R11794 VN.n7522 VN.n7505 0.002
R11795 VN.n6728 VN.n6720 0.002
R11796 VN.n7133 VN.n7116 0.002
R11797 VN.n6283 VN.n6275 0.002
R11798 VN.n5890 VN.n5873 0.002
R11799 VN.n5491 VN.n5483 0.002
R11800 VN.n5098 VN.n5081 0.002
R11801 VN.n4712 VN.n4704 0.002
R11802 VN.n4323 VN.n4306 0.002
R11803 VN.n3955 VN.n3947 0.002
R11804 VN.n11969 VN.n11961 0.002
R11805 VN.n11240 VN.n11232 0.002
R11806 VN.n10922 VN.n10900 0.002
R11807 VN.n10472 VN.n10464 0.002
R11808 VN.n10048 VN.n10031 0.002
R11809 VN.n9596 VN.n9588 0.002
R11810 VN.n9166 VN.n9149 0.002
R11811 VN.n8734 VN.n8726 0.002
R11812 VN.n8304 VN.n8287 0.002
R11813 VN.n7885 VN.n7877 0.002
R11814 VN.n7459 VN.n7442 0.002
R11815 VN.n6694 VN.n6686 0.002
R11816 VN.n7070 VN.n7053 0.002
R11817 VN.n6249 VN.n6241 0.002
R11818 VN.n5827 VN.n5810 0.002
R11819 VN.n5457 VN.n5449 0.002
R11820 VN.n6660 VN.n6652 0.002
R11821 VN.n7396 VN.n7379 0.002
R11822 VN.n7851 VN.n7843 0.002
R11823 VN.n8241 VN.n8224 0.002
R11824 VN.n8700 VN.n8692 0.002
R11825 VN.n9103 VN.n9086 0.002
R11826 VN.n9562 VN.n9554 0.002
R11827 VN.n9985 VN.n9968 0.002
R11828 VN.n10437 VN.n10429 0.002
R11829 VN.n10864 VN.n10847 0.002
R11830 VN.n11273 VN.n11265 0.002
R11831 VN.n11924 VN.n11912 0.002
R11832 VN.n11876 VN.n11868 0.002
R11833 VN.n11307 VN.n11299 0.002
R11834 VN.n10806 VN.n10784 0.002
R11835 VN.n10402 VN.n10394 0.002
R11836 VN.n9922 VN.n9905 0.002
R11837 VN.n9528 VN.n9520 0.002
R11838 VN.n9040 VN.n9023 0.002
R11839 VN.n8666 VN.n8658 0.002
R11840 VN.n11617 VN.n11609 0.002
R11841 VN.n11341 VN.n11333 0.002
R11842 VN.n10748 VN.n10726 0.002
R11843 VN.n10367 VN.n10359 0.002
R11844 VN.n12282 VN.n12266 0.002
R11845 VN.n12314 VN.n12301 0.002
R11846 VN.n12299 VN.n12284 0.002
R11847 VN.n273 VN.n260 0.002
R11848 VN.n542 VN.n533 0.002
R11849 VN.n945 VN.n932 0.002
R11850 VN.n1217 VN.n1208 0.002
R11851 VN.n1632 VN.n1619 0.002
R11852 VN.n1907 VN.n1898 0.002
R11853 VN.n2340 VN.n2327 0.002
R11854 VN.n2616 VN.n2607 0.002
R11855 VN.n3059 VN.n3046 0.002
R11856 VN.n3338 VN.n3329 0.002
R11857 VN.n3802 VN.n3789 0.002
R11858 VN.n4082 VN.n4073 0.002
R11859 VN.n4556 VN.n4543 0.002
R11860 VN.n4839 VN.n4830 0.002
R11861 VN.n5334 VN.n5321 0.002
R11862 VN.n5618 VN.n5609 0.002
R11863 VN.n6123 VN.n6110 0.002
R11864 VN.n6410 VN.n6401 0.002
R11865 VN.n7007 VN.n6994 0.002
R11866 VN.n6855 VN.n6846 0.002
R11867 VN.n7755 VN.n7742 0.002
R11868 VN.n8046 VN.n8037 0.002
R11869 VN.n8603 VN.n8590 0.002
R11870 VN.n8895 VN.n8886 0.002
R11871 VN.n9462 VN.n9449 0.002
R11872 VN.n9757 VN.n9748 0.002
R11873 VN.n10676 VN.n10663 0.002
R11874 VN.n10662 VN.n10335 0.002
R11875 VN.n11506 VN.n11497 0.002
R11876 VN.n12630 VN.n12345 0.002
R11877 VN.n12632 VN.n12321 0.002
R11878 VN.n12343 VN.n12329 0.002
R11879 VN.n288 VN.n280 0.002
R11880 VN.n558 VN.n549 0.002
R11881 VN.n960 VN.n952 0.002
R11882 VN.n1233 VN.n1224 0.002
R11883 VN.n1647 VN.n1639 0.002
R11884 VN.n1923 VN.n1914 0.002
R11885 VN.n2355 VN.n2347 0.002
R11886 VN.n2632 VN.n2623 0.002
R11887 VN.n3074 VN.n3066 0.002
R11888 VN.n3354 VN.n3345 0.002
R11889 VN.n3817 VN.n3809 0.002
R11890 VN.n4098 VN.n4089 0.002
R11891 VN.n4571 VN.n4563 0.002
R11892 VN.n4855 VN.n4846 0.002
R11893 VN.n5349 VN.n5341 0.002
R11894 VN.n5634 VN.n5625 0.002
R11895 VN.n6138 VN.n6130 0.002
R11896 VN.n6426 VN.n6417 0.002
R11897 VN.n6987 VN.n6979 0.002
R11898 VN.n6871 VN.n6862 0.002
R11899 VN.n7770 VN.n7762 0.002
R11900 VN.n8062 VN.n8053 0.002
R11901 VN.n8618 VN.n8610 0.002
R11902 VN.n8911 VN.n8902 0.002
R11903 VN.n9796 VN.n9469 0.002
R11904 VN.n9795 VN.n9477 0.002
R11905 VN.n10691 VN.n10683 0.002
R11906 VN.n10644 VN.n10636 0.002
R11907 VN.n12422 VN.n12413 0.002
R11908 VN.n12663 VN.n12639 0.002
R11909 VN.n12661 VN.n12647 0.002
R11910 VN.n303 VN.n295 0.002
R11911 VN.n574 VN.n565 0.002
R11912 VN.n975 VN.n967 0.002
R11913 VN.n1249 VN.n1240 0.002
R11914 VN.n1662 VN.n1654 0.002
R11915 VN.n1939 VN.n1930 0.002
R11916 VN.n2370 VN.n2362 0.002
R11917 VN.n2648 VN.n2639 0.002
R11918 VN.n3089 VN.n3081 0.002
R11919 VN.n3370 VN.n3361 0.002
R11920 VN.n3832 VN.n3824 0.002
R11921 VN.n4114 VN.n4105 0.002
R11922 VN.n4586 VN.n4578 0.002
R11923 VN.n4871 VN.n4862 0.002
R11924 VN.n5364 VN.n5356 0.002
R11925 VN.n5650 VN.n5641 0.002
R11926 VN.n6153 VN.n6145 0.002
R11927 VN.n6442 VN.n6433 0.002
R11928 VN.n6972 VN.n6964 0.002
R11929 VN.n6887 VN.n6878 0.002
R11930 VN.n7785 VN.n7777 0.002
R11931 VN.n8078 VN.n8069 0.002
R11932 VN.n8950 VN.n8625 0.002
R11933 VN.n8949 VN.n8633 0.002
R11934 VN.n9811 VN.n9803 0.002
R11935 VN.n9779 VN.n9765 0.002
R11936 VN.n12438 VN.n12429 0.002
R11937 VN.n12774 VN.n12670 0.002
R11938 VN.n12772 VN.n12678 0.002
R11939 VN.n318 VN.n310 0.002
R11940 VN.n590 VN.n581 0.002
R11941 VN.n990 VN.n982 0.002
R11942 VN.n1265 VN.n1256 0.002
R11943 VN.n1677 VN.n1669 0.002
R11944 VN.n1955 VN.n1946 0.002
R11945 VN.n2385 VN.n2377 0.002
R11946 VN.n2664 VN.n2655 0.002
R11947 VN.n3104 VN.n3096 0.002
R11948 VN.n3386 VN.n3377 0.002
R11949 VN.n3847 VN.n3839 0.002
R11950 VN.n4130 VN.n4121 0.002
R11951 VN.n4601 VN.n4593 0.002
R11952 VN.n4887 VN.n4878 0.002
R11953 VN.n5379 VN.n5371 0.002
R11954 VN.n5666 VN.n5657 0.002
R11955 VN.n6168 VN.n6160 0.002
R11956 VN.n6458 VN.n6449 0.002
R11957 VN.n6957 VN.n6949 0.002
R11958 VN.n6903 VN.n6894 0.002
R11959 VN.n8117 VN.n7792 0.002
R11960 VN.n8116 VN.n7800 0.002
R11961 VN.n8965 VN.n8957 0.002
R11962 VN.n8933 VN.n8919 0.002
R11963 VN.n12454 VN.n12445 0.002
R11964 VN.n12808 VN.n12781 0.002
R11965 VN.n12806 VN.n12792 0.002
R11966 VN.n333 VN.n325 0.002
R11967 VN.n606 VN.n597 0.002
R11968 VN.n1005 VN.n997 0.002
R11969 VN.n1281 VN.n1272 0.002
R11970 VN.n1692 VN.n1684 0.002
R11971 VN.n1971 VN.n1962 0.002
R11972 VN.n2400 VN.n2392 0.002
R11973 VN.n2680 VN.n2671 0.002
R11974 VN.n3119 VN.n3111 0.002
R11975 VN.n3402 VN.n3393 0.002
R11976 VN.n3862 VN.n3854 0.002
R11977 VN.n4146 VN.n4137 0.002
R11978 VN.n4616 VN.n4608 0.002
R11979 VN.n4903 VN.n4894 0.002
R11980 VN.n5394 VN.n5386 0.002
R11981 VN.n5682 VN.n5673 0.002
R11982 VN.n6183 VN.n6175 0.002
R11983 VN.n6474 VN.n6465 0.002
R11984 VN.n6942 VN.n6619 0.002
R11985 VN.n6941 VN.n6627 0.002
R11986 VN.n8132 VN.n8124 0.002
R11987 VN.n8100 VN.n8086 0.002
R11988 VN.n12470 VN.n12461 0.002
R11989 VN.n12839 VN.n12812 0.002
R11990 VN.n12837 VN.n12823 0.002
R11991 VN.n348 VN.n340 0.002
R11992 VN.n622 VN.n613 0.002
R11993 VN.n1020 VN.n1012 0.002
R11994 VN.n1297 VN.n1288 0.002
R11995 VN.n1707 VN.n1699 0.002
R11996 VN.n1987 VN.n1978 0.002
R11997 VN.n2415 VN.n2407 0.002
R11998 VN.n2696 VN.n2687 0.002
R11999 VN.n3134 VN.n3126 0.002
R12000 VN.n3418 VN.n3409 0.002
R12001 VN.n3877 VN.n3869 0.002
R12002 VN.n4162 VN.n4153 0.002
R12003 VN.n4631 VN.n4623 0.002
R12004 VN.n4919 VN.n4910 0.002
R12005 VN.n5409 VN.n5401 0.002
R12006 VN.n5698 VN.n5689 0.002
R12007 VN.n6513 VN.n6190 0.002
R12008 VN.n6512 VN.n6198 0.002
R12009 VN.n6612 VN.n6604 0.002
R12010 VN.n6925 VN.n6911 0.002
R12011 VN.n12486 VN.n12477 0.002
R12012 VN.n12867 VN.n12843 0.002
R12013 VN.n12865 VN.n12851 0.002
R12014 VN.n363 VN.n355 0.002
R12015 VN.n638 VN.n629 0.002
R12016 VN.n1035 VN.n1027 0.002
R12017 VN.n1313 VN.n1304 0.002
R12018 VN.n1722 VN.n1714 0.002
R12019 VN.n2003 VN.n1994 0.002
R12020 VN.n2430 VN.n2422 0.002
R12021 VN.n2712 VN.n2703 0.002
R12022 VN.n3149 VN.n3141 0.002
R12023 VN.n3434 VN.n3425 0.002
R12024 VN.n3892 VN.n3884 0.002
R12025 VN.n4178 VN.n4169 0.002
R12026 VN.n4646 VN.n4638 0.002
R12027 VN.n4935 VN.n4926 0.002
R12028 VN.n5737 VN.n5416 0.002
R12029 VN.n5736 VN.n5424 0.002
R12030 VN.n6528 VN.n6520 0.002
R12031 VN.n6496 VN.n6482 0.002
R12032 VN.n12502 VN.n12493 0.002
R12033 VN.n12898 VN.n12874 0.002
R12034 VN.n12896 VN.n12882 0.002
R12035 VN.n378 VN.n370 0.002
R12036 VN.n654 VN.n645 0.002
R12037 VN.n1050 VN.n1042 0.002
R12038 VN.n1329 VN.n1320 0.002
R12039 VN.n1737 VN.n1729 0.002
R12040 VN.n2019 VN.n2010 0.002
R12041 VN.n2445 VN.n2437 0.002
R12042 VN.n2728 VN.n2719 0.002
R12043 VN.n3164 VN.n3156 0.002
R12044 VN.n3450 VN.n3441 0.002
R12045 VN.n3907 VN.n3899 0.002
R12046 VN.n4194 VN.n4185 0.002
R12047 VN.n4974 VN.n4653 0.002
R12048 VN.n4973 VN.n4661 0.002
R12049 VN.n5752 VN.n5744 0.002
R12050 VN.n5720 VN.n5706 0.002
R12051 VN.n12518 VN.n12509 0.002
R12052 VN.n12929 VN.n12905 0.002
R12053 VN.n12927 VN.n12913 0.002
R12054 VN.n393 VN.n385 0.002
R12055 VN.n670 VN.n661 0.002
R12056 VN.n1065 VN.n1057 0.002
R12057 VN.n1345 VN.n1336 0.002
R12058 VN.n1752 VN.n1744 0.002
R12059 VN.n2035 VN.n2026 0.002
R12060 VN.n2460 VN.n2452 0.002
R12061 VN.n2744 VN.n2735 0.002
R12062 VN.n3179 VN.n3171 0.002
R12063 VN.n3466 VN.n3457 0.002
R12064 VN.n4233 VN.n3914 0.002
R12065 VN.n4232 VN.n3922 0.002
R12066 VN.n4989 VN.n4981 0.002
R12067 VN.n4957 VN.n4943 0.002
R12068 VN.n12534 VN.n12525 0.002
R12069 VN.n12960 VN.n12936 0.002
R12070 VN.n12958 VN.n12944 0.002
R12071 VN.n408 VN.n400 0.002
R12072 VN.n686 VN.n677 0.002
R12073 VN.n1080 VN.n1072 0.002
R12074 VN.n1361 VN.n1352 0.002
R12075 VN.n1767 VN.n1759 0.002
R12076 VN.n2051 VN.n2042 0.002
R12077 VN.n2475 VN.n2467 0.002
R12078 VN.n2760 VN.n2751 0.002
R12079 VN.n3505 VN.n3186 0.002
R12080 VN.n3504 VN.n3194 0.002
R12081 VN.n4248 VN.n4240 0.002
R12082 VN.n4216 VN.n4202 0.002
R12083 VN.n12550 VN.n12541 0.002
R12084 VN.n12991 VN.n12967 0.002
R12085 VN.n12989 VN.n12975 0.002
R12086 VN.n423 VN.n415 0.002
R12087 VN.n702 VN.n693 0.002
R12088 VN.n1095 VN.n1087 0.002
R12089 VN.n1377 VN.n1368 0.002
R12090 VN.n1782 VN.n1774 0.002
R12091 VN.n2067 VN.n2058 0.002
R12092 VN.n2799 VN.n2482 0.002
R12093 VN.n2798 VN.n2490 0.002
R12094 VN.n3520 VN.n3512 0.002
R12095 VN.n3488 VN.n3474 0.002
R12096 VN.n12566 VN.n12557 0.002
R12097 VN.n13022 VN.n12998 0.002
R12098 VN.n13020 VN.n13006 0.002
R12099 VN.n438 VN.n430 0.002
R12100 VN.n718 VN.n709 0.002
R12101 VN.n1110 VN.n1102 0.002
R12102 VN.n1393 VN.n1384 0.002
R12103 VN.n2106 VN.n1789 0.002
R12104 VN.n2105 VN.n1797 0.002
R12105 VN.n2814 VN.n2806 0.002
R12106 VN.n2782 VN.n2768 0.002
R12107 VN.n12582 VN.n12573 0.002
R12108 VN.n13053 VN.n13029 0.002
R12109 VN.n13051 VN.n13037 0.002
R12110 VN.n453 VN.n445 0.002
R12111 VN.n734 VN.n725 0.002
R12112 VN.n1432 VN.n1117 0.002
R12113 VN.n1431 VN.n1125 0.002
R12114 VN.n2121 VN.n2113 0.002
R12115 VN.n2089 VN.n2075 0.002
R12116 VN.n12598 VN.n12589 0.002
R12117 VN.n13084 VN.n13060 0.002
R12118 VN.n13082 VN.n13068 0.002
R12119 VN.n772 VN.n460 0.002
R12120 VN.n771 VN.n468 0.002
R12121 VN.n1447 VN.n1439 0.002
R12122 VN.n1415 VN.n1401 0.002
R12123 VN.n12756 VN.n12748 0.002
R12124 VN.n13104 VN.n13096 0.002
R12125 VN.n12614 VN.n12606 0.002
R12126 VN.n755 VN.n747 0.002
R12127 VN.n794 VN.n785 0.002
R12128 VN.n12737 VN.n12720 0.002
R12129 VN.n12233 VN.n12225 0.002
R12130 VN.n12385 VN.n12377 0.002
R12131 VN.n14 VN.n12 0.002
R12132 VN.n14 VN.n13 0.002
R12133 VN.n2320 VN.n2305 0.002
R12134 VN.n925 VN.n906 0.002
R12135 VN.n253 VN.n244 0.002
R12136 VN.n3782 VN.n3767 0.002
R12137 VN.n5314 VN.n5299 0.002
R12138 VN.t76 VN.n6593 0.002
R12139 VN.n8583 VN.n8568 0.002
R12140 VN.n10328 VN.n10313 0.002
R12141 VN.n11567 VN.n11561 0.002
R12142 VN.n9843 VN.n9842 0.002
R12143 VN.n8997 VN.n8996 0.002
R12144 VN.n8164 VN.n8163 0.002
R12145 VN.n7353 VN.n7352 0.002
R12146 VN.n6560 VN.n6559 0.002
R12147 VN.n5784 VN.n5783 0.002
R12148 VN.n5021 VN.n5020 0.002
R12149 VN.n4280 VN.n4279 0.002
R12150 VN.n3552 VN.n3551 0.002
R12151 VN.n2846 VN.n2845 0.002
R12152 VN.n2153 VN.n2152 0.002
R12153 VN.n1479 VN.n1478 0.002
R12154 VN.n24 VN.n23 0.002
R12155 VN.n90 VN.n89 0.002
R12156 VN.t8 VN.n11681 0.002
R12157 VN.n11506 VN.n11505 0.002
R12158 VN.n12253 VN.n12252 0.002
R12159 VN.n1606 VN.n1605 0.002
R12160 VN.n3033 VN.n3032 0.002
R12161 VN.n4530 VN.n4529 0.002
R12162 VN.n6097 VN.n6096 0.002
R12163 VN.n7729 VN.n7728 0.002
R12164 VN.n9436 VN.n9435 0.002
R12165 VN.n10174 VN.n10173 0.002
R12166 VN.n9664 VN.n9663 0.002
R12167 VN.n9292 VN.n9291 0.002
R12168 VN.n8802 VN.n8801 0.002
R12169 VN.n8430 VN.n8429 0.002
R12170 VN.n7953 VN.n7952 0.002
R12171 VN.n7585 VN.n7584 0.002
R12172 VN.n6762 VN.n6761 0.002
R12173 VN.n7196 VN.n7195 0.002
R12174 VN.n6317 VN.n6316 0.002
R12175 VN.n5953 VN.n5952 0.002
R12176 VN.n5525 VN.n5524 0.002
R12177 VN.n5161 VN.n5160 0.002
R12178 VN.n4746 VN.n4745 0.002
R12179 VN.n4386 VN.n4385 0.002
R12180 VN.n3989 VN.n3988 0.002
R12181 VN.n3629 VN.n3628 0.002
R12182 VN.n3245 VN.n3244 0.002
R12183 VN.n2889 VN.n2888 0.002
R12184 VN.n2523 VN.n2522 0.002
R12185 VN.n10507 VN.n10506 0.002
R12186 VN.n10111 VN.n10110 0.002
R12187 VN.n9630 VN.n9629 0.002
R12188 VN.n9229 VN.n9228 0.002
R12189 VN.n8768 VN.n8767 0.002
R12190 VN.n8367 VN.n8366 0.002
R12191 VN.n7919 VN.n7918 0.002
R12192 VN.n7522 VN.n7521 0.002
R12193 VN.n6728 VN.n6727 0.002
R12194 VN.n7133 VN.n7132 0.002
R12195 VN.n6283 VN.n6282 0.002
R12196 VN.n5890 VN.n5889 0.002
R12197 VN.n5491 VN.n5490 0.002
R12198 VN.n5098 VN.n5097 0.002
R12199 VN.n4712 VN.n4711 0.002
R12200 VN.n4323 VN.n4322 0.002
R12201 VN.n3955 VN.n3954 0.002
R12202 VN.n10472 VN.n10471 0.002
R12203 VN.n10048 VN.n10047 0.002
R12204 VN.n9596 VN.n9595 0.002
R12205 VN.n9166 VN.n9165 0.002
R12206 VN.n8734 VN.n8733 0.002
R12207 VN.n8304 VN.n8303 0.002
R12208 VN.n7885 VN.n7884 0.002
R12209 VN.n7459 VN.n7458 0.002
R12210 VN.n6694 VN.n6693 0.002
R12211 VN.n7070 VN.n7069 0.002
R12212 VN.n6249 VN.n6248 0.002
R12213 VN.n5827 VN.n5826 0.002
R12214 VN.n5457 VN.n5456 0.002
R12215 VN.n11273 VN.n11272 0.002
R12216 VN.n10864 VN.n10863 0.002
R12217 VN.n10437 VN.n10436 0.002
R12218 VN.n9985 VN.n9984 0.002
R12219 VN.n9562 VN.n9561 0.002
R12220 VN.n9103 VN.n9102 0.002
R12221 VN.n8700 VN.n8699 0.002
R12222 VN.n8241 VN.n8240 0.002
R12223 VN.n7851 VN.n7850 0.002
R12224 VN.n7396 VN.n7395 0.002
R12225 VN.n6660 VN.n6659 0.002
R12226 VN.n10402 VN.n10401 0.002
R12227 VN.n9922 VN.n9921 0.002
R12228 VN.n9528 VN.n9527 0.002
R12229 VN.n9040 VN.n9039 0.002
R12230 VN.n8666 VN.n8665 0.002
R12231 VN.n10367 VN.n10366 0.002
R12232 VN.n10691 VN.n10684 0.002
R12233 VN.n9811 VN.n9804 0.002
R12234 VN.n8965 VN.n8958 0.002
R12235 VN.n8132 VN.n8125 0.002
R12236 VN.n6612 VN.n6605 0.002
R12237 VN.n6528 VN.n6521 0.002
R12238 VN.n5752 VN.n5745 0.002
R12239 VN.n4989 VN.n4982 0.002
R12240 VN.n4248 VN.n4241 0.002
R12241 VN.n3520 VN.n3513 0.002
R12242 VN.n2814 VN.n2807 0.002
R12243 VN.n2121 VN.n2114 0.002
R12244 VN.n1447 VN.n1440 0.002
R12245 VN.n12756 VN.n12755 0.002
R12246 VN.n13104 VN.n13103 0.002
R12247 VN.n12614 VN.n12613 0.002
R12248 VN.n12233 VN.n12232 0.002
R12249 VN.n12385 VN.n12384 0.002
R12250 VN.n2304 VN.n2303 0.002
R12251 VN.n3766 VN.n3765 0.002
R12252 VN.n5298 VN.n5297 0.002
R12253 VN.n8567 VN.n8566 0.002
R12254 VN.n10312 VN.n10311 0.002
R12255 VN.n12713 VN.n12704 0.002
R12256 VN.n227 VN.n210 0.002
R12257 VN.n524 VN.n515 0.002
R12258 VN.n898 VN.n881 0.002
R12259 VN.n1199 VN.n1190 0.002
R12260 VN.n1581 VN.n1564 0.002
R12261 VN.n1889 VN.n1880 0.002
R12262 VN.n2289 VN.n2272 0.002
R12263 VN.n2598 VN.n2589 0.002
R12264 VN.n3011 VN.n2994 0.002
R12265 VN.n3320 VN.n3311 0.002
R12266 VN.n3751 VN.n3734 0.002
R12267 VN.n4064 VN.n4055 0.002
R12268 VN.n4508 VN.n4491 0.002
R12269 VN.n4821 VN.n4812 0.002
R12270 VN.n5283 VN.n5266 0.002
R12271 VN.n5600 VN.n5591 0.002
R12272 VN.n6075 VN.n6058 0.002
R12273 VN.n6392 VN.n6383 0.002
R12274 VN.n7318 VN.n7301 0.002
R12275 VN.n6837 VN.n6828 0.002
R12276 VN.n7707 VN.n7690 0.002
R12277 VN.n8028 VN.n8019 0.002
R12278 VN.n8552 VN.n8535 0.002
R12279 VN.n8877 VN.n8868 0.002
R12280 VN.n9414 VN.n9397 0.002
R12281 VN.n9739 VN.n9730 0.002
R12282 VN.n10297 VN.n10280 0.002
R12283 VN.n10627 VN.n10617 0.002
R12284 VN.n11465 VN.n11449 0.002
R12285 VN.n11118 VN.n11109 0.002
R12286 VN.n3228 VN.n3219 0.002
R12287 VN.n3600 VN.n3583 0.002
R12288 VN.n3972 VN.n3963 0.002
R12289 VN.n4357 VN.n4340 0.002
R12290 VN.n4729 VN.n4720 0.002
R12291 VN.n5132 VN.n5115 0.002
R12292 VN.n5508 VN.n5499 0.002
R12293 VN.n5924 VN.n5907 0.002
R12294 VN.n6300 VN.n6291 0.002
R12295 VN.n7167 VN.n7150 0.002
R12296 VN.n6745 VN.n6736 0.002
R12297 VN.n7556 VN.n7539 0.002
R12298 VN.n7936 VN.n7927 0.002
R12299 VN.n8401 VN.n8384 0.002
R12300 VN.n8785 VN.n8776 0.002
R12301 VN.n9263 VN.n9246 0.002
R12302 VN.n9647 VN.n9638 0.002
R12303 VN.n10145 VN.n10128 0.002
R12304 VN.n10525 VN.n10515 0.002
R12305 VN.n11009 VN.n10997 0.002
R12306 VN.n11188 VN.n11179 0.002
R12307 VN.n11036 VN.n11035 0.002
R12308 VN.n11172 VN.n11171 0.002
R12309 VN.n4695 VN.n4686 0.002
R12310 VN.n5069 VN.n5052 0.002
R12311 VN.n5474 VN.n5465 0.002
R12312 VN.n5861 VN.n5844 0.002
R12313 VN.n6266 VN.n6257 0.002
R12314 VN.n7104 VN.n7087 0.002
R12315 VN.n6711 VN.n6702 0.002
R12316 VN.n7493 VN.n7476 0.002
R12317 VN.n7902 VN.n7893 0.002
R12318 VN.n8338 VN.n8321 0.002
R12319 VN.n8751 VN.n8742 0.002
R12320 VN.n9200 VN.n9183 0.002
R12321 VN.n9613 VN.n9604 0.002
R12322 VN.n10082 VN.n10065 0.002
R12323 VN.n10490 VN.n10480 0.002
R12324 VN.n10951 VN.n10939 0.002
R12325 VN.n11222 VN.n11213 0.002
R12326 VN.n10980 VN.n10979 0.002
R12327 VN.n11206 VN.n11205 0.002
R12328 VN.n6232 VN.n6223 0.002
R12329 VN.n7041 VN.n7024 0.002
R12330 VN.n6677 VN.n6668 0.002
R12331 VN.n7430 VN.n7413 0.002
R12332 VN.n7868 VN.n7859 0.002
R12333 VN.n8275 VN.n8258 0.002
R12334 VN.n8717 VN.n8708 0.002
R12335 VN.n9137 VN.n9120 0.002
R12336 VN.n9579 VN.n9570 0.002
R12337 VN.n10019 VN.n10002 0.002
R12338 VN.n10455 VN.n10445 0.002
R12339 VN.n10893 VN.n10881 0.002
R12340 VN.n11256 VN.n11247 0.002
R12341 VN.n10922 VN.n10921 0.002
R12342 VN.n11240 VN.n11239 0.002
R12343 VN.n7834 VN.n7825 0.002
R12344 VN.n8212 VN.n8195 0.002
R12345 VN.n8683 VN.n8674 0.002
R12346 VN.n9074 VN.n9057 0.002
R12347 VN.n9545 VN.n9536 0.002
R12348 VN.n9956 VN.n9939 0.002
R12349 VN.n10420 VN.n10410 0.002
R12350 VN.n10835 VN.n10823 0.002
R12351 VN.n11289 VN.n11281 0.002
R12352 VN.n9511 VN.n9502 0.002
R12353 VN.n9893 VN.n9876 0.002
R12354 VN.n10385 VN.n10375 0.002
R12355 VN.n10777 VN.n10765 0.002
R12356 VN.n11323 VN.n11314 0.002
R12357 VN.n10806 VN.n10805 0.002
R12358 VN.n11307 VN.n11306 0.002
R12359 VN.n11357 VN.n11348 0.002
R12360 VN.n10748 VN.n10747 0.002
R12361 VN.n11341 VN.n11340 0.002
R12362 VN.n12630 VN.n12346 0.002
R12363 VN.n12632 VN.n12322 0.002
R12364 VN.n12343 VN.n12330 0.002
R12365 VN.n288 VN.n281 0.002
R12366 VN.n558 VN.n550 0.002
R12367 VN.n960 VN.n953 0.002
R12368 VN.n1233 VN.n1225 0.002
R12369 VN.n1647 VN.n1640 0.002
R12370 VN.n1923 VN.n1915 0.002
R12371 VN.n2355 VN.n2348 0.002
R12372 VN.n2632 VN.n2624 0.002
R12373 VN.n3074 VN.n3067 0.002
R12374 VN.n3354 VN.n3346 0.002
R12375 VN.n3817 VN.n3810 0.002
R12376 VN.n4098 VN.n4090 0.002
R12377 VN.n4571 VN.n4564 0.002
R12378 VN.n4855 VN.n4847 0.002
R12379 VN.n5349 VN.n5342 0.002
R12380 VN.n5634 VN.n5626 0.002
R12381 VN.n6138 VN.n6131 0.002
R12382 VN.n6426 VN.n6418 0.002
R12383 VN.n6987 VN.n6980 0.002
R12384 VN.n6871 VN.n6863 0.002
R12385 VN.n7770 VN.n7763 0.002
R12386 VN.n8062 VN.n8054 0.002
R12387 VN.n8618 VN.n8611 0.002
R12388 VN.n8911 VN.n8903 0.002
R12389 VN.n9796 VN.n9470 0.002
R12390 VN.n9795 VN.n9478 0.002
R12391 VN.n10644 VN.n10643 0.002
R12392 VN.n12422 VN.n12414 0.002
R12393 VN.n12663 VN.n12640 0.002
R12394 VN.n12661 VN.n12648 0.002
R12395 VN.n303 VN.n296 0.002
R12396 VN.n574 VN.n566 0.002
R12397 VN.n975 VN.n968 0.002
R12398 VN.n1249 VN.n1241 0.002
R12399 VN.n1662 VN.n1655 0.002
R12400 VN.n1939 VN.n1931 0.002
R12401 VN.n2370 VN.n2363 0.002
R12402 VN.n2648 VN.n2640 0.002
R12403 VN.n3089 VN.n3082 0.002
R12404 VN.n3370 VN.n3362 0.002
R12405 VN.n3832 VN.n3825 0.002
R12406 VN.n4114 VN.n4106 0.002
R12407 VN.n4586 VN.n4579 0.002
R12408 VN.n4871 VN.n4863 0.002
R12409 VN.n5364 VN.n5357 0.002
R12410 VN.n5650 VN.n5642 0.002
R12411 VN.n6153 VN.n6146 0.002
R12412 VN.n6442 VN.n6434 0.002
R12413 VN.n6972 VN.n6965 0.002
R12414 VN.n6887 VN.n6879 0.002
R12415 VN.n7785 VN.n7778 0.002
R12416 VN.n8078 VN.n8070 0.002
R12417 VN.n8950 VN.n8626 0.002
R12418 VN.n8949 VN.n8634 0.002
R12419 VN.n9779 VN.n9778 0.002
R12420 VN.n12438 VN.n12430 0.002
R12421 VN.n12774 VN.n12671 0.002
R12422 VN.n12772 VN.n12679 0.002
R12423 VN.n318 VN.n311 0.002
R12424 VN.n590 VN.n582 0.002
R12425 VN.n990 VN.n983 0.002
R12426 VN.n1265 VN.n1257 0.002
R12427 VN.n1677 VN.n1670 0.002
R12428 VN.n1955 VN.n1947 0.002
R12429 VN.n2385 VN.n2378 0.002
R12430 VN.n2664 VN.n2656 0.002
R12431 VN.n3104 VN.n3097 0.002
R12432 VN.n3386 VN.n3378 0.002
R12433 VN.n3847 VN.n3840 0.002
R12434 VN.n4130 VN.n4122 0.002
R12435 VN.n4601 VN.n4594 0.002
R12436 VN.n4887 VN.n4879 0.002
R12437 VN.n5379 VN.n5372 0.002
R12438 VN.n5666 VN.n5658 0.002
R12439 VN.n6168 VN.n6161 0.002
R12440 VN.n6458 VN.n6450 0.002
R12441 VN.n6957 VN.n6950 0.002
R12442 VN.n6903 VN.n6895 0.002
R12443 VN.n8117 VN.n7793 0.002
R12444 VN.n8116 VN.n7801 0.002
R12445 VN.n8933 VN.n8932 0.002
R12446 VN.n12454 VN.n12446 0.002
R12447 VN.n12808 VN.n12782 0.002
R12448 VN.n12806 VN.n12793 0.002
R12449 VN.n333 VN.n326 0.002
R12450 VN.n606 VN.n598 0.002
R12451 VN.n1005 VN.n998 0.002
R12452 VN.n1281 VN.n1273 0.002
R12453 VN.n1692 VN.n1685 0.002
R12454 VN.n1971 VN.n1963 0.002
R12455 VN.n2400 VN.n2393 0.002
R12456 VN.n2680 VN.n2672 0.002
R12457 VN.n3119 VN.n3112 0.002
R12458 VN.n3402 VN.n3394 0.002
R12459 VN.n3862 VN.n3855 0.002
R12460 VN.n4146 VN.n4138 0.002
R12461 VN.n4616 VN.n4609 0.002
R12462 VN.n4903 VN.n4895 0.002
R12463 VN.n5394 VN.n5387 0.002
R12464 VN.n5682 VN.n5674 0.002
R12465 VN.n6183 VN.n6176 0.002
R12466 VN.n6474 VN.n6466 0.002
R12467 VN.n6942 VN.n6620 0.002
R12468 VN.n6941 VN.n6628 0.002
R12469 VN.n8100 VN.n8099 0.002
R12470 VN.n12470 VN.n12462 0.002
R12471 VN.n12839 VN.n12813 0.002
R12472 VN.n12837 VN.n12824 0.002
R12473 VN.n348 VN.n341 0.002
R12474 VN.n622 VN.n614 0.002
R12475 VN.n1020 VN.n1013 0.002
R12476 VN.n1297 VN.n1289 0.002
R12477 VN.n1707 VN.n1700 0.002
R12478 VN.n1987 VN.n1979 0.002
R12479 VN.n2415 VN.n2408 0.002
R12480 VN.n2696 VN.n2688 0.002
R12481 VN.n3134 VN.n3127 0.002
R12482 VN.n3418 VN.n3410 0.002
R12483 VN.n3877 VN.n3870 0.002
R12484 VN.n4162 VN.n4154 0.002
R12485 VN.n4631 VN.n4624 0.002
R12486 VN.n4919 VN.n4911 0.002
R12487 VN.n5409 VN.n5402 0.002
R12488 VN.n5698 VN.n5690 0.002
R12489 VN.n6513 VN.n6191 0.002
R12490 VN.n6512 VN.n6199 0.002
R12491 VN.n6925 VN.n6924 0.002
R12492 VN.n12486 VN.n12478 0.002
R12493 VN.n12867 VN.n12844 0.002
R12494 VN.n12865 VN.n12852 0.002
R12495 VN.n363 VN.n356 0.002
R12496 VN.n638 VN.n630 0.002
R12497 VN.n1035 VN.n1028 0.002
R12498 VN.n1313 VN.n1305 0.002
R12499 VN.n1722 VN.n1715 0.002
R12500 VN.n2003 VN.n1995 0.002
R12501 VN.n2430 VN.n2423 0.002
R12502 VN.n2712 VN.n2704 0.002
R12503 VN.n3149 VN.n3142 0.002
R12504 VN.n3434 VN.n3426 0.002
R12505 VN.n3892 VN.n3885 0.002
R12506 VN.n4178 VN.n4170 0.002
R12507 VN.n4646 VN.n4639 0.002
R12508 VN.n4935 VN.n4927 0.002
R12509 VN.n5737 VN.n5417 0.002
R12510 VN.n5736 VN.n5425 0.002
R12511 VN.n6496 VN.n6495 0.002
R12512 VN.n12502 VN.n12494 0.002
R12513 VN.n12898 VN.n12875 0.002
R12514 VN.n12896 VN.n12883 0.002
R12515 VN.n378 VN.n371 0.002
R12516 VN.n654 VN.n646 0.002
R12517 VN.n1050 VN.n1043 0.002
R12518 VN.n1329 VN.n1321 0.002
R12519 VN.n1737 VN.n1730 0.002
R12520 VN.n2019 VN.n2011 0.002
R12521 VN.n2445 VN.n2438 0.002
R12522 VN.n2728 VN.n2720 0.002
R12523 VN.n3164 VN.n3157 0.002
R12524 VN.n3450 VN.n3442 0.002
R12525 VN.n3907 VN.n3900 0.002
R12526 VN.n4194 VN.n4186 0.002
R12527 VN.n4974 VN.n4654 0.002
R12528 VN.n4973 VN.n4662 0.002
R12529 VN.n5720 VN.n5719 0.002
R12530 VN.n12518 VN.n12510 0.002
R12531 VN.n12929 VN.n12906 0.002
R12532 VN.n12927 VN.n12914 0.002
R12533 VN.n393 VN.n386 0.002
R12534 VN.n670 VN.n662 0.002
R12535 VN.n1065 VN.n1058 0.002
R12536 VN.n1345 VN.n1337 0.002
R12537 VN.n1752 VN.n1745 0.002
R12538 VN.n2035 VN.n2027 0.002
R12539 VN.n2460 VN.n2453 0.002
R12540 VN.n2744 VN.n2736 0.002
R12541 VN.n3179 VN.n3172 0.002
R12542 VN.n3466 VN.n3458 0.002
R12543 VN.n4233 VN.n3915 0.002
R12544 VN.n4232 VN.n3923 0.002
R12545 VN.n4957 VN.n4956 0.002
R12546 VN.n12534 VN.n12526 0.002
R12547 VN.n12960 VN.n12937 0.002
R12548 VN.n12958 VN.n12945 0.002
R12549 VN.n408 VN.n401 0.002
R12550 VN.n686 VN.n678 0.002
R12551 VN.n1080 VN.n1073 0.002
R12552 VN.n1361 VN.n1353 0.002
R12553 VN.n1767 VN.n1760 0.002
R12554 VN.n2051 VN.n2043 0.002
R12555 VN.n2475 VN.n2468 0.002
R12556 VN.n2760 VN.n2752 0.002
R12557 VN.n3505 VN.n3187 0.002
R12558 VN.n3504 VN.n3195 0.002
R12559 VN.n4216 VN.n4215 0.002
R12560 VN.n12550 VN.n12542 0.002
R12561 VN.n12991 VN.n12968 0.002
R12562 VN.n12989 VN.n12976 0.002
R12563 VN.n423 VN.n416 0.002
R12564 VN.n702 VN.n694 0.002
R12565 VN.n1095 VN.n1088 0.002
R12566 VN.n1377 VN.n1369 0.002
R12567 VN.n1782 VN.n1775 0.002
R12568 VN.n2067 VN.n2059 0.002
R12569 VN.n2799 VN.n2483 0.002
R12570 VN.n2798 VN.n2491 0.002
R12571 VN.n3488 VN.n3487 0.002
R12572 VN.n12566 VN.n12558 0.002
R12573 VN.n13022 VN.n12999 0.002
R12574 VN.n13020 VN.n13007 0.002
R12575 VN.n438 VN.n431 0.002
R12576 VN.n718 VN.n710 0.002
R12577 VN.n1110 VN.n1103 0.002
R12578 VN.n1393 VN.n1385 0.002
R12579 VN.n2106 VN.n1790 0.002
R12580 VN.n2105 VN.n1798 0.002
R12581 VN.n2782 VN.n2781 0.002
R12582 VN.n12582 VN.n12574 0.002
R12583 VN.n13053 VN.n13030 0.002
R12584 VN.n13051 VN.n13038 0.002
R12585 VN.n453 VN.n446 0.002
R12586 VN.n734 VN.n726 0.002
R12587 VN.n1432 VN.n1118 0.002
R12588 VN.n1431 VN.n1126 0.002
R12589 VN.n2089 VN.n2088 0.002
R12590 VN.n12598 VN.n12590 0.002
R12591 VN.n13084 VN.n13061 0.002
R12592 VN.n13082 VN.n13069 0.002
R12593 VN.n772 VN.n461 0.002
R12594 VN.n771 VN.n469 0.002
R12595 VN.n1415 VN.n1414 0.002
R12596 VN.n794 VN.n793 0.002
R12597 VN.n12737 VN.n12736 0.002
R12598 VN.n12405 VN.n12392 0.002
R12599 VN.n12115 VN.n12100 0.002
R12600 VN.n12144 VN.n12141 0.002
R12601 VN.n755 VN.n751 0.002
R12602 VN.n11852 VN.n11849 0.002
R12603 VN.t51 VN.n31 0.002
R12604 VN.t51 VN.n98 0.002
R12605 VN.n12259 VN.n12239 0.002
R12606 VN.n3039 VN.n3020 0.002
R12607 VN.n4536 VN.n4517 0.002
R12608 VN.n6103 VN.n6084 0.002
R12609 VN.n7735 VN.n7716 0.002
R12610 VN.n9442 VN.n9423 0.002
R12611 VN.n11489 VN.n11474 0.002
R12612 VN.n11789 VN.n11788 0.002
R12613 VN.n253 VN.n252 0.002
R12614 VN.n864 VN.n863 0.002
R12615 VN.n1550 VN.n1549 0.002
R12616 VN.n2255 VN.n2254 0.002
R12617 VN.n2977 VN.n2976 0.002
R12618 VN.n3717 VN.n3716 0.002
R12619 VN.n4474 VN.n4473 0.002
R12620 VN.n5249 VN.n5248 0.002
R12621 VN.n6041 VN.n6040 0.002
R12622 VN.n7284 VN.n7283 0.002
R12623 VN.n7673 VN.n7672 0.002
R12624 VN.n8518 VN.n8517 0.002
R12625 VN.n9380 VN.n9379 0.002
R12626 VN.n10263 VN.n10262 0.002
R12627 VN.n9779 VN.n9764 0.002
R12628 VN.n8078 VN.n8077 0.002
R12629 VN.n6887 VN.n6886 0.002
R12630 VN.n6442 VN.n6441 0.002
R12631 VN.n5650 VN.n5649 0.002
R12632 VN.n4871 VN.n4870 0.002
R12633 VN.n4114 VN.n4113 0.002
R12634 VN.n3370 VN.n3369 0.002
R12635 VN.n2648 VN.n2647 0.002
R12636 VN.n1939 VN.n1938 0.002
R12637 VN.n1249 VN.n1248 0.002
R12638 VN.n574 VN.n573 0.002
R12639 VN.n12662 VN.n12661 0.002
R12640 VN.n12422 VN.n12421 0.002
R12641 VN.n8933 VN.n8918 0.002
R12642 VN.n6903 VN.n6902 0.002
R12643 VN.n6458 VN.n6457 0.002
R12644 VN.n5666 VN.n5665 0.002
R12645 VN.n4887 VN.n4886 0.002
R12646 VN.n4130 VN.n4129 0.002
R12647 VN.n3386 VN.n3385 0.002
R12648 VN.n2664 VN.n2663 0.002
R12649 VN.n1955 VN.n1954 0.002
R12650 VN.n1265 VN.n1264 0.002
R12651 VN.n590 VN.n589 0.002
R12652 VN.n12773 VN.n12772 0.002
R12653 VN.n12438 VN.n12437 0.002
R12654 VN.n8100 VN.n8085 0.002
R12655 VN.n6474 VN.n6473 0.002
R12656 VN.n5682 VN.n5681 0.002
R12657 VN.n4903 VN.n4902 0.002
R12658 VN.n4146 VN.n4145 0.002
R12659 VN.n3402 VN.n3401 0.002
R12660 VN.n2680 VN.n2679 0.002
R12661 VN.n1971 VN.n1970 0.002
R12662 VN.n1281 VN.n1280 0.002
R12663 VN.n606 VN.n605 0.002
R12664 VN.n12807 VN.n12806 0.002
R12665 VN.n12454 VN.n12453 0.002
R12666 VN.n6925 VN.n6910 0.002
R12667 VN.n5698 VN.n5697 0.002
R12668 VN.n4919 VN.n4918 0.002
R12669 VN.n4162 VN.n4161 0.002
R12670 VN.n3418 VN.n3417 0.002
R12671 VN.n2696 VN.n2695 0.002
R12672 VN.n1987 VN.n1986 0.002
R12673 VN.n1297 VN.n1296 0.002
R12674 VN.n622 VN.n621 0.002
R12675 VN.n12838 VN.n12837 0.002
R12676 VN.n12470 VN.n12469 0.002
R12677 VN.n6496 VN.n6481 0.002
R12678 VN.n4935 VN.n4934 0.002
R12679 VN.n4178 VN.n4177 0.002
R12680 VN.n3434 VN.n3433 0.002
R12681 VN.n2712 VN.n2711 0.002
R12682 VN.n2003 VN.n2002 0.002
R12683 VN.n1313 VN.n1312 0.002
R12684 VN.n638 VN.n637 0.002
R12685 VN.n12866 VN.n12865 0.002
R12686 VN.n12486 VN.n12485 0.002
R12687 VN.n5720 VN.n5705 0.002
R12688 VN.n4194 VN.n4193 0.002
R12689 VN.n3450 VN.n3449 0.002
R12690 VN.n2728 VN.n2727 0.002
R12691 VN.n2019 VN.n2018 0.002
R12692 VN.n1329 VN.n1328 0.002
R12693 VN.n654 VN.n653 0.002
R12694 VN.n12897 VN.n12896 0.002
R12695 VN.n12502 VN.n12501 0.002
R12696 VN.n4957 VN.n4942 0.002
R12697 VN.n3466 VN.n3465 0.002
R12698 VN.n2744 VN.n2743 0.002
R12699 VN.n2035 VN.n2034 0.002
R12700 VN.n1345 VN.n1344 0.002
R12701 VN.n670 VN.n669 0.002
R12702 VN.n12928 VN.n12927 0.002
R12703 VN.n12518 VN.n12517 0.002
R12704 VN.n4216 VN.n4201 0.002
R12705 VN.n2760 VN.n2759 0.002
R12706 VN.n2051 VN.n2050 0.002
R12707 VN.n1361 VN.n1360 0.002
R12708 VN.n686 VN.n685 0.002
R12709 VN.n12959 VN.n12958 0.002
R12710 VN.n12534 VN.n12533 0.002
R12711 VN.n3488 VN.n3473 0.002
R12712 VN.n2067 VN.n2066 0.002
R12713 VN.n1377 VN.n1376 0.002
R12714 VN.n702 VN.n701 0.002
R12715 VN.n12990 VN.n12989 0.002
R12716 VN.n12550 VN.n12549 0.002
R12717 VN.n2782 VN.n2767 0.002
R12718 VN.n1393 VN.n1392 0.002
R12719 VN.n718 VN.n717 0.002
R12720 VN.n13021 VN.n13020 0.002
R12721 VN.n12566 VN.n12565 0.002
R12722 VN.n2089 VN.n2074 0.002
R12723 VN.n734 VN.n733 0.002
R12724 VN.n13052 VN.n13051 0.002
R12725 VN.n12582 VN.n12581 0.002
R12726 VN.n1415 VN.n1400 0.002
R12727 VN.n13083 VN.n13082 0.002
R12728 VN.n12598 VN.n12597 0.002
R12729 VN.n12614 VN.n12605 0.002
R12730 VN.n1163 VN.n1162 0.002
R12731 VN.n1853 VN.n1852 0.002
R12732 VN.n2562 VN.n2561 0.002
R12733 VN.n3284 VN.n3283 0.002
R12734 VN.n4028 VN.n4027 0.002
R12735 VN.n4785 VN.n4784 0.002
R12736 VN.n5564 VN.n5563 0.002
R12737 VN.n6356 VN.n6355 0.002
R12738 VN.n6801 VN.n6800 0.002
R12739 VN.n7992 VN.n7991 0.002
R12740 VN.n8841 VN.n8840 0.002
R12741 VN.n9703 VN.n9702 0.002
R12742 VN.n10588 VN.n10587 0.002
R12743 VN.n11398 VN.n11397 0.002
R12744 VN.n9757 VN.n9747 0.002
R12745 VN.n8895 VN.n8885 0.002
R12746 VN.n8046 VN.n8036 0.002
R12747 VN.n6855 VN.n6845 0.002
R12748 VN.n6410 VN.n6400 0.002
R12749 VN.n5618 VN.n5608 0.002
R12750 VN.n4839 VN.n4829 0.002
R12751 VN.n4082 VN.n4072 0.002
R12752 VN.n3338 VN.n3328 0.002
R12753 VN.n2616 VN.n2606 0.002
R12754 VN.n1907 VN.n1897 0.002
R12755 VN.n1217 VN.n1207 0.002
R12756 VN.n542 VN.n532 0.002
R12757 VN.n12300 VN.n12299 0.002
R12758 VN.n12283 VN.n12282 0.002
R12759 VN.n10644 VN.n10635 0.002
R12760 VN.n8911 VN.n8910 0.002
R12761 VN.n8062 VN.n8061 0.002
R12762 VN.n6871 VN.n6870 0.002
R12763 VN.n6426 VN.n6425 0.002
R12764 VN.n5634 VN.n5633 0.002
R12765 VN.n4855 VN.n4854 0.002
R12766 VN.n4098 VN.n4097 0.002
R12767 VN.n3354 VN.n3353 0.002
R12768 VN.n2632 VN.n2631 0.002
R12769 VN.n1923 VN.n1922 0.002
R12770 VN.n1233 VN.n1232 0.002
R12771 VN.n558 VN.n557 0.002
R12772 VN.n12344 VN.n12343 0.002
R12773 VN.n12631 VN.n12630 0.002
R12774 VN.n12259 VN.n12238 0.002
R12775 VN.n12713 VN.n12703 0.002
R12776 VN.n227 VN.n200 0.002
R12777 VN.n524 VN.n514 0.002
R12778 VN.n898 VN.n871 0.002
R12779 VN.n1199 VN.n1189 0.002
R12780 VN.n1581 VN.n1554 0.002
R12781 VN.n1889 VN.n1879 0.002
R12782 VN.n2289 VN.n2262 0.002
R12783 VN.n2598 VN.n2588 0.002
R12784 VN.n3011 VN.n2984 0.002
R12785 VN.n3320 VN.n3310 0.002
R12786 VN.n3751 VN.n3724 0.002
R12787 VN.n4064 VN.n4054 0.002
R12788 VN.n4508 VN.n4481 0.002
R12789 VN.n4821 VN.n4811 0.002
R12790 VN.n5283 VN.n5256 0.002
R12791 VN.n5600 VN.n5590 0.002
R12792 VN.n6075 VN.n6048 0.002
R12793 VN.n6392 VN.n6382 0.002
R12794 VN.n7318 VN.n7291 0.002
R12795 VN.n6837 VN.n6827 0.002
R12796 VN.n7707 VN.n7680 0.002
R12797 VN.n8028 VN.n8018 0.002
R12798 VN.n8552 VN.n8525 0.002
R12799 VN.n8877 VN.n8867 0.002
R12800 VN.n9414 VN.n9387 0.002
R12801 VN.n9739 VN.n9729 0.002
R12802 VN.n10297 VN.n10270 0.002
R12803 VN.n10627 VN.n10616 0.002
R12804 VN.n11465 VN.n11448 0.002
R12805 VN.n11118 VN.n11108 0.002
R12806 VN.n12165 VN.n12151 0.002
R12807 VN.n1612 VN.n1589 0.002
R12808 VN.n1831 VN.n1821 0.002
R12809 VN.n2201 VN.n2174 0.002
R12810 VN.n2540 VN.n2530 0.002
R12811 VN.n2923 VN.n2896 0.002
R12812 VN.n3262 VN.n3252 0.002
R12813 VN.n3663 VN.n3636 0.002
R12814 VN.n4006 VN.n3996 0.002
R12815 VN.n4420 VN.n4393 0.002
R12816 VN.n4763 VN.n4753 0.002
R12817 VN.n5195 VN.n5168 0.002
R12818 VN.n5542 VN.n5532 0.002
R12819 VN.n5987 VN.n5960 0.002
R12820 VN.n6334 VN.n6324 0.002
R12821 VN.n7230 VN.n7203 0.002
R12822 VN.n6779 VN.n6769 0.002
R12823 VN.n7619 VN.n7592 0.002
R12824 VN.n7970 VN.n7960 0.002
R12825 VN.n8464 VN.n8437 0.002
R12826 VN.n8819 VN.n8809 0.002
R12827 VN.n9326 VN.n9299 0.002
R12828 VN.n9681 VN.n9671 0.002
R12829 VN.n10209 VN.n10181 0.002
R12830 VN.n10566 VN.n10555 0.002
R12831 VN.n11069 VN.n11048 0.002
R12832 VN.n12081 VN.n12068 0.002
R12833 VN.n11154 VN.n11146 0.002
R12834 VN.n3039 VN.n3019 0.002
R12835 VN.n3228 VN.n3218 0.002
R12836 VN.n3600 VN.n3573 0.002
R12837 VN.n3972 VN.n3962 0.002
R12838 VN.n4357 VN.n4330 0.002
R12839 VN.n4729 VN.n4719 0.002
R12840 VN.n5132 VN.n5105 0.002
R12841 VN.n5508 VN.n5498 0.002
R12842 VN.n5924 VN.n5897 0.002
R12843 VN.n6300 VN.n6290 0.002
R12844 VN.n7167 VN.n7140 0.002
R12845 VN.n6745 VN.n6735 0.002
R12846 VN.n7556 VN.n7529 0.002
R12847 VN.n7936 VN.n7926 0.002
R12848 VN.n8401 VN.n8374 0.002
R12849 VN.n8785 VN.n8775 0.002
R12850 VN.n9263 VN.n9236 0.002
R12851 VN.n9647 VN.n9637 0.002
R12852 VN.n10145 VN.n10118 0.002
R12853 VN.n10525 VN.n10514 0.002
R12854 VN.n11009 VN.n10987 0.002
R12855 VN.n11188 VN.n11187 0.002
R12856 VN.n12036 VN.n12028 0.002
R12857 VN.n4536 VN.n4516 0.002
R12858 VN.n4695 VN.n4685 0.002
R12859 VN.n5069 VN.n5042 0.002
R12860 VN.n5474 VN.n5464 0.002
R12861 VN.n5861 VN.n5834 0.002
R12862 VN.n6266 VN.n6256 0.002
R12863 VN.n7104 VN.n7077 0.002
R12864 VN.n6711 VN.n6701 0.002
R12865 VN.n7493 VN.n7466 0.002
R12866 VN.n7902 VN.n7892 0.002
R12867 VN.n8338 VN.n8311 0.002
R12868 VN.n8751 VN.n8741 0.002
R12869 VN.n9200 VN.n9173 0.002
R12870 VN.n9613 VN.n9603 0.002
R12871 VN.n10082 VN.n10055 0.002
R12872 VN.n10490 VN.n10479 0.002
R12873 VN.n10951 VN.n10929 0.002
R12874 VN.n11222 VN.n11221 0.002
R12875 VN.n11991 VN.n11983 0.002
R12876 VN.n6103 VN.n6083 0.002
R12877 VN.n6232 VN.n6222 0.002
R12878 VN.n7041 VN.n7014 0.002
R12879 VN.n6677 VN.n6667 0.002
R12880 VN.n7430 VN.n7403 0.002
R12881 VN.n7868 VN.n7858 0.002
R12882 VN.n8275 VN.n8248 0.002
R12883 VN.n8717 VN.n8707 0.002
R12884 VN.n9137 VN.n9110 0.002
R12885 VN.n9579 VN.n9569 0.002
R12886 VN.n10019 VN.n9992 0.002
R12887 VN.n10455 VN.n10444 0.002
R12888 VN.n10893 VN.n10871 0.002
R12889 VN.n11256 VN.n11255 0.002
R12890 VN.n11946 VN.n11938 0.002
R12891 VN.n7735 VN.n7715 0.002
R12892 VN.n7834 VN.n7824 0.002
R12893 VN.n8212 VN.n8185 0.002
R12894 VN.n8683 VN.n8673 0.002
R12895 VN.n9074 VN.n9047 0.002
R12896 VN.n9545 VN.n9535 0.002
R12897 VN.n9956 VN.n9929 0.002
R12898 VN.n10420 VN.n10409 0.002
R12899 VN.n10835 VN.n10813 0.002
R12900 VN.n11289 VN.n11280 0.002
R12901 VN.n11897 VN.n11889 0.002
R12902 VN.n9442 VN.n9422 0.002
R12903 VN.n9511 VN.n9501 0.002
R12904 VN.n9893 VN.n9866 0.002
R12905 VN.n10385 VN.n10374 0.002
R12906 VN.n10777 VN.n10755 0.002
R12907 VN.n11323 VN.n11322 0.002
R12908 VN.n11639 VN.n11631 0.002
R12909 VN.n11489 VN.n11473 0.002
R12910 VN.n11357 VN.n11356 0.002
R12911 VN.n11594 VN.n11586 0.002
R12912 VN.n12405 VN.n12393 0.002
R12913 VN.n12128 VN.n12127 0.002
R12914 VN.n11791 VN.n11789 0.002
R12915 VN.n11047 VN.n11046 0.001
R12916 VN.t8 VN.n11791 0.001
R12917 VN.n7378 VN.n7377 0.001
R12918 VN.n8223 VN.n8222 0.001
R12919 VN.n9085 VN.n9084 0.001
R12920 VN.n9967 VN.n9966 0.001
R12921 VN.n10846 VN.n10845 0.001
R12922 VN.n854 VN.n853 0.001
R12923 VN.n1540 VN.n1539 0.001
R12924 VN.n2245 VN.n2244 0.001
R12925 VN.n2967 VN.n2966 0.001
R12926 VN.n3707 VN.n3706 0.001
R12927 VN.n4464 VN.n4463 0.001
R12928 VN.n5239 VN.n5238 0.001
R12929 VN.n6031 VN.n6030 0.001
R12930 VN.n7274 VN.n7273 0.001
R12931 VN.n7663 VN.n7662 0.001
R12932 VN.n8508 VN.n8507 0.001
R12933 VN.n9370 VN.n9369 0.001
R12934 VN.n10253 VN.n10252 0.001
R12935 VN.n11425 VN.n11424 0.001
R12936 VN.n175 VN.n174 0.001
R12937 VN.n11539 VN.n11538 0.001
R12938 VN.n10719 VN.n10718 0.001
R12939 VN.n9859 VN.n9858 0.001
R12940 VN.n9011 VN.n9010 0.001
R12941 VN.n8178 VN.n8177 0.001
R12942 VN.n7367 VN.n7366 0.001
R12943 VN.n6574 VN.n6573 0.001
R12944 VN.n5798 VN.n5797 0.001
R12945 VN.n5035 VN.n5034 0.001
R12946 VN.n4294 VN.n4293 0.001
R12947 VN.n3566 VN.n3565 0.001
R12948 VN.n2860 VN.n2859 0.001
R12949 VN.n2167 VN.n2166 0.001
R12950 VN.n1493 VN.n1492 0.001
R12951 VN.n843 VN.n842 0.001
R12952 VN.n816 VN.n815 0.001
R12953 VN.n13132 VN.n13131 0.001
R12954 VN.n11006 VN.n11005 0.001
R12955 VN.n10948 VN.n10947 0.001
R12956 VN.n10890 VN.n10889 0.001
R12957 VN.n10832 VN.n10831 0.001
R12958 VN.n10774 VN.n10773 0.001
R12959 VN.n828 VN.n827 0.001
R12960 VN.n12722 VN.n12721 0.001
R12961 VN.n10209 VN.n10192 0.001
R12962 VN.n2319 VN.n2318 0.001
R12963 VN.n3781 VN.n3780 0.001
R12964 VN.n5313 VN.n5312 0.001
R12965 VN.n6601 VN.n6600 0.001
R12966 VN.n8582 VN.n8581 0.001
R12967 VN.n10327 VN.n10326 0.001
R12968 VN.n11852 VN.n11843 0.001
R12969 VN.n9 VN.n8 0.001
R12970 VN.n11 VN.n10 0.001
R12971 VN.n11564 VN.n11563 0.001
R12972 VN.n11117 VN.n11116 0.001
R12973 VN.n11462 VN.n11461 0.001
R12974 VN.n10626 VN.n10625 0.001
R12975 VN.n10294 VN.n10293 0.001
R12976 VN.n9738 VN.n9737 0.001
R12977 VN.n9411 VN.n9410 0.001
R12978 VN.n8876 VN.n8875 0.001
R12979 VN.n8549 VN.n8548 0.001
R12980 VN.n8027 VN.n8026 0.001
R12981 VN.n7704 VN.n7703 0.001
R12982 VN.n6836 VN.n6835 0.001
R12983 VN.n7315 VN.n7314 0.001
R12984 VN.n6391 VN.n6390 0.001
R12985 VN.n6072 VN.n6071 0.001
R12986 VN.n5599 VN.n5598 0.001
R12987 VN.n5280 VN.n5279 0.001
R12988 VN.n4820 VN.n4819 0.001
R12989 VN.n4505 VN.n4504 0.001
R12990 VN.n4063 VN.n4062 0.001
R12991 VN.n3748 VN.n3747 0.001
R12992 VN.n3319 VN.n3318 0.001
R12993 VN.n3008 VN.n3007 0.001
R12994 VN.n2597 VN.n2596 0.001
R12995 VN.n2286 VN.n2285 0.001
R12996 VN.n1888 VN.n1887 0.001
R12997 VN.n1578 VN.n1577 0.001
R12998 VN.n1198 VN.n1197 0.001
R12999 VN.n895 VN.n894 0.001
R13000 VN.n523 VN.n522 0.001
R13001 VN.n224 VN.n223 0.001
R13002 VN.n12712 VN.n12711 0.001
R13003 VN.n10554 VN.n10553 0.001
R13004 VN.n10206 VN.n10205 0.001
R13005 VN.n9680 VN.n9679 0.001
R13006 VN.n9323 VN.n9322 0.001
R13007 VN.n8818 VN.n8817 0.001
R13008 VN.n8461 VN.n8460 0.001
R13009 VN.n7969 VN.n7968 0.001
R13010 VN.n7616 VN.n7615 0.001
R13011 VN.n6778 VN.n6777 0.001
R13012 VN.n7227 VN.n7226 0.001
R13013 VN.n6333 VN.n6332 0.001
R13014 VN.n5984 VN.n5983 0.001
R13015 VN.n5541 VN.n5540 0.001
R13016 VN.n5192 VN.n5191 0.001
R13017 VN.n4762 VN.n4761 0.001
R13018 VN.n4417 VN.n4416 0.001
R13019 VN.n4005 VN.n4004 0.001
R13020 VN.n3660 VN.n3659 0.001
R13021 VN.n3261 VN.n3260 0.001
R13022 VN.n2920 VN.n2919 0.001
R13023 VN.n2539 VN.n2538 0.001
R13024 VN.n2198 VN.n2197 0.001
R13025 VN.n1830 VN.n1829 0.001
R13026 VN.n10524 VN.n10523 0.001
R13027 VN.n10142 VN.n10141 0.001
R13028 VN.n9646 VN.n9645 0.001
R13029 VN.n9260 VN.n9259 0.001
R13030 VN.n8784 VN.n8783 0.001
R13031 VN.n8398 VN.n8397 0.001
R13032 VN.n7935 VN.n7934 0.001
R13033 VN.n7553 VN.n7552 0.001
R13034 VN.n6744 VN.n6743 0.001
R13035 VN.n7164 VN.n7163 0.001
R13036 VN.n6299 VN.n6298 0.001
R13037 VN.n5921 VN.n5920 0.001
R13038 VN.n5507 VN.n5506 0.001
R13039 VN.n5129 VN.n5128 0.001
R13040 VN.n4728 VN.n4727 0.001
R13041 VN.n4354 VN.n4353 0.001
R13042 VN.n3971 VN.n3970 0.001
R13043 VN.n3597 VN.n3596 0.001
R13044 VN.n3227 VN.n3226 0.001
R13045 VN.n10489 VN.n10488 0.001
R13046 VN.n10079 VN.n10078 0.001
R13047 VN.n9612 VN.n9611 0.001
R13048 VN.n9197 VN.n9196 0.001
R13049 VN.n8750 VN.n8749 0.001
R13050 VN.n8335 VN.n8334 0.001
R13051 VN.n7901 VN.n7900 0.001
R13052 VN.n7490 VN.n7489 0.001
R13053 VN.n6710 VN.n6709 0.001
R13054 VN.n7101 VN.n7100 0.001
R13055 VN.n6265 VN.n6264 0.001
R13056 VN.n5858 VN.n5857 0.001
R13057 VN.n5473 VN.n5472 0.001
R13058 VN.n5066 VN.n5065 0.001
R13059 VN.n4694 VN.n4693 0.001
R13060 VN.n10454 VN.n10453 0.001
R13061 VN.n10016 VN.n10015 0.001
R13062 VN.n9578 VN.n9577 0.001
R13063 VN.n9134 VN.n9133 0.001
R13064 VN.n8716 VN.n8715 0.001
R13065 VN.n8272 VN.n8271 0.001
R13066 VN.n7867 VN.n7866 0.001
R13067 VN.n7427 VN.n7426 0.001
R13068 VN.n6676 VN.n6675 0.001
R13069 VN.n7038 VN.n7037 0.001
R13070 VN.n6231 VN.n6230 0.001
R13071 VN.n10419 VN.n10418 0.001
R13072 VN.n9953 VN.n9952 0.001
R13073 VN.n9544 VN.n9543 0.001
R13074 VN.n9071 VN.n9070 0.001
R13075 VN.n8682 VN.n8681 0.001
R13076 VN.n8209 VN.n8208 0.001
R13077 VN.n7833 VN.n7832 0.001
R13078 VN.n10384 VN.n10383 0.001
R13079 VN.n9890 VN.n9889 0.001
R13080 VN.n9510 VN.n9509 0.001
R13081 VN.n12395 VN.n12394 0.001
R13082 VN.n11852 VN.n11846 0.001
R13083 VN.n2871 VN.n2870 0.001
R13084 VN.n3611 VN.n3610 0.001
R13085 VN.n4368 VN.n4367 0.001
R13086 VN.n5143 VN.n5142 0.001
R13087 VN.n5935 VN.n5934 0.001
R13088 VN.n7178 VN.n7177 0.001
R13089 VN.n7567 VN.n7566 0.001
R13090 VN.n8412 VN.n8411 0.001
R13091 VN.n9274 VN.n9273 0.001
R13092 VN.n10156 VN.n10155 0.001
R13093 VN.n11021 VN.n11020 0.001
R13094 VN.n4305 VN.n4304 0.001
R13095 VN.n5080 VN.n5079 0.001
R13096 VN.n5872 VN.n5871 0.001
R13097 VN.n7115 VN.n7114 0.001
R13098 VN.n7504 VN.n7503 0.001
R13099 VN.n8349 VN.n8348 0.001
R13100 VN.n9211 VN.n9210 0.001
R13101 VN.n10093 VN.n10092 0.001
R13102 VN.n10963 VN.n10962 0.001
R13103 VN.n5809 VN.n5808 0.001
R13104 VN.n7052 VN.n7051 0.001
R13105 VN.n7441 VN.n7440 0.001
R13106 VN.n8286 VN.n8285 0.001
R13107 VN.n9148 VN.n9147 0.001
R13108 VN.n10030 VN.n10029 0.001
R13109 VN.n10905 VN.n10904 0.001
R13110 VN.n9022 VN.n9021 0.001
R13111 VN.n9904 VN.n9903 0.001
R13112 VN.n10789 VN.n10788 0.001
R13113 VN.n10731 VN.n10730 0.001
R13114 VN.n11100 VN.n11091 0.001
R13115 VN.n11373 VN.n11372 0.001
R13116 VN.n10346 VN.n10345 0.001
R13117 VN.n9491 VN.n9490 0.001
R13118 VN.n8645 VN.n8644 0.001
R13119 VN.n7814 VN.n7813 0.001
R13120 VN.n6639 VN.n6638 0.001
R13121 VN.n6210 VN.n6209 0.001
R13122 VN.n5436 VN.n5435 0.001
R13123 VN.n4675 VN.n4674 0.001
R13124 VN.n3934 VN.n3933 0.001
R13125 VN.n3208 VN.n3207 0.001
R13126 VN.n2502 VN.n2501 0.001
R13127 VN.n1811 VN.n1810 0.001
R13128 VN.n1137 VN.n1136 0.001
R13129 VN.n485 VN.n484 0.001
R13130 VN.n12692 VN.n12691 0.001
R13131 VN.n12362 VN.n12361 0.001
R13132 VN.n176 VN.n175 0.001
R13133 VN.t8 VN.n11703 0.001
R13134 VN.n11867 VN.t8 0.001
R13135 VN.t8 VN.n11669 0.001
R13136 VN.t8 VN.n11717 0.001
R13137 VN.t8 VN.n11728 0.001
R13138 VN.t8 VN.n11739 0.001
R13139 VN.t8 VN.n11750 0.001
R13140 VN.t8 VN.n11761 0.001
R13141 VN.t8 VN.n11770 0.001
R13142 VN.n2201 VN.n2184 0.001
R13143 VN.n2923 VN.n2906 0.001
R13144 VN.n3663 VN.n3646 0.001
R13145 VN.n4420 VN.n4403 0.001
R13146 VN.n5195 VN.n5178 0.001
R13147 VN.n5987 VN.n5970 0.001
R13148 VN.n7230 VN.n7213 0.001
R13149 VN.n7619 VN.n7602 0.001
R13150 VN.n8464 VN.n8447 0.001
R13151 VN.n9326 VN.n9309 0.001
R13152 VN.n182 VN.n170 0.001
R13153 VN.n12367 VN.n12366 0.001
R13154 VN.n2508 VN.n2507 0.001
R13155 VN.n1143 VN.n1142 0.001
R13156 VN.n490 VN.n489 0.001
R13157 VN.n12698 VN.n12697 0.001
R13158 VN.n1816 VN.n1815 0.001
R13159 VN.n3940 VN.n3939 0.001
R13160 VN.n3213 VN.n3212 0.001
R13161 VN.n5442 VN.n5441 0.001
R13162 VN.n4680 VN.n4679 0.001
R13163 VN.n6217 VN.n6216 0.001
R13164 VN.n6645 VN.n6644 0.001
R13165 VN.n8651 VN.n8650 0.001
R13166 VN.n7819 VN.n7818 0.001
R13167 VN.n10352 VN.n10351 0.001
R13168 VN.n9496 VN.n9495 0.001
R13169 VN.n11380 VN.n11379 0.001
R13170 VN.n11852 VN.n11851 0.001
R13171 VN.n1612 VN.n1591 0.001
R13172 VN.n12282 VN.n12281 0.001
R13173 VN.n12314 VN.n12313 0.001
R13174 VN.n12299 VN.n12298 0.001
R13175 VN.n273 VN.n272 0.001
R13176 VN.n542 VN.n541 0.001
R13177 VN.n945 VN.n944 0.001
R13178 VN.n1217 VN.n1216 0.001
R13179 VN.n1632 VN.n1631 0.001
R13180 VN.n1907 VN.n1906 0.001
R13181 VN.n2340 VN.n2339 0.001
R13182 VN.n2616 VN.n2615 0.001
R13183 VN.n3059 VN.n3058 0.001
R13184 VN.n3338 VN.n3337 0.001
R13185 VN.n3802 VN.n3801 0.001
R13186 VN.n4082 VN.n4081 0.001
R13187 VN.n4556 VN.n4555 0.001
R13188 VN.n4839 VN.n4838 0.001
R13189 VN.n5334 VN.n5333 0.001
R13190 VN.n5618 VN.n5617 0.001
R13191 VN.n6123 VN.n6122 0.001
R13192 VN.n6410 VN.n6409 0.001
R13193 VN.n7007 VN.n7006 0.001
R13194 VN.n6855 VN.n6854 0.001
R13195 VN.n7755 VN.n7754 0.001
R13196 VN.n8046 VN.n8045 0.001
R13197 VN.n8603 VN.n8602 0.001
R13198 VN.n8895 VN.n8894 0.001
R13199 VN.n9462 VN.n9461 0.001
R13200 VN.n9757 VN.n9756 0.001
R13201 VN.n10676 VN.n10675 0.001
R13202 VN.n10662 VN.n10661 0.001
R13203 VN.n12375 VN.n12374 0.001
R13204 VN.n11575 VN.n11572 0.001
R13205 VN.t160 VN.n11575 0.001
R13206 VN.t35 VN.n11380 0.001
R13207 VN.t82 VN.n12367 0.001
R13208 VN.t57 VN.n2508 0.001
R13209 VN.t108 VN.n1816 0.001
R13210 VN.t94 VN.n1143 0.001
R13211 VN.t41 VN.n490 0.001
R13212 VN.t101 VN.n12698 0.001
R13213 VN.t28 VN.n3940 0.001
R13214 VN.t183 VN.n3213 0.001
R13215 VN.t176 VN.n5442 0.001
R13216 VN.t32 VN.n4680 0.001
R13217 VN.t146 VN.n6217 0.001
R13218 VN.t253 VN.n6645 0.001
R13219 VN.t39 VN.n8651 0.001
R13220 VN.t73 VN.n7819 0.001
R13221 VN.t241 VN.n10352 0.001
R13222 VN.t0 VN.n9496 0.001
R13223 VN.n170 VN.t51 0.001
R13224 VN.n11852 VN.n11850 0.001
R13225 VN.n14 VN.n3 0.001
R13226 VN.n11525 VN.n11524 0.001
R13227 VN.n11372 VN.n11371 0.001
R13228 VN.n10345 VN.n10344 0.001
R13229 VN.n9490 VN.n9489 0.001
R13230 VN.n8644 VN.n8643 0.001
R13231 VN.n7813 VN.n7812 0.001
R13232 VN.n6638 VN.n6637 0.001
R13233 VN.n6209 VN.n6208 0.001
R13234 VN.n5435 VN.n5434 0.001
R13235 VN.n4674 VN.n4673 0.001
R13236 VN.n3933 VN.n3932 0.001
R13237 VN.n3207 VN.n3206 0.001
R13238 VN.n2501 VN.n2500 0.001
R13239 VN.n1810 VN.n1809 0.001
R13240 VN.n1136 VN.n1135 0.001
R13241 VN.n484 VN.n483 0.001
R13242 VN.n12691 VN.n12690 0.001
R13243 VN.n12361 VN.n12360 0.001
R13244 VN.n11154 VN.n11145 0.001
R13245 VN.n11852 VN.n11845 0.001
R13246 VN.n11852 VN.n11844 0.001
R13247 VN.n11852 VN.n11842 0.001
R13248 VN.n11852 VN.n11841 0.001
R13249 VN.n11852 VN.n11848 0.001
R13250 VN.n11188 VN.n11186 0.001
R13251 VN.n11222 VN.n11220 0.001
R13252 VN.n11256 VN.n11254 0.001
R13253 VN.n11323 VN.n11321 0.001
R13254 VN.n11357 VN.n11355 0.001
R13255 VN.n14 VN.n11 0.001
R13256 VN.n14 VN.n9 0.001
R13257 VN.n11289 VN.n11288 0.001
R13258 VN.n12110 VN.n12109 0.001
R13259 VN.n173 VN.n172 0.001
R13260 VN.n11538 VN.n11537 0.001
R13261 VN.n10718 VN.n10717 0.001
R13262 VN.n9858 VN.n9857 0.001
R13263 VN.n9010 VN.n9009 0.001
R13264 VN.n8177 VN.n8176 0.001
R13265 VN.n7366 VN.n7365 0.001
R13266 VN.n6573 VN.n6572 0.001
R13267 VN.n5797 VN.n5796 0.001
R13268 VN.n5034 VN.n5033 0.001
R13269 VN.n4293 VN.n4292 0.001
R13270 VN.n3565 VN.n3564 0.001
R13271 VN.n2859 VN.n2858 0.001
R13272 VN.n2166 VN.n2165 0.001
R13273 VN.n1492 VN.n1491 0.001
R13274 VN.n842 VN.n841 0.001
R13275 VN.n815 VN.n814 0.001
R13276 VN.n13131 VN.n13130 0.001
R13277 VN.n12158 VN.n12157 0.001
R13278 VN.n12245 VN.n12244 0.001
R13279 VN.n12710 VN.n12709 0.001
R13280 VN.n216 VN.n215 0.001
R13281 VN.n521 VN.n520 0.001
R13282 VN.n887 VN.n886 0.001
R13283 VN.n1196 VN.n1195 0.001
R13284 VN.n1570 VN.n1569 0.001
R13285 VN.n1886 VN.n1885 0.001
R13286 VN.n2278 VN.n2277 0.001
R13287 VN.n2595 VN.n2594 0.001
R13288 VN.n3000 VN.n2999 0.001
R13289 VN.n3317 VN.n3316 0.001
R13290 VN.n3740 VN.n3739 0.001
R13291 VN.n4061 VN.n4060 0.001
R13292 VN.n4497 VN.n4496 0.001
R13293 VN.n4818 VN.n4817 0.001
R13294 VN.n5272 VN.n5271 0.001
R13295 VN.n5597 VN.n5596 0.001
R13296 VN.n6064 VN.n6063 0.001
R13297 VN.n6389 VN.n6388 0.001
R13298 VN.n7307 VN.n7306 0.001
R13299 VN.n6834 VN.n6833 0.001
R13300 VN.n7696 VN.n7695 0.001
R13301 VN.n8025 VN.n8024 0.001
R13302 VN.n8541 VN.n8540 0.001
R13303 VN.n8874 VN.n8873 0.001
R13304 VN.n9403 VN.n9402 0.001
R13305 VN.n9736 VN.n9735 0.001
R13306 VN.n10286 VN.n10285 0.001
R13307 VN.n10623 VN.n10622 0.001
R13308 VN.n11455 VN.n11454 0.001
R13309 VN.n11115 VN.n11114 0.001
R13310 VN.n12031 VN.n12030 0.001
R13311 VN.n3026 VN.n3025 0.001
R13312 VN.n3225 VN.n3224 0.001
R13313 VN.n3589 VN.n3588 0.001
R13314 VN.n3969 VN.n3968 0.001
R13315 VN.n4346 VN.n4345 0.001
R13316 VN.n4726 VN.n4725 0.001
R13317 VN.n5121 VN.n5120 0.001
R13318 VN.n5505 VN.n5504 0.001
R13319 VN.n5913 VN.n5912 0.001
R13320 VN.n6297 VN.n6296 0.001
R13321 VN.n7156 VN.n7155 0.001
R13322 VN.n6742 VN.n6741 0.001
R13323 VN.n7545 VN.n7544 0.001
R13324 VN.n7933 VN.n7932 0.001
R13325 VN.n8390 VN.n8389 0.001
R13326 VN.n8782 VN.n8781 0.001
R13327 VN.n9252 VN.n9251 0.001
R13328 VN.n9644 VN.n9643 0.001
R13329 VN.n10134 VN.n10133 0.001
R13330 VN.n10521 VN.n10520 0.001
R13331 VN.n11003 VN.n11002 0.001
R13332 VN.n11185 VN.n11184 0.001
R13333 VN.n12054 VN.n12053 0.001
R13334 VN.n2308 VN.n2307 0.001
R13335 VN.n2518 VN.n2517 0.001
R13336 VN.n2875 VN.n2874 0.001
R13337 VN.n3240 VN.n3239 0.001
R13338 VN.n3615 VN.n3614 0.001
R13339 VN.n3984 VN.n3983 0.001
R13340 VN.n4372 VN.n4371 0.001
R13341 VN.n4741 VN.n4740 0.001
R13342 VN.n5147 VN.n5146 0.001
R13343 VN.n5520 VN.n5519 0.001
R13344 VN.n5939 VN.n5938 0.001
R13345 VN.n6312 VN.n6311 0.001
R13346 VN.n7182 VN.n7181 0.001
R13347 VN.n6757 VN.n6756 0.001
R13348 VN.n7571 VN.n7570 0.001
R13349 VN.n7948 VN.n7947 0.001
R13350 VN.n8416 VN.n8415 0.001
R13351 VN.n8797 VN.n8796 0.001
R13352 VN.n9278 VN.n9277 0.001
R13353 VN.n9659 VN.n9658 0.001
R13354 VN.n10160 VN.n10159 0.001
R13355 VN.n10537 VN.n10536 0.001
R13356 VN.n10558 VN.n10557 0.001
R13357 VN.n11051 VN.n11050 0.001
R13358 VN.n11149 VN.n11148 0.001
R13359 VN.n12071 VN.n12070 0.001
R13360 VN.n10198 VN.n10197 0.001
R13361 VN.n9315 VN.n9314 0.001
R13362 VN.n8453 VN.n8452 0.001
R13363 VN.n7608 VN.n7607 0.001
R13364 VN.n7219 VN.n7218 0.001
R13365 VN.n5976 VN.n5975 0.001
R13366 VN.n5184 VN.n5183 0.001
R13367 VN.n4409 VN.n4408 0.001
R13368 VN.n3652 VN.n3651 0.001
R13369 VN.n2912 VN.n2911 0.001
R13370 VN.n2190 VN.n2189 0.001
R13371 VN.n1599 VN.n1598 0.001
R13372 VN.n1828 VN.n1827 0.001
R13373 VN.n2537 VN.n2536 0.001
R13374 VN.n3259 VN.n3258 0.001
R13375 VN.n4003 VN.n4002 0.001
R13376 VN.n4760 VN.n4759 0.001
R13377 VN.n5539 VN.n5538 0.001
R13378 VN.n6331 VN.n6330 0.001
R13379 VN.n6776 VN.n6775 0.001
R13380 VN.n7967 VN.n7966 0.001
R13381 VN.n8816 VN.n8815 0.001
R13382 VN.n9678 VN.n9677 0.001
R13383 VN.n11402 VN.n11401 0.001
R13384 VN.n11090 VN.n11089 0.001
R13385 VN.n12105 VN.n12104 0.001
R13386 VN.n920 VN.n919 0.001
R13387 VN.n1161 VN.n1160 0.001
R13388 VN.n1514 VN.n1513 0.001
R13389 VN.n1851 VN.n1850 0.001
R13390 VN.n2222 VN.n2221 0.001
R13391 VN.n2560 VN.n2559 0.001
R13392 VN.n2944 VN.n2943 0.001
R13393 VN.n3282 VN.n3281 0.001
R13394 VN.n3684 VN.n3683 0.001
R13395 VN.n4026 VN.n4025 0.001
R13396 VN.n4441 VN.n4440 0.001
R13397 VN.n4783 VN.n4782 0.001
R13398 VN.n5216 VN.n5215 0.001
R13399 VN.n5562 VN.n5561 0.001
R13400 VN.n6008 VN.n6007 0.001
R13401 VN.n6354 VN.n6353 0.001
R13402 VN.n7251 VN.n7250 0.001
R13403 VN.n6799 VN.n6798 0.001
R13404 VN.n7640 VN.n7639 0.001
R13405 VN.n7990 VN.n7989 0.001
R13406 VN.n8485 VN.n8484 0.001
R13407 VN.n8839 VN.n8838 0.001
R13408 VN.n9347 VN.n9346 0.001
R13409 VN.n9701 VN.n9700 0.001
R13410 VN.n10230 VN.n10229 0.001
R13411 VN.n10586 VN.n10585 0.001
R13412 VN.n11429 VN.n11428 0.001
R13413 VN.n11130 VN.n11129 0.001
R13414 VN.n10606 VN.n10605 0.001
R13415 VN.n10257 VN.n10256 0.001
R13416 VN.n9715 VN.n9714 0.001
R13417 VN.n9374 VN.n9373 0.001
R13418 VN.n8853 VN.n8852 0.001
R13419 VN.n8512 VN.n8511 0.001
R13420 VN.n8004 VN.n8003 0.001
R13421 VN.n7667 VN.n7666 0.001
R13422 VN.n6813 VN.n6812 0.001
R13423 VN.n7278 VN.n7277 0.001
R13424 VN.n6368 VN.n6367 0.001
R13425 VN.n6035 VN.n6034 0.001
R13426 VN.n5576 VN.n5575 0.001
R13427 VN.n5243 VN.n5242 0.001
R13428 VN.n4797 VN.n4796 0.001
R13429 VN.n4468 VN.n4467 0.001
R13430 VN.n4040 VN.n4039 0.001
R13431 VN.n3711 VN.n3710 0.001
R13432 VN.n3296 VN.n3295 0.001
R13433 VN.n2971 VN.n2970 0.001
R13434 VN.n2574 VN.n2573 0.001
R13435 VN.n2249 VN.n2248 0.001
R13436 VN.n1865 VN.n1864 0.001
R13437 VN.n1544 VN.n1543 0.001
R13438 VN.n1175 VN.n1174 0.001
R13439 VN.n858 VN.n857 0.001
R13440 VN.n500 VN.n499 0.001
R13441 VN.n247 VN.n246 0.001
R13442 VN.n12131 VN.n12130 0.001
R13443 VN.n11024 VN.n11023 0.001
R13444 VN.n11167 VN.n11166 0.001
R13445 VN.n11986 VN.n11985 0.001
R13446 VN.n4523 VN.n4522 0.001
R13447 VN.n4692 VN.n4691 0.001
R13448 VN.n5058 VN.n5057 0.001
R13449 VN.n5471 VN.n5470 0.001
R13450 VN.n5850 VN.n5849 0.001
R13451 VN.n6263 VN.n6262 0.001
R13452 VN.n7093 VN.n7092 0.001
R13453 VN.n6708 VN.n6707 0.001
R13454 VN.n7482 VN.n7481 0.001
R13455 VN.n7899 VN.n7898 0.001
R13456 VN.n8327 VN.n8326 0.001
R13457 VN.n8748 VN.n8747 0.001
R13458 VN.n9189 VN.n9188 0.001
R13459 VN.n9610 VN.n9609 0.001
R13460 VN.n10071 VN.n10070 0.001
R13461 VN.n10486 VN.n10485 0.001
R13462 VN.n10945 VN.n10944 0.001
R13463 VN.n11219 VN.n11218 0.001
R13464 VN.n12009 VN.n12008 0.001
R13465 VN.n3770 VN.n3769 0.001
R13466 VN.n3950 VN.n3949 0.001
R13467 VN.n4309 VN.n4308 0.001
R13468 VN.n4707 VN.n4706 0.001
R13469 VN.n5084 VN.n5083 0.001
R13470 VN.n5486 VN.n5485 0.001
R13471 VN.n5876 VN.n5875 0.001
R13472 VN.n6278 VN.n6277 0.001
R13473 VN.n7119 VN.n7118 0.001
R13474 VN.n6723 VN.n6722 0.001
R13475 VN.n7508 VN.n7507 0.001
R13476 VN.n7914 VN.n7913 0.001
R13477 VN.n8353 VN.n8352 0.001
R13478 VN.n8763 VN.n8762 0.001
R13479 VN.n9215 VN.n9214 0.001
R13480 VN.n9625 VN.n9624 0.001
R13481 VN.n10097 VN.n10096 0.001
R13482 VN.n10502 VN.n10501 0.001
R13483 VN.n10966 VN.n10965 0.001
R13484 VN.n11201 VN.n11200 0.001
R13485 VN.n11941 VN.n11940 0.001
R13486 VN.n6090 VN.n6089 0.001
R13487 VN.n6229 VN.n6228 0.001
R13488 VN.n7030 VN.n7029 0.001
R13489 VN.n6674 VN.n6673 0.001
R13490 VN.n7419 VN.n7418 0.001
R13491 VN.n7865 VN.n7864 0.001
R13492 VN.n8264 VN.n8263 0.001
R13493 VN.n8714 VN.n8713 0.001
R13494 VN.n9126 VN.n9125 0.001
R13495 VN.n9576 VN.n9575 0.001
R13496 VN.n10008 VN.n10007 0.001
R13497 VN.n10451 VN.n10450 0.001
R13498 VN.n10887 VN.n10886 0.001
R13499 VN.n11253 VN.n11252 0.001
R13500 VN.n11964 VN.n11963 0.001
R13501 VN.n5302 VN.n5301 0.001
R13502 VN.n5452 VN.n5451 0.001
R13503 VN.n5813 VN.n5812 0.001
R13504 VN.n6244 VN.n6243 0.001
R13505 VN.n7056 VN.n7055 0.001
R13506 VN.n6689 VN.n6688 0.001
R13507 VN.n7445 VN.n7444 0.001
R13508 VN.n7880 VN.n7879 0.001
R13509 VN.n8290 VN.n8289 0.001
R13510 VN.n8729 VN.n8728 0.001
R13511 VN.n9152 VN.n9151 0.001
R13512 VN.n9591 VN.n9590 0.001
R13513 VN.n10034 VN.n10033 0.001
R13514 VN.n10467 VN.n10466 0.001
R13515 VN.n10908 VN.n10907 0.001
R13516 VN.n11235 VN.n11234 0.001
R13517 VN.n6655 VN.n6654 0.001
R13518 VN.n7382 VN.n7381 0.001
R13519 VN.n7846 VN.n7845 0.001
R13520 VN.n8227 VN.n8226 0.001
R13521 VN.n8695 VN.n8694 0.001
R13522 VN.n9089 VN.n9088 0.001
R13523 VN.n9557 VN.n9556 0.001
R13524 VN.n9971 VN.n9970 0.001
R13525 VN.n10432 VN.n10431 0.001
R13526 VN.n10850 VN.n10849 0.001
R13527 VN.n11268 VN.n11267 0.001
R13528 VN.n11915 VN.n11914 0.001
R13529 VN.n11892 VN.n11891 0.001
R13530 VN.n7722 VN.n7721 0.001
R13531 VN.n7831 VN.n7830 0.001
R13532 VN.n8201 VN.n8200 0.001
R13533 VN.n8680 VN.n8679 0.001
R13534 VN.n9063 VN.n9062 0.001
R13535 VN.n9542 VN.n9541 0.001
R13536 VN.n9945 VN.n9944 0.001
R13537 VN.n10416 VN.n10415 0.001
R13538 VN.n10829 VN.n10828 0.001
R13539 VN.n11287 VN.n11286 0.001
R13540 VN.n11634 VN.n11633 0.001
R13541 VN.n9429 VN.n9428 0.001
R13542 VN.n9508 VN.n9507 0.001
R13543 VN.n9882 VN.n9881 0.001
R13544 VN.n10381 VN.n10380 0.001
R13545 VN.n10771 VN.n10770 0.001
R13546 VN.n11320 VN.n11319 0.001
R13547 VN.n11871 VN.n11870 0.001
R13548 VN.n8571 VN.n8570 0.001
R13549 VN.n8661 VN.n8660 0.001
R13550 VN.n9026 VN.n9025 0.001
R13551 VN.n9523 VN.n9522 0.001
R13552 VN.n9908 VN.n9907 0.001
R13553 VN.n10397 VN.n10396 0.001
R13554 VN.n10792 VN.n10791 0.001
R13555 VN.n11302 VN.n11301 0.001
R13556 VN.n11589 VN.n11588 0.001
R13557 VN.n11480 VN.n11479 0.001
R13558 VN.n11354 VN.n11353 0.001
R13559 VN.n11612 VN.n11611 0.001
R13560 VN.n10316 VN.n10315 0.001
R13561 VN.n10362 VN.n10361 0.001
R13562 VN.n10734 VN.n10733 0.001
R13563 VN.n11336 VN.n11335 0.001
R13564 VN.n11094 VN.n11093 0.001
R13565 VN.n11500 VN.n11499 0.001
R13566 VN.n10338 VN.n10337 0.001
R13567 VN.n10666 VN.n10665 0.001
R13568 VN.n9751 VN.n9750 0.001
R13569 VN.n9452 VN.n9451 0.001
R13570 VN.n8889 VN.n8888 0.001
R13571 VN.n8593 VN.n8592 0.001
R13572 VN.n8040 VN.n8039 0.001
R13573 VN.n7745 VN.n7744 0.001
R13574 VN.n6849 VN.n6848 0.001
R13575 VN.n6997 VN.n6996 0.001
R13576 VN.n6404 VN.n6403 0.001
R13577 VN.n6113 VN.n6112 0.001
R13578 VN.n5612 VN.n5611 0.001
R13579 VN.n5324 VN.n5323 0.001
R13580 VN.n4833 VN.n4832 0.001
R13581 VN.n4546 VN.n4545 0.001
R13582 VN.n4076 VN.n4075 0.001
R13583 VN.n3792 VN.n3791 0.001
R13584 VN.n3332 VN.n3331 0.001
R13585 VN.n3049 VN.n3048 0.001
R13586 VN.n2610 VN.n2609 0.001
R13587 VN.n2330 VN.n2329 0.001
R13588 VN.n1901 VN.n1900 0.001
R13589 VN.n1622 VN.n1621 0.001
R13590 VN.n1211 VN.n1210 0.001
R13591 VN.n935 VN.n934 0.001
R13592 VN.n536 VN.n535 0.001
R13593 VN.n263 VN.n262 0.001
R13594 VN.n12287 VN.n12286 0.001
R13595 VN.n12304 VN.n12303 0.001
R13596 VN.n12269 VN.n12268 0.001
R13597 VN.n10639 VN.n10638 0.001
R13598 VN.n10690 VN.n10689 0.001
R13599 VN.n12629 VN.n12628 0.001
R13600 VN.n12328 VN.n12327 0.001
R13601 VN.n12342 VN.n12341 0.001
R13602 VN.n287 VN.n286 0.001
R13603 VN.n556 VN.n555 0.001
R13604 VN.n959 VN.n958 0.001
R13605 VN.n1231 VN.n1230 0.001
R13606 VN.n1646 VN.n1645 0.001
R13607 VN.n1921 VN.n1920 0.001
R13608 VN.n2354 VN.n2353 0.001
R13609 VN.n2630 VN.n2629 0.001
R13610 VN.n3073 VN.n3072 0.001
R13611 VN.n3352 VN.n3351 0.001
R13612 VN.n3816 VN.n3815 0.001
R13613 VN.n4096 VN.n4095 0.001
R13614 VN.n4570 VN.n4569 0.001
R13615 VN.n4853 VN.n4852 0.001
R13616 VN.n5348 VN.n5347 0.001
R13617 VN.n5632 VN.n5631 0.001
R13618 VN.n6137 VN.n6136 0.001
R13619 VN.n6424 VN.n6423 0.001
R13620 VN.n6986 VN.n6985 0.001
R13621 VN.n6869 VN.n6868 0.001
R13622 VN.n7769 VN.n7768 0.001
R13623 VN.n8060 VN.n8059 0.001
R13624 VN.n8617 VN.n8616 0.001
R13625 VN.n8909 VN.n8908 0.001
R13626 VN.n9476 VN.n9475 0.001
R13627 VN.n9794 VN.n9793 0.001
R13628 VN.n9768 VN.n9767 0.001
R13629 VN.n9810 VN.n9809 0.001
R13630 VN.n12420 VN.n12419 0.001
R13631 VN.n12646 VN.n12645 0.001
R13632 VN.n12660 VN.n12659 0.001
R13633 VN.n302 VN.n301 0.001
R13634 VN.n572 VN.n571 0.001
R13635 VN.n974 VN.n973 0.001
R13636 VN.n1247 VN.n1246 0.001
R13637 VN.n1661 VN.n1660 0.001
R13638 VN.n1937 VN.n1936 0.001
R13639 VN.n2369 VN.n2368 0.001
R13640 VN.n2646 VN.n2645 0.001
R13641 VN.n3088 VN.n3087 0.001
R13642 VN.n3368 VN.n3367 0.001
R13643 VN.n3831 VN.n3830 0.001
R13644 VN.n4112 VN.n4111 0.001
R13645 VN.n4585 VN.n4584 0.001
R13646 VN.n4869 VN.n4868 0.001
R13647 VN.n5363 VN.n5362 0.001
R13648 VN.n5648 VN.n5647 0.001
R13649 VN.n6152 VN.n6151 0.001
R13650 VN.n6440 VN.n6439 0.001
R13651 VN.n6971 VN.n6970 0.001
R13652 VN.n6885 VN.n6884 0.001
R13653 VN.n7784 VN.n7783 0.001
R13654 VN.n8076 VN.n8075 0.001
R13655 VN.n8632 VN.n8631 0.001
R13656 VN.n8948 VN.n8947 0.001
R13657 VN.n8922 VN.n8921 0.001
R13658 VN.n8964 VN.n8963 0.001
R13659 VN.n12436 VN.n12435 0.001
R13660 VN.n12677 VN.n12676 0.001
R13661 VN.n12771 VN.n12770 0.001
R13662 VN.n317 VN.n316 0.001
R13663 VN.n588 VN.n587 0.001
R13664 VN.n989 VN.n988 0.001
R13665 VN.n1263 VN.n1262 0.001
R13666 VN.n1676 VN.n1675 0.001
R13667 VN.n1953 VN.n1952 0.001
R13668 VN.n2384 VN.n2383 0.001
R13669 VN.n2662 VN.n2661 0.001
R13670 VN.n3103 VN.n3102 0.001
R13671 VN.n3384 VN.n3383 0.001
R13672 VN.n3846 VN.n3845 0.001
R13673 VN.n4128 VN.n4127 0.001
R13674 VN.n4600 VN.n4599 0.001
R13675 VN.n4885 VN.n4884 0.001
R13676 VN.n5378 VN.n5377 0.001
R13677 VN.n5664 VN.n5663 0.001
R13678 VN.n6167 VN.n6166 0.001
R13679 VN.n6456 VN.n6455 0.001
R13680 VN.n6956 VN.n6955 0.001
R13681 VN.n6901 VN.n6900 0.001
R13682 VN.n7799 VN.n7798 0.001
R13683 VN.n8115 VN.n8114 0.001
R13684 VN.n8089 VN.n8088 0.001
R13685 VN.n8131 VN.n8130 0.001
R13686 VN.n12452 VN.n12451 0.001
R13687 VN.n12791 VN.n12790 0.001
R13688 VN.n12805 VN.n12804 0.001
R13689 VN.n332 VN.n331 0.001
R13690 VN.n604 VN.n603 0.001
R13691 VN.n1004 VN.n1003 0.001
R13692 VN.n1279 VN.n1278 0.001
R13693 VN.n1691 VN.n1690 0.001
R13694 VN.n1969 VN.n1968 0.001
R13695 VN.n2399 VN.n2398 0.001
R13696 VN.n2678 VN.n2677 0.001
R13697 VN.n3118 VN.n3117 0.001
R13698 VN.n3400 VN.n3399 0.001
R13699 VN.n3861 VN.n3860 0.001
R13700 VN.n4144 VN.n4143 0.001
R13701 VN.n4615 VN.n4614 0.001
R13702 VN.n4901 VN.n4900 0.001
R13703 VN.n5393 VN.n5392 0.001
R13704 VN.n5680 VN.n5679 0.001
R13705 VN.n6182 VN.n6181 0.001
R13706 VN.n6472 VN.n6471 0.001
R13707 VN.n6626 VN.n6625 0.001
R13708 VN.n6940 VN.n6939 0.001
R13709 VN.n6914 VN.n6913 0.001
R13710 VN.n6611 VN.n6610 0.001
R13711 VN.n12468 VN.n12467 0.001
R13712 VN.n12822 VN.n12821 0.001
R13713 VN.n12836 VN.n12835 0.001
R13714 VN.n347 VN.n346 0.001
R13715 VN.n620 VN.n619 0.001
R13716 VN.n1019 VN.n1018 0.001
R13717 VN.n1295 VN.n1294 0.001
R13718 VN.n1706 VN.n1705 0.001
R13719 VN.n1985 VN.n1984 0.001
R13720 VN.n2414 VN.n2413 0.001
R13721 VN.n2694 VN.n2693 0.001
R13722 VN.n3133 VN.n3132 0.001
R13723 VN.n3416 VN.n3415 0.001
R13724 VN.n3876 VN.n3875 0.001
R13725 VN.n4160 VN.n4159 0.001
R13726 VN.n4630 VN.n4629 0.001
R13727 VN.n4917 VN.n4916 0.001
R13728 VN.n5408 VN.n5407 0.001
R13729 VN.n5696 VN.n5695 0.001
R13730 VN.n6197 VN.n6196 0.001
R13731 VN.n6511 VN.n6510 0.001
R13732 VN.n6485 VN.n6484 0.001
R13733 VN.n6527 VN.n6526 0.001
R13734 VN.n12484 VN.n12483 0.001
R13735 VN.n12850 VN.n12849 0.001
R13736 VN.n12864 VN.n12863 0.001
R13737 VN.n362 VN.n361 0.001
R13738 VN.n636 VN.n635 0.001
R13739 VN.n1034 VN.n1033 0.001
R13740 VN.n1311 VN.n1310 0.001
R13741 VN.n1721 VN.n1720 0.001
R13742 VN.n2001 VN.n2000 0.001
R13743 VN.n2429 VN.n2428 0.001
R13744 VN.n2710 VN.n2709 0.001
R13745 VN.n3148 VN.n3147 0.001
R13746 VN.n3432 VN.n3431 0.001
R13747 VN.n3891 VN.n3890 0.001
R13748 VN.n4176 VN.n4175 0.001
R13749 VN.n4645 VN.n4644 0.001
R13750 VN.n4933 VN.n4932 0.001
R13751 VN.n5423 VN.n5422 0.001
R13752 VN.n5735 VN.n5734 0.001
R13753 VN.n5709 VN.n5708 0.001
R13754 VN.n5751 VN.n5750 0.001
R13755 VN.n12500 VN.n12499 0.001
R13756 VN.n12881 VN.n12880 0.001
R13757 VN.n12895 VN.n12894 0.001
R13758 VN.n377 VN.n376 0.001
R13759 VN.n652 VN.n651 0.001
R13760 VN.n1049 VN.n1048 0.001
R13761 VN.n1327 VN.n1326 0.001
R13762 VN.n1736 VN.n1735 0.001
R13763 VN.n2017 VN.n2016 0.001
R13764 VN.n2444 VN.n2443 0.001
R13765 VN.n2726 VN.n2725 0.001
R13766 VN.n3163 VN.n3162 0.001
R13767 VN.n3448 VN.n3447 0.001
R13768 VN.n3906 VN.n3905 0.001
R13769 VN.n4192 VN.n4191 0.001
R13770 VN.n4660 VN.n4659 0.001
R13771 VN.n4972 VN.n4971 0.001
R13772 VN.n4946 VN.n4945 0.001
R13773 VN.n4988 VN.n4987 0.001
R13774 VN.n12516 VN.n12515 0.001
R13775 VN.n12912 VN.n12911 0.001
R13776 VN.n12926 VN.n12925 0.001
R13777 VN.n392 VN.n391 0.001
R13778 VN.n668 VN.n667 0.001
R13779 VN.n1064 VN.n1063 0.001
R13780 VN.n1343 VN.n1342 0.001
R13781 VN.n1751 VN.n1750 0.001
R13782 VN.n2033 VN.n2032 0.001
R13783 VN.n2459 VN.n2458 0.001
R13784 VN.n2742 VN.n2741 0.001
R13785 VN.n3178 VN.n3177 0.001
R13786 VN.n3464 VN.n3463 0.001
R13787 VN.n3921 VN.n3920 0.001
R13788 VN.n4231 VN.n4230 0.001
R13789 VN.n4205 VN.n4204 0.001
R13790 VN.n4247 VN.n4246 0.001
R13791 VN.n12532 VN.n12531 0.001
R13792 VN.n12943 VN.n12942 0.001
R13793 VN.n12957 VN.n12956 0.001
R13794 VN.n407 VN.n406 0.001
R13795 VN.n684 VN.n683 0.001
R13796 VN.n1079 VN.n1078 0.001
R13797 VN.n1359 VN.n1358 0.001
R13798 VN.n1766 VN.n1765 0.001
R13799 VN.n2049 VN.n2048 0.001
R13800 VN.n2474 VN.n2473 0.001
R13801 VN.n2758 VN.n2757 0.001
R13802 VN.n3193 VN.n3192 0.001
R13803 VN.n3503 VN.n3502 0.001
R13804 VN.n3477 VN.n3476 0.001
R13805 VN.n3519 VN.n3518 0.001
R13806 VN.n12548 VN.n12547 0.001
R13807 VN.n12974 VN.n12973 0.001
R13808 VN.n12988 VN.n12987 0.001
R13809 VN.n422 VN.n421 0.001
R13810 VN.n700 VN.n699 0.001
R13811 VN.n1094 VN.n1093 0.001
R13812 VN.n1375 VN.n1374 0.001
R13813 VN.n1781 VN.n1780 0.001
R13814 VN.n2065 VN.n2064 0.001
R13815 VN.n2489 VN.n2488 0.001
R13816 VN.n2797 VN.n2796 0.001
R13817 VN.n2771 VN.n2770 0.001
R13818 VN.n2813 VN.n2812 0.001
R13819 VN.n12564 VN.n12563 0.001
R13820 VN.n13005 VN.n13004 0.001
R13821 VN.n13019 VN.n13018 0.001
R13822 VN.n437 VN.n436 0.001
R13823 VN.n716 VN.n715 0.001
R13824 VN.n1109 VN.n1108 0.001
R13825 VN.n1391 VN.n1390 0.001
R13826 VN.n1796 VN.n1795 0.001
R13827 VN.n2104 VN.n2103 0.001
R13828 VN.n2078 VN.n2077 0.001
R13829 VN.n2120 VN.n2119 0.001
R13830 VN.n12580 VN.n12579 0.001
R13831 VN.n13036 VN.n13035 0.001
R13832 VN.n13050 VN.n13049 0.001
R13833 VN.n452 VN.n451 0.001
R13834 VN.n732 VN.n731 0.001
R13835 VN.n1124 VN.n1123 0.001
R13836 VN.n1430 VN.n1429 0.001
R13837 VN.n1404 VN.n1403 0.001
R13838 VN.n1446 VN.n1445 0.001
R13839 VN.n12596 VN.n12595 0.001
R13840 VN.n13067 VN.n13066 0.001
R13841 VN.n13081 VN.n13080 0.001
R13842 VN.n467 VN.n466 0.001
R13843 VN.n770 VN.n769 0.001
R13844 VN.n743 VN.n742 0.001
R13845 VN.n788 VN.n787 0.001
R13846 VN.n12609 VN.n12608 0.001
R13847 VN.n13099 VN.n13098 0.001
R13848 VN.n12751 VN.n12750 0.001
R13849 VN.n12380 VN.n12379 0.001
R13850 VN.n12228 VN.n12227 0.001
R13851 VN.n12725 VN.n12724 0.001
R13852 VN.n11853 VN.n11852 0.001
R13853 VN.n11852 VN.n11847 0.001
R13854 VN.n12364 VN.n12363 0.001
R13855 VN.n12694 VN.n12693 0.001
R13856 VN.n487 VN.n486 0.001
R13857 VN.n1139 VN.n1138 0.001
R13858 VN.n1813 VN.n1812 0.001
R13859 VN.n2504 VN.n2503 0.001
R13860 VN.n3210 VN.n3209 0.001
R13861 VN.n3936 VN.n3935 0.001
R13862 VN.n4677 VN.n4676 0.001
R13863 VN.n5438 VN.n5437 0.001
R13864 VN.n6212 VN.n6211 0.001
R13865 VN.n6641 VN.n6640 0.001
R13866 VN.n7816 VN.n7815 0.001
R13867 VN.n8647 VN.n8646 0.001
R13868 VN.n9493 VN.n9492 0.001
R13869 VN.n10348 VN.n10347 0.001
R13870 VN.n11375 VN.n11374 0.001
R13871 VN.t160 VN.n11578 0.001
R13872 VN.n11572 VN.n11571 0.001
R13873 VN.n12408 VN.n12405 0.001
R13874 VN.t82 VN.n12411 0.001
R13875 VN.n13113 VN.t236 0.001
R13876 VN.n13137 VN.n13115 0.001
R13877 VN.t160 VN.n12171 0.001
R13878 VN.t160 VN.n12168 0.001
R13879 VN.n12168 VN.n12165 0.001
R13880 VN.t236 VN.n12262 0.001
R13881 VN.t236 VN.n12265 0.001
R13882 VN.t101 VN.n12719 0.001
R13883 VN.t101 VN.n12716 0.001
R13884 VN.n12716 VN.n12713 0.001
R13885 VN.t12 VN.n233 0.001
R13886 VN.t12 VN.n230 0.001
R13887 VN.n230 VN.n227 0.001
R13888 VN.t41 VN.n530 0.001
R13889 VN.t41 VN.n527 0.001
R13890 VN.n527 VN.n524 0.001
R13891 VN.t24 VN.n904 0.001
R13892 VN.t24 VN.n901 0.001
R13893 VN.n901 VN.n898 0.001
R13894 VN.t94 VN.n1205 0.001
R13895 VN.t94 VN.n1202 0.001
R13896 VN.n1202 VN.n1199 0.001
R13897 VN.t224 VN.n1587 0.001
R13898 VN.t224 VN.n1584 0.001
R13899 VN.n1584 VN.n1581 0.001
R13900 VN.t108 VN.n1895 0.001
R13901 VN.t108 VN.n1892 0.001
R13902 VN.n1892 VN.n1889 0.001
R13903 VN.t49 VN.n2295 0.001
R13904 VN.t49 VN.n2292 0.001
R13905 VN.n2292 VN.n2289 0.001
R13906 VN.t57 VN.n2604 0.001
R13907 VN.t57 VN.n2601 0.001
R13908 VN.n2601 VN.n2598 0.001
R13909 VN.t63 VN.n3017 0.001
R13910 VN.t63 VN.n3014 0.001
R13911 VN.n3014 VN.n3011 0.001
R13912 VN.t183 VN.n3326 0.001
R13913 VN.t183 VN.n3323 0.001
R13914 VN.n3323 VN.n3320 0.001
R13915 VN.t14 VN.n3757 0.001
R13916 VN.t14 VN.n3754 0.001
R13917 VN.n3754 VN.n3751 0.001
R13918 VN.t28 VN.n4070 0.001
R13919 VN.t28 VN.n4067 0.001
R13920 VN.n4067 VN.n4064 0.001
R13921 VN.t99 VN.n4514 0.001
R13922 VN.t99 VN.n4511 0.001
R13923 VN.n4511 VN.n4508 0.001
R13924 VN.t32 VN.n4827 0.001
R13925 VN.t32 VN.n4824 0.001
R13926 VN.n4824 VN.n4821 0.001
R13927 VN.t71 VN.n5289 0.001
R13928 VN.t71 VN.n5286 0.001
R13929 VN.n5286 VN.n5283 0.001
R13930 VN.t176 VN.n5606 0.001
R13931 VN.t176 VN.n5603 0.001
R13932 VN.n5603 VN.n5600 0.001
R13933 VN.t10 VN.n6081 0.001
R13934 VN.t10 VN.n6078 0.001
R13935 VN.n6078 VN.n6075 0.001
R13936 VN.t146 VN.n6398 0.001
R13937 VN.t146 VN.n6395 0.001
R13938 VN.n6395 VN.n6392 0.001
R13939 VN.t76 VN.n7324 0.001
R13940 VN.t76 VN.n7321 0.001
R13941 VN.n7321 VN.n7318 0.001
R13942 VN.t253 VN.n6843 0.001
R13943 VN.t253 VN.n6840 0.001
R13944 VN.n6840 VN.n6837 0.001
R13945 VN.t80 VN.n7713 0.001
R13946 VN.t80 VN.n7710 0.001
R13947 VN.n7710 VN.n7707 0.001
R13948 VN.t73 VN.n8034 0.001
R13949 VN.t73 VN.n8031 0.001
R13950 VN.n8031 VN.n8028 0.001
R13951 VN.t26 VN.n8558 0.001
R13952 VN.t26 VN.n8555 0.001
R13953 VN.n8555 VN.n8552 0.001
R13954 VN.t39 VN.n8883 0.001
R13955 VN.t39 VN.n8880 0.001
R13956 VN.n8880 VN.n8877 0.001
R13957 VN.t125 VN.n9420 0.001
R13958 VN.t125 VN.n9417 0.001
R13959 VN.n9417 VN.n9414 0.001
R13960 VN.t0 VN.n9745 0.001
R13961 VN.t0 VN.n9742 0.001
R13962 VN.n9742 VN.n9739 0.001
R13963 VN.t120 VN.n10303 0.001
R13964 VN.t120 VN.n10300 0.001
R13965 VN.n10300 VN.n10297 0.001
R13966 VN.t241 VN.n10633 0.001
R13967 VN.t241 VN.n10630 0.001
R13968 VN.n10630 VN.n10627 0.001
R13969 VN.t106 VN.n11471 0.001
R13970 VN.t106 VN.n11468 0.001
R13971 VN.n11468 VN.n11465 0.001
R13972 VN.t35 VN.n11121 0.001
R13973 VN.t35 VN.n11124 0.001
R13974 VN.t160 VN.n12042 0.001
R13975 VN.t160 VN.n12039 0.001
R13976 VN.n12039 VN.n12036 0.001
R13977 VN.t63 VN.n3042 0.001
R13978 VN.t63 VN.n3045 0.001
R13979 VN.t183 VN.n3234 0.001
R13980 VN.t183 VN.n3231 0.001
R13981 VN.n3231 VN.n3228 0.001
R13982 VN.t14 VN.n3606 0.001
R13983 VN.t14 VN.n3603 0.001
R13984 VN.n3603 VN.n3600 0.001
R13985 VN.t28 VN.n3978 0.001
R13986 VN.t28 VN.n3975 0.001
R13987 VN.n3975 VN.n3972 0.001
R13988 VN.t99 VN.n4363 0.001
R13989 VN.t99 VN.n4360 0.001
R13990 VN.n4360 VN.n4357 0.001
R13991 VN.t32 VN.n4735 0.001
R13992 VN.t32 VN.n4732 0.001
R13993 VN.n4732 VN.n4729 0.001
R13994 VN.t71 VN.n5138 0.001
R13995 VN.t71 VN.n5135 0.001
R13996 VN.n5135 VN.n5132 0.001
R13997 VN.t176 VN.n5514 0.001
R13998 VN.t176 VN.n5511 0.001
R13999 VN.n5511 VN.n5508 0.001
R14000 VN.t10 VN.n5930 0.001
R14001 VN.t10 VN.n5927 0.001
R14002 VN.n5927 VN.n5924 0.001
R14003 VN.t146 VN.n6306 0.001
R14004 VN.t146 VN.n6303 0.001
R14005 VN.n6303 VN.n6300 0.001
R14006 VN.t76 VN.n7173 0.001
R14007 VN.t76 VN.n7170 0.001
R14008 VN.n7170 VN.n7167 0.001
R14009 VN.t253 VN.n6751 0.001
R14010 VN.t253 VN.n6748 0.001
R14011 VN.n6748 VN.n6745 0.001
R14012 VN.t80 VN.n7562 0.001
R14013 VN.t80 VN.n7559 0.001
R14014 VN.n7559 VN.n7556 0.001
R14015 VN.t73 VN.n7942 0.001
R14016 VN.t73 VN.n7939 0.001
R14017 VN.n7939 VN.n7936 0.001
R14018 VN.t26 VN.n8407 0.001
R14019 VN.t26 VN.n8404 0.001
R14020 VN.n8404 VN.n8401 0.001
R14021 VN.t39 VN.n8791 0.001
R14022 VN.t39 VN.n8788 0.001
R14023 VN.n8788 VN.n8785 0.001
R14024 VN.t125 VN.n9269 0.001
R14025 VN.t125 VN.n9266 0.001
R14026 VN.n9266 VN.n9263 0.001
R14027 VN.t0 VN.n9653 0.001
R14028 VN.t0 VN.n9650 0.001
R14029 VN.n9650 VN.n9647 0.001
R14030 VN.t120 VN.n10151 0.001
R14031 VN.t120 VN.n10148 0.001
R14032 VN.n10148 VN.n10145 0.001
R14033 VN.t241 VN.n10531 0.001
R14034 VN.t241 VN.n10528 0.001
R14035 VN.n10528 VN.n10525 0.001
R14036 VN.t106 VN.n11015 0.001
R14037 VN.t106 VN.n11012 0.001
R14038 VN.n11012 VN.n11009 0.001
R14039 VN.t35 VN.n11191 0.001
R14040 VN.t35 VN.n11194 0.001
R14041 VN.t160 VN.n12065 0.001
R14042 VN.t160 VN.n12062 0.001
R14043 VN.n12062 VN.n12059 0.001
R14044 VN.t49 VN.n2323 0.001
R14045 VN.t49 VN.n2326 0.001
R14046 VN.t57 VN.n2529 0.001
R14047 VN.t57 VN.n2526 0.001
R14048 VN.n2526 VN.n2523 0.001
R14049 VN.t63 VN.n2895 0.001
R14050 VN.t63 VN.n2892 0.001
R14051 VN.n2892 VN.n2889 0.001
R14052 VN.t183 VN.n3251 0.001
R14053 VN.t183 VN.n3248 0.001
R14054 VN.n3248 VN.n3245 0.001
R14055 VN.t14 VN.n3635 0.001
R14056 VN.t14 VN.n3632 0.001
R14057 VN.n3632 VN.n3629 0.001
R14058 VN.t28 VN.n3995 0.001
R14059 VN.t28 VN.n3992 0.001
R14060 VN.n3992 VN.n3989 0.001
R14061 VN.t99 VN.n4392 0.001
R14062 VN.t99 VN.n4389 0.001
R14063 VN.n4389 VN.n4386 0.001
R14064 VN.t32 VN.n4752 0.001
R14065 VN.t32 VN.n4749 0.001
R14066 VN.n4749 VN.n4746 0.001
R14067 VN.t71 VN.n5167 0.001
R14068 VN.t71 VN.n5164 0.001
R14069 VN.n5164 VN.n5161 0.001
R14070 VN.t176 VN.n5531 0.001
R14071 VN.t176 VN.n5528 0.001
R14072 VN.n5528 VN.n5525 0.001
R14073 VN.t10 VN.n5959 0.001
R14074 VN.t10 VN.n5956 0.001
R14075 VN.n5956 VN.n5953 0.001
R14076 VN.t146 VN.n6323 0.001
R14077 VN.t146 VN.n6320 0.001
R14078 VN.n6320 VN.n6317 0.001
R14079 VN.t76 VN.n7202 0.001
R14080 VN.t76 VN.n7199 0.001
R14081 VN.n7199 VN.n7196 0.001
R14082 VN.t253 VN.n6768 0.001
R14083 VN.t253 VN.n6765 0.001
R14084 VN.n6765 VN.n6762 0.001
R14085 VN.t80 VN.n7591 0.001
R14086 VN.t80 VN.n7588 0.001
R14087 VN.n7588 VN.n7585 0.001
R14088 VN.t73 VN.n7959 0.001
R14089 VN.t73 VN.n7956 0.001
R14090 VN.n7956 VN.n7953 0.001
R14091 VN.t26 VN.n8436 0.001
R14092 VN.t26 VN.n8433 0.001
R14093 VN.n8433 VN.n8430 0.001
R14094 VN.t39 VN.n8808 0.001
R14095 VN.t39 VN.n8805 0.001
R14096 VN.n8805 VN.n8802 0.001
R14097 VN.t125 VN.n9298 0.001
R14098 VN.t125 VN.n9295 0.001
R14099 VN.n9295 VN.n9292 0.001
R14100 VN.t0 VN.n9670 0.001
R14101 VN.t0 VN.n9667 0.001
R14102 VN.n9667 VN.n9664 0.001
R14103 VN.t120 VN.n10180 0.001
R14104 VN.t120 VN.n10177 0.001
R14105 VN.n10177 VN.n10174 0.001
R14106 VN.t241 VN.n10551 0.001
R14107 VN.t241 VN.n10548 0.001
R14108 VN.n10548 VN.n10545 0.001
R14109 VN.t241 VN.n10572 0.001
R14110 VN.t241 VN.n10569 0.001
R14111 VN.n10569 VN.n10566 0.001
R14112 VN.t106 VN.n11075 0.001
R14113 VN.t106 VN.n11072 0.001
R14114 VN.n11072 VN.n11069 0.001
R14115 VN.t35 VN.n11157 0.001
R14116 VN.t35 VN.n11160 0.001
R14117 VN.t160 VN.n12087 0.001
R14118 VN.t160 VN.n12084 0.001
R14119 VN.n12084 VN.n12081 0.001
R14120 VN.t120 VN.n10215 0.001
R14121 VN.t120 VN.n10212 0.001
R14122 VN.n10212 VN.n10209 0.001
R14123 VN.t125 VN.n9332 0.001
R14124 VN.t125 VN.n9329 0.001
R14125 VN.n9329 VN.n9326 0.001
R14126 VN.t26 VN.n8470 0.001
R14127 VN.t26 VN.n8467 0.001
R14128 VN.n8467 VN.n8464 0.001
R14129 VN.t80 VN.n7625 0.001
R14130 VN.t80 VN.n7622 0.001
R14131 VN.n7622 VN.n7619 0.001
R14132 VN.t76 VN.n7236 0.001
R14133 VN.t76 VN.n7233 0.001
R14134 VN.n7233 VN.n7230 0.001
R14135 VN.t10 VN.n5993 0.001
R14136 VN.t10 VN.n5990 0.001
R14137 VN.n5990 VN.n5987 0.001
R14138 VN.t71 VN.n5201 0.001
R14139 VN.t71 VN.n5198 0.001
R14140 VN.n5198 VN.n5195 0.001
R14141 VN.t99 VN.n4426 0.001
R14142 VN.t99 VN.n4423 0.001
R14143 VN.n4423 VN.n4420 0.001
R14144 VN.t14 VN.n3669 0.001
R14145 VN.t14 VN.n3666 0.001
R14146 VN.n3666 VN.n3663 0.001
R14147 VN.t63 VN.n2929 0.001
R14148 VN.t63 VN.n2926 0.001
R14149 VN.n2926 VN.n2923 0.001
R14150 VN.t49 VN.n2207 0.001
R14151 VN.t49 VN.n2204 0.001
R14152 VN.n2204 VN.n2201 0.001
R14153 VN.t224 VN.n1615 0.001
R14154 VN.t224 VN.n1618 0.001
R14155 VN.t108 VN.n1837 0.001
R14156 VN.t108 VN.n1834 0.001
R14157 VN.n1834 VN.n1831 0.001
R14158 VN.t57 VN.n2546 0.001
R14159 VN.t57 VN.n2543 0.001
R14160 VN.n2543 VN.n2540 0.001
R14161 VN.t183 VN.n3268 0.001
R14162 VN.t183 VN.n3265 0.001
R14163 VN.n3265 VN.n3262 0.001
R14164 VN.t28 VN.n4012 0.001
R14165 VN.t28 VN.n4009 0.001
R14166 VN.n4009 VN.n4006 0.001
R14167 VN.t32 VN.n4769 0.001
R14168 VN.t32 VN.n4766 0.001
R14169 VN.n4766 VN.n4763 0.001
R14170 VN.t176 VN.n5548 0.001
R14171 VN.t176 VN.n5545 0.001
R14172 VN.n5545 VN.n5542 0.001
R14173 VN.t146 VN.n6340 0.001
R14174 VN.t146 VN.n6337 0.001
R14175 VN.n6337 VN.n6334 0.001
R14176 VN.t253 VN.n6785 0.001
R14177 VN.t253 VN.n6782 0.001
R14178 VN.n6782 VN.n6779 0.001
R14179 VN.t73 VN.n7976 0.001
R14180 VN.t73 VN.n7973 0.001
R14181 VN.n7973 VN.n7970 0.001
R14182 VN.t39 VN.n8825 0.001
R14183 VN.t39 VN.n8822 0.001
R14184 VN.n8822 VN.n8819 0.001
R14185 VN.t0 VN.n9687 0.001
R14186 VN.t0 VN.n9684 0.001
R14187 VN.n9684 VN.n9681 0.001
R14188 VN.t106 VN.n11420 0.001
R14189 VN.t106 VN.n11417 0.001
R14190 VN.n11417 VN.n11414 0.001
R14191 VN.n11385 VN.t35 0.001
R14192 VN.n11397 VN.n11388 0.001
R14193 VN.t160 VN.n12121 0.001
R14194 VN.t160 VN.n12118 0.001
R14195 VN.n12118 VN.n12115 0.001
R14196 VN.t24 VN.n928 0.001
R14197 VN.t24 VN.n931 0.001
R14198 VN.t94 VN.n1169 0.001
R14199 VN.t94 VN.n1166 0.001
R14200 VN.n1166 VN.n1163 0.001
R14201 VN.t224 VN.n1532 0.001
R14202 VN.t224 VN.n1529 0.001
R14203 VN.n1529 VN.n1526 0.001
R14204 VN.t108 VN.n1859 0.001
R14205 VN.t108 VN.n1856 0.001
R14206 VN.n1856 VN.n1853 0.001
R14207 VN.t49 VN.n2240 0.001
R14208 VN.t49 VN.n2237 0.001
R14209 VN.n2237 VN.n2234 0.001
R14210 VN.t57 VN.n2568 0.001
R14211 VN.t57 VN.n2565 0.001
R14212 VN.n2565 VN.n2562 0.001
R14213 VN.t63 VN.n2962 0.001
R14214 VN.t63 VN.n2959 0.001
R14215 VN.n2959 VN.n2956 0.001
R14216 VN.t183 VN.n3290 0.001
R14217 VN.t183 VN.n3287 0.001
R14218 VN.n3287 VN.n3284 0.001
R14219 VN.t14 VN.n3702 0.001
R14220 VN.t14 VN.n3699 0.001
R14221 VN.n3699 VN.n3696 0.001
R14222 VN.t28 VN.n4034 0.001
R14223 VN.t28 VN.n4031 0.001
R14224 VN.n4031 VN.n4028 0.001
R14225 VN.t99 VN.n4459 0.001
R14226 VN.t99 VN.n4456 0.001
R14227 VN.n4456 VN.n4453 0.001
R14228 VN.t32 VN.n4791 0.001
R14229 VN.t32 VN.n4788 0.001
R14230 VN.n4788 VN.n4785 0.001
R14231 VN.t71 VN.n5234 0.001
R14232 VN.t71 VN.n5231 0.001
R14233 VN.n5231 VN.n5228 0.001
R14234 VN.t176 VN.n5570 0.001
R14235 VN.t176 VN.n5567 0.001
R14236 VN.n5567 VN.n5564 0.001
R14237 VN.t10 VN.n6026 0.001
R14238 VN.t10 VN.n6023 0.001
R14239 VN.n6023 VN.n6020 0.001
R14240 VN.t146 VN.n6362 0.001
R14241 VN.t146 VN.n6359 0.001
R14242 VN.n6359 VN.n6356 0.001
R14243 VN.t76 VN.n7269 0.001
R14244 VN.t76 VN.n7266 0.001
R14245 VN.n7266 VN.n7263 0.001
R14246 VN.t253 VN.n6807 0.001
R14247 VN.t253 VN.n6804 0.001
R14248 VN.n6804 VN.n6801 0.001
R14249 VN.t80 VN.n7658 0.001
R14250 VN.t80 VN.n7655 0.001
R14251 VN.n7655 VN.n7652 0.001
R14252 VN.t73 VN.n7998 0.001
R14253 VN.t73 VN.n7995 0.001
R14254 VN.n7995 VN.n7992 0.001
R14255 VN.t26 VN.n8503 0.001
R14256 VN.t26 VN.n8500 0.001
R14257 VN.n8500 VN.n8497 0.001
R14258 VN.t39 VN.n8847 0.001
R14259 VN.t39 VN.n8844 0.001
R14260 VN.n8844 VN.n8841 0.001
R14261 VN.t125 VN.n9365 0.001
R14262 VN.t125 VN.n9362 0.001
R14263 VN.n9362 VN.n9359 0.001
R14264 VN.t0 VN.n9709 0.001
R14265 VN.t0 VN.n9706 0.001
R14266 VN.n9706 VN.n9703 0.001
R14267 VN.t120 VN.n10248 0.001
R14268 VN.t120 VN.n10245 0.001
R14269 VN.n10245 VN.n10242 0.001
R14270 VN.t241 VN.n10594 0.001
R14271 VN.t241 VN.n10591 0.001
R14272 VN.n10591 VN.n10588 0.001
R14273 VN.t106 VN.n11447 0.001
R14274 VN.t106 VN.n11444 0.001
R14275 VN.n11444 VN.n11441 0.001
R14276 VN.t35 VN.n11141 0.001
R14277 VN.t35 VN.n11144 0.001
R14278 VN.t241 VN.n10615 0.001
R14279 VN.t241 VN.n10612 0.001
R14280 VN.n10612 VN.n10609 0.001
R14281 VN.t120 VN.n10269 0.001
R14282 VN.t120 VN.n10266 0.001
R14283 VN.n10266 VN.n10263 0.001
R14284 VN.t0 VN.n9728 0.001
R14285 VN.t0 VN.n9725 0.001
R14286 VN.n9725 VN.n9722 0.001
R14287 VN.t125 VN.n9386 0.001
R14288 VN.t125 VN.n9383 0.001
R14289 VN.n9383 VN.n9380 0.001
R14290 VN.t39 VN.n8866 0.001
R14291 VN.t39 VN.n8863 0.001
R14292 VN.n8863 VN.n8860 0.001
R14293 VN.t26 VN.n8524 0.001
R14294 VN.t26 VN.n8521 0.001
R14295 VN.n8521 VN.n8518 0.001
R14296 VN.t73 VN.n8017 0.001
R14297 VN.t73 VN.n8014 0.001
R14298 VN.n8014 VN.n8011 0.001
R14299 VN.t80 VN.n7679 0.001
R14300 VN.t80 VN.n7676 0.001
R14301 VN.n7676 VN.n7673 0.001
R14302 VN.t253 VN.n6826 0.001
R14303 VN.t253 VN.n6823 0.001
R14304 VN.n6823 VN.n6820 0.001
R14305 VN.t76 VN.n7290 0.001
R14306 VN.t76 VN.n7287 0.001
R14307 VN.n7287 VN.n7284 0.001
R14308 VN.t146 VN.n6381 0.001
R14309 VN.t146 VN.n6378 0.001
R14310 VN.n6378 VN.n6375 0.001
R14311 VN.t10 VN.n6047 0.001
R14312 VN.t10 VN.n6044 0.001
R14313 VN.n6044 VN.n6041 0.001
R14314 VN.t176 VN.n5589 0.001
R14315 VN.t176 VN.n5586 0.001
R14316 VN.n5586 VN.n5583 0.001
R14317 VN.t71 VN.n5255 0.001
R14318 VN.t71 VN.n5252 0.001
R14319 VN.n5252 VN.n5249 0.001
R14320 VN.t32 VN.n4810 0.001
R14321 VN.t32 VN.n4807 0.001
R14322 VN.n4807 VN.n4804 0.001
R14323 VN.t99 VN.n4480 0.001
R14324 VN.t99 VN.n4477 0.001
R14325 VN.n4477 VN.n4474 0.001
R14326 VN.t28 VN.n4053 0.001
R14327 VN.t28 VN.n4050 0.001
R14328 VN.n4050 VN.n4047 0.001
R14329 VN.t14 VN.n3723 0.001
R14330 VN.t14 VN.n3720 0.001
R14331 VN.n3720 VN.n3717 0.001
R14332 VN.t183 VN.n3309 0.001
R14333 VN.t183 VN.n3306 0.001
R14334 VN.n3306 VN.n3303 0.001
R14335 VN.t63 VN.n2983 0.001
R14336 VN.t63 VN.n2980 0.001
R14337 VN.n2980 VN.n2977 0.001
R14338 VN.t57 VN.n2587 0.001
R14339 VN.t57 VN.n2584 0.001
R14340 VN.n2584 VN.n2581 0.001
R14341 VN.t49 VN.n2261 0.001
R14342 VN.t49 VN.n2258 0.001
R14343 VN.n2258 VN.n2255 0.001
R14344 VN.t108 VN.n1878 0.001
R14345 VN.t108 VN.n1875 0.001
R14346 VN.n1875 VN.n1872 0.001
R14347 VN.t224 VN.n1553 0.001
R14348 VN.t224 VN.n1535 0.001
R14349 VN.t94 VN.n1188 0.001
R14350 VN.t94 VN.n1185 0.001
R14351 VN.n1185 VN.n1182 0.001
R14352 VN.t24 VN.n870 0.001
R14353 VN.t24 VN.n867 0.001
R14354 VN.n867 VN.n864 0.001
R14355 VN.t41 VN.n513 0.001
R14356 VN.t41 VN.n510 0.001
R14357 VN.n510 VN.n507 0.001
R14358 VN.t12 VN.n256 0.001
R14359 VN.t12 VN.n259 0.001
R14360 VN.t160 VN.n12150 0.001
R14361 VN.t160 VN.n12147 0.001
R14362 VN.n12147 VN.n12144 0.001
R14363 VN.t106 VN.n11042 0.001
R14364 VN.t106 VN.n11039 0.001
R14365 VN.n11039 VN.n11036 0.001
R14366 VN.t35 VN.n11175 0.001
R14367 VN.t35 VN.n11178 0.001
R14368 VN.t160 VN.n11997 0.001
R14369 VN.t160 VN.n11994 0.001
R14370 VN.n11994 VN.n11991 0.001
R14371 VN.t99 VN.n4539 0.001
R14372 VN.t99 VN.n4542 0.001
R14373 VN.t32 VN.n4701 0.001
R14374 VN.t32 VN.n4698 0.001
R14375 VN.n4698 VN.n4695 0.001
R14376 VN.t71 VN.n5075 0.001
R14377 VN.t71 VN.n5072 0.001
R14378 VN.n5072 VN.n5069 0.001
R14379 VN.t176 VN.n5480 0.001
R14380 VN.t176 VN.n5477 0.001
R14381 VN.n5477 VN.n5474 0.001
R14382 VN.t10 VN.n5867 0.001
R14383 VN.t10 VN.n5864 0.001
R14384 VN.n5864 VN.n5861 0.001
R14385 VN.t146 VN.n6272 0.001
R14386 VN.t146 VN.n6269 0.001
R14387 VN.n6269 VN.n6266 0.001
R14388 VN.t76 VN.n7110 0.001
R14389 VN.t76 VN.n7107 0.001
R14390 VN.n7107 VN.n7104 0.001
R14391 VN.t253 VN.n6717 0.001
R14392 VN.t253 VN.n6714 0.001
R14393 VN.n6714 VN.n6711 0.001
R14394 VN.t80 VN.n7499 0.001
R14395 VN.t80 VN.n7496 0.001
R14396 VN.n7496 VN.n7493 0.001
R14397 VN.t73 VN.n7908 0.001
R14398 VN.t73 VN.n7905 0.001
R14399 VN.n7905 VN.n7902 0.001
R14400 VN.t26 VN.n8344 0.001
R14401 VN.t26 VN.n8341 0.001
R14402 VN.n8341 VN.n8338 0.001
R14403 VN.t39 VN.n8757 0.001
R14404 VN.t39 VN.n8754 0.001
R14405 VN.n8754 VN.n8751 0.001
R14406 VN.t125 VN.n9206 0.001
R14407 VN.t125 VN.n9203 0.001
R14408 VN.n9203 VN.n9200 0.001
R14409 VN.t0 VN.n9619 0.001
R14410 VN.t0 VN.n9616 0.001
R14411 VN.n9616 VN.n9613 0.001
R14412 VN.t120 VN.n10088 0.001
R14413 VN.t120 VN.n10085 0.001
R14414 VN.n10085 VN.n10082 0.001
R14415 VN.t241 VN.n10496 0.001
R14416 VN.t241 VN.n10493 0.001
R14417 VN.n10493 VN.n10490 0.001
R14418 VN.t106 VN.n10957 0.001
R14419 VN.t106 VN.n10954 0.001
R14420 VN.n10954 VN.n10951 0.001
R14421 VN.t35 VN.n11225 0.001
R14422 VN.t35 VN.n11228 0.001
R14423 VN.t160 VN.n12020 0.001
R14424 VN.t160 VN.n12017 0.001
R14425 VN.n12017 VN.n12014 0.001
R14426 VN.t14 VN.n3785 0.001
R14427 VN.t14 VN.n3788 0.001
R14428 VN.t28 VN.n3961 0.001
R14429 VN.t28 VN.n3958 0.001
R14430 VN.n3958 VN.n3955 0.001
R14431 VN.t99 VN.n4329 0.001
R14432 VN.t99 VN.n4326 0.001
R14433 VN.n4326 VN.n4323 0.001
R14434 VN.t32 VN.n4718 0.001
R14435 VN.t32 VN.n4715 0.001
R14436 VN.n4715 VN.n4712 0.001
R14437 VN.t71 VN.n5104 0.001
R14438 VN.t71 VN.n5101 0.001
R14439 VN.n5101 VN.n5098 0.001
R14440 VN.t176 VN.n5497 0.001
R14441 VN.t176 VN.n5494 0.001
R14442 VN.n5494 VN.n5491 0.001
R14443 VN.t10 VN.n5896 0.001
R14444 VN.t10 VN.n5893 0.001
R14445 VN.n5893 VN.n5890 0.001
R14446 VN.t146 VN.n6289 0.001
R14447 VN.t146 VN.n6286 0.001
R14448 VN.n6286 VN.n6283 0.001
R14449 VN.t76 VN.n7139 0.001
R14450 VN.t76 VN.n7136 0.001
R14451 VN.n7136 VN.n7133 0.001
R14452 VN.t253 VN.n6734 0.001
R14453 VN.t253 VN.n6731 0.001
R14454 VN.n6731 VN.n6728 0.001
R14455 VN.t80 VN.n7528 0.001
R14456 VN.t80 VN.n7525 0.001
R14457 VN.n7525 VN.n7522 0.001
R14458 VN.t73 VN.n7925 0.001
R14459 VN.t73 VN.n7922 0.001
R14460 VN.n7922 VN.n7919 0.001
R14461 VN.t26 VN.n8373 0.001
R14462 VN.t26 VN.n8370 0.001
R14463 VN.n8370 VN.n8367 0.001
R14464 VN.t39 VN.n8774 0.001
R14465 VN.t39 VN.n8771 0.001
R14466 VN.n8771 VN.n8768 0.001
R14467 VN.t125 VN.n9235 0.001
R14468 VN.t125 VN.n9232 0.001
R14469 VN.n9232 VN.n9229 0.001
R14470 VN.t0 VN.n9636 0.001
R14471 VN.t0 VN.n9633 0.001
R14472 VN.n9633 VN.n9630 0.001
R14473 VN.t120 VN.n10117 0.001
R14474 VN.t120 VN.n10114 0.001
R14475 VN.n10114 VN.n10111 0.001
R14476 VN.t241 VN.n10513 0.001
R14477 VN.t241 VN.n10510 0.001
R14478 VN.n10510 VN.n10507 0.001
R14479 VN.t106 VN.n10986 0.001
R14480 VN.t106 VN.n10983 0.001
R14481 VN.n10983 VN.n10980 0.001
R14482 VN.t35 VN.n11209 0.001
R14483 VN.t35 VN.n11212 0.001
R14484 VN.t160 VN.n11952 0.001
R14485 VN.t160 VN.n11949 0.001
R14486 VN.n11949 VN.n11946 0.001
R14487 VN.t10 VN.n6106 0.001
R14488 VN.t10 VN.n6109 0.001
R14489 VN.t146 VN.n6238 0.001
R14490 VN.t146 VN.n6235 0.001
R14491 VN.n6235 VN.n6232 0.001
R14492 VN.t76 VN.n7047 0.001
R14493 VN.t76 VN.n7044 0.001
R14494 VN.n7044 VN.n7041 0.001
R14495 VN.t253 VN.n6683 0.001
R14496 VN.t253 VN.n6680 0.001
R14497 VN.n6680 VN.n6677 0.001
R14498 VN.t80 VN.n7436 0.001
R14499 VN.t80 VN.n7433 0.001
R14500 VN.n7433 VN.n7430 0.001
R14501 VN.t73 VN.n7874 0.001
R14502 VN.t73 VN.n7871 0.001
R14503 VN.n7871 VN.n7868 0.001
R14504 VN.t26 VN.n8281 0.001
R14505 VN.t26 VN.n8278 0.001
R14506 VN.n8278 VN.n8275 0.001
R14507 VN.t39 VN.n8723 0.001
R14508 VN.t39 VN.n8720 0.001
R14509 VN.n8720 VN.n8717 0.001
R14510 VN.t125 VN.n9143 0.001
R14511 VN.t125 VN.n9140 0.001
R14512 VN.n9140 VN.n9137 0.001
R14513 VN.t0 VN.n9585 0.001
R14514 VN.t0 VN.n9582 0.001
R14515 VN.n9582 VN.n9579 0.001
R14516 VN.t120 VN.n10025 0.001
R14517 VN.t120 VN.n10022 0.001
R14518 VN.n10022 VN.n10019 0.001
R14519 VN.t241 VN.n10461 0.001
R14520 VN.t241 VN.n10458 0.001
R14521 VN.n10458 VN.n10455 0.001
R14522 VN.t106 VN.n10899 0.001
R14523 VN.t106 VN.n10896 0.001
R14524 VN.n10896 VN.n10893 0.001
R14525 VN.t35 VN.n11259 0.001
R14526 VN.t35 VN.n11262 0.001
R14527 VN.t160 VN.n11975 0.001
R14528 VN.t160 VN.n11972 0.001
R14529 VN.n11972 VN.n11969 0.001
R14530 VN.t71 VN.n5317 0.001
R14531 VN.t71 VN.n5320 0.001
R14532 VN.t176 VN.n5463 0.001
R14533 VN.t176 VN.n5460 0.001
R14534 VN.n5460 VN.n5457 0.001
R14535 VN.t10 VN.n5833 0.001
R14536 VN.t10 VN.n5830 0.001
R14537 VN.n5830 VN.n5827 0.001
R14538 VN.t146 VN.n6255 0.001
R14539 VN.t146 VN.n6252 0.001
R14540 VN.n6252 VN.n6249 0.001
R14541 VN.t76 VN.n7076 0.001
R14542 VN.t76 VN.n7073 0.001
R14543 VN.n7073 VN.n7070 0.001
R14544 VN.t253 VN.n6700 0.001
R14545 VN.t253 VN.n6697 0.001
R14546 VN.n6697 VN.n6694 0.001
R14547 VN.t80 VN.n7465 0.001
R14548 VN.t80 VN.n7462 0.001
R14549 VN.n7462 VN.n7459 0.001
R14550 VN.t73 VN.n7891 0.001
R14551 VN.t73 VN.n7888 0.001
R14552 VN.n7888 VN.n7885 0.001
R14553 VN.t26 VN.n8310 0.001
R14554 VN.t26 VN.n8307 0.001
R14555 VN.n8307 VN.n8304 0.001
R14556 VN.t39 VN.n8740 0.001
R14557 VN.t39 VN.n8737 0.001
R14558 VN.n8737 VN.n8734 0.001
R14559 VN.t125 VN.n9172 0.001
R14560 VN.t125 VN.n9169 0.001
R14561 VN.n9169 VN.n9166 0.001
R14562 VN.t0 VN.n9602 0.001
R14563 VN.t0 VN.n9599 0.001
R14564 VN.n9599 VN.n9596 0.001
R14565 VN.t120 VN.n10054 0.001
R14566 VN.t120 VN.n10051 0.001
R14567 VN.n10051 VN.n10048 0.001
R14568 VN.t241 VN.n10478 0.001
R14569 VN.t241 VN.n10475 0.001
R14570 VN.n10475 VN.n10472 0.001
R14571 VN.t106 VN.n10928 0.001
R14572 VN.t106 VN.n10925 0.001
R14573 VN.n10925 VN.n10922 0.001
R14574 VN.t35 VN.n11243 0.001
R14575 VN.t35 VN.n11246 0.001
R14576 VN.t253 VN.n6666 0.001
R14577 VN.t253 VN.n6663 0.001
R14578 VN.n6663 VN.n6660 0.001
R14579 VN.t80 VN.n7402 0.001
R14580 VN.t80 VN.n7399 0.001
R14581 VN.n7399 VN.n7396 0.001
R14582 VN.t73 VN.n7857 0.001
R14583 VN.t73 VN.n7854 0.001
R14584 VN.n7854 VN.n7851 0.001
R14585 VN.t26 VN.n8247 0.001
R14586 VN.t26 VN.n8244 0.001
R14587 VN.n8244 VN.n8241 0.001
R14588 VN.t39 VN.n8706 0.001
R14589 VN.t39 VN.n8703 0.001
R14590 VN.n8703 VN.n8700 0.001
R14591 VN.t125 VN.n9109 0.001
R14592 VN.t125 VN.n9106 0.001
R14593 VN.n9106 VN.n9103 0.001
R14594 VN.t0 VN.n9568 0.001
R14595 VN.t0 VN.n9565 0.001
R14596 VN.n9565 VN.n9562 0.001
R14597 VN.t120 VN.n9991 0.001
R14598 VN.t120 VN.n9988 0.001
R14599 VN.n9988 VN.n9985 0.001
R14600 VN.t241 VN.n10443 0.001
R14601 VN.t241 VN.n10440 0.001
R14602 VN.n10440 VN.n10437 0.001
R14603 VN.t106 VN.n10870 0.001
R14604 VN.t106 VN.n10867 0.001
R14605 VN.n10867 VN.n10864 0.001
R14606 VN.t35 VN.n11276 0.001
R14607 VN.t35 VN.n11279 0.001
R14608 VN.t160 VN.n11930 0.001
R14609 VN.t160 VN.n11927 0.001
R14610 VN.n11927 VN.n11924 0.001
R14611 VN.t160 VN.n11903 0.001
R14612 VN.t160 VN.n11900 0.001
R14613 VN.n11900 VN.n11897 0.001
R14614 VN.t80 VN.n7738 0.001
R14615 VN.t80 VN.n7741 0.001
R14616 VN.t73 VN.n7840 0.001
R14617 VN.t73 VN.n7837 0.001
R14618 VN.n7837 VN.n7834 0.001
R14619 VN.t26 VN.n8218 0.001
R14620 VN.t26 VN.n8215 0.001
R14621 VN.n8215 VN.n8212 0.001
R14622 VN.t39 VN.n8689 0.001
R14623 VN.t39 VN.n8686 0.001
R14624 VN.n8686 VN.n8683 0.001
R14625 VN.t125 VN.n9080 0.001
R14626 VN.t125 VN.n9077 0.001
R14627 VN.n9077 VN.n9074 0.001
R14628 VN.t0 VN.n9551 0.001
R14629 VN.t0 VN.n9548 0.001
R14630 VN.n9548 VN.n9545 0.001
R14631 VN.t120 VN.n9962 0.001
R14632 VN.t120 VN.n9959 0.001
R14633 VN.n9959 VN.n9956 0.001
R14634 VN.t241 VN.n10426 0.001
R14635 VN.t241 VN.n10423 0.001
R14636 VN.n10423 VN.n10420 0.001
R14637 VN.t106 VN.n10841 0.001
R14638 VN.t106 VN.n10838 0.001
R14639 VN.n10838 VN.n10835 0.001
R14640 VN.t35 VN.n11292 0.001
R14641 VN.t35 VN.n11295 0.001
R14642 VN.t160 VN.n11645 0.001
R14643 VN.t160 VN.n11642 0.001
R14644 VN.n11642 VN.n11639 0.001
R14645 VN.t125 VN.n9445 0.001
R14646 VN.t125 VN.n9448 0.001
R14647 VN.t0 VN.n9517 0.001
R14648 VN.t0 VN.n9514 0.001
R14649 VN.n9514 VN.n9511 0.001
R14650 VN.t120 VN.n9899 0.001
R14651 VN.t120 VN.n9896 0.001
R14652 VN.n9896 VN.n9893 0.001
R14653 VN.t241 VN.n10391 0.001
R14654 VN.t241 VN.n10388 0.001
R14655 VN.n10388 VN.n10385 0.001
R14656 VN.t106 VN.n10783 0.001
R14657 VN.t106 VN.n10780 0.001
R14658 VN.n10780 VN.n10777 0.001
R14659 VN.t35 VN.n11326 0.001
R14660 VN.t35 VN.n11329 0.001
R14661 VN.t160 VN.n11882 0.001
R14662 VN.t160 VN.n11879 0.001
R14663 VN.n11879 VN.n11876 0.001
R14664 VN.t26 VN.n8586 0.001
R14665 VN.t26 VN.n8589 0.001
R14666 VN.t39 VN.n8672 0.001
R14667 VN.t39 VN.n8669 0.001
R14668 VN.n8669 VN.n8666 0.001
R14669 VN.t125 VN.n9046 0.001
R14670 VN.t125 VN.n9043 0.001
R14671 VN.n9043 VN.n9040 0.001
R14672 VN.t0 VN.n9534 0.001
R14673 VN.t0 VN.n9531 0.001
R14674 VN.n9531 VN.n9528 0.001
R14675 VN.t120 VN.n9928 0.001
R14676 VN.t120 VN.n9925 0.001
R14677 VN.n9925 VN.n9922 0.001
R14678 VN.t241 VN.n10408 0.001
R14679 VN.t241 VN.n10405 0.001
R14680 VN.n10405 VN.n10402 0.001
R14681 VN.t106 VN.n10812 0.001
R14682 VN.t106 VN.n10809 0.001
R14683 VN.n10809 VN.n10806 0.001
R14684 VN.t35 VN.n11310 0.001
R14685 VN.t35 VN.n11313 0.001
R14686 VN.t160 VN.n11600 0.001
R14687 VN.t160 VN.n11597 0.001
R14688 VN.n11597 VN.n11594 0.001
R14689 VN.t106 VN.n11492 0.001
R14690 VN.t106 VN.n11495 0.001
R14691 VN.t35 VN.n11360 0.001
R14692 VN.t35 VN.n11363 0.001
R14693 VN.t160 VN.n11623 0.001
R14694 VN.t160 VN.n11620 0.001
R14695 VN.n11620 VN.n11617 0.001
R14696 VN.t120 VN.n10331 0.001
R14697 VN.t120 VN.n10334 0.001
R14698 VN.t241 VN.n10373 0.001
R14699 VN.t241 VN.n10370 0.001
R14700 VN.n10370 VN.n10367 0.001
R14701 VN.t106 VN.n10754 0.001
R14702 VN.t106 VN.n10751 0.001
R14703 VN.n10751 VN.n10748 0.001
R14704 VN.t35 VN.n11344 0.001
R14705 VN.t35 VN.n11347 0.001
R14706 VN.n12174 VN.t160 0.001
R14707 VN.n12182 VN.n12174 0.001
R14708 VN.t35 VN.n11106 0.001
R14709 VN.t35 VN.n11103 0.001
R14710 VN.n11103 VN.n11100 0.001
R14711 VN.t106 VN.n11509 0.001
R14712 VN.t106 VN.n11512 0.001
R14713 VN.n10653 VN.t241 0.001
R14714 VN.n10662 VN.n10656 0.001
R14715 VN.t120 VN.n10679 0.001
R14716 VN.t120 VN.n10682 0.001
R14717 VN.t0 VN.n9760 0.001
R14718 VN.t0 VN.n9763 0.001
R14719 VN.t125 VN.n9465 0.001
R14720 VN.t125 VN.n9468 0.001
R14721 VN.t39 VN.n8898 0.001
R14722 VN.t39 VN.n8901 0.001
R14723 VN.t26 VN.n8606 0.001
R14724 VN.t26 VN.n8609 0.001
R14725 VN.t73 VN.n8049 0.001
R14726 VN.t73 VN.n8052 0.001
R14727 VN.t80 VN.n7758 0.001
R14728 VN.t80 VN.n7761 0.001
R14729 VN.t253 VN.n6858 0.001
R14730 VN.t253 VN.n6861 0.001
R14731 VN.t76 VN.n7013 0.001
R14732 VN.t76 VN.n7010 0.001
R14733 VN.n7010 VN.n7007 0.001
R14734 VN.t146 VN.n6413 0.001
R14735 VN.t146 VN.n6416 0.001
R14736 VN.t10 VN.n6126 0.001
R14737 VN.t10 VN.n6129 0.001
R14738 VN.t176 VN.n5621 0.001
R14739 VN.t176 VN.n5624 0.001
R14740 VN.t71 VN.n5337 0.001
R14741 VN.t71 VN.n5340 0.001
R14742 VN.t32 VN.n4842 0.001
R14743 VN.t32 VN.n4845 0.001
R14744 VN.t99 VN.n4559 0.001
R14745 VN.t99 VN.n4562 0.001
R14746 VN.t28 VN.n4085 0.001
R14747 VN.t28 VN.n4088 0.001
R14748 VN.t14 VN.n3805 0.001
R14749 VN.t14 VN.n3808 0.001
R14750 VN.t183 VN.n3341 0.001
R14751 VN.t183 VN.n3344 0.001
R14752 VN.t63 VN.n3062 0.001
R14753 VN.t63 VN.n3065 0.001
R14754 VN.t57 VN.n2619 0.001
R14755 VN.t57 VN.n2622 0.001
R14756 VN.t49 VN.n2343 0.001
R14757 VN.t49 VN.n2346 0.001
R14758 VN.t108 VN.n1910 0.001
R14759 VN.t108 VN.n1913 0.001
R14760 VN.t224 VN.n1635 0.001
R14761 VN.t224 VN.n1638 0.001
R14762 VN.t94 VN.n1220 0.001
R14763 VN.t94 VN.n1223 0.001
R14764 VN.t24 VN.n948 0.001
R14765 VN.t24 VN.n951 0.001
R14766 VN.t41 VN.n545 0.001
R14767 VN.t41 VN.n548 0.001
R14768 VN.t12 VN.n276 0.001
R14769 VN.t12 VN.n279 0.001
R14770 VN.n12299 VN.n12293 0.001
R14771 VN.t236 VN.n12317 0.001
R14772 VN.t236 VN.n12320 0.001
R14773 VN.n12282 VN.n12275 0.001
R14774 VN.n12281 VN.n12280 0.001
R14775 VN.n12313 VN.n12312 0.001
R14776 VN.n12298 VN.n12297 0.001
R14777 VN.n272 VN.n271 0.001
R14778 VN.n541 VN.n540 0.001
R14779 VN.n944 VN.n943 0.001
R14780 VN.n1216 VN.n1215 0.001
R14781 VN.n1631 VN.n1630 0.001
R14782 VN.n1906 VN.n1905 0.001
R14783 VN.n2339 VN.n2338 0.001
R14784 VN.n2615 VN.n2614 0.001
R14785 VN.n3058 VN.n3057 0.001
R14786 VN.n3337 VN.n3336 0.001
R14787 VN.n3801 VN.n3800 0.001
R14788 VN.n4081 VN.n4080 0.001
R14789 VN.n4555 VN.n4554 0.001
R14790 VN.n4838 VN.n4837 0.001
R14791 VN.n5333 VN.n5332 0.001
R14792 VN.n5617 VN.n5616 0.001
R14793 VN.n6122 VN.n6121 0.001
R14794 VN.n6409 VN.n6408 0.001
R14795 VN.n7006 VN.n7005 0.001
R14796 VN.n6854 VN.n6853 0.001
R14797 VN.n7754 VN.n7753 0.001
R14798 VN.n8045 VN.n8044 0.001
R14799 VN.n8602 VN.n8601 0.001
R14800 VN.n8894 VN.n8893 0.001
R14801 VN.n9461 VN.n9460 0.001
R14802 VN.n9756 VN.n9755 0.001
R14803 VN.n10675 VN.n10674 0.001
R14804 VN.n10661 VN.n10660 0.001
R14805 VN.n11515 VN.t106 0.001
R14806 VN.n11524 VN.n11517 0.001
R14807 VN.t241 VN.n10647 0.001
R14808 VN.t241 VN.n10650 0.001
R14809 VN.t120 VN.n10694 0.001
R14810 VN.t120 VN.n10697 0.001
R14811 VN.n12623 VN.t82 0.001
R14812 VN.n12630 VN.n12623 0.001
R14813 VN.t236 VN.n12635 0.001
R14814 VN.t236 VN.n12638 0.001
R14815 VN.n12343 VN.n12336 0.001
R14816 VN.t12 VN.n291 0.001
R14817 VN.t12 VN.n294 0.001
R14818 VN.t41 VN.n561 0.001
R14819 VN.t41 VN.n564 0.001
R14820 VN.t24 VN.n963 0.001
R14821 VN.t24 VN.n966 0.001
R14822 VN.t94 VN.n1236 0.001
R14823 VN.t94 VN.n1239 0.001
R14824 VN.t224 VN.n1650 0.001
R14825 VN.t224 VN.n1653 0.001
R14826 VN.t108 VN.n1926 0.001
R14827 VN.t108 VN.n1929 0.001
R14828 VN.t49 VN.n2358 0.001
R14829 VN.t49 VN.n2361 0.001
R14830 VN.t57 VN.n2635 0.001
R14831 VN.t57 VN.n2638 0.001
R14832 VN.t63 VN.n3077 0.001
R14833 VN.t63 VN.n3080 0.001
R14834 VN.t183 VN.n3357 0.001
R14835 VN.t183 VN.n3360 0.001
R14836 VN.t14 VN.n3820 0.001
R14837 VN.t14 VN.n3823 0.001
R14838 VN.t28 VN.n4101 0.001
R14839 VN.t28 VN.n4104 0.001
R14840 VN.t99 VN.n4574 0.001
R14841 VN.t99 VN.n4577 0.001
R14842 VN.t32 VN.n4858 0.001
R14843 VN.t32 VN.n4861 0.001
R14844 VN.t71 VN.n5352 0.001
R14845 VN.t71 VN.n5355 0.001
R14846 VN.t176 VN.n5637 0.001
R14847 VN.t176 VN.n5640 0.001
R14848 VN.t10 VN.n6141 0.001
R14849 VN.t10 VN.n6144 0.001
R14850 VN.t146 VN.n6429 0.001
R14851 VN.t146 VN.n6432 0.001
R14852 VN.t76 VN.n6993 0.001
R14853 VN.t76 VN.n6990 0.001
R14854 VN.n6990 VN.n6987 0.001
R14855 VN.t253 VN.n6874 0.001
R14856 VN.t253 VN.n6877 0.001
R14857 VN.t80 VN.n7773 0.001
R14858 VN.t80 VN.n7776 0.001
R14859 VN.t73 VN.n8065 0.001
R14860 VN.t73 VN.n8068 0.001
R14861 VN.t26 VN.n8621 0.001
R14862 VN.t26 VN.n8624 0.001
R14863 VN.t39 VN.n8914 0.001
R14864 VN.t39 VN.n8917 0.001
R14865 VN.t125 VN.n9799 0.001
R14866 VN.t125 VN.n9802 0.001
R14867 VN.n9788 VN.t0 0.001
R14868 VN.n9795 VN.n9788 0.001
R14869 VN.n10699 VN.t120 0.001
R14870 VN.n10707 VN.n10699 0.001
R14871 VN.t0 VN.n9782 0.001
R14872 VN.t0 VN.n9785 0.001
R14873 VN.t125 VN.n9814 0.001
R14874 VN.t125 VN.n9817 0.001
R14875 VN.t82 VN.n12425 0.001
R14876 VN.t82 VN.n12428 0.001
R14877 VN.t236 VN.n12666 0.001
R14878 VN.t236 VN.n12669 0.001
R14879 VN.n12661 VN.n12654 0.001
R14880 VN.t12 VN.n306 0.001
R14881 VN.t12 VN.n309 0.001
R14882 VN.t41 VN.n577 0.001
R14883 VN.t41 VN.n580 0.001
R14884 VN.t24 VN.n978 0.001
R14885 VN.t24 VN.n981 0.001
R14886 VN.t94 VN.n1252 0.001
R14887 VN.t94 VN.n1255 0.001
R14888 VN.t224 VN.n1665 0.001
R14889 VN.t224 VN.n1668 0.001
R14890 VN.t108 VN.n1942 0.001
R14891 VN.t108 VN.n1945 0.001
R14892 VN.t49 VN.n2373 0.001
R14893 VN.t49 VN.n2376 0.001
R14894 VN.t57 VN.n2651 0.001
R14895 VN.t57 VN.n2654 0.001
R14896 VN.t63 VN.n3092 0.001
R14897 VN.t63 VN.n3095 0.001
R14898 VN.t183 VN.n3373 0.001
R14899 VN.t183 VN.n3376 0.001
R14900 VN.t14 VN.n3835 0.001
R14901 VN.t14 VN.n3838 0.001
R14902 VN.t28 VN.n4117 0.001
R14903 VN.t28 VN.n4120 0.001
R14904 VN.t99 VN.n4589 0.001
R14905 VN.t99 VN.n4592 0.001
R14906 VN.t32 VN.n4874 0.001
R14907 VN.t32 VN.n4877 0.001
R14908 VN.t71 VN.n5367 0.001
R14909 VN.t71 VN.n5370 0.001
R14910 VN.t176 VN.n5653 0.001
R14911 VN.t176 VN.n5656 0.001
R14912 VN.t10 VN.n6156 0.001
R14913 VN.t10 VN.n6159 0.001
R14914 VN.t146 VN.n6445 0.001
R14915 VN.t146 VN.n6448 0.001
R14916 VN.t76 VN.n6978 0.001
R14917 VN.t76 VN.n6975 0.001
R14918 VN.n6975 VN.n6972 0.001
R14919 VN.t253 VN.n6890 0.001
R14920 VN.t253 VN.n6893 0.001
R14921 VN.t80 VN.n7788 0.001
R14922 VN.t80 VN.n7791 0.001
R14923 VN.t73 VN.n8081 0.001
R14924 VN.t73 VN.n8084 0.001
R14925 VN.t26 VN.n8953 0.001
R14926 VN.t26 VN.n8956 0.001
R14927 VN.n8942 VN.t39 0.001
R14928 VN.n8949 VN.n8942 0.001
R14929 VN.n9819 VN.t125 0.001
R14930 VN.n9827 VN.n9819 0.001
R14931 VN.t39 VN.n8936 0.001
R14932 VN.t39 VN.n8939 0.001
R14933 VN.t26 VN.n8968 0.001
R14934 VN.t26 VN.n8971 0.001
R14935 VN.t82 VN.n12441 0.001
R14936 VN.t82 VN.n12444 0.001
R14937 VN.t236 VN.n12777 0.001
R14938 VN.t236 VN.n12780 0.001
R14939 VN.n12765 VN.t101 0.001
R14940 VN.n12772 VN.n12765 0.001
R14941 VN.t12 VN.n321 0.001
R14942 VN.t12 VN.n324 0.001
R14943 VN.t41 VN.n593 0.001
R14944 VN.t41 VN.n596 0.001
R14945 VN.t24 VN.n993 0.001
R14946 VN.t24 VN.n996 0.001
R14947 VN.t94 VN.n1268 0.001
R14948 VN.t94 VN.n1271 0.001
R14949 VN.t224 VN.n1680 0.001
R14950 VN.t224 VN.n1683 0.001
R14951 VN.t108 VN.n1958 0.001
R14952 VN.t108 VN.n1961 0.001
R14953 VN.t49 VN.n2388 0.001
R14954 VN.t49 VN.n2391 0.001
R14955 VN.t57 VN.n2667 0.001
R14956 VN.t57 VN.n2670 0.001
R14957 VN.t63 VN.n3107 0.001
R14958 VN.t63 VN.n3110 0.001
R14959 VN.t183 VN.n3389 0.001
R14960 VN.t183 VN.n3392 0.001
R14961 VN.t14 VN.n3850 0.001
R14962 VN.t14 VN.n3853 0.001
R14963 VN.t28 VN.n4133 0.001
R14964 VN.t28 VN.n4136 0.001
R14965 VN.t99 VN.n4604 0.001
R14966 VN.t99 VN.n4607 0.001
R14967 VN.t32 VN.n4890 0.001
R14968 VN.t32 VN.n4893 0.001
R14969 VN.t71 VN.n5382 0.001
R14970 VN.t71 VN.n5385 0.001
R14971 VN.t176 VN.n5669 0.001
R14972 VN.t176 VN.n5672 0.001
R14973 VN.t10 VN.n6171 0.001
R14974 VN.t10 VN.n6174 0.001
R14975 VN.t146 VN.n6461 0.001
R14976 VN.t146 VN.n6464 0.001
R14977 VN.t76 VN.n6963 0.001
R14978 VN.t76 VN.n6960 0.001
R14979 VN.n6960 VN.n6957 0.001
R14980 VN.t253 VN.n6906 0.001
R14981 VN.t253 VN.n6909 0.001
R14982 VN.t80 VN.n8120 0.001
R14983 VN.t80 VN.n8123 0.001
R14984 VN.n8109 VN.t73 0.001
R14985 VN.n8116 VN.n8109 0.001
R14986 VN.n8973 VN.t26 0.001
R14987 VN.n8981 VN.n8973 0.001
R14988 VN.t73 VN.n8103 0.001
R14989 VN.t73 VN.n8106 0.001
R14990 VN.t80 VN.n8135 0.001
R14991 VN.t80 VN.n8138 0.001
R14992 VN.t82 VN.n12457 0.001
R14993 VN.t82 VN.n12460 0.001
R14994 VN.t236 VN.n12811 0.001
R14995 VN.n12808 VN.n12788 0.001
R14996 VN.n12806 VN.n12799 0.001
R14997 VN.t12 VN.n336 0.001
R14998 VN.t12 VN.n339 0.001
R14999 VN.t41 VN.n609 0.001
R15000 VN.t41 VN.n612 0.001
R15001 VN.t24 VN.n1008 0.001
R15002 VN.t24 VN.n1011 0.001
R15003 VN.t94 VN.n1284 0.001
R15004 VN.t94 VN.n1287 0.001
R15005 VN.t224 VN.n1695 0.001
R15006 VN.t224 VN.n1698 0.001
R15007 VN.t108 VN.n1974 0.001
R15008 VN.t108 VN.n1977 0.001
R15009 VN.t49 VN.n2403 0.001
R15010 VN.t49 VN.n2406 0.001
R15011 VN.t57 VN.n2683 0.001
R15012 VN.t57 VN.n2686 0.001
R15013 VN.t63 VN.n3122 0.001
R15014 VN.t63 VN.n3125 0.001
R15015 VN.t183 VN.n3405 0.001
R15016 VN.t183 VN.n3408 0.001
R15017 VN.t14 VN.n3865 0.001
R15018 VN.t14 VN.n3868 0.001
R15019 VN.t28 VN.n4149 0.001
R15020 VN.t28 VN.n4152 0.001
R15021 VN.t99 VN.n4619 0.001
R15022 VN.t99 VN.n4622 0.001
R15023 VN.t32 VN.n4906 0.001
R15024 VN.t32 VN.n4909 0.001
R15025 VN.t71 VN.n5397 0.001
R15026 VN.t71 VN.n5400 0.001
R15027 VN.t176 VN.n5685 0.001
R15028 VN.t176 VN.n5688 0.001
R15029 VN.t10 VN.n6186 0.001
R15030 VN.t10 VN.n6189 0.001
R15031 VN.t146 VN.n6477 0.001
R15032 VN.t146 VN.n6480 0.001
R15033 VN.t76 VN.n6948 0.001
R15034 VN.t76 VN.n6945 0.001
R15035 VN.n6945 VN.n6942 0.001
R15036 VN.n6934 VN.t253 0.001
R15037 VN.n6941 VN.n6934 0.001
R15038 VN.n8140 VN.t80 0.001
R15039 VN.n8148 VN.n8140 0.001
R15040 VN.t253 VN.n6928 0.001
R15041 VN.t253 VN.n6931 0.001
R15042 VN.t76 VN.n6618 0.001
R15043 VN.t76 VN.n6615 0.001
R15044 VN.n6615 VN.n6612 0.001
R15045 VN.t82 VN.n12473 0.001
R15046 VN.t82 VN.n12476 0.001
R15047 VN.t236 VN.n12842 0.001
R15048 VN.n12839 VN.n12819 0.001
R15049 VN.n12837 VN.n12830 0.001
R15050 VN.t12 VN.n351 0.001
R15051 VN.t12 VN.n354 0.001
R15052 VN.t41 VN.n625 0.001
R15053 VN.t41 VN.n628 0.001
R15054 VN.t24 VN.n1023 0.001
R15055 VN.t24 VN.n1026 0.001
R15056 VN.t94 VN.n1300 0.001
R15057 VN.t94 VN.n1303 0.001
R15058 VN.t224 VN.n1710 0.001
R15059 VN.t224 VN.n1713 0.001
R15060 VN.t108 VN.n1990 0.001
R15061 VN.t108 VN.n1993 0.001
R15062 VN.t49 VN.n2418 0.001
R15063 VN.t49 VN.n2421 0.001
R15064 VN.t57 VN.n2699 0.001
R15065 VN.t57 VN.n2702 0.001
R15066 VN.t63 VN.n3137 0.001
R15067 VN.t63 VN.n3140 0.001
R15068 VN.t183 VN.n3421 0.001
R15069 VN.t183 VN.n3424 0.001
R15070 VN.t14 VN.n3880 0.001
R15071 VN.t14 VN.n3883 0.001
R15072 VN.t28 VN.n4165 0.001
R15073 VN.t28 VN.n4168 0.001
R15074 VN.t99 VN.n4634 0.001
R15075 VN.t99 VN.n4637 0.001
R15076 VN.t32 VN.n4922 0.001
R15077 VN.t32 VN.n4925 0.001
R15078 VN.t71 VN.n5412 0.001
R15079 VN.t71 VN.n5415 0.001
R15080 VN.t176 VN.n5701 0.001
R15081 VN.t176 VN.n5704 0.001
R15082 VN.t10 VN.n6516 0.001
R15083 VN.t10 VN.n6519 0.001
R15084 VN.n6505 VN.t146 0.001
R15085 VN.n6512 VN.n6505 0.001
R15086 VN.n7329 VN.t76 0.001
R15087 VN.n7337 VN.n7329 0.001
R15088 VN.t146 VN.n6499 0.001
R15089 VN.t146 VN.n6502 0.001
R15090 VN.t10 VN.n6531 0.001
R15091 VN.t10 VN.n6534 0.001
R15092 VN.t82 VN.n12489 0.001
R15093 VN.t82 VN.n12492 0.001
R15094 VN.t236 VN.n12870 0.001
R15095 VN.t236 VN.n12873 0.001
R15096 VN.n12865 VN.n12858 0.001
R15097 VN.t12 VN.n366 0.001
R15098 VN.t12 VN.n369 0.001
R15099 VN.t41 VN.n641 0.001
R15100 VN.t41 VN.n644 0.001
R15101 VN.t24 VN.n1038 0.001
R15102 VN.t24 VN.n1041 0.001
R15103 VN.t94 VN.n1316 0.001
R15104 VN.t94 VN.n1319 0.001
R15105 VN.t224 VN.n1725 0.001
R15106 VN.t224 VN.n1728 0.001
R15107 VN.t108 VN.n2006 0.001
R15108 VN.t108 VN.n2009 0.001
R15109 VN.t49 VN.n2433 0.001
R15110 VN.t49 VN.n2436 0.001
R15111 VN.t57 VN.n2715 0.001
R15112 VN.t57 VN.n2718 0.001
R15113 VN.t63 VN.n3152 0.001
R15114 VN.t63 VN.n3155 0.001
R15115 VN.t183 VN.n3437 0.001
R15116 VN.t183 VN.n3440 0.001
R15117 VN.t14 VN.n3895 0.001
R15118 VN.t14 VN.n3898 0.001
R15119 VN.t28 VN.n4181 0.001
R15120 VN.t28 VN.n4184 0.001
R15121 VN.t99 VN.n4649 0.001
R15122 VN.t99 VN.n4652 0.001
R15123 VN.t32 VN.n4938 0.001
R15124 VN.t32 VN.n4941 0.001
R15125 VN.t71 VN.n5740 0.001
R15126 VN.t71 VN.n5743 0.001
R15127 VN.n5729 VN.t176 0.001
R15128 VN.n5736 VN.n5729 0.001
R15129 VN.n6536 VN.t10 0.001
R15130 VN.n6544 VN.n6536 0.001
R15131 VN.t176 VN.n5723 0.001
R15132 VN.t176 VN.n5726 0.001
R15133 VN.t71 VN.n5755 0.001
R15134 VN.t71 VN.n5758 0.001
R15135 VN.t82 VN.n12505 0.001
R15136 VN.t82 VN.n12508 0.001
R15137 VN.t236 VN.n12901 0.001
R15138 VN.t236 VN.n12904 0.001
R15139 VN.n12896 VN.n12889 0.001
R15140 VN.t12 VN.n381 0.001
R15141 VN.t12 VN.n384 0.001
R15142 VN.t41 VN.n657 0.001
R15143 VN.t41 VN.n660 0.001
R15144 VN.t24 VN.n1053 0.001
R15145 VN.t24 VN.n1056 0.001
R15146 VN.t94 VN.n1332 0.001
R15147 VN.t94 VN.n1335 0.001
R15148 VN.t224 VN.n1740 0.001
R15149 VN.t224 VN.n1743 0.001
R15150 VN.t108 VN.n2022 0.001
R15151 VN.t108 VN.n2025 0.001
R15152 VN.t49 VN.n2448 0.001
R15153 VN.t49 VN.n2451 0.001
R15154 VN.t57 VN.n2731 0.001
R15155 VN.t57 VN.n2734 0.001
R15156 VN.t63 VN.n3167 0.001
R15157 VN.t63 VN.n3170 0.001
R15158 VN.t183 VN.n3453 0.001
R15159 VN.t183 VN.n3456 0.001
R15160 VN.t14 VN.n3910 0.001
R15161 VN.t14 VN.n3913 0.001
R15162 VN.t28 VN.n4197 0.001
R15163 VN.t28 VN.n4200 0.001
R15164 VN.t99 VN.n4977 0.001
R15165 VN.t99 VN.n4980 0.001
R15166 VN.n4966 VN.t32 0.001
R15167 VN.n4973 VN.n4966 0.001
R15168 VN.n5760 VN.t71 0.001
R15169 VN.n5768 VN.n5760 0.001
R15170 VN.t32 VN.n4960 0.001
R15171 VN.t32 VN.n4963 0.001
R15172 VN.t99 VN.n4992 0.001
R15173 VN.t99 VN.n4995 0.001
R15174 VN.t82 VN.n12521 0.001
R15175 VN.t82 VN.n12524 0.001
R15176 VN.t236 VN.n12932 0.001
R15177 VN.t236 VN.n12935 0.001
R15178 VN.n12927 VN.n12920 0.001
R15179 VN.t12 VN.n396 0.001
R15180 VN.t12 VN.n399 0.001
R15181 VN.t41 VN.n673 0.001
R15182 VN.t41 VN.n676 0.001
R15183 VN.t24 VN.n1068 0.001
R15184 VN.t24 VN.n1071 0.001
R15185 VN.t94 VN.n1348 0.001
R15186 VN.t94 VN.n1351 0.001
R15187 VN.t224 VN.n1755 0.001
R15188 VN.t224 VN.n1758 0.001
R15189 VN.t108 VN.n2038 0.001
R15190 VN.t108 VN.n2041 0.001
R15191 VN.t49 VN.n2463 0.001
R15192 VN.t49 VN.n2466 0.001
R15193 VN.t57 VN.n2747 0.001
R15194 VN.t57 VN.n2750 0.001
R15195 VN.t63 VN.n3182 0.001
R15196 VN.t63 VN.n3185 0.001
R15197 VN.t183 VN.n3469 0.001
R15198 VN.t183 VN.n3472 0.001
R15199 VN.t14 VN.n4236 0.001
R15200 VN.t14 VN.n4239 0.001
R15201 VN.n4225 VN.t28 0.001
R15202 VN.n4232 VN.n4225 0.001
R15203 VN.n4997 VN.t99 0.001
R15204 VN.n5005 VN.n4997 0.001
R15205 VN.t28 VN.n4219 0.001
R15206 VN.t28 VN.n4222 0.001
R15207 VN.t14 VN.n4251 0.001
R15208 VN.t14 VN.n4254 0.001
R15209 VN.t82 VN.n12537 0.001
R15210 VN.t82 VN.n12540 0.001
R15211 VN.t236 VN.n12963 0.001
R15212 VN.t236 VN.n12966 0.001
R15213 VN.n12958 VN.n12951 0.001
R15214 VN.t12 VN.n411 0.001
R15215 VN.t12 VN.n414 0.001
R15216 VN.t41 VN.n689 0.001
R15217 VN.t41 VN.n692 0.001
R15218 VN.t24 VN.n1083 0.001
R15219 VN.t24 VN.n1086 0.001
R15220 VN.t94 VN.n1364 0.001
R15221 VN.t94 VN.n1367 0.001
R15222 VN.t224 VN.n1770 0.001
R15223 VN.t224 VN.n1773 0.001
R15224 VN.t108 VN.n2054 0.001
R15225 VN.t108 VN.n2057 0.001
R15226 VN.t49 VN.n2478 0.001
R15227 VN.t49 VN.n2481 0.001
R15228 VN.t57 VN.n2763 0.001
R15229 VN.t57 VN.n2766 0.001
R15230 VN.t63 VN.n3508 0.001
R15231 VN.t63 VN.n3511 0.001
R15232 VN.n3497 VN.t183 0.001
R15233 VN.n3504 VN.n3497 0.001
R15234 VN.n4256 VN.t14 0.001
R15235 VN.n4264 VN.n4256 0.001
R15236 VN.t183 VN.n3491 0.001
R15237 VN.t183 VN.n3494 0.001
R15238 VN.t63 VN.n3523 0.001
R15239 VN.t63 VN.n3526 0.001
R15240 VN.t82 VN.n12553 0.001
R15241 VN.t82 VN.n12556 0.001
R15242 VN.t236 VN.n12994 0.001
R15243 VN.t236 VN.n12997 0.001
R15244 VN.n12989 VN.n12982 0.001
R15245 VN.t12 VN.n426 0.001
R15246 VN.t12 VN.n429 0.001
R15247 VN.t41 VN.n705 0.001
R15248 VN.t41 VN.n708 0.001
R15249 VN.t24 VN.n1098 0.001
R15250 VN.t24 VN.n1101 0.001
R15251 VN.t94 VN.n1380 0.001
R15252 VN.t94 VN.n1383 0.001
R15253 VN.t224 VN.n1785 0.001
R15254 VN.t224 VN.n1788 0.001
R15255 VN.t108 VN.n2070 0.001
R15256 VN.t108 VN.n2073 0.001
R15257 VN.t49 VN.n2802 0.001
R15258 VN.t49 VN.n2805 0.001
R15259 VN.n2791 VN.t57 0.001
R15260 VN.n2798 VN.n2791 0.001
R15261 VN.n3528 VN.t63 0.001
R15262 VN.n3536 VN.n3528 0.001
R15263 VN.t57 VN.n2785 0.001
R15264 VN.t57 VN.n2788 0.001
R15265 VN.t49 VN.n2817 0.001
R15266 VN.t49 VN.n2820 0.001
R15267 VN.t82 VN.n12569 0.001
R15268 VN.t82 VN.n12572 0.001
R15269 VN.t236 VN.n13025 0.001
R15270 VN.t236 VN.n13028 0.001
R15271 VN.n13020 VN.n13013 0.001
R15272 VN.t12 VN.n441 0.001
R15273 VN.t12 VN.n444 0.001
R15274 VN.t41 VN.n721 0.001
R15275 VN.t41 VN.n724 0.001
R15276 VN.t24 VN.n1113 0.001
R15277 VN.t24 VN.n1116 0.001
R15278 VN.t94 VN.n1396 0.001
R15279 VN.t94 VN.n1399 0.001
R15280 VN.t224 VN.n2109 0.001
R15281 VN.t224 VN.n2112 0.001
R15282 VN.n2098 VN.t108 0.001
R15283 VN.n2105 VN.n2098 0.001
R15284 VN.n2822 VN.t49 0.001
R15285 VN.n2830 VN.n2822 0.001
R15286 VN.t108 VN.n2092 0.001
R15287 VN.t108 VN.n2095 0.001
R15288 VN.t224 VN.n2124 0.001
R15289 VN.t224 VN.n2127 0.001
R15290 VN.t82 VN.n12585 0.001
R15291 VN.t82 VN.n12588 0.001
R15292 VN.t236 VN.n13056 0.001
R15293 VN.t236 VN.n13059 0.001
R15294 VN.n13051 VN.n13044 0.001
R15295 VN.t12 VN.n456 0.001
R15296 VN.t12 VN.n459 0.001
R15297 VN.t41 VN.n737 0.001
R15298 VN.t41 VN.n740 0.001
R15299 VN.t24 VN.n1435 0.001
R15300 VN.t24 VN.n1438 0.001
R15301 VN.n1424 VN.t94 0.001
R15302 VN.n1431 VN.n1424 0.001
R15303 VN.n2129 VN.t224 0.001
R15304 VN.n2137 VN.n2129 0.001
R15305 VN.t94 VN.n1418 0.001
R15306 VN.t94 VN.n1421 0.001
R15307 VN.t24 VN.n1450 0.001
R15308 VN.t24 VN.n1453 0.001
R15309 VN.t82 VN.n12601 0.001
R15310 VN.t82 VN.n12604 0.001
R15311 VN.t236 VN.n13087 0.001
R15312 VN.t236 VN.n13090 0.001
R15313 VN.n13082 VN.n13075 0.001
R15314 VN.t12 VN.n775 0.001
R15315 VN.t12 VN.n778 0.001
R15316 VN.n764 VN.t41 0.001
R15317 VN.n771 VN.n764 0.001
R15318 VN.n1455 VN.t24 0.001
R15319 VN.n1463 VN.n1455 0.001
R15320 VN.t41 VN.n758 0.001
R15321 VN.t41 VN.n761 0.001
R15322 VN.t12 VN.n797 0.001
R15323 VN.t12 VN.n800 0.001
R15324 VN.t82 VN.n12617 0.001
R15325 VN.t82 VN.n12620 0.001
R15326 VN.t236 VN.n13107 0.001
R15327 VN.t236 VN.n13110 0.001
R15328 VN.t101 VN.n12759 0.001
R15329 VN.t101 VN.n12762 0.001
R15330 VN.n802 VN.t12 0.001
R15331 VN.n821 VN.n802 0.001
R15332 VN.t82 VN.n12391 0.001
R15333 VN.t82 VN.n12388 0.001
R15334 VN.n12388 VN.n12385 0.001
R15335 VN.t236 VN.n12236 0.001
R15336 VN.t236 VN.n12219 0.001
R15337 VN.t101 VN.n12743 0.001
R15338 VN.t101 VN.n12740 0.001
R15339 VN.n12740 VN.n12737 0.001
R15340 VN.t82 VN.n12408 0.001
R15341 VN.n12236 VN.n12233 0.001
R15342 VN.n821 VN.n805 0.001
R15343 VN.n11121 VN.n11118 0.001
R15344 VN.n12262 VN.n12259 0.001
R15345 VN.n256 VN.n253 0.001
R15346 VN.n1553 VN.n1550 0.001
R15347 VN.n11141 VN.n11138 0.001
R15348 VN.n928 VN.n925 0.001
R15349 VN.n11397 VN.n11385 0.001
R15350 VN.n11157 VN.n11154 0.001
R15351 VN.n1615 VN.n1612 0.001
R15352 VN.n2323 VN.n2320 0.001
R15353 VN.n11175 VN.n11172 0.001
R15354 VN.n11191 VN.n11188 0.001
R15355 VN.n3042 VN.n3039 0.001
R15356 VN.n3785 VN.n3782 0.001
R15357 VN.n11209 VN.n11206 0.001
R15358 VN.n11225 VN.n11222 0.001
R15359 VN.n4539 VN.n4536 0.001
R15360 VN.n5317 VN.n5314 0.001
R15361 VN.n11243 VN.n11240 0.001
R15362 VN.n11259 VN.n11256 0.001
R15363 VN.n6106 VN.n6103 0.001
R15364 VN.n11276 VN.n11273 0.001
R15365 VN.n11292 VN.n11289 0.001
R15366 VN.n7738 VN.n7735 0.001
R15367 VN.n8586 VN.n8583 0.001
R15368 VN.n11310 VN.n11307 0.001
R15369 VN.n11326 VN.n11323 0.001
R15370 VN.n9445 VN.n9442 0.001
R15371 VN.n10331 VN.n10328 0.001
R15372 VN.n11344 VN.n11341 0.001
R15373 VN.n11360 VN.n11357 0.001
R15374 VN.n11492 VN.n11489 0.001
R15375 VN.n13137 VN.n13113 0.001
R15376 VN.n12182 VN.n12177 0.001
R15377 VN.n12282 VN.n12272 0.001
R15378 VN.n12317 VN.n12314 0.001
R15379 VN.n12299 VN.n12290 0.001
R15380 VN.n276 VN.n273 0.001
R15381 VN.n545 VN.n542 0.001
R15382 VN.n948 VN.n945 0.001
R15383 VN.n1220 VN.n1217 0.001
R15384 VN.n1635 VN.n1632 0.001
R15385 VN.n1910 VN.n1907 0.001
R15386 VN.n2343 VN.n2340 0.001
R15387 VN.n2619 VN.n2616 0.001
R15388 VN.n3062 VN.n3059 0.001
R15389 VN.n3341 VN.n3338 0.001
R15390 VN.n3805 VN.n3802 0.001
R15391 VN.n4085 VN.n4082 0.001
R15392 VN.n4559 VN.n4556 0.001
R15393 VN.n4842 VN.n4839 0.001
R15394 VN.n5337 VN.n5334 0.001
R15395 VN.n5621 VN.n5618 0.001
R15396 VN.n6126 VN.n6123 0.001
R15397 VN.n6413 VN.n6410 0.001
R15398 VN.n6858 VN.n6855 0.001
R15399 VN.n7758 VN.n7755 0.001
R15400 VN.n8049 VN.n8046 0.001
R15401 VN.n8606 VN.n8603 0.001
R15402 VN.n8898 VN.n8895 0.001
R15403 VN.n9465 VN.n9462 0.001
R15404 VN.n9760 VN.n9757 0.001
R15405 VN.n10679 VN.n10676 0.001
R15406 VN.n10662 VN.n10653 0.001
R15407 VN.n11509 VN.n11506 0.001
R15408 VN.n11524 VN.n11515 0.001
R15409 VN.n12630 VN.n12626 0.001
R15410 VN.n12635 VN.n12632 0.001
R15411 VN.n12343 VN.n12339 0.001
R15412 VN.n291 VN.n288 0.001
R15413 VN.n561 VN.n558 0.001
R15414 VN.n963 VN.n960 0.001
R15415 VN.n1236 VN.n1233 0.001
R15416 VN.n1650 VN.n1647 0.001
R15417 VN.n1926 VN.n1923 0.001
R15418 VN.n2358 VN.n2355 0.001
R15419 VN.n2635 VN.n2632 0.001
R15420 VN.n3077 VN.n3074 0.001
R15421 VN.n3357 VN.n3354 0.001
R15422 VN.n3820 VN.n3817 0.001
R15423 VN.n4101 VN.n4098 0.001
R15424 VN.n4574 VN.n4571 0.001
R15425 VN.n4858 VN.n4855 0.001
R15426 VN.n5352 VN.n5349 0.001
R15427 VN.n5637 VN.n5634 0.001
R15428 VN.n6141 VN.n6138 0.001
R15429 VN.n6429 VN.n6426 0.001
R15430 VN.n6874 VN.n6871 0.001
R15431 VN.n7773 VN.n7770 0.001
R15432 VN.n8065 VN.n8062 0.001
R15433 VN.n8621 VN.n8618 0.001
R15434 VN.n8914 VN.n8911 0.001
R15435 VN.n9799 VN.n9796 0.001
R15436 VN.n9795 VN.n9791 0.001
R15437 VN.n10694 VN.n10691 0.001
R15438 VN.n10647 VN.n10644 0.001
R15439 VN.n10707 VN.n10702 0.001
R15440 VN.n9782 VN.n9779 0.001
R15441 VN.n9814 VN.n9811 0.001
R15442 VN.n8949 VN.n8945 0.001
R15443 VN.n8953 VN.n8950 0.001
R15444 VN.n8081 VN.n8078 0.001
R15445 VN.n7788 VN.n7785 0.001
R15446 VN.n6890 VN.n6887 0.001
R15447 VN.n6445 VN.n6442 0.001
R15448 VN.n6156 VN.n6153 0.001
R15449 VN.n5653 VN.n5650 0.001
R15450 VN.n5367 VN.n5364 0.001
R15451 VN.n4874 VN.n4871 0.001
R15452 VN.n4589 VN.n4586 0.001
R15453 VN.n4117 VN.n4114 0.001
R15454 VN.n3835 VN.n3832 0.001
R15455 VN.n3373 VN.n3370 0.001
R15456 VN.n3092 VN.n3089 0.001
R15457 VN.n2651 VN.n2648 0.001
R15458 VN.n2373 VN.n2370 0.001
R15459 VN.n1942 VN.n1939 0.001
R15460 VN.n1665 VN.n1662 0.001
R15461 VN.n1252 VN.n1249 0.001
R15462 VN.n978 VN.n975 0.001
R15463 VN.n577 VN.n574 0.001
R15464 VN.n306 VN.n303 0.001
R15465 VN.n12661 VN.n12657 0.001
R15466 VN.n12666 VN.n12663 0.001
R15467 VN.n12425 VN.n12422 0.001
R15468 VN.n9827 VN.n9822 0.001
R15469 VN.n8936 VN.n8933 0.001
R15470 VN.n8968 VN.n8965 0.001
R15471 VN.n8116 VN.n8112 0.001
R15472 VN.n8120 VN.n8117 0.001
R15473 VN.n6906 VN.n6903 0.001
R15474 VN.n6461 VN.n6458 0.001
R15475 VN.n6171 VN.n6168 0.001
R15476 VN.n5669 VN.n5666 0.001
R15477 VN.n5382 VN.n5379 0.001
R15478 VN.n4890 VN.n4887 0.001
R15479 VN.n4604 VN.n4601 0.001
R15480 VN.n4133 VN.n4130 0.001
R15481 VN.n3850 VN.n3847 0.001
R15482 VN.n3389 VN.n3386 0.001
R15483 VN.n3107 VN.n3104 0.001
R15484 VN.n2667 VN.n2664 0.001
R15485 VN.n2388 VN.n2385 0.001
R15486 VN.n1958 VN.n1955 0.001
R15487 VN.n1680 VN.n1677 0.001
R15488 VN.n1268 VN.n1265 0.001
R15489 VN.n993 VN.n990 0.001
R15490 VN.n593 VN.n590 0.001
R15491 VN.n321 VN.n318 0.001
R15492 VN.n12772 VN.n12768 0.001
R15493 VN.n12777 VN.n12774 0.001
R15494 VN.n12441 VN.n12438 0.001
R15495 VN.n8981 VN.n8976 0.001
R15496 VN.n8103 VN.n8100 0.001
R15497 VN.n8135 VN.n8132 0.001
R15498 VN.n6941 VN.n6937 0.001
R15499 VN.n6477 VN.n6474 0.001
R15500 VN.n6186 VN.n6183 0.001
R15501 VN.n5685 VN.n5682 0.001
R15502 VN.n5397 VN.n5394 0.001
R15503 VN.n4906 VN.n4903 0.001
R15504 VN.n4619 VN.n4616 0.001
R15505 VN.n4149 VN.n4146 0.001
R15506 VN.n3865 VN.n3862 0.001
R15507 VN.n3405 VN.n3402 0.001
R15508 VN.n3122 VN.n3119 0.001
R15509 VN.n2683 VN.n2680 0.001
R15510 VN.n2403 VN.n2400 0.001
R15511 VN.n1974 VN.n1971 0.001
R15512 VN.n1695 VN.n1692 0.001
R15513 VN.n1284 VN.n1281 0.001
R15514 VN.n1008 VN.n1005 0.001
R15515 VN.n609 VN.n606 0.001
R15516 VN.n336 VN.n333 0.001
R15517 VN.n12806 VN.n12802 0.001
R15518 VN.n12811 VN.n12808 0.001
R15519 VN.n12457 VN.n12454 0.001
R15520 VN.n8148 VN.n8143 0.001
R15521 VN.n6928 VN.n6925 0.001
R15522 VN.n6512 VN.n6508 0.001
R15523 VN.n6516 VN.n6513 0.001
R15524 VN.n5701 VN.n5698 0.001
R15525 VN.n5412 VN.n5409 0.001
R15526 VN.n4922 VN.n4919 0.001
R15527 VN.n4634 VN.n4631 0.001
R15528 VN.n4165 VN.n4162 0.001
R15529 VN.n3880 VN.n3877 0.001
R15530 VN.n3421 VN.n3418 0.001
R15531 VN.n3137 VN.n3134 0.001
R15532 VN.n2699 VN.n2696 0.001
R15533 VN.n2418 VN.n2415 0.001
R15534 VN.n1990 VN.n1987 0.001
R15535 VN.n1710 VN.n1707 0.001
R15536 VN.n1300 VN.n1297 0.001
R15537 VN.n1023 VN.n1020 0.001
R15538 VN.n625 VN.n622 0.001
R15539 VN.n351 VN.n348 0.001
R15540 VN.n12837 VN.n12833 0.001
R15541 VN.n12842 VN.n12839 0.001
R15542 VN.n12473 VN.n12470 0.001
R15543 VN.n7337 VN.n7332 0.001
R15544 VN.n6499 VN.n6496 0.001
R15545 VN.n6531 VN.n6528 0.001
R15546 VN.n5736 VN.n5732 0.001
R15547 VN.n5740 VN.n5737 0.001
R15548 VN.n4938 VN.n4935 0.001
R15549 VN.n4649 VN.n4646 0.001
R15550 VN.n4181 VN.n4178 0.001
R15551 VN.n3895 VN.n3892 0.001
R15552 VN.n3437 VN.n3434 0.001
R15553 VN.n3152 VN.n3149 0.001
R15554 VN.n2715 VN.n2712 0.001
R15555 VN.n2433 VN.n2430 0.001
R15556 VN.n2006 VN.n2003 0.001
R15557 VN.n1725 VN.n1722 0.001
R15558 VN.n1316 VN.n1313 0.001
R15559 VN.n1038 VN.n1035 0.001
R15560 VN.n641 VN.n638 0.001
R15561 VN.n366 VN.n363 0.001
R15562 VN.n12865 VN.n12861 0.001
R15563 VN.n12870 VN.n12867 0.001
R15564 VN.n12489 VN.n12486 0.001
R15565 VN.n6544 VN.n6539 0.001
R15566 VN.n5723 VN.n5720 0.001
R15567 VN.n5755 VN.n5752 0.001
R15568 VN.n4973 VN.n4969 0.001
R15569 VN.n4977 VN.n4974 0.001
R15570 VN.n4197 VN.n4194 0.001
R15571 VN.n3910 VN.n3907 0.001
R15572 VN.n3453 VN.n3450 0.001
R15573 VN.n3167 VN.n3164 0.001
R15574 VN.n2731 VN.n2728 0.001
R15575 VN.n2448 VN.n2445 0.001
R15576 VN.n2022 VN.n2019 0.001
R15577 VN.n1740 VN.n1737 0.001
R15578 VN.n1332 VN.n1329 0.001
R15579 VN.n1053 VN.n1050 0.001
R15580 VN.n657 VN.n654 0.001
R15581 VN.n381 VN.n378 0.001
R15582 VN.n12896 VN.n12892 0.001
R15583 VN.n12901 VN.n12898 0.001
R15584 VN.n12505 VN.n12502 0.001
R15585 VN.n5768 VN.n5763 0.001
R15586 VN.n4960 VN.n4957 0.001
R15587 VN.n4992 VN.n4989 0.001
R15588 VN.n4232 VN.n4228 0.001
R15589 VN.n4236 VN.n4233 0.001
R15590 VN.n3469 VN.n3466 0.001
R15591 VN.n3182 VN.n3179 0.001
R15592 VN.n2747 VN.n2744 0.001
R15593 VN.n2463 VN.n2460 0.001
R15594 VN.n2038 VN.n2035 0.001
R15595 VN.n1755 VN.n1752 0.001
R15596 VN.n1348 VN.n1345 0.001
R15597 VN.n1068 VN.n1065 0.001
R15598 VN.n673 VN.n670 0.001
R15599 VN.n396 VN.n393 0.001
R15600 VN.n12927 VN.n12923 0.001
R15601 VN.n12932 VN.n12929 0.001
R15602 VN.n12521 VN.n12518 0.001
R15603 VN.n5005 VN.n5000 0.001
R15604 VN.n4219 VN.n4216 0.001
R15605 VN.n4251 VN.n4248 0.001
R15606 VN.n3504 VN.n3500 0.001
R15607 VN.n3508 VN.n3505 0.001
R15608 VN.n2763 VN.n2760 0.001
R15609 VN.n2478 VN.n2475 0.001
R15610 VN.n2054 VN.n2051 0.001
R15611 VN.n1770 VN.n1767 0.001
R15612 VN.n1364 VN.n1361 0.001
R15613 VN.n1083 VN.n1080 0.001
R15614 VN.n689 VN.n686 0.001
R15615 VN.n411 VN.n408 0.001
R15616 VN.n12958 VN.n12954 0.001
R15617 VN.n12963 VN.n12960 0.001
R15618 VN.n12537 VN.n12534 0.001
R15619 VN.n4264 VN.n4259 0.001
R15620 VN.n3491 VN.n3488 0.001
R15621 VN.n3523 VN.n3520 0.001
R15622 VN.n2798 VN.n2794 0.001
R15623 VN.n2802 VN.n2799 0.001
R15624 VN.n2070 VN.n2067 0.001
R15625 VN.n1785 VN.n1782 0.001
R15626 VN.n1380 VN.n1377 0.001
R15627 VN.n1098 VN.n1095 0.001
R15628 VN.n705 VN.n702 0.001
R15629 VN.n426 VN.n423 0.001
R15630 VN.n12989 VN.n12985 0.001
R15631 VN.n12994 VN.n12991 0.001
R15632 VN.n12553 VN.n12550 0.001
R15633 VN.n3536 VN.n3531 0.001
R15634 VN.n2785 VN.n2782 0.001
R15635 VN.n2817 VN.n2814 0.001
R15636 VN.n2105 VN.n2101 0.001
R15637 VN.n2109 VN.n2106 0.001
R15638 VN.n1396 VN.n1393 0.001
R15639 VN.n1113 VN.n1110 0.001
R15640 VN.n721 VN.n718 0.001
R15641 VN.n441 VN.n438 0.001
R15642 VN.n13020 VN.n13016 0.001
R15643 VN.n13025 VN.n13022 0.001
R15644 VN.n12569 VN.n12566 0.001
R15645 VN.n2830 VN.n2825 0.001
R15646 VN.n2092 VN.n2089 0.001
R15647 VN.n2124 VN.n2121 0.001
R15648 VN.n1431 VN.n1427 0.001
R15649 VN.n1435 VN.n1432 0.001
R15650 VN.n737 VN.n734 0.001
R15651 VN.n456 VN.n453 0.001
R15652 VN.n13051 VN.n13047 0.001
R15653 VN.n13056 VN.n13053 0.001
R15654 VN.n12585 VN.n12582 0.001
R15655 VN.n2137 VN.n2132 0.001
R15656 VN.n1418 VN.n1415 0.001
R15657 VN.n1450 VN.n1447 0.001
R15658 VN.n771 VN.n767 0.001
R15659 VN.n775 VN.n772 0.001
R15660 VN.n13082 VN.n13078 0.001
R15661 VN.n13087 VN.n13084 0.001
R15662 VN.n12601 VN.n12598 0.001
R15663 VN.n1463 VN.n1458 0.001
R15664 VN.n758 VN.n755 0.001
R15665 VN.n797 VN.n794 0.001
R15666 VN.n12759 VN.n12756 0.001
R15667 VN.n13107 VN.n13104 0.001
R15668 VN.n12617 VN.n12614 0.001
R15669 VN.n15 VN.n14 0.001
R15670 VN.n14 VN.n7 0.001
R15671 VN.n11540 VN.n11539 0.001
R15672 VN.n10720 VN.n10719 0.001
R15673 VN.n9860 VN.n9859 0.001
R15674 VN.n9012 VN.n9011 0.001
R15675 VN.n8179 VN.n8178 0.001
R15676 VN.n7368 VN.n7367 0.001
R15677 VN.n6575 VN.n6574 0.001
R15678 VN.n5799 VN.n5798 0.001
R15679 VN.n5036 VN.n5035 0.001
R15680 VN.n4295 VN.n4294 0.001
R15681 VN.n3567 VN.n3566 0.001
R15682 VN.n2861 VN.n2860 0.001
R15683 VN.n2168 VN.n2167 0.001
R15684 VN.n1494 VN.n1493 0.001
R15685 VN.n844 VN.n843 0.001
R15686 VN.n817 VN.n816 0.001
R15687 VN.n13133 VN.n13132 0.001
R15688 VN.n11779 VN.n11778 0.001
R15689 VN.n12360 VN.n12359 0.001
R15690 VN.n16 VN.n15 0.001
R15691 VN.n7 VN.n6 0.001
R15692 VN.n11541 VN.n11540 0.001
R15693 VN.n10721 VN.n10720 0.001
R15694 VN.n9861 VN.n9860 0.001
R15695 VN.n9013 VN.n9012 0.001
R15696 VN.n8180 VN.n8179 0.001
R15697 VN.n7369 VN.n7368 0.001
R15698 VN.n6576 VN.n6575 0.001
R15699 VN.n5800 VN.n5799 0.001
R15700 VN.n5037 VN.n5036 0.001
R15701 VN.n4296 VN.n4295 0.001
R15702 VN.n3568 VN.n3567 0.001
R15703 VN.n2862 VN.n2861 0.001
R15704 VN.n2169 VN.n2168 0.001
R15705 VN.n1495 VN.n1494 0.001
R15706 VN.n845 VN.n844 0.001
R15707 VN.n818 VN.n817 0.001
R15708 VN.n13135 VN.n13124 0.001
R15709 VN.n819 VN.n808 0.001
R15710 VN.n11542 VN.n11530 0.001
R15711 VN.n10722 VN.n10711 0.001
R15712 VN.n9862 VN.n9851 0.001
R15713 VN.n9014 VN.n9003 0.001
R15714 VN.n8181 VN.n8170 0.001
R15715 VN.n7370 VN.n7359 0.001
R15716 VN.n6577 VN.n6566 0.001
R15717 VN.n5801 VN.n5790 0.001
R15718 VN.n5038 VN.n5027 0.001
R15719 VN.n4297 VN.n4286 0.001
R15720 VN.n3569 VN.n3558 0.001
R15721 VN.n2863 VN.n2852 0.001
R15722 VN.n2170 VN.n2159 0.001
R15723 VN.n1496 VN.n1485 0.001
R15724 VN.n846 VN.n835 0.001
R15725 VN.n179 VN.n178 0.001
R15726 VN.n13134 VN.n13133 0.001
R15727 VN.n11782 VN.n11781 0.001
R15728 VN.n174 VN.n173 0.001
R15729 VN.n11571 VN.n11567 0.001
C0 fc2 s3 12294.20fF
C1 fc2 s4 4037.63fF
C2 s2 out 7185.27fF
C3 VN s4 12347.40fF
C4 VP fc1 5164.57fF
C5 dw_2450_33450# fc2 7202.83fF
C6 out s3 4043.75fF
C7 dw_2450_2450# s4 112.05fF
C8 VP s1 21658.10fF
C9 fc2 VN 2899.38fF
C10 fc1 s1 7117.35fF
C11 dw_2450_33450# out 1677.01fF
C12 fc1 s2 21602.30fF
C13 dw_2450_33450# s3 120.53fF
C14 fc1 out 5543.06fF
C15 dw_2450_2450# fc2 1719.66fF
C16 fc2 out 3189.96fF
C17 dw_2450_2450# VN 7050.43fF
C18 s4 a_400_62400# -1496.16fF
C19 s3 a_400_62400# -1469.96fF
C20 out a_400_62400# 3551.74fF
C21 s2 a_400_62400# -2409.67fF
C22 s1 a_400_62400# -2481.33fF
C23 VN a_400_62400# -5083.38fF
C24 fc2 a_400_62400# -4550.72fF
C25 fc1 a_400_62400# 5423.77fF
C26 VP a_400_62400# 1690.54fF
C27 dw_2450_2450# a_400_62400# 9423.81fF $ **FLOATING
C28 dw_2450_33450# a_400_62400# 9479.45fF $ **FLOATING
C29 VN.n0 a_400_62400# 3.15fF
C30 VN.n1 a_400_62400# 0.75fF
C31 VN.n2 a_400_62400# 1.18fF
C32 VN.n3 a_400_62400# 2.79fF
C33 VN.n4 a_400_62400# 0.75fF
C34 VN.n5 a_400_62400# 1.18fF
C35 VN.n6 a_400_62400# 0.51fF
C36 VN.n8 a_400_62400# 0.52fF
C37 VN.n9 a_400_62400# 0.71fF
C38 VN.n10 a_400_62400# 0.52fF
C39 VN.n11 a_400_62400# 0.71fF
C40 VN.n12 a_400_62400# 2.09fF
C41 VN.n13 a_400_62400# 2.07fF
C42 VN.n14 a_400_62400# 218.10fF
C43 VN.n16 a_400_62400# 0.51fF
C44 VN.n17 a_400_62400# 5.29fF
C45 VN.n18 a_400_62400# 3.68fF
C46 VN.n19 a_400_62400# 0.04fF
C47 VN.n20 a_400_62400# 0.03fF
C48 VN.n21 a_400_62400# 0.02fF
C49 VN.n22 a_400_62400# 0.06fF
C50 VN.n23 a_400_62400# 0.13fF
C51 VN.n24 a_400_62400# 0.39fF
C52 VN.n25 a_400_62400# 0.83fF
C53 VN.n26 a_400_62400# 0.04fF
C54 VN.n27 a_400_62400# 0.04fF
C55 VN.n28 a_400_62400# 0.03fF
C56 VN.n29 a_400_62400# 0.32fF
C57 VN.n30 a_400_62400# 0.20fF
C58 VN.n31 a_400_62400# 0.24fF
C59 VN.n32 a_400_62400# 3.25fF
C60 VN.n33 a_400_62400# 5.87fF
C61 VN.n34 a_400_62400# 3.76fF
C62 VN.n35 a_400_62400# 5.87fF
C63 VN.n36 a_400_62400# 3.74fF
C64 VN.n37 a_400_62400# 3.25fF
C65 VN.n38 a_400_62400# 5.87fF
C66 VN.n39 a_400_62400# 3.74fF
C67 VN.n40 a_400_62400# 3.25fF
C68 VN.n41 a_400_62400# 5.87fF
C69 VN.n42 a_400_62400# 3.74fF
C70 VN.n43 a_400_62400# 3.25fF
C71 VN.n44 a_400_62400# 5.87fF
C72 VN.n45 a_400_62400# 3.74fF
C73 VN.n46 a_400_62400# 3.25fF
C74 VN.n47 a_400_62400# 5.87fF
C75 VN.n48 a_400_62400# 3.74fF
C76 VN.n49 a_400_62400# 3.25fF
C77 VN.n50 a_400_62400# 5.87fF
C78 VN.n51 a_400_62400# 3.74fF
C79 VN.n52 a_400_62400# 3.25fF
C80 VN.n53 a_400_62400# 5.87fF
C81 VN.n54 a_400_62400# 3.74fF
C82 VN.n55 a_400_62400# 3.25fF
C83 VN.n56 a_400_62400# 5.87fF
C84 VN.n57 a_400_62400# 3.74fF
C85 VN.n58 a_400_62400# 3.25fF
C86 VN.n59 a_400_62400# 5.87fF
C87 VN.n60 a_400_62400# 3.74fF
C88 VN.n61 a_400_62400# 3.25fF
C89 VN.n62 a_400_62400# 5.87fF
C90 VN.n63 a_400_62400# 3.74fF
C91 VN.n64 a_400_62400# 3.25fF
C92 VN.n65 a_400_62400# 5.87fF
C93 VN.n66 a_400_62400# 3.74fF
C94 VN.n67 a_400_62400# 3.25fF
C95 VN.n68 a_400_62400# 5.87fF
C96 VN.n69 a_400_62400# 3.74fF
C97 VN.n70 a_400_62400# 3.25fF
C98 VN.n71 a_400_62400# 5.12fF
C99 VN.n72 a_400_62400# 3.74fF
C100 VN.n73 a_400_62400# 0.28fF
C101 VN.n74 a_400_62400# 2.93fF
C102 VN.n75 a_400_62400# 1.71fF
C103 VN.n76 a_400_62400# 0.41fF
C104 VN.n77 a_400_62400# 0.42fF
C105 VN.n78 a_400_62400# 2.84fF
C106 VN.n79 a_400_62400# 1.60fF
C107 VN.n80 a_400_62400# 0.44fF
C108 VN.n81 a_400_62400# 1.24fF
C109 VN.n82 a_400_62400# 5.48fF
C110 VN.n83 a_400_62400# 2.47fF
C111 VN.t408 a_400_62400# 0.03fF
C112 VN.n84 a_400_62400# 1.19fF
C113 VN.t1064 a_400_62400# 0.03fF
C114 VN.n85 a_400_62400# 1.20fF
C115 VN.n86 a_400_62400# 0.04fF
C116 VN.n87 a_400_62400# 0.03fF
C117 VN.n88 a_400_62400# 0.07fF
C118 VN.n89 a_400_62400# 0.13fF
C119 VN.n90 a_400_62400# 0.39fF
C120 VN.n91 a_400_62400# 0.83fF
C121 VN.n92 a_400_62400# 0.04fF
C122 VN.n93 a_400_62400# 0.04fF
C123 VN.n94 a_400_62400# 0.03fF
C124 VN.n95 a_400_62400# 0.32fF
C125 VN.n96 a_400_62400# 0.02fF
C126 VN.n97 a_400_62400# 0.20fF
C127 VN.n98 a_400_62400# 0.24fF
C128 VN.n99 a_400_62400# 5.26fF
C129 VN.n100 a_400_62400# 3.62fF
C130 VN.t1459 a_400_62400# 0.03fF
C131 VN.n101 a_400_62400# 0.02fF
C132 VN.n102 a_400_62400# 0.50fF
C133 VN.n103 a_400_62400# 27.83fF
C134 VN.t478 a_400_62400# 0.03fF
C135 VN.n104 a_400_62400# 1.20fF
C136 VN.t1632 a_400_62400# 0.03fF
C137 VN.n105 a_400_62400# 0.02fF
C138 VN.n106 a_400_62400# 0.50fF
C139 VN.t2198 a_400_62400# 0.03fF
C140 VN.n107 a_400_62400# 1.19fF
C141 VN.t2133 a_400_62400# 0.03fF
C142 VN.n108 a_400_62400# 1.20fF
C143 VN.t761 a_400_62400# 0.03fF
C144 VN.n109 a_400_62400# 0.02fF
C145 VN.n110 a_400_62400# 0.50fF
C146 VN.t1448 a_400_62400# 0.03fF
C147 VN.n111 a_400_62400# 1.19fF
C148 VN.t1259 a_400_62400# 0.03fF
C149 VN.n112 a_400_62400# 1.20fF
C150 VN.t2537 a_400_62400# 0.03fF
C151 VN.n113 a_400_62400# 0.02fF
C152 VN.n114 a_400_62400# 0.50fF
C153 VN.t579 a_400_62400# 0.03fF
C154 VN.n115 a_400_62400# 1.19fF
C155 VN.t389 a_400_62400# 0.03fF
C156 VN.n116 a_400_62400# 1.20fF
C157 VN.t1672 a_400_62400# 0.03fF
C158 VN.n117 a_400_62400# 0.02fF
C159 VN.n118 a_400_62400# 0.50fF
C160 VN.t2237 a_400_62400# 0.03fF
C161 VN.n119 a_400_62400# 1.19fF
C162 VN.t2042 a_400_62400# 0.03fF
C163 VN.n120 a_400_62400# 1.20fF
C164 VN.t2171 a_400_62400# 0.03fF
C165 VN.n121 a_400_62400# 0.02fF
C166 VN.n122 a_400_62400# 0.50fF
C167 VN.t173 a_400_62400# 0.03fF
C168 VN.n123 a_400_62400# 1.19fF
C169 VN.t2511 a_400_62400# 0.03fF
C170 VN.n124 a_400_62400# 1.20fF
C171 VN.t1304 a_400_62400# 0.03fF
C172 VN.n125 a_400_62400# 0.02fF
C173 VN.n126 a_400_62400# 0.50fF
C174 VN.t1834 a_400_62400# 0.03fF
C175 VN.n127 a_400_62400# 1.19fF
C176 VN.t1648 a_400_62400# 0.03fF
C177 VN.n128 a_400_62400# 1.20fF
C178 VN.t440 a_400_62400# 0.03fF
C179 VN.n129 a_400_62400# 0.02fF
C180 VN.n130 a_400_62400# 0.50fF
C181 VN.t960 a_400_62400# 0.03fF
C182 VN.n131 a_400_62400# 1.19fF
C183 VN.t887 a_400_62400# 0.03fF
C184 VN.n132 a_400_62400# 1.20fF
C185 VN.t2085 a_400_62400# 0.03fF
C186 VN.n133 a_400_62400# 0.02fF
C187 VN.n134 a_400_62400# 0.50fF
C188 VN.t52 a_400_62400# 0.03fF
C189 VN.n135 a_400_62400# 1.19fF
C190 VN.t2548 a_400_62400# 0.03fF
C191 VN.n136 a_400_62400# 1.20fF
C192 VN.t1210 a_400_62400# 0.03fF
C193 VN.n137 a_400_62400# 0.02fF
C194 VN.n138 a_400_62400# 0.50fF
C195 VN.t1747 a_400_62400# 0.03fF
C196 VN.n139 a_400_62400# 1.19fF
C197 VN.t1680 a_400_62400# 0.03fF
C198 VN.n140 a_400_62400# 1.20fF
C199 VN.t347 a_400_62400# 0.03fF
C200 VN.n141 a_400_62400# 0.02fF
C201 VN.n142 a_400_62400# 0.50fF
C202 VN.t874 a_400_62400# 0.03fF
C203 VN.n143 a_400_62400# 1.19fF
C204 VN.t814 a_400_62400# 0.03fF
C205 VN.n144 a_400_62400# 1.20fF
C206 VN.t1990 a_400_62400# 0.03fF
C207 VN.n145 a_400_62400# 0.02fF
C208 VN.n146 a_400_62400# 0.50fF
C209 VN.t2535 a_400_62400# 0.03fF
C210 VN.n147 a_400_62400# 1.19fF
C211 VN.t2471 a_400_62400# 0.03fF
C212 VN.n148 a_400_62400# 1.20fF
C213 VN.t1116 a_400_62400# 0.03fF
C214 VN.n149 a_400_62400# 0.02fF
C215 VN.n150 a_400_62400# 0.50fF
C216 VN.t1792 a_400_62400# 0.03fF
C217 VN.n151 a_400_62400# 1.19fF
C218 VN.t1608 a_400_62400# 0.03fF
C219 VN.n152 a_400_62400# 1.20fF
C220 VN.t395 a_400_62400# 0.03fF
C221 VN.n153 a_400_62400# 0.02fF
C222 VN.n154 a_400_62400# 0.50fF
C223 VN.t917 a_400_62400# 0.03fF
C224 VN.n155 a_400_62400# 1.19fF
C225 VN.t742 a_400_62400# 0.03fF
C226 VN.n156 a_400_62400# 1.20fF
C227 VN.t1537 a_400_62400# 0.03fF
C228 VN.n157 a_400_62400# 0.02fF
C229 VN.n158 a_400_62400# 0.50fF
C230 VN.t492 a_400_62400# 0.03fF
C231 VN.n159 a_400_62400# 1.19fF
C232 VN.t285 a_400_62400# 0.03fF
C233 VN.n160 a_400_62400# 1.20fF
C234 VN.t665 a_400_62400# 0.03fF
C235 VN.n161 a_400_62400# 0.02fF
C236 VN.n162 a_400_62400# 0.50fF
C237 VN.t2147 a_400_62400# 0.03fF
C238 VN.n163 a_400_62400# 1.19fF
C239 VN.t1937 a_400_62400# 0.03fF
C240 VN.n164 a_400_62400# 1.20fF
C241 VN.t2325 a_400_62400# 0.03fF
C242 VN.n165 a_400_62400# 0.02fF
C243 VN.n166 a_400_62400# 0.50fF
C244 VN.t1277 a_400_62400# 0.03fF
C245 VN.n167 a_400_62400# 1.19fF
C246 VN.t335 a_400_62400# 0.03fF
C247 VN.n168 a_400_62400# 0.59fF
C248 VN.t51 a_400_62400# 229.46fF
C249 VN.t588 a_400_62400# 0.03fF
C250 VN.n169 a_400_62400# 1.75fF
C251 VN.n170 a_400_62400# 0.33fF
C252 VN.n171 a_400_62400# 28.25fF
C253 VN.n172 a_400_62400# 2.32fF
C254 VN.n173 a_400_62400# 4.41fF
C255 VN.n174 a_400_62400# 24.43fF
C256 VN.n175 a_400_62400# 13.29fF
C257 VN.n176 a_400_62400# 3.21fF
C258 VN.n177 a_400_62400# 1.02fF
C259 VN.n178 a_400_62400# 0.70fF
C260 VN.n179 a_400_62400# 13.15fF
C261 VN.n180 a_400_62400# 5.93fF
C262 VN.n181 a_400_62400# 3.15fF
C263 VN.n182 a_400_62400# 6.92fF
C264 VN.n183 a_400_62400# 0.35fF
C265 VN.n184 a_400_62400# 0.19fF
C266 VN.n185 a_400_62400# 2.01fF
C267 VN.n186 a_400_62400# 0.14fF
C268 VN.n187 a_400_62400# 0.03fF
C269 VN.n188 a_400_62400# 0.01fF
C270 VN.n189 a_400_62400# 0.01fF
C271 VN.n190 a_400_62400# 0.01fF
C272 VN.n191 a_400_62400# 0.02fF
C273 VN.n192 a_400_62400# 0.03fF
C274 VN.n193 a_400_62400# 0.03fF
C275 VN.n194 a_400_62400# 0.14fF
C276 VN.n195 a_400_62400# 0.13fF
C277 VN.n196 a_400_62400# 0.20fF
C278 VN.n197 a_400_62400# 0.37fF
C279 VN.t2366 a_400_62400# 0.03fF
C280 VN.n198 a_400_62400# 0.85fF
C281 VN.n199 a_400_62400# 0.81fF
C282 VN.n200 a_400_62400# 2.53fF
C283 VN.n201 a_400_62400# 0.08fF
C284 VN.n202 a_400_62400# 0.04fF
C285 VN.n203 a_400_62400# 0.05fF
C286 VN.n204 a_400_62400# 1.33fF
C287 VN.n205 a_400_62400# 0.03fF
C288 VN.n206 a_400_62400# 0.01fF
C289 VN.n207 a_400_62400# 0.02fF
C290 VN.n208 a_400_62400# 0.11fF
C291 VN.n209 a_400_62400# 0.48fF
C292 VN.n210 a_400_62400# 2.48fF
C293 VN.t520 a_400_62400# 0.03fF
C294 VN.n211 a_400_62400# 0.32fF
C295 VN.n212 a_400_62400# 0.48fF
C296 VN.n213 a_400_62400# 0.81fF
C297 VN.n214 a_400_62400# 0.16fF
C298 VN.t2018 a_400_62400# 0.03fF
C299 VN.n215 a_400_62400# 0.19fF
C300 VN.n217 a_400_62400# 0.93fF
C301 VN.n218 a_400_62400# 0.30fF
C302 VN.n219 a_400_62400# 0.34fF
C303 VN.n220 a_400_62400# 0.12fF
C304 VN.n221 a_400_62400# 0.30fF
C305 VN.n222 a_400_62400# 0.93fF
C306 VN.n223 a_400_62400# 1.55fF
C307 VN.n224 a_400_62400# 0.29fF
C308 VN.n225 a_400_62400# 0.34fF
C309 VN.n226 a_400_62400# 0.12fF
C310 VN.n227 a_400_62400# 2.52fF
C311 VN.t1622 a_400_62400# 0.03fF
C312 VN.n228 a_400_62400# 0.32fF
C313 VN.n229 a_400_62400# 1.22fF
C314 VN.n230 a_400_62400# 0.07fF
C315 VN.t145 a_400_62400# 0.03fF
C316 VN.n231 a_400_62400# 0.16fF
C317 VN.n232 a_400_62400# 0.19fF
C318 VN.n234 a_400_62400# 27.83fF
C319 VN.n235 a_400_62400# 0.13fF
C320 VN.n236 a_400_62400# 0.28fF
C321 VN.n237 a_400_62400# 0.09fF
C322 VN.n238 a_400_62400# 0.08fF
C323 VN.n239 a_400_62400# 0.09fF
C324 VN.n240 a_400_62400# 0.24fF
C325 VN.n241 a_400_62400# 0.26fF
C326 VN.n242 a_400_62400# 1.39fF
C327 VN.n243 a_400_62400# 0.72fF
C328 VN.n244 a_400_62400# 3.13fF
C329 VN.n245 a_400_62400# 0.16fF
C330 VN.t231 a_400_62400# 0.03fF
C331 VN.n246 a_400_62400# 0.19fF
C332 VN.t1386 a_400_62400# 0.03fF
C333 VN.n248 a_400_62400# 0.32fF
C334 VN.n249 a_400_62400# 0.48fF
C335 VN.n250 a_400_62400# 0.81fF
C336 VN.n251 a_400_62400# 0.95fF
C337 VN.n252 a_400_62400# 2.31fF
C338 VN.n253 a_400_62400# 3.27fF
C339 VN.t1018 a_400_62400# 0.03fF
C340 VN.n254 a_400_62400# 0.16fF
C341 VN.n255 a_400_62400# 0.19fF
C342 VN.t2486 a_400_62400# 0.03fF
C343 VN.n257 a_400_62400# 0.32fF
C344 VN.n258 a_400_62400# 1.22fF
C345 VN.n259 a_400_62400# 0.07fF
C346 VN.n260 a_400_62400# 2.51fF
C347 VN.n261 a_400_62400# 0.16fF
C348 VN.t1145 a_400_62400# 0.03fF
C349 VN.n262 a_400_62400# 0.19fF
C350 VN.t2289 a_400_62400# 0.03fF
C351 VN.n264 a_400_62400# 0.32fF
C352 VN.n265 a_400_62400# 0.48fF
C353 VN.n266 a_400_62400# 0.81fF
C354 VN.n267 a_400_62400# 1.24fF
C355 VN.n268 a_400_62400# 0.43fF
C356 VN.n269 a_400_62400# 0.43fF
C357 VN.n270 a_400_62400# 1.24fF
C358 VN.n271 a_400_62400# 1.46fF
C359 VN.n272 a_400_62400# 0.21fF
C360 VN.n273 a_400_62400# 6.64fF
C361 VN.t1810 a_400_62400# 0.03fF
C362 VN.n274 a_400_62400# 0.16fF
C363 VN.n275 a_400_62400# 0.19fF
C364 VN.t864 a_400_62400# 0.03fF
C365 VN.n277 a_400_62400# 0.32fF
C366 VN.n278 a_400_62400# 1.22fF
C367 VN.n279 a_400_62400# 0.07fF
C368 VN.n280 a_400_62400# 2.51fF
C369 VN.n281 a_400_62400# 3.57fF
C370 VN.t1420 a_400_62400# 0.03fF
C371 VN.n282 a_400_62400# 0.32fF
C372 VN.n283 a_400_62400# 0.48fF
C373 VN.n284 a_400_62400# 0.81fF
C374 VN.n285 a_400_62400# 0.16fF
C375 VN.t282 a_400_62400# 0.03fF
C376 VN.n286 a_400_62400# 0.19fF
C377 VN.n288 a_400_62400# 6.91fF
C378 VN.t935 a_400_62400# 0.03fF
C379 VN.n289 a_400_62400# 0.16fF
C380 VN.n290 a_400_62400# 0.19fF
C381 VN.t2526 a_400_62400# 0.03fF
C382 VN.n292 a_400_62400# 0.32fF
C383 VN.n293 a_400_62400# 1.22fF
C384 VN.n294 a_400_62400# 0.07fF
C385 VN.n295 a_400_62400# 2.51fF
C386 VN.n296 a_400_62400# 3.57fF
C387 VN.t1886 a_400_62400# 0.03fF
C388 VN.n297 a_400_62400# 0.32fF
C389 VN.n298 a_400_62400# 0.48fF
C390 VN.n299 a_400_62400# 0.81fF
C391 VN.n300 a_400_62400# 0.16fF
C392 VN.t752 a_400_62400# 0.03fF
C393 VN.n301 a_400_62400# 0.19fF
C394 VN.n303 a_400_62400# 6.92fF
C395 VN.t13 a_400_62400# 0.03fF
C396 VN.n304 a_400_62400# 0.16fF
C397 VN.n305 a_400_62400# 0.19fF
C398 VN.t507 a_400_62400# 0.03fF
C399 VN.n307 a_400_62400# 0.32fF
C400 VN.n308 a_400_62400# 1.22fF
C401 VN.n309 a_400_62400# 0.07fF
C402 VN.n310 a_400_62400# 2.51fF
C403 VN.n311 a_400_62400# 3.57fF
C404 VN.t1014 a_400_62400# 0.03fF
C405 VN.n312 a_400_62400# 0.32fF
C406 VN.n313 a_400_62400# 0.48fF
C407 VN.n314 a_400_62400# 0.81fF
C408 VN.n315 a_400_62400# 0.16fF
C409 VN.t2410 a_400_62400# 0.03fF
C410 VN.n316 a_400_62400# 0.19fF
C411 VN.n318 a_400_62400# 6.92fF
C412 VN.t566 a_400_62400# 0.03fF
C413 VN.n319 a_400_62400# 0.16fF
C414 VN.n320 a_400_62400# 0.19fF
C415 VN.t2160 a_400_62400# 0.03fF
C416 VN.n322 a_400_62400# 0.32fF
C417 VN.n323 a_400_62400# 1.22fF
C418 VN.n324 a_400_62400# 0.07fF
C419 VN.n325 a_400_62400# 2.51fF
C420 VN.n326 a_400_62400# 3.57fF
C421 VN.t140 a_400_62400# 0.03fF
C422 VN.n327 a_400_62400# 0.32fF
C423 VN.n328 a_400_62400# 0.48fF
C424 VN.n329 a_400_62400# 0.81fF
C425 VN.n330 a_400_62400# 0.16fF
C426 VN.t1545 a_400_62400# 0.03fF
C427 VN.n331 a_400_62400# 0.19fF
C428 VN.n333 a_400_62400# 6.92fF
C429 VN.t2226 a_400_62400# 0.03fF
C430 VN.n334 a_400_62400# 0.16fF
C431 VN.n335 a_400_62400# 0.19fF
C432 VN.t1292 a_400_62400# 0.03fF
C433 VN.n337 a_400_62400# 0.32fF
C434 VN.n338 a_400_62400# 1.22fF
C435 VN.n339 a_400_62400# 0.07fF
C436 VN.n340 a_400_62400# 2.51fF
C437 VN.n341 a_400_62400# 3.57fF
C438 VN.t1804 a_400_62400# 0.03fF
C439 VN.n342 a_400_62400# 0.32fF
C440 VN.n343 a_400_62400# 0.48fF
C441 VN.n344 a_400_62400# 0.81fF
C442 VN.n345 a_400_62400# 0.16fF
C443 VN.t675 a_400_62400# 0.03fF
C444 VN.n346 a_400_62400# 0.19fF
C445 VN.n348 a_400_62400# 6.92fF
C446 VN.t1479 a_400_62400# 0.03fF
C447 VN.n349 a_400_62400# 0.16fF
C448 VN.n350 a_400_62400# 0.19fF
C449 VN.t425 a_400_62400# 0.03fF
C450 VN.n352 a_400_62400# 0.32fF
C451 VN.n353 a_400_62400# 1.22fF
C452 VN.n354 a_400_62400# 0.07fF
C453 VN.n355 a_400_62400# 2.51fF
C454 VN.n356 a_400_62400# 3.57fF
C455 VN.t929 a_400_62400# 0.03fF
C456 VN.n357 a_400_62400# 0.32fF
C457 VN.n358 a_400_62400# 0.48fF
C458 VN.n359 a_400_62400# 0.81fF
C459 VN.n360 a_400_62400# 0.16fF
C460 VN.t2334 a_400_62400# 0.03fF
C461 VN.n361 a_400_62400# 0.19fF
C462 VN.n363 a_400_62400# 6.92fF
C463 VN.t611 a_400_62400# 0.03fF
C464 VN.n364 a_400_62400# 0.16fF
C465 VN.n365 a_400_62400# 0.19fF
C466 VN.t2071 a_400_62400# 0.03fF
C467 VN.n367 a_400_62400# 0.32fF
C468 VN.n368 a_400_62400# 1.22fF
C469 VN.n369 a_400_62400# 0.07fF
C470 VN.n370 a_400_62400# 2.51fF
C471 VN.n371 a_400_62400# 3.57fF
C472 VN.t3 a_400_62400# 0.03fF
C473 VN.n372 a_400_62400# 0.32fF
C474 VN.n373 a_400_62400# 0.48fF
C475 VN.n374 a_400_62400# 0.81fF
C476 VN.n375 a_400_62400# 0.16fF
C477 VN.t1469 a_400_62400# 0.03fF
C478 VN.n376 a_400_62400# 0.19fF
C479 VN.n378 a_400_62400# 6.92fF
C480 VN.t2263 a_400_62400# 0.03fF
C481 VN.n379 a_400_62400# 0.16fF
C482 VN.n380 a_400_62400# 0.19fF
C483 VN.t1200 a_400_62400# 0.03fF
C484 VN.n382 a_400_62400# 0.32fF
C485 VN.n383 a_400_62400# 1.22fF
C486 VN.n384 a_400_62400# 0.07fF
C487 VN.n385 a_400_62400# 2.51fF
C488 VN.n386 a_400_62400# 3.57fF
C489 VN.t1723 a_400_62400# 0.03fF
C490 VN.n387 a_400_62400# 0.32fF
C491 VN.n388 a_400_62400# 0.48fF
C492 VN.n389 a_400_62400# 0.81fF
C493 VN.n390 a_400_62400# 0.16fF
C494 VN.t600 a_400_62400# 0.03fF
C495 VN.n391 a_400_62400# 0.19fF
C496 VN.n393 a_400_62400# 6.92fF
C497 VN.t1398 a_400_62400# 0.03fF
C498 VN.n394 a_400_62400# 0.16fF
C499 VN.n395 a_400_62400# 0.19fF
C500 VN.t332 a_400_62400# 0.03fF
C501 VN.n397 a_400_62400# 0.32fF
C502 VN.n398 a_400_62400# 1.22fF
C503 VN.n399 a_400_62400# 0.07fF
C504 VN.n400 a_400_62400# 2.51fF
C505 VN.n401 a_400_62400# 3.57fF
C506 VN.t850 a_400_62400# 0.03fF
C507 VN.n402 a_400_62400# 0.32fF
C508 VN.n403 a_400_62400# 0.48fF
C509 VN.n404 a_400_62400# 0.81fF
C510 VN.n405 a_400_62400# 0.16fF
C511 VN.t2375 a_400_62400# 0.03fF
C512 VN.n406 a_400_62400# 0.19fF
C513 VN.n408 a_400_62400# 6.92fF
C514 VN.t537 a_400_62400# 0.03fF
C515 VN.n409 a_400_62400# 0.16fF
C516 VN.n410 a_400_62400# 0.19fF
C517 VN.t1978 a_400_62400# 0.03fF
C518 VN.n412 a_400_62400# 0.32fF
C519 VN.n413 a_400_62400# 1.22fF
C520 VN.n414 a_400_62400# 0.07fF
C521 VN.n415 a_400_62400# 2.51fF
C522 VN.n416 a_400_62400# 3.57fF
C523 VN.t84 a_400_62400# 0.03fF
C524 VN.n417 a_400_62400# 0.32fF
C525 VN.n418 a_400_62400# 0.48fF
C526 VN.n419 a_400_62400# 0.81fF
C527 VN.n420 a_400_62400# 0.16fF
C528 VN.t1508 a_400_62400# 0.03fF
C529 VN.n421 a_400_62400# 0.19fF
C530 VN.n423 a_400_62400# 6.92fF
C531 VN.t2192 a_400_62400# 0.03fF
C532 VN.n424 a_400_62400# 0.16fF
C533 VN.n425 a_400_62400# 0.19fF
C534 VN.t1247 a_400_62400# 0.03fF
C535 VN.n427 a_400_62400# 0.32fF
C536 VN.n428 a_400_62400# 1.22fF
C537 VN.n429 a_400_62400# 0.07fF
C538 VN.n430 a_400_62400# 2.51fF
C539 VN.n431 a_400_62400# 3.57fF
C540 VN.t788 a_400_62400# 0.03fF
C541 VN.n432 a_400_62400# 0.32fF
C542 VN.n433 a_400_62400# 0.48fF
C543 VN.n434 a_400_62400# 0.81fF
C544 VN.n435 a_400_62400# 0.16fF
C545 VN.t2178 a_400_62400# 0.03fF
C546 VN.n436 a_400_62400# 0.19fF
C547 VN.n438 a_400_62400# 6.92fF
C548 VN.t1323 a_400_62400# 0.03fF
C549 VN.n439 a_400_62400# 0.16fF
C550 VN.n440 a_400_62400# 0.19fF
C551 VN.t2365 a_400_62400# 0.03fF
C552 VN.n442 a_400_62400# 0.32fF
C553 VN.n443 a_400_62400# 1.22fF
C554 VN.n444 a_400_62400# 0.07fF
C555 VN.n445 a_400_62400# 2.51fF
C556 VN.n446 a_400_62400# 3.57fF
C557 VN.t2440 a_400_62400# 0.03fF
C558 VN.n447 a_400_62400# 0.32fF
C559 VN.n448 a_400_62400# 0.48fF
C560 VN.n449 a_400_62400# 0.81fF
C561 VN.n450 a_400_62400# 0.16fF
C562 VN.t1310 a_400_62400# 0.03fF
C563 VN.n451 a_400_62400# 0.19fF
C564 VN.n453 a_400_62400# 6.92fF
C565 VN.t1966 a_400_62400# 0.03fF
C566 VN.n454 a_400_62400# 0.16fF
C567 VN.n455 a_400_62400# 0.19fF
C568 VN.t1495 a_400_62400# 0.03fF
C569 VN.n457 a_400_62400# 0.32fF
C570 VN.n458 a_400_62400# 1.22fF
C571 VN.n459 a_400_62400# 0.07fF
C572 VN.n460 a_400_62400# 2.51fF
C573 VN.n461 a_400_62400# 3.57fF
C574 VN.t1578 a_400_62400# 0.03fF
C575 VN.n462 a_400_62400# 0.32fF
C576 VN.n463 a_400_62400# 0.48fF
C577 VN.n464 a_400_62400# 0.81fF
C578 VN.n465 a_400_62400# 0.16fF
C579 VN.t449 a_400_62400# 0.03fF
C580 VN.n466 a_400_62400# 0.19fF
C581 VN.n468 a_400_62400# 2.51fF
C582 VN.n469 a_400_62400# 3.59fF
C583 VN.t451 a_400_62400# 0.03fF
C584 VN.n470 a_400_62400# 0.32fF
C585 VN.n471 a_400_62400# 0.48fF
C586 VN.n472 a_400_62400# 0.81fF
C587 VN.t763 a_400_62400# 0.03fF
C588 VN.n473 a_400_62400# 1.63fF
C589 VN.n474 a_400_62400# 0.56fF
C590 VN.n475 a_400_62400# 0.59fF
C591 VN.n476 a_400_62400# 0.49fF
C592 VN.n477 a_400_62400# 0.28fF
C593 VN.n478 a_400_62400# 0.34fF
C594 VN.n479 a_400_62400# 1.71fF
C595 VN.n480 a_400_62400# 1.21fF
C596 VN.n481 a_400_62400# 1.54fF
C597 VN.n482 a_400_62400# 4.06fF
C598 VN.t257 a_400_62400# 28.64fF
C599 VN.n483 a_400_62400# 28.43fF
C600 VN.n485 a_400_62400# 0.50fF
C601 VN.n486 a_400_62400# 0.31fF
C602 VN.n487 a_400_62400# 3.78fF
C603 VN.n488 a_400_62400# 2.68fF
C604 VN.n489 a_400_62400# 5.46fF
C605 VN.n490 a_400_62400# 0.34fF
C606 VN.n491 a_400_62400# 0.02fF
C607 VN.t2165 a_400_62400# 0.03fF
C608 VN.n492 a_400_62400# 0.34fF
C609 VN.t2451 a_400_62400# 0.03fF
C610 VN.n493 a_400_62400# 1.28fF
C611 VN.n494 a_400_62400# 0.94fF
C612 VN.n495 a_400_62400# 1.05fF
C613 VN.n496 a_400_62400# 3.03fF
C614 VN.n497 a_400_62400# 2.51fF
C615 VN.n498 a_400_62400# 0.16fF
C616 VN.t1299 a_400_62400# 0.03fF
C617 VN.n499 a_400_62400# 0.19fF
C618 VN.t2418 a_400_62400# 0.03fF
C619 VN.n501 a_400_62400# 0.32fF
C620 VN.n502 a_400_62400# 0.48fF
C621 VN.n503 a_400_62400# 0.81fF
C622 VN.n504 a_400_62400# 1.86fF
C623 VN.n505 a_400_62400# 1.53fF
C624 VN.n506 a_400_62400# 0.47fF
C625 VN.n507 a_400_62400# 2.71fF
C626 VN.t1587 a_400_62400# 0.03fF
C627 VN.n508 a_400_62400# 0.32fF
C628 VN.n509 a_400_62400# 1.22fF
C629 VN.n510 a_400_62400# 0.07fF
C630 VN.t1363 a_400_62400# 0.03fF
C631 VN.n511 a_400_62400# 0.16fF
C632 VN.n512 a_400_62400# 0.19fF
C633 VN.n514 a_400_62400# 2.53fF
C634 VN.n515 a_400_62400# 2.51fF
C635 VN.t1556 a_400_62400# 0.03fF
C636 VN.n516 a_400_62400# 0.32fF
C637 VN.n517 a_400_62400# 0.48fF
C638 VN.n518 a_400_62400# 0.81fF
C639 VN.n519 a_400_62400# 0.16fF
C640 VN.t433 a_400_62400# 0.03fF
C641 VN.n520 a_400_62400# 0.19fF
C642 VN.n522 a_400_62400# 1.55fF
C643 VN.n523 a_400_62400# 0.29fF
C644 VN.n524 a_400_62400# 2.52fF
C645 VN.t722 a_400_62400# 0.03fF
C646 VN.n525 a_400_62400# 0.32fF
C647 VN.n526 a_400_62400# 1.22fF
C648 VN.n527 a_400_62400# 0.07fF
C649 VN.t615 a_400_62400# 0.03fF
C650 VN.n528 a_400_62400# 0.16fF
C651 VN.n529 a_400_62400# 0.19fF
C652 VN.n531 a_400_62400# 27.83fF
C653 VN.n532 a_400_62400# 3.93fF
C654 VN.n533 a_400_62400# 2.51fF
C655 VN.n534 a_400_62400# 0.16fF
C656 VN.t2080 a_400_62400# 0.03fF
C657 VN.n535 a_400_62400# 0.19fF
C658 VN.t685 a_400_62400# 0.03fF
C659 VN.n537 a_400_62400# 0.32fF
C660 VN.n538 a_400_62400# 0.48fF
C661 VN.n539 a_400_62400# 0.81fF
C662 VN.n540 a_400_62400# 1.46fF
C663 VN.n541 a_400_62400# 0.21fF
C664 VN.n542 a_400_62400# 2.81fF
C665 VN.t2267 a_400_62400# 0.03fF
C666 VN.n543 a_400_62400# 0.16fF
C667 VN.n544 a_400_62400# 0.19fF
C668 VN.t2376 a_400_62400# 0.03fF
C669 VN.n546 a_400_62400# 0.32fF
C670 VN.n547 a_400_62400# 1.22fF
C671 VN.n548 a_400_62400# 0.07fF
C672 VN.n549 a_400_62400# 2.51fF
C673 VN.n550 a_400_62400# 3.57fF
C674 VN.t2344 a_400_62400# 0.03fF
C675 VN.n551 a_400_62400# 0.32fF
C676 VN.n552 a_400_62400# 0.48fF
C677 VN.n553 a_400_62400# 0.81fF
C678 VN.n554 a_400_62400# 0.16fF
C679 VN.t1207 a_400_62400# 0.03fF
C680 VN.n555 a_400_62400# 0.19fF
C681 VN.n557 a_400_62400# 3.93fF
C682 VN.n558 a_400_62400# 3.08fF
C683 VN.t1403 a_400_62400# 0.03fF
C684 VN.n559 a_400_62400# 0.16fF
C685 VN.n560 a_400_62400# 0.19fF
C686 VN.t1509 a_400_62400# 0.03fF
C687 VN.n562 a_400_62400# 0.32fF
C688 VN.n563 a_400_62400# 1.22fF
C689 VN.n564 a_400_62400# 0.07fF
C690 VN.n565 a_400_62400# 2.51fF
C691 VN.n566 a_400_62400# 3.57fF
C692 VN.t302 a_400_62400# 0.03fF
C693 VN.n567 a_400_62400# 0.32fF
C694 VN.n568 a_400_62400# 0.48fF
C695 VN.n569 a_400_62400# 0.81fF
C696 VN.n570 a_400_62400# 0.16fF
C697 VN.t1677 a_400_62400# 0.03fF
C698 VN.n571 a_400_62400# 0.19fF
C699 VN.n573 a_400_62400# 3.75fF
C700 VN.n574 a_400_62400# 3.08fF
C701 VN.t1870 a_400_62400# 0.03fF
C702 VN.n575 a_400_62400# 0.16fF
C703 VN.n576 a_400_62400# 0.19fF
C704 VN.t1983 a_400_62400# 0.03fF
C705 VN.n578 a_400_62400# 0.32fF
C706 VN.n579 a_400_62400# 1.22fF
C707 VN.n580 a_400_62400# 0.07fF
C708 VN.n581 a_400_62400# 2.51fF
C709 VN.n582 a_400_62400# 3.57fF
C710 VN.t1950 a_400_62400# 0.03fF
C711 VN.n583 a_400_62400# 0.32fF
C712 VN.n584 a_400_62400# 0.48fF
C713 VN.n585 a_400_62400# 0.81fF
C714 VN.n586 a_400_62400# 0.16fF
C715 VN.t811 a_400_62400# 0.03fF
C716 VN.n587 a_400_62400# 0.19fF
C717 VN.n589 a_400_62400# 3.75fF
C718 VN.n590 a_400_62400# 3.08fF
C719 VN.t1000 a_400_62400# 0.03fF
C720 VN.n591 a_400_62400# 0.16fF
C721 VN.n592 a_400_62400# 0.19fF
C722 VN.t1110 a_400_62400# 0.03fF
C723 VN.n594 a_400_62400# 0.32fF
C724 VN.n595 a_400_62400# 1.22fF
C725 VN.n596 a_400_62400# 0.07fF
C726 VN.n597 a_400_62400# 2.51fF
C727 VN.n598 a_400_62400# 3.57fF
C728 VN.t1081 a_400_62400# 0.03fF
C729 VN.n599 a_400_62400# 0.32fF
C730 VN.n600 a_400_62400# 0.48fF
C731 VN.n601 a_400_62400# 0.81fF
C732 VN.n602 a_400_62400# 0.16fF
C733 VN.t2587 a_400_62400# 0.03fF
C734 VN.n603 a_400_62400# 0.19fF
C735 VN.n605 a_400_62400# 3.75fF
C736 VN.n606 a_400_62400# 3.08fF
C737 VN.t119 a_400_62400# 0.03fF
C738 VN.n607 a_400_62400# 0.16fF
C739 VN.n608 a_400_62400# 0.19fF
C740 VN.t246 a_400_62400# 0.03fF
C741 VN.n610 a_400_62400# 0.32fF
C742 VN.n611 a_400_62400# 1.22fF
C743 VN.n612 a_400_62400# 0.07fF
C744 VN.n613 a_400_62400# 2.51fF
C745 VN.n614 a_400_62400# 3.57fF
C746 VN.t349 a_400_62400# 0.03fF
C747 VN.n615 a_400_62400# 0.32fF
C748 VN.n616 a_400_62400# 0.48fF
C749 VN.n617 a_400_62400# 0.81fF
C750 VN.n618 a_400_62400# 0.16fF
C751 VN.t1717 a_400_62400# 0.03fF
C752 VN.n619 a_400_62400# 0.19fF
C753 VN.n621 a_400_62400# 3.75fF
C754 VN.n622 a_400_62400# 3.08fF
C755 VN.t1786 a_400_62400# 0.03fF
C756 VN.n623 a_400_62400# 0.16fF
C757 VN.n624 a_400_62400# 0.19fF
C758 VN.t2037 a_400_62400# 0.03fF
C759 VN.n626 a_400_62400# 0.32fF
C760 VN.n627 a_400_62400# 1.22fF
C761 VN.n628 a_400_62400# 0.07fF
C762 VN.n629 a_400_62400# 2.51fF
C763 VN.n630 a_400_62400# 3.57fF
C764 VN.t1993 a_400_62400# 0.03fF
C765 VN.n631 a_400_62400# 0.32fF
C766 VN.n632 a_400_62400# 0.48fF
C767 VN.n633 a_400_62400# 0.81fF
C768 VN.n634 a_400_62400# 0.16fF
C769 VN.t844 a_400_62400# 0.03fF
C770 VN.n635 a_400_62400# 0.19fF
C771 VN.n637 a_400_62400# 3.75fF
C772 VN.n638 a_400_62400# 3.08fF
C773 VN.t909 a_400_62400# 0.03fF
C774 VN.n639 a_400_62400# 0.16fF
C775 VN.n640 a_400_62400# 0.19fF
C776 VN.t1164 a_400_62400# 0.03fF
C777 VN.n642 a_400_62400# 0.32fF
C778 VN.n643 a_400_62400# 1.22fF
C779 VN.n644 a_400_62400# 0.07fF
C780 VN.n645 a_400_62400# 2.51fF
C781 VN.n646 a_400_62400# 3.57fF
C782 VN.t1120 a_400_62400# 0.03fF
C783 VN.n647 a_400_62400# 0.32fF
C784 VN.n648 a_400_62400# 0.48fF
C785 VN.n649 a_400_62400# 0.81fF
C786 VN.n650 a_400_62400# 0.16fF
C787 VN.t2508 a_400_62400# 0.03fF
C788 VN.n651 a_400_62400# 0.19fF
C789 VN.n653 a_400_62400# 3.75fF
C790 VN.n654 a_400_62400# 3.08fF
C791 VN.t2571 a_400_62400# 0.03fF
C792 VN.n655 a_400_62400# 0.16fF
C793 VN.n656 a_400_62400# 0.19fF
C794 VN.t295 a_400_62400# 0.03fF
C795 VN.n658 a_400_62400# 0.32fF
C796 VN.n659 a_400_62400# 1.22fF
C797 VN.n660 a_400_62400# 0.07fF
C798 VN.n661 a_400_62400# 2.51fF
C799 VN.n662 a_400_62400# 3.57fF
C800 VN.t258 a_400_62400# 0.03fF
C801 VN.n663 a_400_62400# 0.32fF
C802 VN.n664 a_400_62400# 0.48fF
C803 VN.n665 a_400_62400# 0.81fF
C804 VN.n666 a_400_62400# 0.16fF
C805 VN.t1646 a_400_62400# 0.03fF
C806 VN.n667 a_400_62400# 0.19fF
C807 VN.n669 a_400_62400# 3.75fF
C808 VN.n670 a_400_62400# 3.08fF
C809 VN.t1700 a_400_62400# 0.03fF
C810 VN.n671 a_400_62400# 0.16fF
C811 VN.n672 a_400_62400# 0.19fF
C812 VN.t1946 a_400_62400# 0.03fF
C813 VN.n674 a_400_62400# 0.32fF
C814 VN.n675 a_400_62400# 1.22fF
C815 VN.n676 a_400_62400# 0.07fF
C816 VN.n677 a_400_62400# 2.51fF
C817 VN.n678 a_400_62400# 3.57fF
C818 VN.t1906 a_400_62400# 0.03fF
C819 VN.n679 a_400_62400# 0.32fF
C820 VN.n680 a_400_62400# 0.48fF
C821 VN.n681 a_400_62400# 0.81fF
C822 VN.n682 a_400_62400# 0.16fF
C823 VN.t775 a_400_62400# 0.03fF
C824 VN.n683 a_400_62400# 0.19fF
C825 VN.n685 a_400_62400# 3.75fF
C826 VN.n686 a_400_62400# 3.08fF
C827 VN.t955 a_400_62400# 0.03fF
C828 VN.n687 a_400_62400# 0.16fF
C829 VN.n688 a_400_62400# 0.19fF
C830 VN.t1076 a_400_62400# 0.03fF
C831 VN.n690 a_400_62400# 0.32fF
C832 VN.n691 a_400_62400# 1.22fF
C833 VN.n692 a_400_62400# 0.07fF
C834 VN.n693 a_400_62400# 2.51fF
C835 VN.n694 a_400_62400# 3.57fF
C836 VN.t1032 a_400_62400# 0.03fF
C837 VN.n695 a_400_62400# 0.32fF
C838 VN.n696 a_400_62400# 0.48fF
C839 VN.n697 a_400_62400# 0.81fF
C840 VN.n698 a_400_62400# 0.16fF
C841 VN.t2425 a_400_62400# 0.03fF
C842 VN.n699 a_400_62400# 0.19fF
C843 VN.n701 a_400_62400# 3.75fF
C844 VN.n702 a_400_62400# 3.08fF
C845 VN.t42 a_400_62400# 0.03fF
C846 VN.n703 a_400_62400# 0.16fF
C847 VN.n704 a_400_62400# 0.19fF
C848 VN.t202 a_400_62400# 0.03fF
C849 VN.n706 a_400_62400# 0.32fF
C850 VN.n707 a_400_62400# 1.22fF
C851 VN.n708 a_400_62400# 0.07fF
C852 VN.n709 a_400_62400# 2.51fF
C853 VN.n710 a_400_62400# 3.57fF
C854 VN.t2180 a_400_62400# 0.03fF
C855 VN.n711 a_400_62400# 0.32fF
C856 VN.n712 a_400_62400# 0.48fF
C857 VN.n713 a_400_62400# 0.81fF
C858 VN.n714 a_400_62400# 0.16fF
C859 VN.t1010 a_400_62400# 0.03fF
C860 VN.n715 a_400_62400# 0.19fF
C861 VN.n717 a_400_62400# 3.75fF
C862 VN.n718 a_400_62400# 3.08fF
C863 VN.t1220 a_400_62400# 0.03fF
C864 VN.n719 a_400_62400# 0.16fF
C865 VN.n720 a_400_62400# 0.19fF
C866 VN.t1441 a_400_62400# 0.03fF
C867 VN.n722 a_400_62400# 0.32fF
C868 VN.n723 a_400_62400# 1.22fF
C869 VN.n724 a_400_62400# 0.07fF
C870 VN.n725 a_400_62400# 2.51fF
C871 VN.n726 a_400_62400# 3.57fF
C872 VN.t1312 a_400_62400# 0.03fF
C873 VN.n727 a_400_62400# 0.32fF
C874 VN.n728 a_400_62400# 0.48fF
C875 VN.n729 a_400_62400# 0.81fF
C876 VN.n730 a_400_62400# 0.16fF
C877 VN.t136 a_400_62400# 0.03fF
C878 VN.n731 a_400_62400# 0.19fF
C879 VN.n733 a_400_62400# 3.75fF
C880 VN.n734 a_400_62400# 3.08fF
C881 VN.t357 a_400_62400# 0.03fF
C882 VN.n735 a_400_62400# 0.16fF
C883 VN.n736 a_400_62400# 0.19fF
C884 VN.t573 a_400_62400# 0.03fF
C885 VN.n738 a_400_62400# 0.32fF
C886 VN.n739 a_400_62400# 1.22fF
C887 VN.n740 a_400_62400# 0.07fF
C888 VN.n741 a_400_62400# 0.16fF
C889 VN.t1057 a_400_62400# 0.03fF
C890 VN.n742 a_400_62400# 0.19fF
C891 VN.t2097 a_400_62400# 0.03fF
C892 VN.n744 a_400_62400# 0.32fF
C893 VN.n745 a_400_62400# 0.48fF
C894 VN.n746 a_400_62400# 0.81fF
C895 VN.n747 a_400_62400# 2.14fF
C896 VN.n748 a_400_62400# 0.19fF
C897 VN.n749 a_400_62400# 0.78fF
C898 VN.n750 a_400_62400# 0.71fF
C899 VN.n751 a_400_62400# 0.55fF
C900 VN.n752 a_400_62400# 0.33fF
C901 VN.n753 a_400_62400# 0.33fF
C902 VN.n754 a_400_62400# 0.91fF
C903 VN.n755 a_400_62400# 2.64fF
C904 VN.t1128 a_400_62400# 0.03fF
C905 VN.n756 a_400_62400# 0.16fF
C906 VN.n757 a_400_62400# 0.19fF
C907 VN.t1366 a_400_62400# 0.03fF
C908 VN.n759 a_400_62400# 0.32fF
C909 VN.n760 a_400_62400# 1.22fF
C910 VN.n761 a_400_62400# 0.07fF
C911 VN.t41 a_400_62400# 64.69fF
C912 VN.t2231 a_400_62400# 0.03fF
C913 VN.n762 a_400_62400# 0.32fF
C914 VN.n763 a_400_62400# 1.22fF
C915 VN.n764 a_400_62400# 0.07fF
C916 VN.t2002 a_400_62400# 0.03fF
C917 VN.n765 a_400_62400# 0.16fF
C918 VN.n766 a_400_62400# 0.19fF
C919 VN.n768 a_400_62400# 0.16fF
C920 VN.t1799 a_400_62400# 0.03fF
C921 VN.n769 a_400_62400# 0.19fF
C922 VN.n771 a_400_62400# 6.92fF
C923 VN.n772 a_400_62400# 6.56fF
C924 VN.t1099 a_400_62400# 0.03fF
C925 VN.n773 a_400_62400# 0.16fF
C926 VN.n774 a_400_62400# 0.19fF
C927 VN.t628 a_400_62400# 0.03fF
C928 VN.n776 a_400_62400# 0.32fF
C929 VN.n777 a_400_62400# 1.22fF
C930 VN.n778 a_400_62400# 0.07fF
C931 VN.n779 a_400_62400# 0.04fF
C932 VN.n780 a_400_62400# 0.16fF
C933 VN.n781 a_400_62400# 0.14fF
C934 VN.n782 a_400_62400# 0.48fF
C935 VN.n783 a_400_62400# 0.62fF
C936 VN.n784 a_400_62400# 1.52fF
C937 VN.n785 a_400_62400# 2.51fF
C938 VN.n786 a_400_62400# 0.16fF
C939 VN.t2095 a_400_62400# 0.03fF
C940 VN.n787 a_400_62400# 0.19fF
C941 VN.t711 a_400_62400# 0.03fF
C942 VN.n789 a_400_62400# 0.32fF
C943 VN.n790 a_400_62400# 0.48fF
C944 VN.n791 a_400_62400# 0.81fF
C945 VN.n792 a_400_62400# 1.70fF
C946 VN.n793 a_400_62400# 3.19fF
C947 VN.n794 a_400_62400# 5.63fF
C948 VN.t232 a_400_62400# 0.03fF
C949 VN.n795 a_400_62400# 0.16fF
C950 VN.n796 a_400_62400# 0.19fF
C951 VN.t2282 a_400_62400# 0.03fF
C952 VN.n798 a_400_62400# 0.32fF
C953 VN.n799 a_400_62400# 1.22fF
C954 VN.n800 a_400_62400# 0.07fF
C955 VN.t12 a_400_62400# 64.17fF
C956 VN.t1413 a_400_62400# 0.03fF
C957 VN.n801 a_400_62400# 1.60fF
C958 VN.n802 a_400_62400# 0.07fF
C959 VN.t2019 a_400_62400# 0.03fF
C960 VN.n803 a_400_62400# 0.02fF
C961 VN.n804 a_400_62400# 0.34fF
C962 VN.n806 a_400_62400# 0.79fF
C963 VN.n807 a_400_62400# 0.23fF
C964 VN.n808 a_400_62400# 1.18fF
C965 VN.t2 a_400_62400# 28.64fF
C966 VN.n809 a_400_62400# 0.79fF
C967 VN.n810 a_400_62400# 0.11fF
C968 VN.n811 a_400_62400# 4.98fF
C969 VN.n812 a_400_62400# 0.80fF
C970 VN.n813 a_400_62400# 0.29fF
C971 VN.n814 a_400_62400# 1.96fF
C972 VN.n816 a_400_62400# 25.18fF
C973 VN.n818 a_400_62400# 1.87fF
C974 VN.n819 a_400_62400# 5.71fF
C975 VN.n820 a_400_62400# 3.66fF
C976 VN.n821 a_400_62400# 6.25fF
C977 VN.n822 a_400_62400# 0.02fF
C978 VN.n823 a_400_62400# 0.04fF
C979 VN.n824 a_400_62400# 0.32fF
C980 VN.n825 a_400_62400# 0.17fF
C981 VN.n826 a_400_62400# 0.75fF
C982 VN.n827 a_400_62400# 0.04fF
C983 VN.n828 a_400_62400# 1.15fF
C984 VN.n829 a_400_62400# 0.30fF
C985 VN.n830 a_400_62400# 0.20fF
C986 VN.n831 a_400_62400# 37.46fF
C987 VN.n832 a_400_62400# 37.46fF
C988 VN.n833 a_400_62400# 0.79fF
C989 VN.n834 a_400_62400# 0.23fF
C990 VN.n835 a_400_62400# 1.18fF
C991 VN.t201 a_400_62400# 28.64fF
C992 VN.n836 a_400_62400# 0.79fF
C993 VN.n837 a_400_62400# 0.11fF
C994 VN.n838 a_400_62400# 4.98fF
C995 VN.n839 a_400_62400# 0.80fF
C996 VN.n840 a_400_62400# 0.29fF
C997 VN.n841 a_400_62400# 1.96fF
C998 VN.n843 a_400_62400# 25.18fF
C999 VN.n845 a_400_62400# 1.87fF
C1000 VN.n846 a_400_62400# 5.36fF
C1001 VN.n847 a_400_62400# 1.52fF
C1002 VN.t679 a_400_62400# 0.03fF
C1003 VN.n848 a_400_62400# 0.85fF
C1004 VN.n849 a_400_62400# 0.81fF
C1005 VN.n850 a_400_62400# 0.33fF
C1006 VN.n851 a_400_62400# 0.12fF
C1007 VN.n852 a_400_62400# 0.28fF
C1008 VN.n853 a_400_62400# 1.72fF
C1009 VN.n854 a_400_62400# 0.71fF
C1010 VN.n855 a_400_62400# 2.51fF
C1011 VN.n856 a_400_62400# 0.16fF
C1012 VN.t2305 a_400_62400# 0.03fF
C1013 VN.n857 a_400_62400# 0.19fF
C1014 VN.t787 a_400_62400# 0.03fF
C1015 VN.n859 a_400_62400# 0.32fF
C1016 VN.n860 a_400_62400# 0.48fF
C1017 VN.n861 a_400_62400# 0.81fF
C1018 VN.n862 a_400_62400# 0.95fF
C1019 VN.n863 a_400_62400# 2.11fF
C1020 VN.n864 a_400_62400# 3.28fF
C1021 VN.t1901 a_400_62400# 0.03fF
C1022 VN.n865 a_400_62400# 0.32fF
C1023 VN.n866 a_400_62400# 1.22fF
C1024 VN.n867 a_400_62400# 0.07fF
C1025 VN.t467 a_400_62400# 0.03fF
C1026 VN.n868 a_400_62400# 0.16fF
C1027 VN.n869 a_400_62400# 0.19fF
C1028 VN.n871 a_400_62400# 2.53fF
C1029 VN.n872 a_400_62400# 0.08fF
C1030 VN.n873 a_400_62400# 0.04fF
C1031 VN.n874 a_400_62400# 0.05fF
C1032 VN.n875 a_400_62400# 1.33fF
C1033 VN.n876 a_400_62400# 0.03fF
C1034 VN.n877 a_400_62400# 0.01fF
C1035 VN.n878 a_400_62400# 0.02fF
C1036 VN.n879 a_400_62400# 0.11fF
C1037 VN.n880 a_400_62400# 0.48fF
C1038 VN.n881 a_400_62400# 2.48fF
C1039 VN.t2562 a_400_62400# 0.03fF
C1040 VN.n882 a_400_62400# 0.32fF
C1041 VN.n883 a_400_62400# 0.48fF
C1042 VN.n884 a_400_62400# 0.81fF
C1043 VN.n885 a_400_62400# 0.16fF
C1044 VN.t1433 a_400_62400# 0.03fF
C1045 VN.n886 a_400_62400# 0.19fF
C1046 VN.n888 a_400_62400# 0.93fF
C1047 VN.n889 a_400_62400# 0.30fF
C1048 VN.n890 a_400_62400# 0.34fF
C1049 VN.n891 a_400_62400# 0.12fF
C1050 VN.n892 a_400_62400# 0.30fF
C1051 VN.n893 a_400_62400# 0.93fF
C1052 VN.n894 a_400_62400# 1.55fF
C1053 VN.n895 a_400_62400# 0.29fF
C1054 VN.n896 a_400_62400# 0.34fF
C1055 VN.n897 a_400_62400# 0.12fF
C1056 VN.n898 a_400_62400# 2.52fF
C1057 VN.t1172 a_400_62400# 0.03fF
C1058 VN.n899 a_400_62400# 0.32fF
C1059 VN.n900 a_400_62400# 1.22fF
C1060 VN.n901 a_400_62400# 0.07fF
C1061 VN.t2117 a_400_62400# 0.03fF
C1062 VN.n902 a_400_62400# 0.16fF
C1063 VN.n903 a_400_62400# 0.19fF
C1064 VN.n905 a_400_62400# 27.83fF
C1065 VN.n906 a_400_62400# 3.19fF
C1066 VN.n907 a_400_62400# 0.61fF
C1067 VN.n908 a_400_62400# 0.30fF
C1068 VN.n909 a_400_62400# 0.51fF
C1069 VN.n910 a_400_62400# 0.21fF
C1070 VN.n911 a_400_62400# 0.38fF
C1071 VN.n912 a_400_62400# 0.29fF
C1072 VN.n913 a_400_62400# 0.40fF
C1073 VN.n914 a_400_62400# 0.28fF
C1074 VN.t1656 a_400_62400# 0.03fF
C1075 VN.n915 a_400_62400# 0.32fF
C1076 VN.n916 a_400_62400# 0.48fF
C1077 VN.n917 a_400_62400# 0.81fF
C1078 VN.n918 a_400_62400# 0.16fF
C1079 VN.t531 a_400_62400# 0.03fF
C1080 VN.n919 a_400_62400# 0.19fF
C1081 VN.n921 a_400_62400# 0.25fF
C1082 VN.n922 a_400_62400# 2.11fF
C1083 VN.n923 a_400_62400# 2.96fF
C1084 VN.n924 a_400_62400# 0.43fF
C1085 VN.n925 a_400_62400# 3.20fF
C1086 VN.t1330 a_400_62400# 0.03fF
C1087 VN.n926 a_400_62400# 0.16fF
C1088 VN.n927 a_400_62400# 0.19fF
C1089 VN.t251 a_400_62400# 0.03fF
C1090 VN.n929 a_400_62400# 0.32fF
C1091 VN.n930 a_400_62400# 1.22fF
C1092 VN.n931 a_400_62400# 0.07fF
C1093 VN.n932 a_400_62400# 2.51fF
C1094 VN.n933 a_400_62400# 0.16fF
C1095 VN.t567 a_400_62400# 0.03fF
C1096 VN.n934 a_400_62400# 0.19fF
C1097 VN.t1692 a_400_62400# 0.03fF
C1098 VN.n936 a_400_62400# 0.32fF
C1099 VN.n937 a_400_62400# 0.48fF
C1100 VN.n938 a_400_62400# 0.81fF
C1101 VN.n939 a_400_62400# 1.24fF
C1102 VN.n940 a_400_62400# 0.43fF
C1103 VN.n941 a_400_62400# 0.43fF
C1104 VN.n942 a_400_62400# 1.24fF
C1105 VN.n943 a_400_62400# 1.46fF
C1106 VN.n944 a_400_62400# 0.21fF
C1107 VN.n945 a_400_62400# 6.64fF
C1108 VN.t1240 a_400_62400# 0.03fF
C1109 VN.n946 a_400_62400# 0.16fF
C1110 VN.n947 a_400_62400# 0.19fF
C1111 VN.t303 a_400_62400# 0.03fF
C1112 VN.n949 a_400_62400# 0.32fF
C1113 VN.n950 a_400_62400# 1.22fF
C1114 VN.n951 a_400_62400# 0.07fF
C1115 VN.n952 a_400_62400# 2.51fF
C1116 VN.n953 a_400_62400# 3.57fF
C1117 VN.t2194 a_400_62400# 0.03fF
C1118 VN.n954 a_400_62400# 0.32fF
C1119 VN.n955 a_400_62400# 0.48fF
C1120 VN.n956 a_400_62400# 0.81fF
C1121 VN.n957 a_400_62400# 0.16fF
C1122 VN.t1028 a_400_62400# 0.03fF
C1123 VN.n958 a_400_62400# 0.19fF
C1124 VN.n960 a_400_62400# 6.91fF
C1125 VN.t375 a_400_62400# 0.03fF
C1126 VN.n961 a_400_62400# 0.16fF
C1127 VN.n962 a_400_62400# 0.19fF
C1128 VN.t778 a_400_62400# 0.03fF
C1129 VN.n964 a_400_62400# 0.32fF
C1130 VN.n965 a_400_62400# 1.22fF
C1131 VN.n966 a_400_62400# 0.07fF
C1132 VN.n967 a_400_62400# 2.51fF
C1133 VN.n968 a_400_62400# 3.57fF
C1134 VN.t1324 a_400_62400# 0.03fF
C1135 VN.n969 a_400_62400# 0.32fF
C1136 VN.n970 a_400_62400# 0.48fF
C1137 VN.n971 a_400_62400# 0.81fF
C1138 VN.n972 a_400_62400# 0.16fF
C1139 VN.t157 a_400_62400# 0.03fF
C1140 VN.n973 a_400_62400# 0.19fF
C1141 VN.n975 a_400_62400# 6.92fF
C1142 VN.t834 a_400_62400# 0.03fF
C1143 VN.n976 a_400_62400# 0.16fF
C1144 VN.n977 a_400_62400# 0.19fF
C1145 VN.t2427 a_400_62400# 0.03fF
C1146 VN.n979 a_400_62400# 0.32fF
C1147 VN.n980 a_400_62400# 1.22fF
C1148 VN.n981 a_400_62400# 0.07fF
C1149 VN.n982 a_400_62400# 2.51fF
C1150 VN.n983 a_400_62400# 3.57fF
C1151 VN.t462 a_400_62400# 0.03fF
C1152 VN.n984 a_400_62400# 0.32fF
C1153 VN.n985 a_400_62400# 0.48fF
C1154 VN.n986 a_400_62400# 0.81fF
C1155 VN.n987 a_400_62400# 0.16fF
C1156 VN.t1820 a_400_62400# 0.03fF
C1157 VN.n988 a_400_62400# 0.19fF
C1158 VN.n990 a_400_62400# 6.92fF
C1159 VN.t2497 a_400_62400# 0.03fF
C1160 VN.n991 a_400_62400# 0.16fF
C1161 VN.n992 a_400_62400# 0.19fF
C1162 VN.t1565 a_400_62400# 0.03fF
C1163 VN.n994 a_400_62400# 0.32fF
C1164 VN.n995 a_400_62400# 1.22fF
C1165 VN.n996 a_400_62400# 0.07fF
C1166 VN.n997 a_400_62400# 2.51fF
C1167 VN.n998 a_400_62400# 3.57fF
C1168 VN.t2111 a_400_62400# 0.03fF
C1169 VN.n999 a_400_62400# 0.32fF
C1170 VN.n1000 a_400_62400# 0.48fF
C1171 VN.n1001 a_400_62400# 0.81fF
C1172 VN.n1002 a_400_62400# 0.16fF
C1173 VN.t947 a_400_62400# 0.03fF
C1174 VN.n1003 a_400_62400# 0.19fF
C1175 VN.n1005 a_400_62400# 6.92fF
C1176 VN.t1752 a_400_62400# 0.03fF
C1177 VN.n1006 a_400_62400# 0.16fF
C1178 VN.n1007 a_400_62400# 0.19fF
C1179 VN.t695 a_400_62400# 0.03fF
C1180 VN.n1009 a_400_62400# 0.32fF
C1181 VN.n1010 a_400_62400# 1.22fF
C1182 VN.n1011 a_400_62400# 0.07fF
C1183 VN.n1012 a_400_62400# 2.51fF
C1184 VN.n1013 a_400_62400# 3.57fF
C1185 VN.t1234 a_400_62400# 0.03fF
C1186 VN.n1014 a_400_62400# 0.32fF
C1187 VN.n1015 a_400_62400# 0.48fF
C1188 VN.n1016 a_400_62400# 0.81fF
C1189 VN.n1017 a_400_62400# 0.16fF
C1190 VN.t25 a_400_62400# 0.03fF
C1191 VN.n1018 a_400_62400# 0.19fF
C1192 VN.n1020 a_400_62400# 6.92fF
C1193 VN.t878 a_400_62400# 0.03fF
C1194 VN.n1021 a_400_62400# 0.16fF
C1195 VN.n1022 a_400_62400# 0.19fF
C1196 VN.t2354 a_400_62400# 0.03fF
C1197 VN.n1024 a_400_62400# 0.32fF
C1198 VN.n1025 a_400_62400# 1.22fF
C1199 VN.n1026 a_400_62400# 0.07fF
C1200 VN.n1027 a_400_62400# 2.51fF
C1201 VN.n1028 a_400_62400# 3.57fF
C1202 VN.t370 a_400_62400# 0.03fF
C1203 VN.n1029 a_400_62400# 0.32fF
C1204 VN.n1030 a_400_62400# 0.48fF
C1205 VN.n1031 a_400_62400# 0.81fF
C1206 VN.n1032 a_400_62400# 0.16fF
C1207 VN.t1736 a_400_62400# 0.03fF
C1208 VN.n1033 a_400_62400# 0.19fF
C1209 VN.n1035 a_400_62400# 6.92fF
C1210 VN.t2538 a_400_62400# 0.03fF
C1211 VN.n1036 a_400_62400# 0.16fF
C1212 VN.n1037 a_400_62400# 0.19fF
C1213 VN.t1486 a_400_62400# 0.03fF
C1214 VN.n1039 a_400_62400# 0.32fF
C1215 VN.n1040 a_400_62400# 1.22fF
C1216 VN.n1041 a_400_62400# 0.07fF
C1217 VN.n1042 a_400_62400# 2.51fF
C1218 VN.n1043 a_400_62400# 3.57fF
C1219 VN.t2022 a_400_62400# 0.03fF
C1220 VN.n1044 a_400_62400# 0.32fF
C1221 VN.n1045 a_400_62400# 0.48fF
C1222 VN.n1046 a_400_62400# 0.81fF
C1223 VN.n1047 a_400_62400# 0.16fF
C1224 VN.t863 a_400_62400# 0.03fF
C1225 VN.n1048 a_400_62400# 0.19fF
C1226 VN.n1050 a_400_62400# 6.92fF
C1227 VN.t1673 a_400_62400# 0.03fF
C1228 VN.n1051 a_400_62400# 0.16fF
C1229 VN.n1052 a_400_62400# 0.19fF
C1230 VN.t619 a_400_62400# 0.03fF
C1231 VN.n1054 a_400_62400# 0.32fF
C1232 VN.n1055 a_400_62400# 1.22fF
C1233 VN.n1056 a_400_62400# 0.07fF
C1234 VN.n1057 a_400_62400# 2.51fF
C1235 VN.n1058 a_400_62400# 3.57fF
C1236 VN.t1148 a_400_62400# 0.03fF
C1237 VN.n1059 a_400_62400# 0.32fF
C1238 VN.n1060 a_400_62400# 0.48fF
C1239 VN.n1061 a_400_62400# 0.81fF
C1240 VN.n1062 a_400_62400# 0.16fF
C1241 VN.t113 a_400_62400# 0.03fF
C1242 VN.n1063 a_400_62400# 0.19fF
C1243 VN.n1065 a_400_62400# 6.92fF
C1244 VN.t806 a_400_62400# 0.03fF
C1245 VN.n1066 a_400_62400# 0.16fF
C1246 VN.n1067 a_400_62400# 0.19fF
C1247 VN.t2271 a_400_62400# 0.03fF
C1248 VN.n1069 a_400_62400# 0.32fF
C1249 VN.n1070 a_400_62400# 1.22fF
C1250 VN.n1071 a_400_62400# 0.07fF
C1251 VN.n1072 a_400_62400# 2.51fF
C1252 VN.n1073 a_400_62400# 3.57fF
C1253 VN.t422 a_400_62400# 0.03fF
C1254 VN.n1074 a_400_62400# 0.32fF
C1255 VN.n1075 a_400_62400# 0.48fF
C1256 VN.n1076 a_400_62400# 0.81fF
C1257 VN.n1077 a_400_62400# 0.16fF
C1258 VN.t1781 a_400_62400# 0.03fF
C1259 VN.n1078 a_400_62400# 0.19fF
C1260 VN.n1080 a_400_62400# 6.92fF
C1261 VN.t2460 a_400_62400# 0.03fF
C1262 VN.n1081 a_400_62400# 0.16fF
C1263 VN.n1082 a_400_62400# 0.19fF
C1264 VN.t1530 a_400_62400# 0.03fF
C1265 VN.n1084 a_400_62400# 0.32fF
C1266 VN.n1085 a_400_62400# 1.22fF
C1267 VN.n1086 a_400_62400# 0.07fF
C1268 VN.n1087 a_400_62400# 2.51fF
C1269 VN.n1088 a_400_62400# 3.57fF
C1270 VN.t1630 a_400_62400# 0.03fF
C1271 VN.n1089 a_400_62400# 0.32fF
C1272 VN.n1090 a_400_62400# 0.48fF
C1273 VN.n1091 a_400_62400# 0.81fF
C1274 VN.n1092 a_400_62400# 0.16fF
C1275 VN.t496 a_400_62400# 0.03fF
C1276 VN.n1093 a_400_62400# 0.19fF
C1277 VN.n1095 a_400_62400# 6.92fF
C1278 VN.t1595 a_400_62400# 0.03fF
C1279 VN.n1096 a_400_62400# 0.16fF
C1280 VN.n1097 a_400_62400# 0.19fF
C1281 VN.t677 a_400_62400# 0.03fF
C1282 VN.n1099 a_400_62400# 0.32fF
C1283 VN.n1100 a_400_62400# 1.22fF
C1284 VN.n1101 a_400_62400# 0.07fF
C1285 VN.n1102 a_400_62400# 2.51fF
C1286 VN.n1103 a_400_62400# 3.57fF
C1287 VN.t757 a_400_62400# 0.03fF
C1288 VN.n1104 a_400_62400# 0.32fF
C1289 VN.n1105 a_400_62400# 0.48fF
C1290 VN.n1106 a_400_62400# 0.81fF
C1291 VN.n1107 a_400_62400# 0.16fF
C1292 VN.t2153 a_400_62400# 0.03fF
C1293 VN.n1108 a_400_62400# 0.19fF
C1294 VN.n1110 a_400_62400# 6.92fF
C1295 VN.t291 a_400_62400# 0.03fF
C1296 VN.n1111 a_400_62400# 0.16fF
C1297 VN.n1112 a_400_62400# 0.19fF
C1298 VN.t2338 a_400_62400# 0.03fF
C1299 VN.n1114 a_400_62400# 0.32fF
C1300 VN.n1115 a_400_62400# 1.22fF
C1301 VN.n1116 a_400_62400# 0.07fF
C1302 VN.n1117 a_400_62400# 2.51fF
C1303 VN.n1118 a_400_62400# 3.57fF
C1304 VN.t2415 a_400_62400# 0.03fF
C1305 VN.n1119 a_400_62400# 0.32fF
C1306 VN.n1120 a_400_62400# 0.48fF
C1307 VN.n1121 a_400_62400# 0.81fF
C1308 VN.n1122 a_400_62400# 0.16fF
C1309 VN.t1284 a_400_62400# 0.03fF
C1310 VN.n1123 a_400_62400# 0.19fF
C1311 VN.n1125 a_400_62400# 2.51fF
C1312 VN.n1126 a_400_62400# 3.59fF
C1313 VN.t1286 a_400_62400# 0.03fF
C1314 VN.n1127 a_400_62400# 0.32fF
C1315 VN.n1128 a_400_62400# 0.48fF
C1316 VN.n1129 a_400_62400# 0.81fF
C1317 VN.t1043 a_400_62400# 0.03fF
C1318 VN.n1130 a_400_62400# 1.63fF
C1319 VN.n1131 a_400_62400# 0.81fF
C1320 VN.n1132 a_400_62400# 1.21fF
C1321 VN.n1133 a_400_62400# 1.54fF
C1322 VN.n1134 a_400_62400# 4.06fF
C1323 VN.t53 a_400_62400# 28.64fF
C1324 VN.n1135 a_400_62400# 28.43fF
C1325 VN.n1137 a_400_62400# 0.50fF
C1326 VN.n1138 a_400_62400# 0.31fF
C1327 VN.n1139 a_400_62400# 3.87fF
C1328 VN.n1140 a_400_62400# 3.29fF
C1329 VN.n1141 a_400_62400# 3.38fF
C1330 VN.n1142 a_400_62400# 5.28fF
C1331 VN.n1143 a_400_62400# 0.34fF
C1332 VN.n1144 a_400_62400# 0.02fF
C1333 VN.t2432 a_400_62400# 0.03fF
C1334 VN.n1145 a_400_62400# 0.34fF
C1335 VN.t215 a_400_62400# 0.03fF
C1336 VN.n1146 a_400_62400# 1.28fF
C1337 VN.n1147 a_400_62400# 0.94fF
C1338 VN.n1148 a_400_62400# 2.51fF
C1339 VN.n1149 a_400_62400# 0.56fF
C1340 VN.n1150 a_400_62400# 0.64fF
C1341 VN.n1151 a_400_62400# 0.12fF
C1342 VN.n1152 a_400_62400# 0.44fF
C1343 VN.n1153 a_400_62400# 0.40fF
C1344 VN.n1154 a_400_62400# 1.03fF
C1345 VN.n1155 a_400_62400# 0.79fF
C1346 VN.t174 a_400_62400# 0.03fF
C1347 VN.n1156 a_400_62400# 0.32fF
C1348 VN.n1157 a_400_62400# 0.48fF
C1349 VN.n1158 a_400_62400# 0.81fF
C1350 VN.n1159 a_400_62400# 0.16fF
C1351 VN.t1572 a_400_62400# 0.03fF
C1352 VN.n1160 a_400_62400# 0.19fF
C1353 VN.n1162 a_400_62400# 1.93fF
C1354 VN.n1163 a_400_62400# 2.89fF
C1355 VN.t1865 a_400_62400# 0.03fF
C1356 VN.n1164 a_400_62400# 0.32fF
C1357 VN.n1165 a_400_62400# 1.22fF
C1358 VN.n1166 a_400_62400# 0.07fF
C1359 VN.t1639 a_400_62400# 0.03fF
C1360 VN.n1167 a_400_62400# 0.16fF
C1361 VN.n1168 a_400_62400# 0.19fF
C1362 VN.n1170 a_400_62400# 1.05fF
C1363 VN.n1171 a_400_62400# 3.07fF
C1364 VN.n1172 a_400_62400# 2.51fF
C1365 VN.n1173 a_400_62400# 0.16fF
C1366 VN.t702 a_400_62400# 0.03fF
C1367 VN.n1174 a_400_62400# 0.19fF
C1368 VN.t1836 a_400_62400# 0.03fF
C1369 VN.n1176 a_400_62400# 0.32fF
C1370 VN.n1177 a_400_62400# 0.48fF
C1371 VN.n1178 a_400_62400# 0.81fF
C1372 VN.n1179 a_400_62400# 1.86fF
C1373 VN.n1180 a_400_62400# 1.53fF
C1374 VN.n1181 a_400_62400# 0.47fF
C1375 VN.n1182 a_400_62400# 2.71fF
C1376 VN.t995 a_400_62400# 0.03fF
C1377 VN.n1183 a_400_62400# 0.32fF
C1378 VN.n1184 a_400_62400# 1.22fF
C1379 VN.n1185 a_400_62400# 0.07fF
C1380 VN.t882 a_400_62400# 0.03fF
C1381 VN.n1186 a_400_62400# 0.16fF
C1382 VN.n1187 a_400_62400# 0.19fF
C1383 VN.n1189 a_400_62400# 2.53fF
C1384 VN.n1190 a_400_62400# 2.51fF
C1385 VN.t961 a_400_62400# 0.03fF
C1386 VN.n1191 a_400_62400# 0.32fF
C1387 VN.n1192 a_400_62400# 0.48fF
C1388 VN.n1193 a_400_62400# 0.81fF
C1389 VN.n1194 a_400_62400# 0.16fF
C1390 VN.t2361 a_400_62400# 0.03fF
C1391 VN.n1195 a_400_62400# 0.19fF
C1392 VN.n1197 a_400_62400# 1.55fF
C1393 VN.n1198 a_400_62400# 0.29fF
C1394 VN.n1199 a_400_62400# 2.52fF
C1395 VN.t115 a_400_62400# 0.03fF
C1396 VN.n1200 a_400_62400# 0.32fF
C1397 VN.n1201 a_400_62400# 1.22fF
C1398 VN.n1202 a_400_62400# 0.07fF
C1399 VN.t2542 a_400_62400# 0.03fF
C1400 VN.n1203 a_400_62400# 0.16fF
C1401 VN.n1204 a_400_62400# 0.19fF
C1402 VN.n1206 a_400_62400# 27.83fF
C1403 VN.n1207 a_400_62400# 3.93fF
C1404 VN.n1208 a_400_62400# 2.51fF
C1405 VN.n1209 a_400_62400# 0.16fF
C1406 VN.t1493 a_400_62400# 0.03fF
C1407 VN.n1210 a_400_62400# 0.19fF
C1408 VN.t54 a_400_62400# 0.03fF
C1409 VN.n1212 a_400_62400# 0.32fF
C1410 VN.n1213 a_400_62400# 0.48fF
C1411 VN.n1214 a_400_62400# 0.81fF
C1412 VN.n1215 a_400_62400# 1.46fF
C1413 VN.n1216 a_400_62400# 0.21fF
C1414 VN.n1217 a_400_62400# 2.81fF
C1415 VN.t1678 a_400_62400# 0.03fF
C1416 VN.n1218 a_400_62400# 0.16fF
C1417 VN.n1219 a_400_62400# 0.19fF
C1418 VN.t1783 a_400_62400# 0.03fF
C1419 VN.n1221 a_400_62400# 0.32fF
C1420 VN.n1222 a_400_62400# 1.22fF
C1421 VN.n1223 a_400_62400# 0.07fF
C1422 VN.n1224 a_400_62400# 2.51fF
C1423 VN.n1225 a_400_62400# 3.57fF
C1424 VN.t593 a_400_62400# 0.03fF
C1425 VN.n1226 a_400_62400# 0.32fF
C1426 VN.n1227 a_400_62400# 0.48fF
C1427 VN.n1228 a_400_62400# 0.81fF
C1428 VN.n1229 a_400_62400# 0.16fF
C1429 VN.t1964 a_400_62400# 0.03fF
C1430 VN.n1230 a_400_62400# 0.19fF
C1431 VN.n1232 a_400_62400# 3.93fF
C1432 VN.n1233 a_400_62400# 3.08fF
C1433 VN.t2176 a_400_62400# 0.03fF
C1434 VN.n1234 a_400_62400# 0.16fF
C1435 VN.n1235 a_400_62400# 0.19fF
C1436 VN.t2275 a_400_62400# 0.03fF
C1437 VN.n1237 a_400_62400# 0.32fF
C1438 VN.n1238 a_400_62400# 1.22fF
C1439 VN.n1239 a_400_62400# 0.07fF
C1440 VN.n1240 a_400_62400# 2.51fF
C1441 VN.n1241 a_400_62400# 3.57fF
C1442 VN.t2246 a_400_62400# 0.03fF
C1443 VN.n1242 a_400_62400# 0.32fF
C1444 VN.n1243 a_400_62400# 0.48fF
C1445 VN.n1244 a_400_62400# 0.81fF
C1446 VN.n1245 a_400_62400# 0.16fF
C1447 VN.t1098 a_400_62400# 0.03fF
C1448 VN.n1246 a_400_62400# 0.19fF
C1449 VN.n1248 a_400_62400# 3.75fF
C1450 VN.n1249 a_400_62400# 3.08fF
C1451 VN.t1309 a_400_62400# 0.03fF
C1452 VN.n1250 a_400_62400# 0.16fF
C1453 VN.n1251 a_400_62400# 0.19fF
C1454 VN.t1406 a_400_62400# 0.03fF
C1455 VN.n1253 a_400_62400# 0.32fF
C1456 VN.n1254 a_400_62400# 1.22fF
C1457 VN.n1255 a_400_62400# 0.07fF
C1458 VN.n1256 a_400_62400# 2.51fF
C1459 VN.n1257 a_400_62400# 3.57fF
C1460 VN.t1384 a_400_62400# 0.03fF
C1461 VN.n1258 a_400_62400# 0.32fF
C1462 VN.n1259 a_400_62400# 0.48fF
C1463 VN.n1260 a_400_62400# 0.81fF
C1464 VN.n1261 a_400_62400# 0.16fF
C1465 VN.t366 a_400_62400# 0.03fF
C1466 VN.n1262 a_400_62400# 0.19fF
C1467 VN.n1264 a_400_62400# 3.75fF
C1468 VN.n1265 a_400_62400# 3.08fF
C1469 VN.t448 a_400_62400# 0.03fF
C1470 VN.n1266 a_400_62400# 0.16fF
C1471 VN.n1267 a_400_62400# 0.19fF
C1472 VN.t546 a_400_62400# 0.03fF
C1473 VN.n1269 a_400_62400# 0.32fF
C1474 VN.n1270 a_400_62400# 1.22fF
C1475 VN.n1271 a_400_62400# 0.07fF
C1476 VN.n1272 a_400_62400# 2.51fF
C1477 VN.n1273 a_400_62400# 3.57fF
C1478 VN.t629 a_400_62400# 0.03fF
C1479 VN.n1274 a_400_62400# 0.32fF
C1480 VN.n1275 a_400_62400# 0.48fF
C1481 VN.n1276 a_400_62400# 0.81fF
C1482 VN.n1277 a_400_62400# 0.16fF
C1483 VN.t2016 a_400_62400# 0.03fF
C1484 VN.n1278 a_400_62400# 0.19fF
C1485 VN.n1280 a_400_62400# 3.75fF
C1486 VN.n1281 a_400_62400# 3.08fF
C1487 VN.t2094 a_400_62400# 0.03fF
C1488 VN.n1282 a_400_62400# 0.16fF
C1489 VN.n1283 a_400_62400# 0.19fF
C1490 VN.t2323 a_400_62400# 0.03fF
C1491 VN.n1285 a_400_62400# 0.32fF
C1492 VN.n1286 a_400_62400# 1.22fF
C1493 VN.n1287 a_400_62400# 0.07fF
C1494 VN.n1288 a_400_62400# 2.51fF
C1495 VN.n1289 a_400_62400# 3.57fF
C1496 VN.t2286 a_400_62400# 0.03fF
C1497 VN.n1290 a_400_62400# 0.32fF
C1498 VN.n1291 a_400_62400# 0.48fF
C1499 VN.n1292 a_400_62400# 0.81fF
C1500 VN.n1293 a_400_62400# 0.16fF
C1501 VN.t1143 a_400_62400# 0.03fF
C1502 VN.n1294 a_400_62400# 0.19fF
C1503 VN.n1296 a_400_62400# 3.75fF
C1504 VN.n1297 a_400_62400# 3.08fF
C1505 VN.t1218 a_400_62400# 0.03fF
C1506 VN.n1298 a_400_62400# 0.16fF
C1507 VN.n1299 a_400_62400# 0.19fF
C1508 VN.t1457 a_400_62400# 0.03fF
C1509 VN.n1301 a_400_62400# 0.32fF
C1510 VN.n1302 a_400_62400# 1.22fF
C1511 VN.n1303 a_400_62400# 0.07fF
C1512 VN.n1304 a_400_62400# 2.51fF
C1513 VN.n1305 a_400_62400# 3.57fF
C1514 VN.t1417 a_400_62400# 0.03fF
C1515 VN.n1306 a_400_62400# 0.32fF
C1516 VN.n1307 a_400_62400# 0.48fF
C1517 VN.n1308 a_400_62400# 0.81fF
C1518 VN.n1309 a_400_62400# 0.16fF
C1519 VN.t279 a_400_62400# 0.03fF
C1520 VN.n1310 a_400_62400# 0.19fF
C1521 VN.n1312 a_400_62400# 3.75fF
C1522 VN.n1313 a_400_62400# 3.08fF
C1523 VN.t355 a_400_62400# 0.03fF
C1524 VN.n1314 a_400_62400# 0.16fF
C1525 VN.n1315 a_400_62400# 0.19fF
C1526 VN.t587 a_400_62400# 0.03fF
C1527 VN.n1317 a_400_62400# 0.32fF
C1528 VN.n1318 a_400_62400# 1.22fF
C1529 VN.n1319 a_400_62400# 0.07fF
C1530 VN.n1320 a_400_62400# 2.51fF
C1531 VN.n1321 a_400_62400# 3.57fF
C1532 VN.t554 a_400_62400# 0.03fF
C1533 VN.n1322 a_400_62400# 0.32fF
C1534 VN.n1323 a_400_62400# 0.48fF
C1535 VN.n1324 a_400_62400# 0.81fF
C1536 VN.n1325 a_400_62400# 0.16fF
C1537 VN.t1930 a_400_62400# 0.03fF
C1538 VN.n1326 a_400_62400# 0.19fF
C1539 VN.n1328 a_400_62400# 3.75fF
C1540 VN.n1329 a_400_62400# 3.08fF
C1541 VN.t2000 a_400_62400# 0.03fF
C1542 VN.n1330 a_400_62400# 0.16fF
C1543 VN.n1331 a_400_62400# 0.19fF
C1544 VN.t2243 a_400_62400# 0.03fF
C1545 VN.n1333 a_400_62400# 0.32fF
C1546 VN.n1334 a_400_62400# 1.22fF
C1547 VN.n1335 a_400_62400# 0.07fF
C1548 VN.n1336 a_400_62400# 2.51fF
C1549 VN.n1337 a_400_62400# 3.57fF
C1550 VN.t2212 a_400_62400# 0.03fF
C1551 VN.n1338 a_400_62400# 0.32fF
C1552 VN.n1339 a_400_62400# 0.48fF
C1553 VN.n1340 a_400_62400# 0.81fF
C1554 VN.n1341 a_400_62400# 0.16fF
C1555 VN.t1055 a_400_62400# 0.03fF
C1556 VN.n1342 a_400_62400# 0.19fF
C1557 VN.n1344 a_400_62400# 3.75fF
C1558 VN.n1345 a_400_62400# 3.08fF
C1559 VN.t1268 a_400_62400# 0.03fF
C1560 VN.n1346 a_400_62400# 0.16fF
C1561 VN.n1347 a_400_62400# 0.19fF
C1562 VN.t1380 a_400_62400# 0.03fF
C1563 VN.n1349 a_400_62400# 0.32fF
C1564 VN.n1350 a_400_62400# 1.22fF
C1565 VN.n1351 a_400_62400# 0.07fF
C1566 VN.n1352 a_400_62400# 2.51fF
C1567 VN.n1353 a_400_62400# 3.57fF
C1568 VN.t1345 a_400_62400# 0.03fF
C1569 VN.n1354 a_400_62400# 0.32fF
C1570 VN.n1355 a_400_62400# 0.48fF
C1571 VN.n1356 a_400_62400# 0.81fF
C1572 VN.n1357 a_400_62400# 0.16fF
C1573 VN.t182 a_400_62400# 0.03fF
C1574 VN.n1358 a_400_62400# 0.19fF
C1575 VN.n1360 a_400_62400# 3.75fF
C1576 VN.n1361 a_400_62400# 3.08fF
C1577 VN.t399 a_400_62400# 0.03fF
C1578 VN.n1362 a_400_62400# 0.16fF
C1579 VN.n1363 a_400_62400# 0.19fF
C1580 VN.t515 a_400_62400# 0.03fF
C1581 VN.n1365 a_400_62400# 0.32fF
C1582 VN.n1366 a_400_62400# 1.22fF
C1583 VN.n1367 a_400_62400# 0.07fF
C1584 VN.n1368 a_400_62400# 2.51fF
C1585 VN.n1369 a_400_62400# 3.57fF
C1586 VN.t499 a_400_62400# 0.03fF
C1587 VN.n1370 a_400_62400# 0.32fF
C1588 VN.n1371 a_400_62400# 0.48fF
C1589 VN.n1372 a_400_62400# 0.81fF
C1590 VN.n1373 a_400_62400# 0.16fF
C1591 VN.t1853 a_400_62400# 0.03fF
C1592 VN.n1374 a_400_62400# 0.19fF
C1593 VN.n1376 a_400_62400# 3.75fF
C1594 VN.n1377 a_400_62400# 3.08fF
C1595 VN.t2064 a_400_62400# 0.03fF
C1596 VN.n1378 a_400_62400# 0.16fF
C1597 VN.n1379 a_400_62400# 0.19fF
C1598 VN.t2284 a_400_62400# 0.03fF
C1599 VN.n1381 a_400_62400# 0.32fF
C1600 VN.n1382 a_400_62400# 1.22fF
C1601 VN.n1383 a_400_62400# 0.07fF
C1602 VN.n1384 a_400_62400# 2.51fF
C1603 VN.n1385 a_400_62400# 3.57fF
C1604 VN.t2154 a_400_62400# 0.03fF
C1605 VN.n1386 a_400_62400# 0.32fF
C1606 VN.n1387 a_400_62400# 0.48fF
C1607 VN.n1388 a_400_62400# 0.81fF
C1608 VN.n1389 a_400_62400# 0.16fF
C1609 VN.t984 a_400_62400# 0.03fF
C1610 VN.n1390 a_400_62400# 0.19fF
C1611 VN.n1392 a_400_62400# 3.75fF
C1612 VN.n1393 a_400_62400# 3.08fF
C1613 VN.t1192 a_400_62400# 0.03fF
C1614 VN.n1394 a_400_62400# 0.16fF
C1615 VN.n1395 a_400_62400# 0.19fF
C1616 VN.t1415 a_400_62400# 0.03fF
C1617 VN.n1397 a_400_62400# 0.32fF
C1618 VN.n1398 a_400_62400# 1.22fF
C1619 VN.n1399 a_400_62400# 0.07fF
C1620 VN.n1400 a_400_62400# 3.65fF
C1621 VN.n1401 a_400_62400# 2.14fF
C1622 VN.n1402 a_400_62400# 0.16fF
C1623 VN.t1895 a_400_62400# 0.03fF
C1624 VN.n1403 a_400_62400# 0.19fF
C1625 VN.t419 a_400_62400# 0.03fF
C1626 VN.n1405 a_400_62400# 0.32fF
C1627 VN.n1406 a_400_62400# 0.48fF
C1628 VN.n1407 a_400_62400# 0.81fF
C1629 VN.n1408 a_400_62400# 0.09fF
C1630 VN.n1409 a_400_62400# 0.01fF
C1631 VN.n1410 a_400_62400# 0.02fF
C1632 VN.n1411 a_400_62400# 0.02fF
C1633 VN.n1412 a_400_62400# 0.32fF
C1634 VN.n1413 a_400_62400# 1.56fF
C1635 VN.n1414 a_400_62400# 1.81fF
C1636 VN.n1415 a_400_62400# 3.08fF
C1637 VN.t1969 a_400_62400# 0.03fF
C1638 VN.n1416 a_400_62400# 0.16fF
C1639 VN.n1417 a_400_62400# 0.19fF
C1640 VN.t2209 a_400_62400# 0.03fF
C1641 VN.n1419 a_400_62400# 0.32fF
C1642 VN.n1420 a_400_62400# 1.22fF
C1643 VN.n1421 a_400_62400# 0.07fF
C1644 VN.t94 a_400_62400# 64.69fF
C1645 VN.t553 a_400_62400# 0.03fF
C1646 VN.n1422 a_400_62400# 0.32fF
C1647 VN.n1423 a_400_62400# 1.22fF
C1648 VN.n1424 a_400_62400# 0.07fF
C1649 VN.t322 a_400_62400# 0.03fF
C1650 VN.n1425 a_400_62400# 0.16fF
C1651 VN.n1426 a_400_62400# 0.19fF
C1652 VN.n1428 a_400_62400# 0.16fF
C1653 VN.t95 a_400_62400# 0.03fF
C1654 VN.n1429 a_400_62400# 0.19fF
C1655 VN.n1431 a_400_62400# 6.92fF
C1656 VN.n1432 a_400_62400# 6.56fF
C1657 VN.t1943 a_400_62400# 0.03fF
C1658 VN.n1433 a_400_62400# 0.16fF
C1659 VN.n1434 a_400_62400# 0.19fF
C1660 VN.t1473 a_400_62400# 0.03fF
C1661 VN.n1436 a_400_62400# 0.32fF
C1662 VN.n1437 a_400_62400# 1.22fF
C1663 VN.n1438 a_400_62400# 0.07fF
C1664 VN.n1439 a_400_62400# 2.51fF
C1665 VN.n1440 a_400_62400# 3.58fF
C1666 VN.t1553 a_400_62400# 0.03fF
C1667 VN.n1441 a_400_62400# 0.32fF
C1668 VN.n1442 a_400_62400# 0.48fF
C1669 VN.n1443 a_400_62400# 0.81fF
C1670 VN.n1444 a_400_62400# 0.16fF
C1671 VN.t416 a_400_62400# 0.03fF
C1672 VN.n1445 a_400_62400# 0.19fF
C1673 VN.n1447 a_400_62400# 7.29fF
C1674 VN.t1072 a_400_62400# 0.03fF
C1675 VN.n1448 a_400_62400# 0.16fF
C1676 VN.n1449 a_400_62400# 0.19fF
C1677 VN.t606 a_400_62400# 0.03fF
C1678 VN.n1451 a_400_62400# 0.32fF
C1679 VN.n1452 a_400_62400# 1.22fF
C1680 VN.n1453 a_400_62400# 0.07fF
C1681 VN.t24 a_400_62400# 64.17fF
C1682 VN.t2258 a_400_62400# 0.03fF
C1683 VN.n1454 a_400_62400# 1.60fF
C1684 VN.n1455 a_400_62400# 0.07fF
C1685 VN.t343 a_400_62400# 0.03fF
C1686 VN.n1456 a_400_62400# 0.02fF
C1687 VN.n1457 a_400_62400# 0.34fF
C1688 VN.n1459 a_400_62400# 2.01fF
C1689 VN.n1460 a_400_62400# 1.68fF
C1690 VN.n1461 a_400_62400# 0.37fF
C1691 VN.n1462 a_400_62400# 0.33fF
C1692 VN.n1463 a_400_62400# 5.87fF
C1693 VN.n1464 a_400_62400# 0.02fF
C1694 VN.n1465 a_400_62400# 0.02fF
C1695 VN.n1466 a_400_62400# 0.03fF
C1696 VN.n1467 a_400_62400# 0.05fF
C1697 VN.n1468 a_400_62400# 0.23fF
C1698 VN.n1469 a_400_62400# 0.02fF
C1699 VN.n1470 a_400_62400# 0.03fF
C1700 VN.n1471 a_400_62400# 0.01fF
C1701 VN.n1472 a_400_62400# 0.01fF
C1702 VN.n1473 a_400_62400# 0.01fF
C1703 VN.n1474 a_400_62400# 0.02fF
C1704 VN.n1475 a_400_62400# 0.03fF
C1705 VN.n1476 a_400_62400# 0.06fF
C1706 VN.n1477 a_400_62400# 0.05fF
C1707 VN.n1478 a_400_62400# 0.15fF
C1708 VN.n1479 a_400_62400# 0.51fF
C1709 VN.n1480 a_400_62400# 0.27fF
C1710 VN.n1481 a_400_62400# 37.46fF
C1711 VN.n1482 a_400_62400# 37.46fF
C1712 VN.n1483 a_400_62400# 0.79fF
C1713 VN.n1484 a_400_62400# 0.23fF
C1714 VN.n1485 a_400_62400# 1.18fF
C1715 VN.t114 a_400_62400# 28.64fF
C1716 VN.n1486 a_400_62400# 0.79fF
C1717 VN.n1487 a_400_62400# 0.11fF
C1718 VN.n1488 a_400_62400# 4.98fF
C1719 VN.n1489 a_400_62400# 0.80fF
C1720 VN.n1490 a_400_62400# 0.29fF
C1721 VN.n1491 a_400_62400# 1.96fF
C1722 VN.n1493 a_400_62400# 25.18fF
C1723 VN.n1495 a_400_62400# 1.87fF
C1724 VN.n1496 a_400_62400# 5.36fF
C1725 VN.n1497 a_400_62400# 1.81fF
C1726 VN.t1528 a_400_62400# 0.03fF
C1727 VN.n1498 a_400_62400# 0.85fF
C1728 VN.n1499 a_400_62400# 0.81fF
C1729 VN.n1500 a_400_62400# 2.51fF
C1730 VN.n1501 a_400_62400# 0.61fF
C1731 VN.n1502 a_400_62400# 0.30fF
C1732 VN.n1503 a_400_62400# 0.51fF
C1733 VN.n1504 a_400_62400# 0.21fF
C1734 VN.n1505 a_400_62400# 0.38fF
C1735 VN.n1506 a_400_62400# 0.29fF
C1736 VN.n1507 a_400_62400# 0.40fF
C1737 VN.n1508 a_400_62400# 0.28fF
C1738 VN.t1070 a_400_62400# 0.03fF
C1739 VN.n1509 a_400_62400# 0.32fF
C1740 VN.n1510 a_400_62400# 0.48fF
C1741 VN.n1511 a_400_62400# 0.81fF
C1742 VN.n1512 a_400_62400# 0.16fF
C1743 VN.t2577 a_400_62400# 0.03fF
C1744 VN.n1513 a_400_62400# 0.19fF
C1745 VN.n1515 a_400_62400# 0.06fF
C1746 VN.n1516 a_400_62400# 0.04fF
C1747 VN.n1517 a_400_62400# 0.04fF
C1748 VN.n1518 a_400_62400# 0.14fF
C1749 VN.n1519 a_400_62400# 0.48fF
C1750 VN.n1520 a_400_62400# 0.50fF
C1751 VN.n1521 a_400_62400# 0.14fF
C1752 VN.n1522 a_400_62400# 0.16fF
C1753 VN.n1523 a_400_62400# 0.09fF
C1754 VN.n1524 a_400_62400# 0.16fF
C1755 VN.n1525 a_400_62400# 0.24fF
C1756 VN.n1526 a_400_62400# 5.35fF
C1757 VN.t1690 a_400_62400# 0.03fF
C1758 VN.n1527 a_400_62400# 0.32fF
C1759 VN.n1528 a_400_62400# 1.22fF
C1760 VN.n1529 a_400_62400# 0.07fF
C1761 VN.t737 a_400_62400# 0.03fF
C1762 VN.n1530 a_400_62400# 0.16fF
C1763 VN.n1531 a_400_62400# 0.19fF
C1764 VN.t942 a_400_62400# 0.03fF
C1765 VN.n1533 a_400_62400# 0.32fF
C1766 VN.n1534 a_400_62400# 1.22fF
C1767 VN.n1535 a_400_62400# 0.07fF
C1768 VN.n1536 a_400_62400# 0.33fF
C1769 VN.n1537 a_400_62400# 0.12fF
C1770 VN.n1538 a_400_62400# 0.28fF
C1771 VN.n1539 a_400_62400# 1.72fF
C1772 VN.n1540 a_400_62400# 0.71fF
C1773 VN.n1541 a_400_62400# 2.51fF
C1774 VN.n1542 a_400_62400# 0.16fF
C1775 VN.t1706 a_400_62400# 0.03fF
C1776 VN.n1543 a_400_62400# 0.19fF
C1777 VN.t340 a_400_62400# 0.03fF
C1778 VN.n1545 a_400_62400# 0.32fF
C1779 VN.n1546 a_400_62400# 0.48fF
C1780 VN.n1547 a_400_62400# 0.81fF
C1781 VN.n1548 a_400_62400# 0.95fF
C1782 VN.n1549 a_400_62400# 2.11fF
C1783 VN.n1550 a_400_62400# 3.28fF
C1784 VN.t2393 a_400_62400# 0.03fF
C1785 VN.n1551 a_400_62400# 0.16fF
C1786 VN.n1552 a_400_62400# 0.19fF
C1787 VN.n1554 a_400_62400# 2.53fF
C1788 VN.n1555 a_400_62400# 0.08fF
C1789 VN.n1556 a_400_62400# 0.04fF
C1790 VN.n1557 a_400_62400# 0.05fF
C1791 VN.n1558 a_400_62400# 1.33fF
C1792 VN.n1559 a_400_62400# 0.03fF
C1793 VN.n1560 a_400_62400# 0.01fF
C1794 VN.n1561 a_400_62400# 0.02fF
C1795 VN.n1562 a_400_62400# 0.11fF
C1796 VN.n1563 a_400_62400# 0.48fF
C1797 VN.n1564 a_400_62400# 2.48fF
C1798 VN.t1984 a_400_62400# 0.03fF
C1799 VN.n1565 a_400_62400# 0.32fF
C1800 VN.n1566 a_400_62400# 0.48fF
C1801 VN.n1567 a_400_62400# 0.81fF
C1802 VN.n1568 a_400_62400# 0.16fF
C1803 VN.t835 a_400_62400# 0.03fF
C1804 VN.n1569 a_400_62400# 0.19fF
C1805 VN.n1571 a_400_62400# 0.93fF
C1806 VN.n1572 a_400_62400# 0.30fF
C1807 VN.n1573 a_400_62400# 0.34fF
C1808 VN.n1574 a_400_62400# 0.12fF
C1809 VN.n1575 a_400_62400# 0.30fF
C1810 VN.n1576 a_400_62400# 0.93fF
C1811 VN.n1577 a_400_62400# 1.55fF
C1812 VN.n1578 a_400_62400# 0.29fF
C1813 VN.n1579 a_400_62400# 0.34fF
C1814 VN.n1580 a_400_62400# 0.12fF
C1815 VN.n1581 a_400_62400# 2.52fF
C1816 VN.t17 a_400_62400# 0.03fF
C1817 VN.n1582 a_400_62400# 0.32fF
C1818 VN.n1583 a_400_62400# 1.22fF
C1819 VN.n1584 a_400_62400# 0.07fF
C1820 VN.t1525 a_400_62400# 0.03fF
C1821 VN.n1585 a_400_62400# 0.16fF
C1822 VN.n1586 a_400_62400# 0.19fF
C1823 VN.n1588 a_400_62400# 27.83fF
C1824 VN.n1589 a_400_62400# 2.30fF
C1825 VN.n1590 a_400_62400# 0.88fF
C1826 VN.n1591 a_400_62400# 0.93fF
C1827 VN.n1592 a_400_62400# 0.97fF
C1828 VN.n1593 a_400_62400# 0.49fF
C1829 VN.t1941 a_400_62400# 0.03fF
C1830 VN.n1594 a_400_62400# 0.32fF
C1831 VN.n1595 a_400_62400# 0.48fF
C1832 VN.n1596 a_400_62400# 0.81fF
C1833 VN.n1597 a_400_62400# 0.16fF
C1834 VN.t801 a_400_62400# 0.03fF
C1835 VN.n1598 a_400_62400# 0.19fF
C1836 VN.n1600 a_400_62400# 0.42fF
C1837 VN.n1601 a_400_62400# 0.34fF
C1838 VN.n1602 a_400_62400# 0.12fF
C1839 VN.n1603 a_400_62400# 0.30fF
C1840 VN.n1604 a_400_62400# 0.88fF
C1841 VN.n1605 a_400_62400# 1.28fF
C1842 VN.n1606 a_400_62400# 0.30fF
C1843 VN.n1607 a_400_62400# 0.28fF
C1844 VN.n1608 a_400_62400# 0.27fF
C1845 VN.n1609 a_400_62400# 0.09fF
C1846 VN.n1610 a_400_62400# 0.12fF
C1847 VN.n1611 a_400_62400# 0.13fF
C1848 VN.n1612 a_400_62400# 2.24fF
C1849 VN.t1604 a_400_62400# 0.03fF
C1850 VN.n1613 a_400_62400# 0.16fF
C1851 VN.n1614 a_400_62400# 0.19fF
C1852 VN.t2560 a_400_62400# 0.03fF
C1853 VN.n1616 a_400_62400# 0.32fF
C1854 VN.n1617 a_400_62400# 1.22fF
C1855 VN.n1618 a_400_62400# 0.07fF
C1856 VN.n1619 a_400_62400# 2.51fF
C1857 VN.n1620 a_400_62400# 0.16fF
C1858 VN.t1342 a_400_62400# 0.03fF
C1859 VN.n1621 a_400_62400# 0.19fF
C1860 VN.t2462 a_400_62400# 0.03fF
C1861 VN.n1623 a_400_62400# 0.32fF
C1862 VN.n1624 a_400_62400# 0.48fF
C1863 VN.n1625 a_400_62400# 0.81fF
C1864 VN.n1626 a_400_62400# 1.24fF
C1865 VN.n1627 a_400_62400# 0.43fF
C1866 VN.n1628 a_400_62400# 0.43fF
C1867 VN.n1629 a_400_62400# 1.24fF
C1868 VN.n1630 a_400_62400# 1.46fF
C1869 VN.n1631 a_400_62400# 0.21fF
C1870 VN.n1632 a_400_62400# 6.64fF
C1871 VN.t656 a_400_62400# 0.03fF
C1872 VN.n1633 a_400_62400# 0.16fF
C1873 VN.n1634 a_400_62400# 0.19fF
C1874 VN.t572 a_400_62400# 0.03fF
C1875 VN.n1636 a_400_62400# 0.32fF
C1876 VN.n1637 a_400_62400# 1.22fF
C1877 VN.n1638 a_400_62400# 0.07fF
C1878 VN.n1639 a_400_62400# 2.51fF
C1879 VN.n1640 a_400_62400# 3.57fF
C1880 VN.t1596 a_400_62400# 0.03fF
C1881 VN.n1641 a_400_62400# 0.32fF
C1882 VN.n1642 a_400_62400# 0.48fF
C1883 VN.n1643 a_400_62400# 0.81fF
C1884 VN.n1644 a_400_62400# 0.16fF
C1885 VN.t479 a_400_62400# 0.03fF
C1886 VN.n1645 a_400_62400# 0.19fF
C1887 VN.n1647 a_400_62400# 6.91fF
C1888 VN.t1131 a_400_62400# 0.03fF
C1889 VN.n1648 a_400_62400# 0.16fF
C1890 VN.n1649 a_400_62400# 0.19fF
C1891 VN.t2230 a_400_62400# 0.03fF
C1892 VN.n1651 a_400_62400# 0.32fF
C1893 VN.n1652 a_400_62400# 1.22fF
C1894 VN.n1653 a_400_62400# 0.07fF
C1895 VN.n1654 a_400_62400# 2.51fF
C1896 VN.n1655 a_400_62400# 3.57fF
C1897 VN.t731 a_400_62400# 0.03fF
C1898 VN.n1656 a_400_62400# 0.32fF
C1899 VN.n1657 a_400_62400# 0.48fF
C1900 VN.n1658 a_400_62400# 0.81fF
C1901 VN.n1659 a_400_62400# 0.16fF
C1902 VN.t2134 a_400_62400# 0.03fF
C1903 VN.n1660 a_400_62400# 0.19fF
C1904 VN.n1662 a_400_62400# 6.92fF
C1905 VN.t267 a_400_62400# 0.03fF
C1906 VN.n1663 a_400_62400# 0.16fF
C1907 VN.n1664 a_400_62400# 0.19fF
C1908 VN.t1365 a_400_62400# 0.03fF
C1909 VN.n1666 a_400_62400# 0.32fF
C1910 VN.n1667 a_400_62400# 1.22fF
C1911 VN.n1668 a_400_62400# 0.07fF
C1912 VN.n1669 a_400_62400# 2.51fF
C1913 VN.n1670 a_400_62400# 3.57fF
C1914 VN.t2385 a_400_62400# 0.03fF
C1915 VN.n1671 a_400_62400# 0.32fF
C1916 VN.n1672 a_400_62400# 0.48fF
C1917 VN.n1673 a_400_62400# 0.81fF
C1918 VN.n1674 a_400_62400# 0.16fF
C1919 VN.t1258 a_400_62400# 0.03fF
C1920 VN.n1675 a_400_62400# 0.19fF
C1921 VN.n1677 a_400_62400# 6.92fF
C1922 VN.t2053 a_400_62400# 0.03fF
C1923 VN.n1678 a_400_62400# 0.16fF
C1924 VN.n1679 a_400_62400# 0.19fF
C1925 VN.t500 a_400_62400# 0.03fF
C1926 VN.n1681 a_400_62400# 0.32fF
C1927 VN.n1682 a_400_62400# 1.22fF
C1928 VN.n1683 a_400_62400# 0.07fF
C1929 VN.n1684 a_400_62400# 2.51fF
C1930 VN.n1685 a_400_62400# 3.57fF
C1931 VN.t1517 a_400_62400# 0.03fF
C1932 VN.n1686 a_400_62400# 0.32fF
C1933 VN.n1687 a_400_62400# 0.48fF
C1934 VN.n1688 a_400_62400# 0.81fF
C1935 VN.n1689 a_400_62400# 0.16fF
C1936 VN.t390 a_400_62400# 0.03fF
C1937 VN.n1690 a_400_62400# 0.19fF
C1938 VN.n1692 a_400_62400# 6.92fF
C1939 VN.t1184 a_400_62400# 0.03fF
C1940 VN.n1693 a_400_62400# 0.16fF
C1941 VN.n1694 a_400_62400# 0.19fF
C1942 VN.t2156 a_400_62400# 0.03fF
C1943 VN.n1696 a_400_62400# 0.32fF
C1944 VN.n1697 a_400_62400# 1.22fF
C1945 VN.n1698 a_400_62400# 0.07fF
C1946 VN.n1699 a_400_62400# 2.51fF
C1947 VN.n1700 a_400_62400# 3.57fF
C1948 VN.t649 a_400_62400# 0.03fF
C1949 VN.n1701 a_400_62400# 0.32fF
C1950 VN.n1702 a_400_62400# 0.48fF
C1951 VN.n1703 a_400_62400# 0.81fF
C1952 VN.n1704 a_400_62400# 0.16fF
C1953 VN.t2043 a_400_62400# 0.03fF
C1954 VN.n1705 a_400_62400# 0.19fF
C1955 VN.n1707 a_400_62400# 6.92fF
C1956 VN.t312 a_400_62400# 0.03fF
C1957 VN.n1708 a_400_62400# 0.16fF
C1958 VN.n1709 a_400_62400# 0.19fF
C1959 VN.t1288 a_400_62400# 0.03fF
C1960 VN.n1711 a_400_62400# 0.32fF
C1961 VN.n1712 a_400_62400# 1.22fF
C1962 VN.n1713 a_400_62400# 0.07fF
C1963 VN.n1714 a_400_62400# 2.51fF
C1964 VN.n1715 a_400_62400# 3.57fF
C1965 VN.t2308 a_400_62400# 0.03fF
C1966 VN.n1716 a_400_62400# 0.32fF
C1967 VN.n1717 a_400_62400# 0.48fF
C1968 VN.n1718 a_400_62400# 0.81fF
C1969 VN.n1719 a_400_62400# 0.16fF
C1970 VN.t1171 a_400_62400# 0.03fF
C1971 VN.n1720 a_400_62400# 0.19fF
C1972 VN.n1722 a_400_62400# 6.92fF
C1973 VN.t1961 a_400_62400# 0.03fF
C1974 VN.n1723 a_400_62400# 0.16fF
C1975 VN.n1724 a_400_62400# 0.19fF
C1976 VN.t421 a_400_62400# 0.03fF
C1977 VN.n1726 a_400_62400# 0.32fF
C1978 VN.n1727 a_400_62400# 1.22fF
C1979 VN.n1728 a_400_62400# 0.07fF
C1980 VN.n1729 a_400_62400# 2.51fF
C1981 VN.n1730 a_400_62400# 3.57fF
C1982 VN.t1438 a_400_62400# 0.03fF
C1983 VN.n1731 a_400_62400# 0.32fF
C1984 VN.n1732 a_400_62400# 0.48fF
C1985 VN.n1733 a_400_62400# 0.81fF
C1986 VN.n1734 a_400_62400# 0.16fF
C1987 VN.t443 a_400_62400# 0.03fF
C1988 VN.n1735 a_400_62400# 0.19fF
C1989 VN.n1737 a_400_62400# 6.92fF
C1990 VN.t1094 a_400_62400# 0.03fF
C1991 VN.n1738 a_400_62400# 0.16fF
C1992 VN.n1739 a_400_62400# 0.19fF
C1993 VN.t2068 a_400_62400# 0.03fF
C1994 VN.n1741 a_400_62400# 0.32fF
C1995 VN.n1742 a_400_62400# 1.22fF
C1996 VN.n1743 a_400_62400# 0.07fF
C1997 VN.n1744 a_400_62400# 2.51fF
C1998 VN.n1745 a_400_62400# 3.57fF
C1999 VN.t693 a_400_62400# 0.03fF
C2000 VN.n1746 a_400_62400# 0.32fF
C2001 VN.n1747 a_400_62400# 0.48fF
C2002 VN.n1748 a_400_62400# 0.81fF
C2003 VN.n1749 a_400_62400# 0.16fF
C2004 VN.t2088 a_400_62400# 0.03fF
C2005 VN.n1750 a_400_62400# 0.19fF
C2006 VN.n1752 a_400_62400# 6.92fF
C2007 VN.t225 a_400_62400# 0.03fF
C2008 VN.n1753 a_400_62400# 0.16fF
C2009 VN.n1754 a_400_62400# 0.19fF
C2010 VN.t1329 a_400_62400# 0.03fF
C2011 VN.n1756 a_400_62400# 0.32fF
C2012 VN.n1757 a_400_62400# 1.22fF
C2013 VN.n1758 a_400_62400# 0.07fF
C2014 VN.n1759 a_400_62400# 2.51fF
C2015 VN.n1760 a_400_62400# 3.57fF
C2016 VN.t2469 a_400_62400# 0.03fF
C2017 VN.n1761 a_400_62400# 0.32fF
C2018 VN.n1762 a_400_62400# 0.48fF
C2019 VN.n1763 a_400_62400# 0.81fF
C2020 VN.n1764 a_400_62400# 0.16fF
C2021 VN.t1341 a_400_62400# 0.03fF
C2022 VN.n1765 a_400_62400# 0.19fF
C2023 VN.n1767 a_400_62400# 6.92fF
C2024 VN.t1873 a_400_62400# 0.03fF
C2025 VN.n1768 a_400_62400# 0.16fF
C2026 VN.n1769 a_400_62400# 0.19fF
C2027 VN.t2003 a_400_62400# 0.03fF
C2028 VN.n1771 a_400_62400# 0.32fF
C2029 VN.n1772 a_400_62400# 1.22fF
C2030 VN.n1773 a_400_62400# 0.07fF
C2031 VN.n1774 a_400_62400# 2.51fF
C2032 VN.n1775 a_400_62400# 3.57fF
C2033 VN.t1605 a_400_62400# 0.03fF
C2034 VN.n1776 a_400_62400# 0.32fF
C2035 VN.n1777 a_400_62400# 0.48fF
C2036 VN.n1778 a_400_62400# 0.81fF
C2037 VN.n1779 a_400_62400# 0.16fF
C2038 VN.t476 a_400_62400# 0.03fF
C2039 VN.n1780 a_400_62400# 0.19fF
C2040 VN.n1782 a_400_62400# 6.92fF
C2041 VN.t1130 a_400_62400# 0.03fF
C2042 VN.n1783 a_400_62400# 0.16fF
C2043 VN.n1784 a_400_62400# 0.19fF
C2044 VN.t1129 a_400_62400# 0.03fF
C2045 VN.n1786 a_400_62400# 0.32fF
C2046 VN.n1787 a_400_62400# 1.22fF
C2047 VN.n1788 a_400_62400# 0.07fF
C2048 VN.n1789 a_400_62400# 2.51fF
C2049 VN.n1790 a_400_62400# 3.57fF
C2050 VN.t740 a_400_62400# 0.03fF
C2051 VN.n1791 a_400_62400# 0.32fF
C2052 VN.n1792 a_400_62400# 0.48fF
C2053 VN.n1793 a_400_62400# 0.81fF
C2054 VN.n1794 a_400_62400# 0.16fF
C2055 VN.t2129 a_400_62400# 0.03fF
C2056 VN.n1795 a_400_62400# 0.19fF
C2057 VN.n1797 a_400_62400# 2.51fF
C2058 VN.n1798 a_400_62400# 3.59fF
C2059 VN.t2585 a_400_62400# 0.03fF
C2060 VN.n1799 a_400_62400# 0.32fF
C2061 VN.n1800 a_400_62400# 0.48fF
C2062 VN.n1801 a_400_62400# 0.81fF
C2063 VN.t831 a_400_62400# 0.03fF
C2064 VN.n1802 a_400_62400# 1.63fF
C2065 VN.n1803 a_400_62400# 0.49fF
C2066 VN.n1804 a_400_62400# 1.64fF
C2067 VN.n1805 a_400_62400# 0.81fF
C2068 VN.n1806 a_400_62400# 1.21fF
C2069 VN.n1807 a_400_62400# 1.54fF
C2070 VN.n1808 a_400_62400# 4.06fF
C2071 VN.t16 a_400_62400# 28.64fF
C2072 VN.n1809 a_400_62400# 28.43fF
C2073 VN.n1811 a_400_62400# 0.50fF
C2074 VN.n1812 a_400_62400# 0.31fF
C2075 VN.n1813 a_400_62400# 3.74fF
C2076 VN.n1814 a_400_62400# 3.29fF
C2077 VN.n1815 a_400_62400# 5.35fF
C2078 VN.n1816 a_400_62400# 0.34fF
C2079 VN.n1817 a_400_62400# 0.02fF
C2080 VN.t2239 a_400_62400# 0.03fF
C2081 VN.n1818 a_400_62400# 0.34fF
C2082 VN.t2527 a_400_62400# 0.03fF
C2083 VN.n1819 a_400_62400# 1.28fF
C2084 VN.n1820 a_400_62400# 0.94fF
C2085 VN.n1821 a_400_62400# 2.53fF
C2086 VN.n1822 a_400_62400# 2.32fF
C2087 VN.t2494 a_400_62400# 0.03fF
C2088 VN.n1823 a_400_62400# 0.32fF
C2089 VN.n1824 a_400_62400# 0.48fF
C2090 VN.n1825 a_400_62400# 0.81fF
C2091 VN.n1826 a_400_62400# 0.16fF
C2092 VN.t1374 a_400_62400# 0.03fF
C2093 VN.n1827 a_400_62400# 0.19fF
C2094 VN.n1829 a_400_62400# 1.55fF
C2095 VN.n1830 a_400_62400# 0.29fF
C2096 VN.n1831 a_400_62400# 3.27fF
C2097 VN.t1663 a_400_62400# 0.03fF
C2098 VN.n1832 a_400_62400# 0.32fF
C2099 VN.n1833 a_400_62400# 1.22fF
C2100 VN.n1834 a_400_62400# 0.07fF
C2101 VN.t1431 a_400_62400# 0.03fF
C2102 VN.n1835 a_400_62400# 0.16fF
C2103 VN.n1836 a_400_62400# 0.19fF
C2104 VN.n1838 a_400_62400# 2.51fF
C2105 VN.n1839 a_400_62400# 0.56fF
C2106 VN.n1840 a_400_62400# 0.64fF
C2107 VN.n1841 a_400_62400# 0.12fF
C2108 VN.n1842 a_400_62400# 0.44fF
C2109 VN.n1843 a_400_62400# 0.40fF
C2110 VN.n1844 a_400_62400# 1.03fF
C2111 VN.n1845 a_400_62400# 0.79fF
C2112 VN.t1628 a_400_62400# 0.03fF
C2113 VN.n1846 a_400_62400# 0.32fF
C2114 VN.n1847 a_400_62400# 0.48fF
C2115 VN.n1848 a_400_62400# 0.81fF
C2116 VN.n1849 a_400_62400# 0.16fF
C2117 VN.t508 a_400_62400# 0.03fF
C2118 VN.n1850 a_400_62400# 0.19fF
C2119 VN.n1852 a_400_62400# 3.50fF
C2120 VN.n1853 a_400_62400# 2.89fF
C2121 VN.t795 a_400_62400# 0.03fF
C2122 VN.n1854 a_400_62400# 0.32fF
C2123 VN.n1855 a_400_62400# 1.22fF
C2124 VN.n1856 a_400_62400# 0.07fF
C2125 VN.t687 a_400_62400# 0.03fF
C2126 VN.n1857 a_400_62400# 0.16fF
C2127 VN.n1858 a_400_62400# 0.19fF
C2128 VN.n1860 a_400_62400# 1.05fF
C2129 VN.n1861 a_400_62400# 3.07fF
C2130 VN.n1862 a_400_62400# 2.51fF
C2131 VN.n1863 a_400_62400# 0.16fF
C2132 VN.t2161 a_400_62400# 0.03fF
C2133 VN.n1864 a_400_62400# 0.19fF
C2134 VN.t756 a_400_62400# 0.03fF
C2135 VN.n1866 a_400_62400# 0.32fF
C2136 VN.n1867 a_400_62400# 0.48fF
C2137 VN.n1868 a_400_62400# 0.81fF
C2138 VN.n1869 a_400_62400# 1.86fF
C2139 VN.n1870 a_400_62400# 1.53fF
C2140 VN.n1871 a_400_62400# 0.47fF
C2141 VN.n1872 a_400_62400# 2.71fF
C2142 VN.t2449 a_400_62400# 0.03fF
C2143 VN.n1873 a_400_62400# 0.32fF
C2144 VN.n1874 a_400_62400# 1.22fF
C2145 VN.n1875 a_400_62400# 0.07fF
C2146 VN.t2345 a_400_62400# 0.03fF
C2147 VN.n1876 a_400_62400# 0.16fF
C2148 VN.n1877 a_400_62400# 0.19fF
C2149 VN.n1879 a_400_62400# 2.53fF
C2150 VN.n1880 a_400_62400# 2.51fF
C2151 VN.t2413 a_400_62400# 0.03fF
C2152 VN.n1881 a_400_62400# 0.32fF
C2153 VN.n1882 a_400_62400# 0.48fF
C2154 VN.n1883 a_400_62400# 0.81fF
C2155 VN.n1884 a_400_62400# 0.16fF
C2156 VN.t1295 a_400_62400# 0.03fF
C2157 VN.n1885 a_400_62400# 0.19fF
C2158 VN.n1887 a_400_62400# 1.55fF
C2159 VN.n1888 a_400_62400# 0.29fF
C2160 VN.n1889 a_400_62400# 2.52fF
C2161 VN.t1585 a_400_62400# 0.03fF
C2162 VN.n1890 a_400_62400# 0.32fF
C2163 VN.n1891 a_400_62400# 1.22fF
C2164 VN.n1892 a_400_62400# 0.07fF
C2165 VN.t1476 a_400_62400# 0.03fF
C2166 VN.n1893 a_400_62400# 0.16fF
C2167 VN.n1894 a_400_62400# 0.19fF
C2168 VN.n1896 a_400_62400# 27.83fF
C2169 VN.n1897 a_400_62400# 3.93fF
C2170 VN.n1898 a_400_62400# 2.51fF
C2171 VN.n1899 a_400_62400# 0.16fF
C2172 VN.t1749 a_400_62400# 0.03fF
C2173 VN.n1900 a_400_62400# 0.19fF
C2174 VN.t382 a_400_62400# 0.03fF
C2175 VN.n1902 a_400_62400# 0.32fF
C2176 VN.n1903 a_400_62400# 0.48fF
C2177 VN.n1904 a_400_62400# 0.81fF
C2178 VN.n1905 a_400_62400# 1.46fF
C2179 VN.n1906 a_400_62400# 0.21fF
C2180 VN.n1907 a_400_62400# 2.81fF
C2181 VN.t1954 a_400_62400# 0.03fF
C2182 VN.n1908 a_400_62400# 0.16fF
C2183 VN.n1909 a_400_62400# 0.19fF
C2184 VN.t2072 a_400_62400# 0.03fF
C2185 VN.n1911 a_400_62400# 0.32fF
C2186 VN.n1912 a_400_62400# 1.22fF
C2187 VN.n1913 a_400_62400# 0.07fF
C2188 VN.n1914 a_400_62400# 2.51fF
C2189 VN.n1915 a_400_62400# 3.57fF
C2190 VN.t2036 a_400_62400# 0.03fF
C2191 VN.n1916 a_400_62400# 0.32fF
C2192 VN.n1917 a_400_62400# 0.48fF
C2193 VN.n1918 a_400_62400# 0.81fF
C2194 VN.n1919 a_400_62400# 0.16fF
C2195 VN.t876 a_400_62400# 0.03fF
C2196 VN.n1920 a_400_62400# 0.19fF
C2197 VN.n1922 a_400_62400# 3.93fF
C2198 VN.n1923 a_400_62400# 3.08fF
C2199 VN.t1086 a_400_62400# 0.03fF
C2200 VN.n1924 a_400_62400# 0.16fF
C2201 VN.n1925 a_400_62400# 0.19fF
C2202 VN.t1201 a_400_62400# 0.03fF
C2203 VN.n1927 a_400_62400# 0.32fF
C2204 VN.n1928 a_400_62400# 1.22fF
C2205 VN.n1929 a_400_62400# 0.07fF
C2206 VN.n1930 a_400_62400# 2.51fF
C2207 VN.n1931 a_400_62400# 3.57fF
C2208 VN.t1162 a_400_62400# 0.03fF
C2209 VN.n1932 a_400_62400# 0.32fF
C2210 VN.n1933 a_400_62400# 0.48fF
C2211 VN.n1934 a_400_62400# 0.81fF
C2212 VN.n1935 a_400_62400# 0.16fF
C2213 VN.t134 a_400_62400# 0.03fF
C2214 VN.n1936 a_400_62400# 0.19fF
C2215 VN.n1938 a_400_62400# 3.75fF
C2216 VN.n1939 a_400_62400# 3.08fF
C2217 VN.t213 a_400_62400# 0.03fF
C2218 VN.n1940 a_400_62400# 0.16fF
C2219 VN.n1941 a_400_62400# 0.19fF
C2220 VN.t333 a_400_62400# 0.03fF
C2221 VN.n1943 a_400_62400# 0.32fF
C2222 VN.n1944 a_400_62400# 1.22fF
C2223 VN.n1945 a_400_62400# 0.07fF
C2224 VN.n1946 a_400_62400# 2.51fF
C2225 VN.n1947 a_400_62400# 3.57fF
C2226 VN.t437 a_400_62400# 0.03fF
C2227 VN.n1948 a_400_62400# 0.32fF
C2228 VN.n1949 a_400_62400# 0.48fF
C2229 VN.n1950 a_400_62400# 0.81fF
C2230 VN.n1951 a_400_62400# 0.16fF
C2231 VN.t1796 a_400_62400# 0.03fF
C2232 VN.n1952 a_400_62400# 0.19fF
C2233 VN.n1954 a_400_62400# 3.75fF
C2234 VN.n1955 a_400_62400# 3.08fF
C2235 VN.t1863 a_400_62400# 0.03fF
C2236 VN.n1956 a_400_62400# 0.16fF
C2237 VN.n1957 a_400_62400# 0.19fF
C2238 VN.t2123 a_400_62400# 0.03fF
C2239 VN.n1959 a_400_62400# 0.32fF
C2240 VN.n1960 a_400_62400# 1.22fF
C2241 VN.n1961 a_400_62400# 0.07fF
C2242 VN.n1962 a_400_62400# 2.51fF
C2243 VN.n1963 a_400_62400# 3.57fF
C2244 VN.t2082 a_400_62400# 0.03fF
C2245 VN.n1964 a_400_62400# 0.32fF
C2246 VN.n1965 a_400_62400# 0.48fF
C2247 VN.n1966 a_400_62400# 0.81fF
C2248 VN.n1967 a_400_62400# 0.16fF
C2249 VN.t921 a_400_62400# 0.03fF
C2250 VN.n1968 a_400_62400# 0.19fF
C2251 VN.n1970 a_400_62400# 3.75fF
C2252 VN.n1971 a_400_62400# 3.08fF
C2253 VN.t993 a_400_62400# 0.03fF
C2254 VN.n1972 a_400_62400# 0.16fF
C2255 VN.n1973 a_400_62400# 0.19fF
C2256 VN.t1248 a_400_62400# 0.03fF
C2257 VN.n1975 a_400_62400# 0.32fF
C2258 VN.n1976 a_400_62400# 1.22fF
C2259 VN.n1977 a_400_62400# 0.07fF
C2260 VN.n1978 a_400_62400# 2.51fF
C2261 VN.n1979 a_400_62400# 3.57fF
C2262 VN.t1208 a_400_62400# 0.03fF
C2263 VN.n1980 a_400_62400# 0.32fF
C2264 VN.n1981 a_400_62400# 0.48fF
C2265 VN.n1982 a_400_62400# 0.81fF
C2266 VN.n1983 a_400_62400# 0.16fF
C2267 VN.t2582 a_400_62400# 0.03fF
C2268 VN.n1984 a_400_62400# 0.19fF
C2269 VN.n1986 a_400_62400# 3.75fF
C2270 VN.n1987 a_400_62400# 3.08fF
C2271 VN.t109 a_400_62400# 0.03fF
C2272 VN.n1988 a_400_62400# 0.16fF
C2273 VN.n1989 a_400_62400# 0.19fF
C2274 VN.t380 a_400_62400# 0.03fF
C2275 VN.n1991 a_400_62400# 0.32fF
C2276 VN.n1992 a_400_62400# 1.22fF
C2277 VN.n1993 a_400_62400# 0.07fF
C2278 VN.n1994 a_400_62400# 2.51fF
C2279 VN.n1995 a_400_62400# 3.57fF
C2280 VN.t345 a_400_62400# 0.03fF
C2281 VN.n1996 a_400_62400# 0.32fF
C2282 VN.n1997 a_400_62400# 0.48fF
C2283 VN.n1998 a_400_62400# 0.81fF
C2284 VN.n1999 a_400_62400# 0.16fF
C2285 VN.t1713 a_400_62400# 0.03fF
C2286 VN.n2000 a_400_62400# 0.19fF
C2287 VN.n2002 a_400_62400# 3.75fF
C2288 VN.n2003 a_400_62400# 3.08fF
C2289 VN.t1778 a_400_62400# 0.03fF
C2290 VN.n2004 a_400_62400# 0.16fF
C2291 VN.n2005 a_400_62400# 0.19fF
C2292 VN.t2034 a_400_62400# 0.03fF
C2293 VN.n2007 a_400_62400# 0.32fF
C2294 VN.n2008 a_400_62400# 1.22fF
C2295 VN.n2009 a_400_62400# 0.07fF
C2296 VN.n2010 a_400_62400# 2.51fF
C2297 VN.n2011 a_400_62400# 3.57fF
C2298 VN.t1988 a_400_62400# 0.03fF
C2299 VN.n2012 a_400_62400# 0.32fF
C2300 VN.n2013 a_400_62400# 0.48fF
C2301 VN.n2014 a_400_62400# 0.81fF
C2302 VN.n2015 a_400_62400# 0.16fF
C2303 VN.t841 a_400_62400# 0.03fF
C2304 VN.n2016 a_400_62400# 0.19fF
C2305 VN.n2018 a_400_62400# 3.75fF
C2306 VN.n2019 a_400_62400# 3.08fF
C2307 VN.t1036 a_400_62400# 0.03fF
C2308 VN.n2020 a_400_62400# 0.16fF
C2309 VN.n2021 a_400_62400# 0.19fF
C2310 VN.t1159 a_400_62400# 0.03fF
C2311 VN.n2023 a_400_62400# 0.32fF
C2312 VN.n2024 a_400_62400# 1.22fF
C2313 VN.n2025 a_400_62400# 0.07fF
C2314 VN.n2026 a_400_62400# 2.51fF
C2315 VN.n2027 a_400_62400# 3.57fF
C2316 VN.t1115 a_400_62400# 0.03fF
C2317 VN.n2028 a_400_62400# 0.32fF
C2318 VN.n2029 a_400_62400# 0.48fF
C2319 VN.n2030 a_400_62400# 0.81fF
C2320 VN.n2031 a_400_62400# 0.16fF
C2321 VN.t2504 a_400_62400# 0.03fF
C2322 VN.n2032 a_400_62400# 0.19fF
C2323 VN.n2034 a_400_62400# 3.75fF
C2324 VN.n2035 a_400_62400# 3.08fF
C2325 VN.t164 a_400_62400# 0.03fF
C2326 VN.n2036 a_400_62400# 0.16fF
C2327 VN.n2037 a_400_62400# 0.19fF
C2328 VN.t292 a_400_62400# 0.03fF
C2329 VN.n2039 a_400_62400# 0.32fF
C2330 VN.n2040 a_400_62400# 1.22fF
C2331 VN.n2041 a_400_62400# 0.07fF
C2332 VN.n2042 a_400_62400# 2.51fF
C2333 VN.n2043 a_400_62400# 3.57fF
C2334 VN.t1800 a_400_62400# 0.03fF
C2335 VN.n2044 a_400_62400# 0.32fF
C2336 VN.n2045 a_400_62400# 0.48fF
C2337 VN.n2046 a_400_62400# 0.81fF
C2338 VN.n2047 a_400_62400# 0.16fF
C2339 VN.t659 a_400_62400# 0.03fF
C2340 VN.n2048 a_400_62400# 0.19fF
C2341 VN.n2050 a_400_62400# 3.75fF
C2342 VN.n2051 a_400_62400# 3.08fF
C2343 VN.t840 a_400_62400# 0.03fF
C2344 VN.n2052 a_400_62400# 0.16fF
C2345 VN.n2053 a_400_62400# 0.19fF
C2346 VN.t1073 a_400_62400# 0.03fF
C2347 VN.n2055 a_400_62400# 0.32fF
C2348 VN.n2056 a_400_62400# 1.22fF
C2349 VN.n2057 a_400_62400# 0.07fF
C2350 VN.n2058 a_400_62400# 2.51fF
C2351 VN.n2059 a_400_62400# 3.57fF
C2352 VN.t923 a_400_62400# 0.03fF
C2353 VN.n2060 a_400_62400# 0.32fF
C2354 VN.n2061 a_400_62400# 0.48fF
C2355 VN.n2062 a_400_62400# 0.81fF
C2356 VN.n2063 a_400_62400# 0.16fF
C2357 VN.t2319 a_400_62400# 0.03fF
C2358 VN.n2064 a_400_62400# 0.19fF
C2359 VN.n2066 a_400_62400# 3.75fF
C2360 VN.n2067 a_400_62400# 3.08fF
C2361 VN.t2503 a_400_62400# 0.03fF
C2362 VN.n2068 a_400_62400# 0.16fF
C2363 VN.n2069 a_400_62400# 0.19fF
C2364 VN.t198 a_400_62400# 0.03fF
C2365 VN.n2071 a_400_62400# 0.32fF
C2366 VN.n2072 a_400_62400# 1.22fF
C2367 VN.n2073 a_400_62400# 0.07fF
C2368 VN.n2074 a_400_62400# 3.65fF
C2369 VN.n2075 a_400_62400# 2.14fF
C2370 VN.n2076 a_400_62400# 0.16fF
C2371 VN.t704 a_400_62400# 0.03fF
C2372 VN.n2077 a_400_62400# 0.19fF
C2373 VN.t1715 a_400_62400# 0.03fF
C2374 VN.n2079 a_400_62400# 0.32fF
C2375 VN.n2080 a_400_62400# 0.48fF
C2376 VN.n2081 a_400_62400# 0.81fF
C2377 VN.n2082 a_400_62400# 0.09fF
C2378 VN.n2083 a_400_62400# 0.01fF
C2379 VN.n2084 a_400_62400# 0.02fF
C2380 VN.n2085 a_400_62400# 0.02fF
C2381 VN.n2086 a_400_62400# 0.32fF
C2382 VN.n2087 a_400_62400# 1.56fF
C2383 VN.n2088 a_400_62400# 1.81fF
C2384 VN.n2089 a_400_62400# 3.08fF
C2385 VN.t769 a_400_62400# 0.03fF
C2386 VN.n2090 a_400_62400# 0.16fF
C2387 VN.n2091 a_400_62400# 0.19fF
C2388 VN.t986 a_400_62400# 0.03fF
C2389 VN.n2093 a_400_62400# 0.32fF
C2390 VN.n2094 a_400_62400# 1.22fF
C2391 VN.n2095 a_400_62400# 0.07fF
C2392 VN.t108 a_400_62400# 64.69fF
C2393 VN.t1855 a_400_62400# 0.03fF
C2394 VN.n2096 a_400_62400# 0.32fF
C2395 VN.n2097 a_400_62400# 1.22fF
C2396 VN.n2098 a_400_62400# 0.07fF
C2397 VN.t1641 a_400_62400# 0.03fF
C2398 VN.n2099 a_400_62400# 0.16fF
C2399 VN.n2100 a_400_62400# 0.19fF
C2400 VN.n2102 a_400_62400# 0.16fF
C2401 VN.t1451 a_400_62400# 0.03fF
C2402 VN.n2103 a_400_62400# 0.19fF
C2403 VN.n2105 a_400_62400# 6.92fF
C2404 VN.n2106 a_400_62400# 6.56fF
C2405 VN.t264 a_400_62400# 0.03fF
C2406 VN.n2107 a_400_62400# 0.16fF
C2407 VN.n2108 a_400_62400# 0.19fF
C2408 VN.t263 a_400_62400# 0.03fF
C2409 VN.n2110 a_400_62400# 0.32fF
C2410 VN.n2111 a_400_62400# 1.22fF
C2411 VN.n2112 a_400_62400# 0.07fF
C2412 VN.n2113 a_400_62400# 2.51fF
C2413 VN.n2114 a_400_62400# 3.58fF
C2414 VN.t2397 a_400_62400# 0.03fF
C2415 VN.n2115 a_400_62400# 0.32fF
C2416 VN.n2116 a_400_62400# 0.48fF
C2417 VN.n2117 a_400_62400# 0.81fF
C2418 VN.n2118 a_400_62400# 0.16fF
C2419 VN.t1253 a_400_62400# 0.03fF
C2420 VN.n2119 a_400_62400# 0.19fF
C2421 VN.n2121 a_400_62400# 7.29fF
C2422 VN.t1914 a_400_62400# 0.03fF
C2423 VN.n2122 a_400_62400# 0.16fF
C2424 VN.n2123 a_400_62400# 0.19fF
C2425 VN.t1913 a_400_62400# 0.03fF
C2426 VN.n2125 a_400_62400# 0.32fF
C2427 VN.n2126 a_400_62400# 1.22fF
C2428 VN.n2127 a_400_62400# 0.07fF
C2429 VN.t224 a_400_62400# 64.17fF
C2430 VN.t1039 a_400_62400# 0.03fF
C2431 VN.n2128 a_400_62400# 1.60fF
C2432 VN.n2129 a_400_62400# 0.07fF
C2433 VN.t1182 a_400_62400# 0.03fF
C2434 VN.n2130 a_400_62400# 0.02fF
C2435 VN.n2131 a_400_62400# 0.34fF
C2436 VN.n2133 a_400_62400# 2.01fF
C2437 VN.n2134 a_400_62400# 1.75fF
C2438 VN.n2135 a_400_62400# 0.37fF
C2439 VN.n2136 a_400_62400# 0.33fF
C2440 VN.n2137 a_400_62400# 5.88fF
C2441 VN.n2138 a_400_62400# 0.02fF
C2442 VN.n2139 a_400_62400# 0.02fF
C2443 VN.n2140 a_400_62400# 0.03fF
C2444 VN.n2141 a_400_62400# 0.05fF
C2445 VN.n2142 a_400_62400# 0.23fF
C2446 VN.n2143 a_400_62400# 0.02fF
C2447 VN.n2144 a_400_62400# 0.03fF
C2448 VN.n2145 a_400_62400# 0.01fF
C2449 VN.n2146 a_400_62400# 0.01fF
C2450 VN.n2147 a_400_62400# 0.01fF
C2451 VN.n2148 a_400_62400# 0.02fF
C2452 VN.n2149 a_400_62400# 0.03fF
C2453 VN.n2150 a_400_62400# 0.06fF
C2454 VN.n2151 a_400_62400# 0.05fF
C2455 VN.n2152 a_400_62400# 0.15fF
C2456 VN.n2153 a_400_62400# 0.51fF
C2457 VN.n2154 a_400_62400# 0.27fF
C2458 VN.n2155 a_400_62400# 37.46fF
C2459 VN.n2156 a_400_62400# 37.46fF
C2460 VN.n2157 a_400_62400# 0.79fF
C2461 VN.n2158 a_400_62400# 0.23fF
C2462 VN.n2159 a_400_62400# 1.18fF
C2463 VN.t92 a_400_62400# 28.64fF
C2464 VN.n2160 a_400_62400# 0.79fF
C2465 VN.n2161 a_400_62400# 0.11fF
C2466 VN.n2162 a_400_62400# 4.98fF
C2467 VN.n2163 a_400_62400# 0.80fF
C2468 VN.n2164 a_400_62400# 0.29fF
C2469 VN.n2165 a_400_62400# 1.96fF
C2470 VN.n2167 a_400_62400# 25.18fF
C2471 VN.n2169 a_400_62400# 1.87fF
C2472 VN.n2170 a_400_62400# 5.36fF
C2473 VN.n2171 a_400_62400# 1.81fF
C2474 VN.t324 a_400_62400# 0.03fF
C2475 VN.n2172 a_400_62400# 0.85fF
C2476 VN.n2173 a_400_62400# 0.81fF
C2477 VN.n2174 a_400_62400# 2.53fF
C2478 VN.n2175 a_400_62400# 0.09fF
C2479 VN.n2176 a_400_62400# 0.05fF
C2480 VN.n2177 a_400_62400# 0.07fF
C2481 VN.n2178 a_400_62400# 1.16fF
C2482 VN.n2179 a_400_62400# 0.01fF
C2483 VN.n2180 a_400_62400# 0.01fF
C2484 VN.n2181 a_400_62400# 0.01fF
C2485 VN.n2182 a_400_62400# 0.09fF
C2486 VN.n2183 a_400_62400# 0.91fF
C2487 VN.n2184 a_400_62400# 0.96fF
C2488 VN.t851 a_400_62400# 0.03fF
C2489 VN.n2185 a_400_62400# 0.32fF
C2490 VN.n2186 a_400_62400# 0.48fF
C2491 VN.n2187 a_400_62400# 0.81fF
C2492 VN.n2188 a_400_62400# 0.16fF
C2493 VN.t2381 a_400_62400# 0.03fF
C2494 VN.n2189 a_400_62400# 0.19fF
C2495 VN.n2191 a_400_62400# 0.93fF
C2496 VN.n2192 a_400_62400# 0.30fF
C2497 VN.n2193 a_400_62400# 0.34fF
C2498 VN.n2194 a_400_62400# 0.12fF
C2499 VN.n2195 a_400_62400# 0.30fF
C2500 VN.n2196 a_400_62400# 0.93fF
C2501 VN.n2197 a_400_62400# 1.55fF
C2502 VN.n2198 a_400_62400# 0.29fF
C2503 VN.n2199 a_400_62400# 0.34fF
C2504 VN.n2200 a_400_62400# 0.12fF
C2505 VN.n2201 a_400_62400# 3.10fF
C2506 VN.t1981 a_400_62400# 0.03fF
C2507 VN.n2202 a_400_62400# 0.32fF
C2508 VN.n2203 a_400_62400# 1.22fF
C2509 VN.n2204 a_400_62400# 0.07fF
C2510 VN.t542 a_400_62400# 0.03fF
C2511 VN.n2205 a_400_62400# 0.16fF
C2512 VN.n2206 a_400_62400# 0.19fF
C2513 VN.n2208 a_400_62400# 2.51fF
C2514 VN.n2209 a_400_62400# 0.61fF
C2515 VN.n2210 a_400_62400# 0.30fF
C2516 VN.n2211 a_400_62400# 0.51fF
C2517 VN.n2212 a_400_62400# 0.21fF
C2518 VN.n2213 a_400_62400# 0.38fF
C2519 VN.n2214 a_400_62400# 0.29fF
C2520 VN.n2215 a_400_62400# 0.40fF
C2521 VN.n2216 a_400_62400# 0.28fF
C2522 VN.t93 a_400_62400# 0.03fF
C2523 VN.n2217 a_400_62400# 0.32fF
C2524 VN.n2218 a_400_62400# 0.48fF
C2525 VN.n2219 a_400_62400# 0.81fF
C2526 VN.n2220 a_400_62400# 0.16fF
C2527 VN.t1512 a_400_62400# 0.03fF
C2528 VN.n2221 a_400_62400# 0.19fF
C2529 VN.n2223 a_400_62400# 0.06fF
C2530 VN.n2224 a_400_62400# 0.04fF
C2531 VN.n2225 a_400_62400# 0.04fF
C2532 VN.n2226 a_400_62400# 0.14fF
C2533 VN.n2227 a_400_62400# 0.48fF
C2534 VN.n2228 a_400_62400# 0.50fF
C2535 VN.n2229 a_400_62400# 0.14fF
C2536 VN.n2230 a_400_62400# 0.16fF
C2537 VN.n2231 a_400_62400# 0.09fF
C2538 VN.n2232 a_400_62400# 0.16fF
C2539 VN.n2233 a_400_62400# 0.24fF
C2540 VN.n2234 a_400_62400# 5.35fF
C2541 VN.t1252 a_400_62400# 0.03fF
C2542 VN.n2235 a_400_62400# 0.32fF
C2543 VN.n2236 a_400_62400# 1.22fF
C2544 VN.n2237 a_400_62400# 0.07fF
C2545 VN.t2197 a_400_62400# 0.03fF
C2546 VN.n2238 a_400_62400# 0.16fF
C2547 VN.n2239 a_400_62400# 0.19fF
C2548 VN.n2241 a_400_62400# 0.33fF
C2549 VN.n2242 a_400_62400# 0.12fF
C2550 VN.n2243 a_400_62400# 0.28fF
C2551 VN.n2244 a_400_62400# 1.72fF
C2552 VN.n2245 a_400_62400# 0.71fF
C2553 VN.n2246 a_400_62400# 2.51fF
C2554 VN.n2247 a_400_62400# 0.16fF
C2555 VN.t644 a_400_62400# 0.03fF
C2556 VN.n2248 a_400_62400# 0.19fF
C2557 VN.t1768 a_400_62400# 0.03fF
C2558 VN.n2250 a_400_62400# 0.32fF
C2559 VN.n2251 a_400_62400# 0.48fF
C2560 VN.n2252 a_400_62400# 0.81fF
C2561 VN.n2253 a_400_62400# 0.95fF
C2562 VN.n2254 a_400_62400# 2.11fF
C2563 VN.n2255 a_400_62400# 3.28fF
C2564 VN.t383 a_400_62400# 0.03fF
C2565 VN.n2256 a_400_62400# 0.32fF
C2566 VN.n2257 a_400_62400# 1.22fF
C2567 VN.n2258 a_400_62400# 0.07fF
C2568 VN.t1326 a_400_62400# 0.03fF
C2569 VN.n2259 a_400_62400# 0.16fF
C2570 VN.n2260 a_400_62400# 0.19fF
C2571 VN.n2262 a_400_62400# 2.53fF
C2572 VN.n2263 a_400_62400# 0.08fF
C2573 VN.n2264 a_400_62400# 0.04fF
C2574 VN.n2265 a_400_62400# 0.05fF
C2575 VN.n2266 a_400_62400# 1.33fF
C2576 VN.n2267 a_400_62400# 0.03fF
C2577 VN.n2268 a_400_62400# 0.01fF
C2578 VN.n2269 a_400_62400# 0.02fF
C2579 VN.n2270 a_400_62400# 0.11fF
C2580 VN.n2271 a_400_62400# 0.48fF
C2581 VN.n2272 a_400_62400# 2.48fF
C2582 VN.t2261 a_400_62400# 0.03fF
C2583 VN.n2273 a_400_62400# 0.32fF
C2584 VN.n2274 a_400_62400# 0.48fF
C2585 VN.n2275 a_400_62400# 0.81fF
C2586 VN.n2276 a_400_62400# 0.16fF
C2587 VN.t1113 a_400_62400# 0.03fF
C2588 VN.n2277 a_400_62400# 0.19fF
C2589 VN.n2279 a_400_62400# 0.93fF
C2590 VN.n2280 a_400_62400# 0.30fF
C2591 VN.n2281 a_400_62400# 0.34fF
C2592 VN.n2282 a_400_62400# 0.12fF
C2593 VN.n2283 a_400_62400# 0.30fF
C2594 VN.n2284 a_400_62400# 0.93fF
C2595 VN.n2285 a_400_62400# 1.55fF
C2596 VN.n2286 a_400_62400# 0.29fF
C2597 VN.n2287 a_400_62400# 0.34fF
C2598 VN.n2288 a_400_62400# 0.12fF
C2599 VN.n2289 a_400_62400# 2.52fF
C2600 VN.t842 a_400_62400# 0.03fF
C2601 VN.n2290 a_400_62400# 0.32fF
C2602 VN.n2291 a_400_62400# 1.22fF
C2603 VN.n2292 a_400_62400# 0.07fF
C2604 VN.t465 a_400_62400# 0.03fF
C2605 VN.n2293 a_400_62400# 0.16fF
C2606 VN.n2294 a_400_62400# 0.19fF
C2607 VN.n2296 a_400_62400# 27.83fF
C2608 VN.n2297 a_400_62400# 0.09fF
C2609 VN.n2298 a_400_62400# 0.27fF
C2610 VN.n2299 a_400_62400# 0.12fF
C2611 VN.n2300 a_400_62400# 0.28fF
C2612 VN.n2301 a_400_62400# 0.13fF
C2613 VN.n2302 a_400_62400# 0.40fF
C2614 VN.n2303 a_400_62400# 0.93fF
C2615 VN.n2304 a_400_62400# 0.60fF
C2616 VN.n2305 a_400_62400# 3.12fF
C2617 VN.n2306 a_400_62400# 0.16fF
C2618 VN.t603 a_400_62400# 0.03fF
C2619 VN.n2307 a_400_62400# 0.19fF
C2620 VN.t1726 a_400_62400# 0.03fF
C2621 VN.n2309 a_400_62400# 0.32fF
C2622 VN.n2310 a_400_62400# 0.48fF
C2623 VN.n2311 a_400_62400# 0.81fF
C2624 VN.n2312 a_400_62400# 2.54fF
C2625 VN.n2313 a_400_62400# 0.23fF
C2626 VN.n2314 a_400_62400# 1.02fF
C2627 VN.n2315 a_400_62400# 0.42fF
C2628 VN.n2316 a_400_62400# 0.34fF
C2629 VN.n2317 a_400_62400# 0.40fF
C2630 VN.n2318 a_400_62400# 0.63fF
C2631 VN.n2319 a_400_62400# 0.21fF
C2632 VN.n2320 a_400_62400# 2.58fF
C2633 VN.t1404 a_400_62400# 0.03fF
C2634 VN.n2321 a_400_62400# 0.16fF
C2635 VN.n2322 a_400_62400# 0.19fF
C2636 VN.t338 a_400_62400# 0.03fF
C2637 VN.n2324 a_400_62400# 0.32fF
C2638 VN.n2325 a_400_62400# 1.22fF
C2639 VN.n2326 a_400_62400# 0.07fF
C2640 VN.n2327 a_400_62400# 2.51fF
C2641 VN.n2328 a_400_62400# 0.16fF
C2642 VN.t249 a_400_62400# 0.03fF
C2643 VN.n2329 a_400_62400# 0.19fF
C2644 VN.t1396 a_400_62400# 0.03fF
C2645 VN.n2331 a_400_62400# 0.32fF
C2646 VN.n2332 a_400_62400# 0.48fF
C2647 VN.n2333 a_400_62400# 0.81fF
C2648 VN.n2334 a_400_62400# 1.24fF
C2649 VN.n2335 a_400_62400# 0.43fF
C2650 VN.n2336 a_400_62400# 0.43fF
C2651 VN.n2337 a_400_62400# 1.24fF
C2652 VN.n2338 a_400_62400# 1.46fF
C2653 VN.n2339 a_400_62400# 0.21fF
C2654 VN.n2340 a_400_62400# 6.64fF
C2655 VN.t910 a_400_62400# 0.03fF
C2656 VN.n2341 a_400_62400# 0.16fF
C2657 VN.n2342 a_400_62400# 0.19fF
C2658 VN.t2506 a_400_62400# 0.03fF
C2659 VN.n2344 a_400_62400# 0.32fF
C2660 VN.n2345 a_400_62400# 1.22fF
C2661 VN.n2346 a_400_62400# 0.07fF
C2662 VN.n2347 a_400_62400# 2.51fF
C2663 VN.n2348 a_400_62400# 3.57fF
C2664 VN.t534 a_400_62400# 0.03fF
C2665 VN.n2349 a_400_62400# 0.32fF
C2666 VN.n2350 a_400_62400# 0.48fF
C2667 VN.n2351 a_400_62400# 0.81fF
C2668 VN.n2352 a_400_62400# 0.16fF
C2669 VN.t1899 a_400_62400# 0.03fF
C2670 VN.n2353 a_400_62400# 0.19fF
C2671 VN.n2355 a_400_62400# 6.91fF
C2672 VN.t2572 a_400_62400# 0.03fF
C2673 VN.n2356 a_400_62400# 0.16fF
C2674 VN.n2357 a_400_62400# 0.19fF
C2675 VN.t1643 a_400_62400# 0.03fF
C2676 VN.n2359 a_400_62400# 0.32fF
C2677 VN.n2360 a_400_62400# 1.22fF
C2678 VN.n2361 a_400_62400# 0.07fF
C2679 VN.n2362 a_400_62400# 2.51fF
C2680 VN.n2363 a_400_62400# 3.57fF
C2681 VN.t2189 a_400_62400# 0.03fF
C2682 VN.n2364 a_400_62400# 0.32fF
C2683 VN.n2365 a_400_62400# 0.48fF
C2684 VN.n2366 a_400_62400# 0.81fF
C2685 VN.n2367 a_400_62400# 0.16fF
C2686 VN.t1024 a_400_62400# 0.03fF
C2687 VN.n2368 a_400_62400# 0.19fF
C2688 VN.n2370 a_400_62400# 6.92fF
C2689 VN.t1833 a_400_62400# 0.03fF
C2690 VN.n2371 a_400_62400# 0.16fF
C2691 VN.n2372 a_400_62400# 0.19fF
C2692 VN.t772 a_400_62400# 0.03fF
C2693 VN.n2374 a_400_62400# 0.32fF
C2694 VN.n2375 a_400_62400# 1.22fF
C2695 VN.n2376 a_400_62400# 0.07fF
C2696 VN.n2377 a_400_62400# 2.51fF
C2697 VN.n2378 a_400_62400# 3.57fF
C2698 VN.t1322 a_400_62400# 0.03fF
C2699 VN.n2379 a_400_62400# 0.32fF
C2700 VN.n2380 a_400_62400# 0.48fF
C2701 VN.n2381 a_400_62400# 0.81fF
C2702 VN.n2382 a_400_62400# 0.16fF
C2703 VN.t152 a_400_62400# 0.03fF
C2704 VN.n2383 a_400_62400# 0.19fF
C2705 VN.n2385 a_400_62400# 6.92fF
C2706 VN.t958 a_400_62400# 0.03fF
C2707 VN.n2386 a_400_62400# 0.16fF
C2708 VN.n2387 a_400_62400# 0.19fF
C2709 VN.t2424 a_400_62400# 0.03fF
C2710 VN.n2389 a_400_62400# 0.32fF
C2711 VN.n2390 a_400_62400# 1.22fF
C2712 VN.n2391 a_400_62400# 0.07fF
C2713 VN.n2392 a_400_62400# 2.51fF
C2714 VN.n2393 a_400_62400# 3.57fF
C2715 VN.t460 a_400_62400# 0.03fF
C2716 VN.n2394 a_400_62400# 0.32fF
C2717 VN.n2395 a_400_62400# 0.48fF
C2718 VN.n2396 a_400_62400# 0.81fF
C2719 VN.n2397 a_400_62400# 0.16fF
C2720 VN.t1816 a_400_62400# 0.03fF
C2721 VN.n2398 a_400_62400# 0.19fF
C2722 VN.n2400 a_400_62400# 6.92fF
C2723 VN.t50 a_400_62400# 0.03fF
C2724 VN.n2401 a_400_62400# 0.16fF
C2725 VN.n2402 a_400_62400# 0.19fF
C2726 VN.t1562 a_400_62400# 0.03fF
C2727 VN.n2404 a_400_62400# 0.32fF
C2728 VN.n2405 a_400_62400# 1.22fF
C2729 VN.n2406 a_400_62400# 0.07fF
C2730 VN.n2407 a_400_62400# 2.51fF
C2731 VN.n2408 a_400_62400# 3.57fF
C2732 VN.t2108 a_400_62400# 0.03fF
C2733 VN.n2409 a_400_62400# 0.32fF
C2734 VN.n2410 a_400_62400# 0.48fF
C2735 VN.n2411 a_400_62400# 0.81fF
C2736 VN.n2412 a_400_62400# 0.16fF
C2737 VN.t941 a_400_62400# 0.03fF
C2738 VN.n2413 a_400_62400# 0.19fF
C2739 VN.n2415 a_400_62400# 6.92fF
C2740 VN.t1746 a_400_62400# 0.03fF
C2741 VN.n2416 a_400_62400# 0.16fF
C2742 VN.n2417 a_400_62400# 0.19fF
C2743 VN.t692 a_400_62400# 0.03fF
C2744 VN.n2419 a_400_62400# 0.32fF
C2745 VN.n2420 a_400_62400# 1.22fF
C2746 VN.n2421 a_400_62400# 0.07fF
C2747 VN.n2422 a_400_62400# 2.51fF
C2748 VN.n2423 a_400_62400# 3.57fF
C2749 VN.t1231 a_400_62400# 0.03fF
C2750 VN.n2424 a_400_62400# 0.32fF
C2751 VN.n2425 a_400_62400# 0.48fF
C2752 VN.n2426 a_400_62400# 0.81fF
C2753 VN.n2427 a_400_62400# 0.16fF
C2754 VN.t208 a_400_62400# 0.03fF
C2755 VN.n2428 a_400_62400# 0.19fF
C2756 VN.n2430 a_400_62400# 6.92fF
C2757 VN.t872 a_400_62400# 0.03fF
C2758 VN.n2431 a_400_62400# 0.16fF
C2759 VN.n2432 a_400_62400# 0.19fF
C2760 VN.t2350 a_400_62400# 0.03fF
C2761 VN.n2434 a_400_62400# 0.32fF
C2762 VN.n2435 a_400_62400# 1.22fF
C2763 VN.n2436 a_400_62400# 0.07fF
C2764 VN.n2437 a_400_62400# 2.51fF
C2765 VN.n2438 a_400_62400# 3.57fF
C2766 VN.t498 a_400_62400# 0.03fF
C2767 VN.n2439 a_400_62400# 0.32fF
C2768 VN.n2440 a_400_62400# 0.48fF
C2769 VN.n2441 a_400_62400# 0.81fF
C2770 VN.n2442 a_400_62400# 0.16fF
C2771 VN.t1858 a_400_62400# 0.03fF
C2772 VN.n2443 a_400_62400# 0.19fF
C2773 VN.n2445 a_400_62400# 6.92fF
C2774 VN.t2534 a_400_62400# 0.03fF
C2775 VN.n2446 a_400_62400# 0.16fF
C2776 VN.n2447 a_400_62400# 0.19fF
C2777 VN.t1603 a_400_62400# 0.03fF
C2778 VN.n2449 a_400_62400# 0.32fF
C2779 VN.n2450 a_400_62400# 1.22fF
C2780 VN.n2451 a_400_62400# 0.07fF
C2781 VN.n2452 a_400_62400# 2.51fF
C2782 VN.n2453 a_400_62400# 3.57fF
C2783 VN.t1285 a_400_62400# 0.03fF
C2784 VN.n2454 a_400_62400# 0.32fF
C2785 VN.n2455 a_400_62400# 0.48fF
C2786 VN.n2456 a_400_62400# 0.81fF
C2787 VN.n2457 a_400_62400# 0.16fF
C2788 VN.t86 a_400_62400# 0.03fF
C2789 VN.n2458 a_400_62400# 0.19fF
C2790 VN.n2460 a_400_62400# 6.92fF
C2791 VN.t1670 a_400_62400# 0.03fF
C2792 VN.n2461 a_400_62400# 0.16fF
C2793 VN.n2462 a_400_62400# 0.19fF
C2794 VN.t323 a_400_62400# 0.03fF
C2795 VN.n2464 a_400_62400# 0.32fF
C2796 VN.n2465 a_400_62400# 1.22fF
C2797 VN.n2466 a_400_62400# 0.07fF
C2798 VN.n2467 a_400_62400# 2.51fF
C2799 VN.n2468 a_400_62400# 3.57fF
C2800 VN.t417 a_400_62400# 0.03fF
C2801 VN.n2469 a_400_62400# 0.32fF
C2802 VN.n2470 a_400_62400# 0.48fF
C2803 VN.n2471 a_400_62400# 0.81fF
C2804 VN.n2472 a_400_62400# 0.16fF
C2805 VN.t1766 a_400_62400# 0.03fF
C2806 VN.n2473 a_400_62400# 0.19fF
C2807 VN.n2475 a_400_62400# 6.92fF
C2808 VN.t2447 a_400_62400# 0.03fF
C2809 VN.n2476 a_400_62400# 0.16fF
C2810 VN.n2477 a_400_62400# 0.19fF
C2811 VN.t1970 a_400_62400# 0.03fF
C2812 VN.n2479 a_400_62400# 0.32fF
C2813 VN.n2480 a_400_62400# 1.22fF
C2814 VN.n2481 a_400_62400# 0.07fF
C2815 VN.n2482 a_400_62400# 2.51fF
C2816 VN.n2483 a_400_62400# 3.57fF
C2817 VN.t2065 a_400_62400# 0.03fF
C2818 VN.n2484 a_400_62400# 0.32fF
C2819 VN.n2485 a_400_62400# 0.48fF
C2820 VN.n2486 a_400_62400# 0.81fF
C2821 VN.n2487 a_400_62400# 0.16fF
C2822 VN.t895 a_400_62400# 0.03fF
C2823 VN.n2488 a_400_62400# 0.19fF
C2824 VN.n2490 a_400_62400# 2.51fF
C2825 VN.n2491 a_400_62400# 3.59fF
C2826 VN.t897 a_400_62400# 0.03fF
C2827 VN.n2492 a_400_62400# 0.32fF
C2828 VN.n2493 a_400_62400# 0.48fF
C2829 VN.n2494 a_400_62400# 0.81fF
C2830 VN.t1127 a_400_62400# 0.03fF
C2831 VN.n2495 a_400_62400# 1.63fF
C2832 VN.n2496 a_400_62400# 0.81fF
C2833 VN.n2497 a_400_62400# 1.21fF
C2834 VN.n2498 a_400_62400# 1.54fF
C2835 VN.n2499 a_400_62400# 4.06fF
C2836 VN.t97 a_400_62400# 28.64fF
C2837 VN.n2500 a_400_62400# 28.43fF
C2838 VN.n2502 a_400_62400# 0.50fF
C2839 VN.n2503 a_400_62400# 0.31fF
C2840 VN.n2504 a_400_62400# 3.88fF
C2841 VN.n2505 a_400_62400# 3.29fF
C2842 VN.n2506 a_400_62400# 2.62fF
C2843 VN.n2507 a_400_62400# 5.27fF
C2844 VN.n2508 a_400_62400# 0.34fF
C2845 VN.n2509 a_400_62400# 0.02fF
C2846 VN.t2514 a_400_62400# 0.03fF
C2847 VN.n2510 a_400_62400# 0.34fF
C2848 VN.t304 a_400_62400# 0.03fF
C2849 VN.n2511 a_400_62400# 1.28fF
C2850 VN.n2512 a_400_62400# 0.94fF
C2851 VN.n2513 a_400_62400# 1.04fF
C2852 VN.n2514 a_400_62400# 2.58fF
C2853 VN.n2515 a_400_62400# 2.51fF
C2854 VN.n2516 a_400_62400# 0.16fF
C2855 VN.t1651 a_400_62400# 0.03fF
C2856 VN.n2517 a_400_62400# 0.19fF
C2857 VN.t261 a_400_62400# 0.03fF
C2858 VN.n2519 a_400_62400# 0.32fF
C2859 VN.n2520 a_400_62400# 0.48fF
C2860 VN.n2521 a_400_62400# 0.81fF
C2861 VN.n2522 a_400_62400# 2.03fF
C2862 VN.n2523 a_400_62400# 4.01fF
C2863 VN.t1951 a_400_62400# 0.03fF
C2864 VN.n2524 a_400_62400# 0.32fF
C2865 VN.n2525 a_400_62400# 1.22fF
C2866 VN.n2526 a_400_62400# 0.07fF
C2867 VN.t1704 a_400_62400# 0.03fF
C2868 VN.n2527 a_400_62400# 0.16fF
C2869 VN.n2528 a_400_62400# 0.19fF
C2870 VN.n2530 a_400_62400# 2.53fF
C2871 VN.n2531 a_400_62400# 2.34fF
C2872 VN.t1911 a_400_62400# 0.03fF
C2873 VN.n2532 a_400_62400# 0.32fF
C2874 VN.n2533 a_400_62400# 0.48fF
C2875 VN.n2534 a_400_62400# 0.81fF
C2876 VN.n2535 a_400_62400# 0.16fF
C2877 VN.t779 a_400_62400# 0.03fF
C2878 VN.n2536 a_400_62400# 0.19fF
C2879 VN.n2538 a_400_62400# 1.55fF
C2880 VN.n2539 a_400_62400# 0.29fF
C2881 VN.n2540 a_400_62400# 3.27fF
C2882 VN.t1082 a_400_62400# 0.03fF
C2883 VN.n2541 a_400_62400# 0.32fF
C2884 VN.n2542 a_400_62400# 1.22fF
C2885 VN.n2543 a_400_62400# 0.07fF
C2886 VN.t964 a_400_62400# 0.03fF
C2887 VN.n2544 a_400_62400# 0.16fF
C2888 VN.n2545 a_400_62400# 0.19fF
C2889 VN.n2547 a_400_62400# 2.51fF
C2890 VN.n2548 a_400_62400# 0.56fF
C2891 VN.n2549 a_400_62400# 0.64fF
C2892 VN.n2550 a_400_62400# 0.12fF
C2893 VN.n2551 a_400_62400# 0.44fF
C2894 VN.n2552 a_400_62400# 0.40fF
C2895 VN.n2553 a_400_62400# 1.03fF
C2896 VN.n2554 a_400_62400# 0.79fF
C2897 VN.t1038 a_400_62400# 0.03fF
C2898 VN.n2555 a_400_62400# 0.32fF
C2899 VN.n2556 a_400_62400# 0.48fF
C2900 VN.n2557 a_400_62400# 0.81fF
C2901 VN.n2558 a_400_62400# 0.16fF
C2902 VN.t2430 a_400_62400# 0.03fF
C2903 VN.n2559 a_400_62400# 0.19fF
C2904 VN.n2561 a_400_62400# 3.50fF
C2905 VN.n2562 a_400_62400# 2.89fF
C2906 VN.t210 a_400_62400# 0.03fF
C2907 VN.n2563 a_400_62400# 0.32fF
C2908 VN.n2564 a_400_62400# 1.22fF
C2909 VN.n2565 a_400_62400# 0.07fF
C2910 VN.t58 a_400_62400# 0.03fF
C2911 VN.n2566 a_400_62400# 0.16fF
C2912 VN.n2567 a_400_62400# 0.19fF
C2913 VN.n2569 a_400_62400# 1.05fF
C2914 VN.n2570 a_400_62400# 3.07fF
C2915 VN.n2571 a_400_62400# 2.51fF
C2916 VN.n2572 a_400_62400# 0.16fF
C2917 VN.t1569 a_400_62400# 0.03fF
C2918 VN.n2573 a_400_62400# 0.19fF
C2919 VN.t166 a_400_62400# 0.03fF
C2920 VN.n2575 a_400_62400# 0.32fF
C2921 VN.n2576 a_400_62400# 0.48fF
C2922 VN.n2577 a_400_62400# 0.81fF
C2923 VN.n2578 a_400_62400# 1.86fF
C2924 VN.n2579 a_400_62400# 1.53fF
C2925 VN.n2580 a_400_62400# 0.47fF
C2926 VN.n2581 a_400_62400# 2.71fF
C2927 VN.t1861 a_400_62400# 0.03fF
C2928 VN.n2582 a_400_62400# 0.32fF
C2929 VN.n2583 a_400_62400# 1.22fF
C2930 VN.n2584 a_400_62400# 0.07fF
C2931 VN.t1750 a_400_62400# 0.03fF
C2932 VN.n2585 a_400_62400# 0.16fF
C2933 VN.n2586 a_400_62400# 0.19fF
C2934 VN.n2588 a_400_62400# 2.53fF
C2935 VN.n2589 a_400_62400# 2.51fF
C2936 VN.t662 a_400_62400# 0.03fF
C2937 VN.n2590 a_400_62400# 0.32fF
C2938 VN.n2591 a_400_62400# 0.48fF
C2939 VN.n2592 a_400_62400# 0.81fF
C2940 VN.n2593 a_400_62400# 0.16fF
C2941 VN.t2051 a_400_62400# 0.03fF
C2942 VN.n2594 a_400_62400# 0.19fF
C2943 VN.n2596 a_400_62400# 1.55fF
C2944 VN.n2597 a_400_62400# 0.29fF
C2945 VN.n2598 a_400_62400# 2.52fF
C2946 VN.t2355 a_400_62400# 0.03fF
C2947 VN.n2599 a_400_62400# 0.32fF
C2948 VN.n2600 a_400_62400# 1.22fF
C2949 VN.n2601 a_400_62400# 0.07fF
C2950 VN.t2248 a_400_62400# 0.03fF
C2951 VN.n2602 a_400_62400# 0.16fF
C2952 VN.n2603 a_400_62400# 0.19fF
C2953 VN.n2605 a_400_62400# 27.83fF
C2954 VN.n2606 a_400_62400# 3.93fF
C2955 VN.n2607 a_400_62400# 2.51fF
C2956 VN.n2608 a_400_62400# 0.16fF
C2957 VN.t1183 a_400_62400# 0.03fF
C2958 VN.n2609 a_400_62400# 0.19fF
C2959 VN.t2322 a_400_62400# 0.03fF
C2960 VN.n2611 a_400_62400# 0.32fF
C2961 VN.n2612 a_400_62400# 0.48fF
C2962 VN.n2613 a_400_62400# 0.81fF
C2963 VN.n2614 a_400_62400# 1.46fF
C2964 VN.n2615 a_400_62400# 0.21fF
C2965 VN.n2616 a_400_62400# 2.81fF
C2966 VN.t1387 a_400_62400# 0.03fF
C2967 VN.n2617 a_400_62400# 0.16fF
C2968 VN.n2618 a_400_62400# 0.19fF
C2969 VN.t1487 a_400_62400# 0.03fF
C2970 VN.n2620 a_400_62400# 0.32fF
C2971 VN.n2621 a_400_62400# 1.22fF
C2972 VN.n2622 a_400_62400# 0.07fF
C2973 VN.n2623 a_400_62400# 2.51fF
C2974 VN.n2624 a_400_62400# 3.57fF
C2975 VN.t1455 a_400_62400# 0.03fF
C2976 VN.n2625 a_400_62400# 0.32fF
C2977 VN.n2626 a_400_62400# 0.48fF
C2978 VN.n2627 a_400_62400# 0.81fF
C2979 VN.n2628 a_400_62400# 0.16fF
C2980 VN.t458 a_400_62400# 0.03fF
C2981 VN.n2629 a_400_62400# 0.19fF
C2982 VN.n2631 a_400_62400# 3.93fF
C2983 VN.n2632 a_400_62400# 3.08fF
C2984 VN.t521 a_400_62400# 0.03fF
C2985 VN.n2633 a_400_62400# 0.16fF
C2986 VN.n2634 a_400_62400# 0.19fF
C2987 VN.t620 a_400_62400# 0.03fF
C2988 VN.n2636 a_400_62400# 0.32fF
C2989 VN.n2637 a_400_62400# 1.22fF
C2990 VN.n2638 a_400_62400# 0.07fF
C2991 VN.n2639 a_400_62400# 2.51fF
C2992 VN.n2640 a_400_62400# 3.57fF
C2993 VN.t708 a_400_62400# 0.03fF
C2994 VN.n2641 a_400_62400# 0.32fF
C2995 VN.n2642 a_400_62400# 0.48fF
C2996 VN.n2643 a_400_62400# 0.81fF
C2997 VN.n2644 a_400_62400# 0.16fF
C2998 VN.t2104 a_400_62400# 0.03fF
C2999 VN.n2645 a_400_62400# 0.19fF
C3000 VN.n2647 a_400_62400# 3.75fF
C3001 VN.n2648 a_400_62400# 3.08fF
C3002 VN.t2172 a_400_62400# 0.03fF
C3003 VN.n2649 a_400_62400# 0.16fF
C3004 VN.n2650 a_400_62400# 0.19fF
C3005 VN.t2400 a_400_62400# 0.03fF
C3006 VN.n2652 a_400_62400# 0.32fF
C3007 VN.n2653 a_400_62400# 1.22fF
C3008 VN.n2654 a_400_62400# 0.07fF
C3009 VN.n2655 a_400_62400# 2.51fF
C3010 VN.n2656 a_400_62400# 3.57fF
C3011 VN.t2364 a_400_62400# 0.03fF
C3012 VN.n2657 a_400_62400# 0.32fF
C3013 VN.n2658 a_400_62400# 0.48fF
C3014 VN.n2659 a_400_62400# 0.81fF
C3015 VN.n2660 a_400_62400# 0.16fF
C3016 VN.t1227 a_400_62400# 0.03fF
C3017 VN.n2661 a_400_62400# 0.19fF
C3018 VN.n2663 a_400_62400# 3.75fF
C3019 VN.n2664 a_400_62400# 3.08fF
C3020 VN.t1305 a_400_62400# 0.03fF
C3021 VN.n2665 a_400_62400# 0.16fF
C3022 VN.n2666 a_400_62400# 0.19fF
C3023 VN.t1531 a_400_62400# 0.03fF
C3024 VN.n2668 a_400_62400# 0.32fF
C3025 VN.n2669 a_400_62400# 1.22fF
C3026 VN.n2670 a_400_62400# 0.07fF
C3027 VN.n2671 a_400_62400# 2.51fF
C3028 VN.n2672 a_400_62400# 3.57fF
C3029 VN.t1494 a_400_62400# 0.03fF
C3030 VN.n2673 a_400_62400# 0.32fF
C3031 VN.n2674 a_400_62400# 0.48fF
C3032 VN.n2675 a_400_62400# 0.81fF
C3033 VN.n2676 a_400_62400# 0.16fF
C3034 VN.t361 a_400_62400# 0.03fF
C3035 VN.n2677 a_400_62400# 0.19fF
C3036 VN.n2679 a_400_62400# 3.75fF
C3037 VN.n2680 a_400_62400# 3.08fF
C3038 VN.t441 a_400_62400# 0.03fF
C3039 VN.n2681 a_400_62400# 0.16fF
C3040 VN.n2682 a_400_62400# 0.19fF
C3041 VN.t660 a_400_62400# 0.03fF
C3042 VN.n2684 a_400_62400# 0.32fF
C3043 VN.n2685 a_400_62400# 1.22fF
C3044 VN.n2686 a_400_62400# 0.07fF
C3045 VN.n2687 a_400_62400# 2.51fF
C3046 VN.n2688 a_400_62400# 3.57fF
C3047 VN.t627 a_400_62400# 0.03fF
C3048 VN.n2689 a_400_62400# 0.32fF
C3049 VN.n2690 a_400_62400# 0.48fF
C3050 VN.n2691 a_400_62400# 0.81fF
C3051 VN.n2692 a_400_62400# 0.16fF
C3052 VN.t2011 a_400_62400# 0.03fF
C3053 VN.n2693 a_400_62400# 0.19fF
C3054 VN.n2695 a_400_62400# 3.75fF
C3055 VN.n2696 a_400_62400# 3.08fF
C3056 VN.t2086 a_400_62400# 0.03fF
C3057 VN.n2697 a_400_62400# 0.16fF
C3058 VN.n2698 a_400_62400# 0.19fF
C3059 VN.t2320 a_400_62400# 0.03fF
C3060 VN.n2700 a_400_62400# 0.32fF
C3061 VN.n2701 a_400_62400# 1.22fF
C3062 VN.n2702 a_400_62400# 0.07fF
C3063 VN.n2703 a_400_62400# 2.51fF
C3064 VN.n2704 a_400_62400# 3.57fF
C3065 VN.t2281 a_400_62400# 0.03fF
C3066 VN.n2705 a_400_62400# 0.32fF
C3067 VN.n2706 a_400_62400# 0.48fF
C3068 VN.n2707 a_400_62400# 0.81fF
C3069 VN.n2708 a_400_62400# 0.16fF
C3070 VN.t1138 a_400_62400# 0.03fF
C3071 VN.n2709 a_400_62400# 0.19fF
C3072 VN.n2711 a_400_62400# 3.75fF
C3073 VN.n2712 a_400_62400# 3.08fF
C3074 VN.t1347 a_400_62400# 0.03fF
C3075 VN.n2713 a_400_62400# 0.16fF
C3076 VN.n2714 a_400_62400# 0.19fF
C3077 VN.t1452 a_400_62400# 0.03fF
C3078 VN.n2716 a_400_62400# 0.32fF
C3079 VN.n2717 a_400_62400# 1.22fF
C3080 VN.n2718 a_400_62400# 0.07fF
C3081 VN.n2719 a_400_62400# 2.51fF
C3082 VN.n2720 a_400_62400# 3.57fF
C3083 VN.t1412 a_400_62400# 0.03fF
C3084 VN.n2721 a_400_62400# 0.32fF
C3085 VN.n2722 a_400_62400# 0.48fF
C3086 VN.n2723 a_400_62400# 0.81fF
C3087 VN.n2724 a_400_62400# 0.16fF
C3088 VN.t275 a_400_62400# 0.03fF
C3089 VN.n2725 a_400_62400# 0.19fF
C3090 VN.n2727 a_400_62400# 3.75fF
C3091 VN.n2728 a_400_62400# 3.08fF
C3092 VN.t481 a_400_62400# 0.03fF
C3093 VN.n2729 a_400_62400# 0.16fF
C3094 VN.n2730 a_400_62400# 0.19fF
C3095 VN.t583 a_400_62400# 0.03fF
C3096 VN.n2732 a_400_62400# 0.32fF
C3097 VN.n2733 a_400_62400# 1.22fF
C3098 VN.n2734 a_400_62400# 0.07fF
C3099 VN.n2735 a_400_62400# 2.51fF
C3100 VN.n2736 a_400_62400# 3.57fF
C3101 VN.t98 a_400_62400# 0.03fF
C3102 VN.n2737 a_400_62400# 0.32fF
C3103 VN.n2738 a_400_62400# 0.48fF
C3104 VN.n2739 a_400_62400# 0.81fF
C3105 VN.n2740 a_400_62400# 0.16fF
C3106 VN.t1505 a_400_62400# 0.03fF
C3107 VN.n2741 a_400_62400# 0.19fF
C3108 VN.n2743 a_400_62400# 3.75fF
C3109 VN.n2744 a_400_62400# 3.08fF
C3110 VN.t1686 a_400_62400# 0.03fF
C3111 VN.n2745 a_400_62400# 0.16fF
C3112 VN.n2746 a_400_62400# 0.19fF
C3113 VN.t1915 a_400_62400# 0.03fF
C3114 VN.n2748 a_400_62400# 0.32fF
C3115 VN.n2749 a_400_62400# 1.22fF
C3116 VN.n2750 a_400_62400# 0.07fF
C3117 VN.n2751 a_400_62400# 2.51fF
C3118 VN.n2752 a_400_62400# 3.57fF
C3119 VN.t1769 a_400_62400# 0.03fF
C3120 VN.n2753 a_400_62400# 0.32fF
C3121 VN.n2754 a_400_62400# 0.48fF
C3122 VN.n2755 a_400_62400# 0.81fF
C3123 VN.n2756 a_400_62400# 0.16fF
C3124 VN.t637 a_400_62400# 0.03fF
C3125 VN.n2757 a_400_62400# 0.19fF
C3126 VN.n2759 a_400_62400# 3.75fF
C3127 VN.n2760 a_400_62400# 3.08fF
C3128 VN.t820 a_400_62400# 0.03fF
C3129 VN.n2761 a_400_62400# 0.16fF
C3130 VN.n2762 a_400_62400# 0.19fF
C3131 VN.t1040 a_400_62400# 0.03fF
C3132 VN.n2764 a_400_62400# 0.32fF
C3133 VN.n2765 a_400_62400# 1.22fF
C3134 VN.n2766 a_400_62400# 0.07fF
C3135 VN.n2767 a_400_62400# 3.65fF
C3136 VN.n2768 a_400_62400# 2.14fF
C3137 VN.n2769 a_400_62400# 0.16fF
C3138 VN.t1547 a_400_62400# 0.03fF
C3139 VN.n2770 a_400_62400# 0.19fF
C3140 VN.t2559 a_400_62400# 0.03fF
C3141 VN.n2772 a_400_62400# 0.32fF
C3142 VN.n2773 a_400_62400# 0.48fF
C3143 VN.n2774 a_400_62400# 0.81fF
C3144 VN.n2775 a_400_62400# 0.09fF
C3145 VN.n2776 a_400_62400# 0.01fF
C3146 VN.n2777 a_400_62400# 0.02fF
C3147 VN.n2778 a_400_62400# 0.02fF
C3148 VN.n2779 a_400_62400# 0.32fF
C3149 VN.n2780 a_400_62400# 1.56fF
C3150 VN.n2781 a_400_62400# 1.81fF
C3151 VN.n2782 a_400_62400# 3.08fF
C3152 VN.t1616 a_400_62400# 0.03fF
C3153 VN.n2783 a_400_62400# 0.16fF
C3154 VN.n2784 a_400_62400# 0.19fF
C3155 VN.t1829 a_400_62400# 0.03fF
C3156 VN.n2786 a_400_62400# 0.32fF
C3157 VN.n2787 a_400_62400# 1.22fF
C3158 VN.n2788 a_400_62400# 0.07fF
C3159 VN.t57 a_400_62400# 64.69fF
C3160 VN.t168 a_400_62400# 0.03fF
C3161 VN.n2789 a_400_62400# 0.32fF
C3162 VN.n2790 a_400_62400# 1.22fF
C3163 VN.n2791 a_400_62400# 0.07fF
C3164 VN.t2477 a_400_62400# 0.03fF
C3165 VN.n2792 a_400_62400# 0.16fF
C3166 VN.n2793 a_400_62400# 0.19fF
C3167 VN.n2795 a_400_62400# 0.16fF
C3168 VN.t2294 a_400_62400# 0.03fF
C3169 VN.n2796 a_400_62400# 0.19fF
C3170 VN.n2798 a_400_62400# 6.92fF
C3171 VN.n2799 a_400_62400# 6.56fF
C3172 VN.t1584 a_400_62400# 0.03fF
C3173 VN.n2800 a_400_62400# 0.16fF
C3174 VN.n2801 a_400_62400# 0.19fF
C3175 VN.t1102 a_400_62400# 0.03fF
C3176 VN.n2803 a_400_62400# 0.32fF
C3177 VN.n2804 a_400_62400# 1.22fF
C3178 VN.n2805 a_400_62400# 0.07fF
C3179 VN.n2806 a_400_62400# 2.51fF
C3180 VN.n2807 a_400_62400# 3.58fF
C3181 VN.t1193 a_400_62400# 0.03fF
C3182 VN.n2808 a_400_62400# 0.32fF
C3183 VN.n2809 a_400_62400# 0.48fF
C3184 VN.n2810 a_400_62400# 0.81fF
C3185 VN.n2811 a_400_62400# 0.16fF
C3186 VN.t2556 a_400_62400# 0.03fF
C3187 VN.n2812 a_400_62400# 0.19fF
C3188 VN.n2814 a_400_62400# 7.29fF
C3189 VN.t720 a_400_62400# 0.03fF
C3190 VN.n2815 a_400_62400# 0.16fF
C3191 VN.n2816 a_400_62400# 0.19fF
C3192 VN.t235 a_400_62400# 0.03fF
C3193 VN.n2818 a_400_62400# 0.32fF
C3194 VN.n2819 a_400_62400# 1.22fF
C3195 VN.n2820 a_400_62400# 0.07fF
C3196 VN.t49 a_400_62400# 64.17fF
C3197 VN.t1883 a_400_62400# 0.03fF
C3198 VN.n2821 a_400_62400# 1.60fF
C3199 VN.n2822 a_400_62400# 0.07fF
C3200 VN.t2491 a_400_62400# 0.03fF
C3201 VN.n2823 a_400_62400# 0.02fF
C3202 VN.n2824 a_400_62400# 0.34fF
C3203 VN.n2826 a_400_62400# 2.01fF
C3204 VN.n2827 a_400_62400# 1.75fF
C3205 VN.n2828 a_400_62400# 0.37fF
C3206 VN.n2829 a_400_62400# 0.33fF
C3207 VN.n2830 a_400_62400# 5.88fF
C3208 VN.n2831 a_400_62400# 0.02fF
C3209 VN.n2832 a_400_62400# 0.02fF
C3210 VN.n2833 a_400_62400# 0.03fF
C3211 VN.n2834 a_400_62400# 0.05fF
C3212 VN.n2835 a_400_62400# 0.23fF
C3213 VN.n2836 a_400_62400# 0.02fF
C3214 VN.n2837 a_400_62400# 0.03fF
C3215 VN.n2838 a_400_62400# 0.01fF
C3216 VN.n2839 a_400_62400# 0.01fF
C3217 VN.n2840 a_400_62400# 0.01fF
C3218 VN.n2841 a_400_62400# 0.02fF
C3219 VN.n2842 a_400_62400# 0.03fF
C3220 VN.n2843 a_400_62400# 0.06fF
C3221 VN.n2844 a_400_62400# 0.05fF
C3222 VN.n2845 a_400_62400# 0.15fF
C3223 VN.n2846 a_400_62400# 0.51fF
C3224 VN.n2847 a_400_62400# 0.27fF
C3225 VN.n2848 a_400_62400# 37.46fF
C3226 VN.n2849 a_400_62400# 37.46fF
C3227 VN.n2850 a_400_62400# 0.79fF
C3228 VN.n2851 a_400_62400# 0.23fF
C3229 VN.n2852 a_400_62400# 1.18fF
C3230 VN.t167 a_400_62400# 28.64fF
C3231 VN.n2853 a_400_62400# 0.79fF
C3232 VN.n2854 a_400_62400# 0.11fF
C3233 VN.n2855 a_400_62400# 4.98fF
C3234 VN.n2856 a_400_62400# 0.80fF
C3235 VN.n2857 a_400_62400# 0.29fF
C3236 VN.n2858 a_400_62400# 1.96fF
C3237 VN.n2860 a_400_62400# 25.18fF
C3238 VN.n2862 a_400_62400# 1.87fF
C3239 VN.n2863 a_400_62400# 5.36fF
C3240 VN.n2864 a_400_62400# 1.81fF
C3241 VN.t1165 a_400_62400# 0.03fF
C3242 VN.n2865 a_400_62400# 0.85fF
C3243 VN.n2866 a_400_62400# 0.81fF
C3244 VN.n2867 a_400_62400# 0.33fF
C3245 VN.n2868 a_400_62400# 0.12fF
C3246 VN.n2869 a_400_62400# 0.28fF
C3247 VN.n2870 a_400_62400# 1.23fF
C3248 VN.n2871 a_400_62400# 0.59fF
C3249 VN.n2872 a_400_62400# 2.51fF
C3250 VN.n2873 a_400_62400# 0.16fF
C3251 VN.t446 a_400_62400# 0.03fF
C3252 VN.n2874 a_400_62400# 0.19fF
C3253 VN.t1150 a_400_62400# 0.03fF
C3254 VN.n2876 a_400_62400# 0.32fF
C3255 VN.n2877 a_400_62400# 0.48fF
C3256 VN.n2878 a_400_62400# 0.81fF
C3257 VN.n2879 a_400_62400# 0.03fF
C3258 VN.n2880 a_400_62400# 0.01fF
C3259 VN.n2881 a_400_62400# 0.02fF
C3260 VN.n2882 a_400_62400# 0.11fF
C3261 VN.n2883 a_400_62400# 0.08fF
C3262 VN.n2884 a_400_62400# 0.04fF
C3263 VN.n2885 a_400_62400# 0.05fF
C3264 VN.n2886 a_400_62400# 1.34fF
C3265 VN.n2887 a_400_62400# 0.48fF
C3266 VN.n2888 a_400_62400# 2.51fF
C3267 VN.n2889 a_400_62400# 2.67fF
C3268 VN.t2273 a_400_62400# 0.03fF
C3269 VN.n2890 a_400_62400# 0.32fF
C3270 VN.n2891 a_400_62400# 1.22fF
C3271 VN.n2892 a_400_62400# 0.07fF
C3272 VN.t1096 a_400_62400# 0.03fF
C3273 VN.n2893 a_400_62400# 0.16fF
C3274 VN.n2894 a_400_62400# 0.19fF
C3275 VN.n2896 a_400_62400# 2.53fF
C3276 VN.n2897 a_400_62400# 0.09fF
C3277 VN.n2898 a_400_62400# 0.05fF
C3278 VN.n2899 a_400_62400# 0.07fF
C3279 VN.n2900 a_400_62400# 1.16fF
C3280 VN.n2901 a_400_62400# 0.01fF
C3281 VN.n2902 a_400_62400# 0.01fF
C3282 VN.n2903 a_400_62400# 0.01fF
C3283 VN.n2904 a_400_62400# 0.09fF
C3284 VN.n2905 a_400_62400# 0.91fF
C3285 VN.n2906 a_400_62400# 0.96fF
C3286 VN.t427 a_400_62400# 0.03fF
C3287 VN.n2907 a_400_62400# 0.32fF
C3288 VN.n2908 a_400_62400# 0.48fF
C3289 VN.n2909 a_400_62400# 0.81fF
C3290 VN.n2910 a_400_62400# 0.16fF
C3291 VN.t2090 a_400_62400# 0.03fF
C3292 VN.n2911 a_400_62400# 0.19fF
C3293 VN.n2913 a_400_62400# 0.93fF
C3294 VN.n2914 a_400_62400# 0.30fF
C3295 VN.n2915 a_400_62400# 0.34fF
C3296 VN.n2916 a_400_62400# 0.12fF
C3297 VN.n2917 a_400_62400# 0.30fF
C3298 VN.n2918 a_400_62400# 0.93fF
C3299 VN.n2919 a_400_62400# 1.55fF
C3300 VN.n2920 a_400_62400# 0.29fF
C3301 VN.n2921 a_400_62400# 0.34fF
C3302 VN.n2922 a_400_62400# 0.12fF
C3303 VN.n2923 a_400_62400# 3.10fF
C3304 VN.t1535 a_400_62400# 0.03fF
C3305 VN.n2924 a_400_62400# 0.32fF
C3306 VN.n2925 a_400_62400# 1.22fF
C3307 VN.n2926 a_400_62400# 0.07fF
C3308 VN.t228 a_400_62400# 0.03fF
C3309 VN.n2927 a_400_62400# 0.16fF
C3310 VN.n2928 a_400_62400# 0.19fF
C3311 VN.n2930 a_400_62400# 2.51fF
C3312 VN.n2931 a_400_62400# 0.61fF
C3313 VN.n2932 a_400_62400# 0.30fF
C3314 VN.n2933 a_400_62400# 0.51fF
C3315 VN.n2934 a_400_62400# 0.21fF
C3316 VN.n2935 a_400_62400# 0.38fF
C3317 VN.n2936 a_400_62400# 0.29fF
C3318 VN.n2937 a_400_62400# 0.40fF
C3319 VN.n2938 a_400_62400# 0.28fF
C3320 VN.t2073 a_400_62400# 0.03fF
C3321 VN.n2939 a_400_62400# 0.32fF
C3322 VN.n2940 a_400_62400# 0.48fF
C3323 VN.n2941 a_400_62400# 0.81fF
C3324 VN.n2942 a_400_62400# 0.16fF
C3325 VN.t1214 a_400_62400# 0.03fF
C3326 VN.n2943 a_400_62400# 0.19fF
C3327 VN.n2945 a_400_62400# 0.06fF
C3328 VN.n2946 a_400_62400# 0.04fF
C3329 VN.n2947 a_400_62400# 0.04fF
C3330 VN.n2948 a_400_62400# 0.14fF
C3331 VN.n2949 a_400_62400# 0.48fF
C3332 VN.n2950 a_400_62400# 0.50fF
C3333 VN.n2951 a_400_62400# 0.14fF
C3334 VN.n2952 a_400_62400# 0.16fF
C3335 VN.n2953 a_400_62400# 0.09fF
C3336 VN.n2954 a_400_62400# 0.16fF
C3337 VN.n2955 a_400_62400# 0.24fF
C3338 VN.n2956 a_400_62400# 5.35fF
C3339 VN.t663 a_400_62400# 0.03fF
C3340 VN.n2957 a_400_62400# 0.32fF
C3341 VN.n2958 a_400_62400# 1.22fF
C3342 VN.n2959 a_400_62400# 0.07fF
C3343 VN.t1878 a_400_62400# 0.03fF
C3344 VN.n2960 a_400_62400# 0.16fF
C3345 VN.n2961 a_400_62400# 0.19fF
C3346 VN.n2963 a_400_62400# 0.33fF
C3347 VN.n2964 a_400_62400# 0.12fF
C3348 VN.n2965 a_400_62400# 0.28fF
C3349 VN.n2966 a_400_62400# 1.72fF
C3350 VN.n2967 a_400_62400# 0.71fF
C3351 VN.n2968 a_400_62400# 2.51fF
C3352 VN.n2969 a_400_62400# 0.16fF
C3353 VN.t1682 a_400_62400# 0.03fF
C3354 VN.n2970 a_400_62400# 0.19fF
C3355 VN.t2536 a_400_62400# 0.03fF
C3356 VN.n2972 a_400_62400# 0.32fF
C3357 VN.n2973 a_400_62400# 0.48fF
C3358 VN.n2974 a_400_62400# 0.81fF
C3359 VN.n2975 a_400_62400# 0.95fF
C3360 VN.n2976 a_400_62400# 2.11fF
C3361 VN.n2977 a_400_62400# 3.28fF
C3362 VN.t1140 a_400_62400# 0.03fF
C3363 VN.n2978 a_400_62400# 0.32fF
C3364 VN.n2979 a_400_62400# 1.22fF
C3365 VN.n2980 a_400_62400# 0.07fF
C3366 VN.t1009 a_400_62400# 0.03fF
C3367 VN.n2981 a_400_62400# 0.16fF
C3368 VN.n2982 a_400_62400# 0.19fF
C3369 VN.n2984 a_400_62400# 2.53fF
C3370 VN.n2985 a_400_62400# 0.08fF
C3371 VN.n2986 a_400_62400# 0.04fF
C3372 VN.n2987 a_400_62400# 0.05fF
C3373 VN.n2988 a_400_62400# 1.33fF
C3374 VN.n2989 a_400_62400# 0.03fF
C3375 VN.n2990 a_400_62400# 0.01fF
C3376 VN.n2991 a_400_62400# 0.02fF
C3377 VN.n2992 a_400_62400# 0.11fF
C3378 VN.n2993 a_400_62400# 0.48fF
C3379 VN.n2994 a_400_62400# 2.48fF
C3380 VN.t1671 a_400_62400# 0.03fF
C3381 VN.n2995 a_400_62400# 0.32fF
C3382 VN.n2996 a_400_62400# 0.48fF
C3383 VN.n2997 a_400_62400# 0.81fF
C3384 VN.n2998 a_400_62400# 0.16fF
C3385 VN.t816 a_400_62400# 0.03fF
C3386 VN.n2999 a_400_62400# 0.19fF
C3387 VN.n3001 a_400_62400# 0.93fF
C3388 VN.n3002 a_400_62400# 0.30fF
C3389 VN.n3003 a_400_62400# 0.34fF
C3390 VN.n3004 a_400_62400# 0.12fF
C3391 VN.n3005 a_400_62400# 0.30fF
C3392 VN.n3006 a_400_62400# 0.93fF
C3393 VN.n3007 a_400_62400# 1.55fF
C3394 VN.n3008 a_400_62400# 0.29fF
C3395 VN.n3009 a_400_62400# 0.34fF
C3396 VN.n3010 a_400_62400# 0.12fF
C3397 VN.n3011 a_400_62400# 2.52fF
C3398 VN.t277 a_400_62400# 0.03fF
C3399 VN.n3012 a_400_62400# 0.32fF
C3400 VN.n3013 a_400_62400# 1.22fF
C3401 VN.n3014 a_400_62400# 0.07fF
C3402 VN.t1498 a_400_62400# 0.03fF
C3403 VN.n3015 a_400_62400# 0.16fF
C3404 VN.n3016 a_400_62400# 0.19fF
C3405 VN.n3018 a_400_62400# 27.83fF
C3406 VN.n3019 a_400_62400# 2.30fF
C3407 VN.n3020 a_400_62400# 4.08fF
C3408 VN.t2025 a_400_62400# 0.03fF
C3409 VN.n3021 a_400_62400# 0.32fF
C3410 VN.n3022 a_400_62400# 0.48fF
C3411 VN.n3023 a_400_62400# 0.81fF
C3412 VN.n3024 a_400_62400# 0.16fF
C3413 VN.t1174 a_400_62400# 0.03fF
C3414 VN.n3025 a_400_62400# 0.19fF
C3415 VN.n3027 a_400_62400# 0.42fF
C3416 VN.n3028 a_400_62400# 0.34fF
C3417 VN.n3029 a_400_62400# 0.12fF
C3418 VN.n3030 a_400_62400# 0.30fF
C3419 VN.n3031 a_400_62400# 0.88fF
C3420 VN.n3032 a_400_62400# 1.28fF
C3421 VN.n3033 a_400_62400# 0.30fF
C3422 VN.n3034 a_400_62400# 0.28fF
C3423 VN.n3035 a_400_62400# 0.27fF
C3424 VN.n3036 a_400_62400# 0.09fF
C3425 VN.n3037 a_400_62400# 0.12fF
C3426 VN.n3038 a_400_62400# 0.13fF
C3427 VN.n3039 a_400_62400# 2.66fF
C3428 VN.t1963 a_400_62400# 0.03fF
C3429 VN.n3040 a_400_62400# 0.16fF
C3430 VN.n3041 a_400_62400# 0.19fF
C3431 VN.t622 a_400_62400# 0.03fF
C3432 VN.n3043 a_400_62400# 0.32fF
C3433 VN.n3044 a_400_62400# 1.22fF
C3434 VN.n3045 a_400_62400# 0.07fF
C3435 VN.n3046 a_400_62400# 2.51fF
C3436 VN.n3047 a_400_62400# 0.16fF
C3437 VN.t2473 a_400_62400# 0.03fF
C3438 VN.n3048 a_400_62400# 0.19fF
C3439 VN.t805 a_400_62400# 0.03fF
C3440 VN.n3050 a_400_62400# 0.32fF
C3441 VN.n3051 a_400_62400# 0.48fF
C3442 VN.n3052 a_400_62400# 0.81fF
C3443 VN.n3053 a_400_62400# 1.24fF
C3444 VN.n3054 a_400_62400# 0.43fF
C3445 VN.n3055 a_400_62400# 0.43fF
C3446 VN.n3056 a_400_62400# 1.24fF
C3447 VN.n3057 a_400_62400# 1.46fF
C3448 VN.n3058 a_400_62400# 0.21fF
C3449 VN.n3059 a_400_62400# 6.64fF
C3450 VN.t632 a_400_62400# 0.03fF
C3451 VN.n3060 a_400_62400# 0.16fF
C3452 VN.n3061 a_400_62400# 0.19fF
C3453 VN.t1925 a_400_62400# 0.03fF
C3454 VN.n3063 a_400_62400# 0.32fF
C3455 VN.n3064 a_400_62400# 1.22fF
C3456 VN.n3065 a_400_62400# 0.07fF
C3457 VN.n3066 a_400_62400# 2.51fF
C3458 VN.n3067 a_400_62400# 3.57fF
C3459 VN.t2458 a_400_62400# 0.03fF
C3460 VN.n3068 a_400_62400# 0.32fF
C3461 VN.n3069 a_400_62400# 0.48fF
C3462 VN.n3070 a_400_62400# 0.81fF
C3463 VN.n3071 a_400_62400# 0.16fF
C3464 VN.t1612 a_400_62400# 0.03fF
C3465 VN.n3072 a_400_62400# 0.19fF
C3466 VN.n3074 a_400_62400# 6.91fF
C3467 VN.t2408 a_400_62400# 0.03fF
C3468 VN.n3075 a_400_62400# 0.16fF
C3469 VN.n3076 a_400_62400# 0.19fF
C3470 VN.t1051 a_400_62400# 0.03fF
C3471 VN.n3078 a_400_62400# 0.32fF
C3472 VN.n3079 a_400_62400# 1.22fF
C3473 VN.n3080 a_400_62400# 0.07fF
C3474 VN.n3081 a_400_62400# 2.51fF
C3475 VN.n3082 a_400_62400# 3.57fF
C3476 VN.t1593 a_400_62400# 0.03fF
C3477 VN.n3083 a_400_62400# 0.32fF
C3478 VN.n3084 a_400_62400# 0.48fF
C3479 VN.n3085 a_400_62400# 0.81fF
C3480 VN.n3086 a_400_62400# 0.16fF
C3481 VN.t745 a_400_62400# 0.03fF
C3482 VN.n3087 a_400_62400# 0.19fF
C3483 VN.n3089 a_400_62400# 6.92fF
C3484 VN.t1541 a_400_62400# 0.03fF
C3485 VN.n3090 a_400_62400# 0.16fF
C3486 VN.n3091 a_400_62400# 0.19fF
C3487 VN.t180 a_400_62400# 0.03fF
C3488 VN.n3093 a_400_62400# 0.32fF
C3489 VN.n3094 a_400_62400# 1.22fF
C3490 VN.n3095 a_400_62400# 0.07fF
C3491 VN.n3096 a_400_62400# 2.51fF
C3492 VN.n3097 a_400_62400# 3.57fF
C3493 VN.t728 a_400_62400# 0.03fF
C3494 VN.n3098 a_400_62400# 0.32fF
C3495 VN.n3099 a_400_62400# 0.48fF
C3496 VN.n3100 a_400_62400# 0.81fF
C3497 VN.n3101 a_400_62400# 0.16fF
C3498 VN.t2402 a_400_62400# 0.03fF
C3499 VN.n3102 a_400_62400# 0.19fF
C3500 VN.n3104 a_400_62400# 6.92fF
C3501 VN.t672 a_400_62400# 0.03fF
C3502 VN.n3105 a_400_62400# 0.16fF
C3503 VN.n3106 a_400_62400# 0.19fF
C3504 VN.t1838 a_400_62400# 0.03fF
C3505 VN.n3108 a_400_62400# 0.32fF
C3506 VN.n3109 a_400_62400# 1.22fF
C3507 VN.n3110 a_400_62400# 0.07fF
C3508 VN.n3111 a_400_62400# 2.51fF
C3509 VN.n3112 a_400_62400# 3.57fF
C3510 VN.t2383 a_400_62400# 0.03fF
C3511 VN.n3113 a_400_62400# 0.32fF
C3512 VN.n3114 a_400_62400# 0.48fF
C3513 VN.n3115 a_400_62400# 0.81fF
C3514 VN.n3116 a_400_62400# 0.16fF
C3515 VN.t1533 a_400_62400# 0.03fF
C3516 VN.n3117 a_400_62400# 0.19fF
C3517 VN.n3119 a_400_62400# 6.92fF
C3518 VN.t2331 a_400_62400# 0.03fF
C3519 VN.n3120 a_400_62400# 0.16fF
C3520 VN.n3121 a_400_62400# 0.19fF
C3521 VN.t966 a_400_62400# 0.03fF
C3522 VN.n3123 a_400_62400# 0.32fF
C3523 VN.n3124 a_400_62400# 1.22fF
C3524 VN.n3125 a_400_62400# 0.07fF
C3525 VN.n3126 a_400_62400# 2.51fF
C3526 VN.n3127 a_400_62400# 3.57fF
C3527 VN.t1514 a_400_62400# 0.03fF
C3528 VN.n3128 a_400_62400# 0.32fF
C3529 VN.n3129 a_400_62400# 0.48fF
C3530 VN.n3130 a_400_62400# 0.81fF
C3531 VN.n3131 a_400_62400# 0.16fF
C3532 VN.t783 a_400_62400# 0.03fF
C3533 VN.n3132 a_400_62400# 0.19fF
C3534 VN.n3134 a_400_62400# 6.92fF
C3535 VN.t1467 a_400_62400# 0.03fF
C3536 VN.n3135 a_400_62400# 0.16fF
C3537 VN.n3136 a_400_62400# 0.19fF
C3538 VN.t62 a_400_62400# 0.03fF
C3539 VN.n3138 a_400_62400# 0.32fF
C3540 VN.n3139 a_400_62400# 1.22fF
C3541 VN.n3140 a_400_62400# 0.07fF
C3542 VN.n3141 a_400_62400# 2.51fF
C3543 VN.n3142 a_400_62400# 3.57fF
C3544 VN.t770 a_400_62400# 0.03fF
C3545 VN.n3143 a_400_62400# 0.32fF
C3546 VN.n3144 a_400_62400# 0.48fF
C3547 VN.n3145 a_400_62400# 0.81fF
C3548 VN.n3146 a_400_62400# 0.16fF
C3549 VN.t2435 a_400_62400# 0.03fF
C3550 VN.n3147 a_400_62400# 0.19fF
C3551 VN.n3149 a_400_62400# 6.92fF
C3552 VN.t597 a_400_62400# 0.03fF
C3553 VN.n3150 a_400_62400# 0.16fF
C3554 VN.n3151 a_400_62400# 0.19fF
C3555 VN.t1882 a_400_62400# 0.03fF
C3556 VN.n3153 a_400_62400# 0.32fF
C3557 VN.n3154 a_400_62400# 1.22fF
C3558 VN.n3155 a_400_62400# 0.07fF
C3559 VN.n3156 a_400_62400# 2.51fF
C3560 VN.n3157 a_400_62400# 3.57fF
C3561 VN.t2130 a_400_62400# 0.03fF
C3562 VN.n3158 a_400_62400# 0.32fF
C3563 VN.n3159 a_400_62400# 0.48fF
C3564 VN.n3160 a_400_62400# 0.81fF
C3565 VN.n3161 a_400_62400# 0.16fF
C3566 VN.t64 a_400_62400# 0.03fF
C3567 VN.n3162 a_400_62400# 0.19fF
C3568 VN.n3164 a_400_62400# 6.92fF
C3569 VN.t2252 a_400_62400# 0.03fF
C3570 VN.n3165 a_400_62400# 0.16fF
C3571 VN.n3166 a_400_62400# 0.19fF
C3572 VN.t1163 a_400_62400# 0.03fF
C3573 VN.n3168 a_400_62400# 0.32fF
C3574 VN.n3169 a_400_62400# 1.22fF
C3575 VN.n3170 a_400_62400# 0.07fF
C3576 VN.n3171 a_400_62400# 2.51fF
C3577 VN.n3172 a_400_62400# 3.57fF
C3578 VN.t1254 a_400_62400# 0.03fF
C3579 VN.n3173 a_400_62400# 0.32fF
C3580 VN.n3174 a_400_62400# 0.48fF
C3581 VN.n3175 a_400_62400# 0.81fF
C3582 VN.n3176 a_400_62400# 0.16fF
C3583 VN.t1755 a_400_62400# 0.03fF
C3584 VN.n3177 a_400_62400# 0.19fF
C3585 VN.n3179 a_400_62400# 6.92fF
C3586 VN.t2434 a_400_62400# 0.03fF
C3587 VN.n3180 a_400_62400# 0.16fF
C3588 VN.n3181 a_400_62400# 0.19fF
C3589 VN.t294 a_400_62400# 0.03fF
C3590 VN.n3183 a_400_62400# 0.32fF
C3591 VN.n3184 a_400_62400# 1.22fF
C3592 VN.n3185 a_400_62400# 0.07fF
C3593 VN.n3186 a_400_62400# 2.51fF
C3594 VN.n3187 a_400_62400# 3.57fF
C3595 VN.t384 a_400_62400# 0.03fF
C3596 VN.n3188 a_400_62400# 0.32fF
C3597 VN.n3189 a_400_62400# 0.48fF
C3598 VN.n3190 a_400_62400# 0.81fF
C3599 VN.n3191 a_400_62400# 0.16fF
C3600 VN.t883 a_400_62400# 0.03fF
C3601 VN.n3192 a_400_62400# 0.19fF
C3602 VN.n3194 a_400_62400# 2.51fF
C3603 VN.n3195 a_400_62400# 3.59fF
C3604 VN.t1740 a_400_62400# 0.03fF
C3605 VN.n3196 a_400_62400# 0.32fF
C3606 VN.n3197 a_400_62400# 0.48fF
C3607 VN.n3198 a_400_62400# 0.81fF
C3608 VN.t1424 a_400_62400# 0.03fF
C3609 VN.n3199 a_400_62400# 1.63fF
C3610 VN.n3200 a_400_62400# 0.49fF
C3611 VN.n3201 a_400_62400# 1.64fF
C3612 VN.n3202 a_400_62400# 0.81fF
C3613 VN.n3203 a_400_62400# 1.21fF
C3614 VN.n3204 a_400_62400# 1.54fF
C3615 VN.n3205 a_400_62400# 4.06fF
C3616 VN.t4 a_400_62400# 28.64fF
C3617 VN.n3206 a_400_62400# 28.43fF
C3618 VN.n3208 a_400_62400# 0.50fF
C3619 VN.n3209 a_400_62400# 0.31fF
C3620 VN.n3210 a_400_62400# 3.74fF
C3621 VN.n3211 a_400_62400# 3.29fF
C3622 VN.n3212 a_400_62400# 5.35fF
C3623 VN.n3213 a_400_62400# 0.34fF
C3624 VN.n3214 a_400_62400# 0.02fF
C3625 VN.t283 a_400_62400# 0.03fF
C3626 VN.n3215 a_400_62400# 0.34fF
C3627 VN.t853 a_400_62400# 0.03fF
C3628 VN.n3216 a_400_62400# 1.28fF
C3629 VN.n3217 a_400_62400# 0.94fF
C3630 VN.n3218 a_400_62400# 2.53fF
C3631 VN.n3219 a_400_62400# 2.51fF
C3632 VN.t557 a_400_62400# 0.03fF
C3633 VN.n3220 a_400_62400# 0.32fF
C3634 VN.n3221 a_400_62400# 0.48fF
C3635 VN.n3222 a_400_62400# 0.81fF
C3636 VN.n3223 a_400_62400# 0.16fF
C3637 VN.t1933 a_400_62400# 0.03fF
C3638 VN.n3224 a_400_62400# 0.19fF
C3639 VN.n3226 a_400_62400# 1.55fF
C3640 VN.n3227 a_400_62400# 0.29fF
C3641 VN.n3228 a_400_62400# 2.52fF
C3642 VN.t2515 a_400_62400# 0.03fF
C3643 VN.n3229 a_400_62400# 0.32fF
C3644 VN.n3230 a_400_62400# 1.22fF
C3645 VN.n3231 a_400_62400# 0.07fF
C3646 VN.t2004 a_400_62400# 0.03fF
C3647 VN.n3232 a_400_62400# 0.16fF
C3648 VN.n3233 a_400_62400# 0.19fF
C3649 VN.n3235 a_400_62400# 1.04fF
C3650 VN.n3236 a_400_62400# 2.60fF
C3651 VN.n3237 a_400_62400# 2.51fF
C3652 VN.n3238 a_400_62400# 0.16fF
C3653 VN.t1058 a_400_62400# 0.03fF
C3654 VN.n3239 a_400_62400# 0.19fF
C3655 VN.t2216 a_400_62400# 0.03fF
C3656 VN.n3241 a_400_62400# 0.32fF
C3657 VN.n3242 a_400_62400# 0.48fF
C3658 VN.n3243 a_400_62400# 0.81fF
C3659 VN.n3244 a_400_62400# 2.46fF
C3660 VN.n3245 a_400_62400# 4.01fF
C3661 VN.t1655 a_400_62400# 0.03fF
C3662 VN.n3246 a_400_62400# 0.32fF
C3663 VN.n3247 a_400_62400# 1.22fF
C3664 VN.n3248 a_400_62400# 0.07fF
C3665 VN.t1273 a_400_62400# 0.03fF
C3666 VN.n3249 a_400_62400# 0.16fF
C3667 VN.n3250 a_400_62400# 0.19fF
C3668 VN.n3252 a_400_62400# 2.53fF
C3669 VN.n3253 a_400_62400# 2.34fF
C3670 VN.t1349 a_400_62400# 0.03fF
C3671 VN.n3254 a_400_62400# 0.32fF
C3672 VN.n3255 a_400_62400# 0.48fF
C3673 VN.n3256 a_400_62400# 0.81fF
C3674 VN.n3257 a_400_62400# 0.16fF
C3675 VN.t184 a_400_62400# 0.03fF
C3676 VN.n3258 a_400_62400# 0.19fF
C3677 VN.n3260 a_400_62400# 1.55fF
C3678 VN.n3261 a_400_62400# 0.29fF
C3679 VN.n3262 a_400_62400# 3.27fF
C3680 VN.t786 a_400_62400# 0.03fF
C3681 VN.n3263 a_400_62400# 0.32fF
C3682 VN.n3264 a_400_62400# 1.22fF
C3683 VN.n3265 a_400_62400# 0.07fF
C3684 VN.t403 a_400_62400# 0.03fF
C3685 VN.n3266 a_400_62400# 0.16fF
C3686 VN.n3267 a_400_62400# 0.19fF
C3687 VN.n3269 a_400_62400# 2.51fF
C3688 VN.n3270 a_400_62400# 0.56fF
C3689 VN.n3271 a_400_62400# 0.64fF
C3690 VN.n3272 a_400_62400# 0.12fF
C3691 VN.n3273 a_400_62400# 0.44fF
C3692 VN.n3274 a_400_62400# 0.40fF
C3693 VN.n3275 a_400_62400# 1.03fF
C3694 VN.n3276 a_400_62400# 0.79fF
C3695 VN.t482 a_400_62400# 0.03fF
C3696 VN.n3277 a_400_62400# 0.32fF
C3697 VN.n3278 a_400_62400# 0.48fF
C3698 VN.n3279 a_400_62400# 0.81fF
C3699 VN.n3280 a_400_62400# 0.16fF
C3700 VN.t1841 a_400_62400# 0.03fF
C3701 VN.n3281 a_400_62400# 0.19fF
C3702 VN.n3283 a_400_62400# 3.50fF
C3703 VN.n3284 a_400_62400# 2.89fF
C3704 VN.t2438 a_400_62400# 0.03fF
C3705 VN.n3285 a_400_62400# 0.32fF
C3706 VN.n3286 a_400_62400# 1.22fF
C3707 VN.n3287 a_400_62400# 0.07fF
C3708 VN.t2052 a_400_62400# 0.03fF
C3709 VN.n3288 a_400_62400# 0.16fF
C3710 VN.n3289 a_400_62400# 0.19fF
C3711 VN.n3291 a_400_62400# 1.05fF
C3712 VN.n3292 a_400_62400# 3.07fF
C3713 VN.n3293 a_400_62400# 2.51fF
C3714 VN.n3294 a_400_62400# 0.16fF
C3715 VN.t2335 a_400_62400# 0.03fF
C3716 VN.n3295 a_400_62400# 0.19fF
C3717 VN.t930 a_400_62400# 0.03fF
C3718 VN.n3297 a_400_62400# 0.32fF
C3719 VN.n3298 a_400_62400# 0.48fF
C3720 VN.n3299 a_400_62400# 0.81fF
C3721 VN.n3300 a_400_62400# 1.86fF
C3722 VN.n3301 a_400_62400# 1.53fF
C3723 VN.n3302 a_400_62400# 0.47fF
C3724 VN.n3303 a_400_62400# 2.71fF
C3725 VN.t411 a_400_62400# 0.03fF
C3726 VN.n3304 a_400_62400# 0.32fF
C3727 VN.n3305 a_400_62400# 1.22fF
C3728 VN.n3306 a_400_62400# 0.07fF
C3729 VN.t2517 a_400_62400# 0.03fF
C3730 VN.n3307 a_400_62400# 0.16fF
C3731 VN.n3308 a_400_62400# 0.19fF
C3732 VN.n3310 a_400_62400# 2.53fF
C3733 VN.n3311 a_400_62400# 2.51fF
C3734 VN.t5 a_400_62400# 0.03fF
C3735 VN.n3312 a_400_62400# 0.32fF
C3736 VN.n3313 a_400_62400# 0.48fF
C3737 VN.n3314 a_400_62400# 0.81fF
C3738 VN.n3315 a_400_62400# 0.16fF
C3739 VN.t1470 a_400_62400# 0.03fF
C3740 VN.n3316 a_400_62400# 0.19fF
C3741 VN.n3318 a_400_62400# 1.55fF
C3742 VN.n3319 a_400_62400# 0.29fF
C3743 VN.n3320 a_400_62400# 2.52fF
C3744 VN.t2060 a_400_62400# 0.03fF
C3745 VN.n3321 a_400_62400# 0.32fF
C3746 VN.n3322 a_400_62400# 1.22fF
C3747 VN.n3323 a_400_62400# 0.07fF
C3748 VN.t1657 a_400_62400# 0.03fF
C3749 VN.n3324 a_400_62400# 0.16fF
C3750 VN.n3325 a_400_62400# 0.19fF
C3751 VN.n3327 a_400_62400# 27.83fF
C3752 VN.n3328 a_400_62400# 3.93fF
C3753 VN.n3329 a_400_62400# 2.51fF
C3754 VN.n3330 a_400_62400# 0.16fF
C3755 VN.t725 a_400_62400# 0.03fF
C3756 VN.n3331 a_400_62400# 0.19fF
C3757 VN.t1725 a_400_62400# 0.03fF
C3758 VN.n3333 a_400_62400# 0.32fF
C3759 VN.n3334 a_400_62400# 0.48fF
C3760 VN.n3335 a_400_62400# 0.81fF
C3761 VN.n3336 a_400_62400# 1.46fF
C3762 VN.n3337 a_400_62400# 0.21fF
C3763 VN.n3338 a_400_62400# 2.81fF
C3764 VN.t789 a_400_62400# 0.03fF
C3765 VN.n3339 a_400_62400# 0.16fF
C3766 VN.n3340 a_400_62400# 0.19fF
C3767 VN.t1189 a_400_62400# 0.03fF
C3768 VN.n3342 a_400_62400# 0.32fF
C3769 VN.n3343 a_400_62400# 1.22fF
C3770 VN.n3344 a_400_62400# 0.07fF
C3771 VN.n3345 a_400_62400# 2.51fF
C3772 VN.n3346 a_400_62400# 3.57fF
C3773 VN.t979 a_400_62400# 0.03fF
C3774 VN.n3347 a_400_62400# 0.32fF
C3775 VN.n3348 a_400_62400# 0.48fF
C3776 VN.n3349 a_400_62400# 0.81fF
C3777 VN.n3350 a_400_62400# 0.16fF
C3778 VN.t2377 a_400_62400# 0.03fF
C3779 VN.n3351 a_400_62400# 0.19fF
C3780 VN.n3353 a_400_62400# 3.93fF
C3781 VN.n3354 a_400_62400# 3.08fF
C3782 VN.t2442 a_400_62400# 0.03fF
C3783 VN.n3355 a_400_62400# 0.16fF
C3784 VN.n3356 a_400_62400# 0.19fF
C3785 VN.t461 a_400_62400# 0.03fF
C3786 VN.n3358 a_400_62400# 0.32fF
C3787 VN.n3359 a_400_62400# 1.22fF
C3788 VN.n3360 a_400_62400# 0.07fF
C3789 VN.n3361 a_400_62400# 2.51fF
C3790 VN.n3362 a_400_62400# 3.57fF
C3791 VN.t87 a_400_62400# 0.03fF
C3792 VN.n3363 a_400_62400# 0.32fF
C3793 VN.n3364 a_400_62400# 0.48fF
C3794 VN.n3365 a_400_62400# 0.81fF
C3795 VN.n3366 a_400_62400# 0.16fF
C3796 VN.t1510 a_400_62400# 0.03fF
C3797 VN.n3367 a_400_62400# 0.19fF
C3798 VN.n3369 a_400_62400# 3.75fF
C3799 VN.n3370 a_400_62400# 3.08fF
C3800 VN.t1579 a_400_62400# 0.03fF
C3801 VN.n3371 a_400_62400# 0.16fF
C3802 VN.n3372 a_400_62400# 0.19fF
C3803 VN.t2110 a_400_62400# 0.03fF
C3804 VN.n3374 a_400_62400# 0.32fF
C3805 VN.n3375 a_400_62400# 1.22fF
C3806 VN.n3376 a_400_62400# 0.07fF
C3807 VN.n3377 a_400_62400# 2.51fF
C3808 VN.n3378 a_400_62400# 3.57fF
C3809 VN.t1765 a_400_62400# 0.03fF
C3810 VN.n3379 a_400_62400# 0.32fF
C3811 VN.n3380 a_400_62400# 0.48fF
C3812 VN.n3381 a_400_62400# 0.81fF
C3813 VN.n3382 a_400_62400# 0.16fF
C3814 VN.t641 a_400_62400# 0.03fF
C3815 VN.n3383 a_400_62400# 0.19fF
C3816 VN.n3385 a_400_62400# 3.75fF
C3817 VN.n3386 a_400_62400# 3.08fF
C3818 VN.t712 a_400_62400# 0.03fF
C3819 VN.n3387 a_400_62400# 0.16fF
C3820 VN.n3388 a_400_62400# 0.19fF
C3821 VN.t1233 a_400_62400# 0.03fF
C3822 VN.n3390 a_400_62400# 0.32fF
C3823 VN.n3391 a_400_62400# 1.22fF
C3824 VN.n3392 a_400_62400# 0.07fF
C3825 VN.n3393 a_400_62400# 2.51fF
C3826 VN.n3394 a_400_62400# 3.57fF
C3827 VN.t894 a_400_62400# 0.03fF
C3828 VN.n3395 a_400_62400# 0.32fF
C3829 VN.n3396 a_400_62400# 0.48fF
C3830 VN.n3397 a_400_62400# 0.81fF
C3831 VN.n3398 a_400_62400# 0.16fF
C3832 VN.t2300 a_400_62400# 0.03fF
C3833 VN.n3399 a_400_62400# 0.19fF
C3834 VN.n3401 a_400_62400# 3.75fF
C3835 VN.n3402 a_400_62400# 3.08fF
C3836 VN.t2367 a_400_62400# 0.03fF
C3837 VN.n3403 a_400_62400# 0.16fF
C3838 VN.n3404 a_400_62400# 0.19fF
C3839 VN.t369 a_400_62400# 0.03fF
C3840 VN.n3406 a_400_62400# 0.32fF
C3841 VN.n3407 a_400_62400# 1.22fF
C3842 VN.n3408 a_400_62400# 0.07fF
C3843 VN.n3409 a_400_62400# 2.51fF
C3844 VN.n3410 a_400_62400# 3.57fF
C3845 VN.t2557 a_400_62400# 0.03fF
C3846 VN.n3411 a_400_62400# 0.32fF
C3847 VN.n3412 a_400_62400# 0.48fF
C3848 VN.n3413 a_400_62400# 0.81fF
C3849 VN.n3414 a_400_62400# 0.16fF
C3850 VN.t1427 a_400_62400# 0.03fF
C3851 VN.n3415 a_400_62400# 0.19fF
C3852 VN.n3417 a_400_62400# 3.75fF
C3853 VN.n3418 a_400_62400# 3.08fF
C3854 VN.t1620 a_400_62400# 0.03fF
C3855 VN.n3419 a_400_62400# 0.16fF
C3856 VN.n3420 a_400_62400# 0.19fF
C3857 VN.t2021 a_400_62400# 0.03fF
C3858 VN.n3422 a_400_62400# 0.32fF
C3859 VN.n3423 a_400_62400# 1.22fF
C3860 VN.n3424 a_400_62400# 0.07fF
C3861 VN.n3425 a_400_62400# 2.51fF
C3862 VN.n3426 a_400_62400# 3.57fF
C3863 VN.t1687 a_400_62400# 0.03fF
C3864 VN.n3427 a_400_62400# 0.32fF
C3865 VN.n3428 a_400_62400# 0.48fF
C3866 VN.n3429 a_400_62400# 0.81fF
C3867 VN.n3430 a_400_62400# 0.16fF
C3868 VN.t562 a_400_62400# 0.03fF
C3869 VN.n3431 a_400_62400# 0.19fF
C3870 VN.n3433 a_400_62400# 3.75fF
C3871 VN.n3434 a_400_62400# 3.08fF
C3872 VN.t749 a_400_62400# 0.03fF
C3873 VN.n3435 a_400_62400# 0.16fF
C3874 VN.n3436 a_400_62400# 0.19fF
C3875 VN.t1146 a_400_62400# 0.03fF
C3876 VN.n3438 a_400_62400# 0.32fF
C3877 VN.n3439 a_400_62400# 1.22fF
C3878 VN.n3440 a_400_62400# 0.07fF
C3879 VN.n3441 a_400_62400# 2.51fF
C3880 VN.n3442 a_400_62400# 3.57fF
C3881 VN.t952 a_400_62400# 0.03fF
C3882 VN.n3443 a_400_62400# 0.32fF
C3883 VN.n3444 a_400_62400# 0.48fF
C3884 VN.n3445 a_400_62400# 0.81fF
C3885 VN.n3446 a_400_62400# 0.16fF
C3886 VN.t2347 a_400_62400# 0.03fF
C3887 VN.n3447 a_400_62400# 0.19fF
C3888 VN.n3449 a_400_62400# 3.75fF
C3889 VN.n3450 a_400_62400# 3.08fF
C3890 VN.t2528 a_400_62400# 0.03fF
C3891 VN.n3451 a_400_62400# 0.16fF
C3892 VN.n3452 a_400_62400# 0.19fF
C3893 VN.t1898 a_400_62400# 0.03fF
C3894 VN.n3454 a_400_62400# 0.32fF
C3895 VN.n3455 a_400_62400# 1.22fF
C3896 VN.n3456 a_400_62400# 0.07fF
C3897 VN.n3457 a_400_62400# 2.51fF
C3898 VN.n3458 a_400_62400# 3.57fF
C3899 VN.t34 a_400_62400# 0.03fF
C3900 VN.n3459 a_400_62400# 0.32fF
C3901 VN.n3460 a_400_62400# 0.48fF
C3902 VN.n3461 a_400_62400# 0.81fF
C3903 VN.n3462 a_400_62400# 0.16fF
C3904 VN.t1477 a_400_62400# 0.03fF
C3905 VN.n3463 a_400_62400# 0.19fF
C3906 VN.n3465 a_400_62400# 3.75fF
C3907 VN.n3466 a_400_62400# 3.08fF
C3908 VN.t1664 a_400_62400# 0.03fF
C3909 VN.n3467 a_400_62400# 0.16fF
C3910 VN.n3468 a_400_62400# 0.19fF
C3911 VN.t1023 a_400_62400# 0.03fF
C3912 VN.n3470 a_400_62400# 0.32fF
C3913 VN.n3471 a_400_62400# 1.22fF
C3914 VN.n3472 a_400_62400# 0.07fF
C3915 VN.n3473 a_400_62400# 3.65fF
C3916 VN.n3474 a_400_62400# 2.14fF
C3917 VN.n3475 a_400_62400# 0.16fF
C3918 VN.t2388 a_400_62400# 0.03fF
C3919 VN.n3476 a_400_62400# 0.19fF
C3920 VN.t868 a_400_62400# 0.03fF
C3921 VN.n3478 a_400_62400# 0.32fF
C3922 VN.n3479 a_400_62400# 0.48fF
C3923 VN.n3480 a_400_62400# 0.81fF
C3924 VN.n3481 a_400_62400# 0.09fF
C3925 VN.n3482 a_400_62400# 0.01fF
C3926 VN.n3483 a_400_62400# 0.02fF
C3927 VN.n3484 a_400_62400# 0.02fF
C3928 VN.n3485 a_400_62400# 0.32fF
C3929 VN.n3486 a_400_62400# 1.56fF
C3930 VN.n3487 a_400_62400# 1.81fF
C3931 VN.n3488 a_400_62400# 3.08fF
C3932 VN.t2450 a_400_62400# 0.03fF
C3933 VN.n3489 a_400_62400# 0.16fF
C3934 VN.n3490 a_400_62400# 0.19fF
C3935 VN.t1814 a_400_62400# 0.03fF
C3936 VN.n3492 a_400_62400# 0.32fF
C3937 VN.n3493 a_400_62400# 1.22fF
C3938 VN.n3494 a_400_62400# 0.07fF
C3939 VN.t183 a_400_62400# 64.69fF
C3940 VN.t151 a_400_62400# 0.03fF
C3941 VN.n3495 a_400_62400# 0.32fF
C3942 VN.n3496 a_400_62400# 1.22fF
C3943 VN.n3497 a_400_62400# 0.07fF
C3944 VN.t796 a_400_62400# 0.03fF
C3945 VN.n3498 a_400_62400# 0.16fF
C3946 VN.n3499 a_400_62400# 0.19fF
C3947 VN.n3501 a_400_62400# 0.16fF
C3948 VN.t609 a_400_62400# 0.03fF
C3949 VN.n3502 a_400_62400# 0.19fF
C3950 VN.n3504 a_400_62400# 6.92fF
C3951 VN.n3505 a_400_62400# 6.56fF
C3952 VN.t1574 a_400_62400# 0.03fF
C3953 VN.n3506 a_400_62400# 0.16fF
C3954 VN.n3507 a_400_62400# 0.19fF
C3955 VN.t1945 a_400_62400# 0.03fF
C3956 VN.n3509 a_400_62400# 0.32fF
C3957 VN.n3510 a_400_62400# 1.22fF
C3958 VN.n3511 a_400_62400# 0.07fF
C3959 VN.n3512 a_400_62400# 2.51fF
C3960 VN.n3513 a_400_62400# 3.58fF
C3961 VN.t2038 a_400_62400# 0.03fF
C3962 VN.n3514 a_400_62400# 0.32fF
C3963 VN.n3515 a_400_62400# 0.48fF
C3964 VN.n3516 a_400_62400# 0.81fF
C3965 VN.n3517 a_400_62400# 0.16fF
C3966 VN.t2544 a_400_62400# 0.03fF
C3967 VN.n3518 a_400_62400# 0.19fF
C3968 VN.n3520 a_400_62400# 7.29fF
C3969 VN.t705 a_400_62400# 0.03fF
C3970 VN.n3521 a_400_62400# 0.16fF
C3971 VN.n3522 a_400_62400# 0.19fF
C3972 VN.t1075 a_400_62400# 0.03fF
C3973 VN.n3524 a_400_62400# 0.32fF
C3974 VN.n3525 a_400_62400# 1.22fF
C3975 VN.n3526 a_400_62400# 0.07fF
C3976 VN.t63 a_400_62400# 64.17fF
C3977 VN.t200 a_400_62400# 0.03fF
C3978 VN.n3527 a_400_62400# 1.60fF
C3979 VN.n3528 a_400_62400# 0.07fF
C3980 VN.t2478 a_400_62400# 0.03fF
C3981 VN.n3529 a_400_62400# 0.02fF
C3982 VN.n3530 a_400_62400# 0.34fF
C3983 VN.n3532 a_400_62400# 2.01fF
C3984 VN.n3533 a_400_62400# 1.75fF
C3985 VN.n3534 a_400_62400# 0.37fF
C3986 VN.n3535 a_400_62400# 0.33fF
C3987 VN.n3536 a_400_62400# 5.88fF
C3988 VN.n3537 a_400_62400# 0.02fF
C3989 VN.n3538 a_400_62400# 0.02fF
C3990 VN.n3539 a_400_62400# 0.03fF
C3991 VN.n3540 a_400_62400# 0.05fF
C3992 VN.n3541 a_400_62400# 0.23fF
C3993 VN.n3542 a_400_62400# 0.02fF
C3994 VN.n3543 a_400_62400# 0.03fF
C3995 VN.n3544 a_400_62400# 0.01fF
C3996 VN.n3545 a_400_62400# 0.01fF
C3997 VN.n3546 a_400_62400# 0.01fF
C3998 VN.n3547 a_400_62400# 0.02fF
C3999 VN.n3548 a_400_62400# 0.03fF
C4000 VN.n3549 a_400_62400# 0.06fF
C4001 VN.n3550 a_400_62400# 0.05fF
C4002 VN.n3551 a_400_62400# 0.15fF
C4003 VN.n3552 a_400_62400# 0.51fF
C4004 VN.n3553 a_400_62400# 0.27fF
C4005 VN.n3554 a_400_62400# 37.46fF
C4006 VN.n3555 a_400_62400# 37.46fF
C4007 VN.n3556 a_400_62400# 0.79fF
C4008 VN.n3557 a_400_62400# 0.23fF
C4009 VN.n3558 a_400_62400# 1.18fF
C4010 VN.t68 a_400_62400# 28.64fF
C4011 VN.n3559 a_400_62400# 0.79fF
C4012 VN.n3560 a_400_62400# 0.11fF
C4013 VN.n3561 a_400_62400# 4.98fF
C4014 VN.n3562 a_400_62400# 0.80fF
C4015 VN.n3563 a_400_62400# 0.29fF
C4016 VN.n3564 a_400_62400# 1.96fF
C4017 VN.n3566 a_400_62400# 25.18fF
C4018 VN.n3568 a_400_62400# 1.87fF
C4019 VN.n3569 a_400_62400# 5.36fF
C4020 VN.n3570 a_400_62400# 1.81fF
C4021 VN.t1149 a_400_62400# 0.03fF
C4022 VN.n3571 a_400_62400# 0.85fF
C4023 VN.n3572 a_400_62400# 0.81fF
C4024 VN.n3573 a_400_62400# 2.53fF
C4025 VN.n3574 a_400_62400# 0.08fF
C4026 VN.n3575 a_400_62400# 0.04fF
C4027 VN.n3576 a_400_62400# 0.05fF
C4028 VN.n3577 a_400_62400# 1.33fF
C4029 VN.n3578 a_400_62400# 0.03fF
C4030 VN.n3579 a_400_62400# 0.01fF
C4031 VN.n3580 a_400_62400# 0.02fF
C4032 VN.n3581 a_400_62400# 0.11fF
C4033 VN.n3582 a_400_62400# 0.48fF
C4034 VN.n3583 a_400_62400# 2.48fF
C4035 VN.t1714 a_400_62400# 0.03fF
C4036 VN.n3584 a_400_62400# 0.32fF
C4037 VN.n3585 a_400_62400# 0.48fF
C4038 VN.n3586 a_400_62400# 0.81fF
C4039 VN.n3587 a_400_62400# 0.16fF
C4040 VN.t714 a_400_62400# 0.03fF
C4041 VN.n3588 a_400_62400# 0.19fF
C4042 VN.n3590 a_400_62400# 0.93fF
C4043 VN.n3591 a_400_62400# 0.30fF
C4044 VN.n3592 a_400_62400# 0.34fF
C4045 VN.n3593 a_400_62400# 0.12fF
C4046 VN.n3594 a_400_62400# 0.30fF
C4047 VN.n3595 a_400_62400# 0.93fF
C4048 VN.n3596 a_400_62400# 1.55fF
C4049 VN.n3597 a_400_62400# 0.29fF
C4050 VN.n3598 a_400_62400# 0.34fF
C4051 VN.n3599 a_400_62400# 0.12fF
C4052 VN.n3600 a_400_62400# 2.52fF
C4053 VN.t2549 a_400_62400# 0.03fF
C4054 VN.n3601 a_400_62400# 0.32fF
C4055 VN.n3602 a_400_62400# 1.22fF
C4056 VN.n3603 a_400_62400# 0.07fF
C4057 VN.t1393 a_400_62400# 0.03fF
C4058 VN.n3604 a_400_62400# 0.16fF
C4059 VN.n3605 a_400_62400# 0.19fF
C4060 VN.n3607 a_400_62400# 0.33fF
C4061 VN.n3608 a_400_62400# 0.12fF
C4062 VN.n3609 a_400_62400# 0.28fF
C4063 VN.n3610 a_400_62400# 1.23fF
C4064 VN.n3611 a_400_62400# 0.59fF
C4065 VN.n3612 a_400_62400# 2.51fF
C4066 VN.n3613 a_400_62400# 0.16fF
C4067 VN.t2369 a_400_62400# 0.03fF
C4068 VN.n3614 a_400_62400# 0.19fF
C4069 VN.t968 a_400_62400# 0.03fF
C4070 VN.n3616 a_400_62400# 0.32fF
C4071 VN.n3617 a_400_62400# 0.48fF
C4072 VN.n3618 a_400_62400# 0.81fF
C4073 VN.n3619 a_400_62400# 0.03fF
C4074 VN.n3620 a_400_62400# 0.01fF
C4075 VN.n3621 a_400_62400# 0.02fF
C4076 VN.n3622 a_400_62400# 0.11fF
C4077 VN.n3623 a_400_62400# 0.08fF
C4078 VN.n3624 a_400_62400# 0.04fF
C4079 VN.n3625 a_400_62400# 0.05fF
C4080 VN.n3626 a_400_62400# 1.34fF
C4081 VN.n3627 a_400_62400# 0.48fF
C4082 VN.n3628 a_400_62400# 2.51fF
C4083 VN.n3629 a_400_62400# 2.67fF
C4084 VN.t1808 a_400_62400# 0.03fF
C4085 VN.n3630 a_400_62400# 0.32fF
C4086 VN.n3631 a_400_62400# 1.22fF
C4087 VN.n3632 a_400_62400# 0.07fF
C4088 VN.t530 a_400_62400# 0.03fF
C4089 VN.n3633 a_400_62400# 0.16fF
C4090 VN.n3634 a_400_62400# 0.19fF
C4091 VN.n3636 a_400_62400# 2.53fF
C4092 VN.n3637 a_400_62400# 0.09fF
C4093 VN.n3638 a_400_62400# 0.05fF
C4094 VN.n3639 a_400_62400# 0.07fF
C4095 VN.n3640 a_400_62400# 1.16fF
C4096 VN.n3641 a_400_62400# 0.01fF
C4097 VN.n3642 a_400_62400# 0.01fF
C4098 VN.n3643 a_400_62400# 0.01fF
C4099 VN.n3644 a_400_62400# 0.09fF
C4100 VN.n3645 a_400_62400# 0.91fF
C4101 VN.n3646 a_400_62400# 0.96fF
C4102 VN.t69 a_400_62400# 0.03fF
C4103 VN.n3647 a_400_62400# 0.32fF
C4104 VN.n3648 a_400_62400# 0.48fF
C4105 VN.n3649 a_400_62400# 0.81fF
C4106 VN.n3650 a_400_62400# 0.16fF
C4107 VN.t1500 a_400_62400# 0.03fF
C4108 VN.n3651 a_400_62400# 0.19fF
C4109 VN.n3653 a_400_62400# 0.93fF
C4110 VN.n3654 a_400_62400# 0.30fF
C4111 VN.n3655 a_400_62400# 0.34fF
C4112 VN.n3656 a_400_62400# 0.12fF
C4113 VN.n3657 a_400_62400# 0.30fF
C4114 VN.n3658 a_400_62400# 0.93fF
C4115 VN.n3659 a_400_62400# 1.55fF
C4116 VN.n3660 a_400_62400# 0.29fF
C4117 VN.n3661 a_400_62400# 0.34fF
C4118 VN.n3662 a_400_62400# 0.12fF
C4119 VN.n3663 a_400_62400# 3.10fF
C4120 VN.t932 a_400_62400# 0.03fF
C4121 VN.n3664 a_400_62400# 0.32fF
C4122 VN.n3665 a_400_62400# 1.22fF
C4123 VN.n3666 a_400_62400# 0.07fF
C4124 VN.t2185 a_400_62400# 0.03fF
C4125 VN.n3667 a_400_62400# 0.16fF
C4126 VN.n3668 a_400_62400# 0.19fF
C4127 VN.n3670 a_400_62400# 2.51fF
C4128 VN.n3671 a_400_62400# 0.61fF
C4129 VN.n3672 a_400_62400# 0.30fF
C4130 VN.n3673 a_400_62400# 0.51fF
C4131 VN.n3674 a_400_62400# 0.21fF
C4132 VN.n3675 a_400_62400# 0.38fF
C4133 VN.n3676 a_400_62400# 0.29fF
C4134 VN.n3677 a_400_62400# 0.40fF
C4135 VN.n3678 a_400_62400# 0.28fF
C4136 VN.t599 a_400_62400# 0.03fF
C4137 VN.n3679 a_400_62400# 0.32fF
C4138 VN.n3680 a_400_62400# 0.48fF
C4139 VN.n3681 a_400_62400# 0.81fF
C4140 VN.n3682 a_400_62400# 0.16fF
C4141 VN.t1973 a_400_62400# 0.03fF
C4142 VN.n3683 a_400_62400# 0.19fF
C4143 VN.n3685 a_400_62400# 0.06fF
C4144 VN.n3686 a_400_62400# 0.04fF
C4145 VN.n3687 a_400_62400# 0.04fF
C4146 VN.n3688 a_400_62400# 0.14fF
C4147 VN.n3689 a_400_62400# 0.48fF
C4148 VN.n3690 a_400_62400# 0.50fF
C4149 VN.n3691 a_400_62400# 0.14fF
C4150 VN.n3692 a_400_62400# 0.16fF
C4151 VN.n3693 a_400_62400# 0.09fF
C4152 VN.n3694 a_400_62400# 0.16fF
C4153 VN.n3695 a_400_62400# 0.24fF
C4154 VN.n3696 a_400_62400# 5.35fF
C4155 VN.t1429 a_400_62400# 0.03fF
C4156 VN.n3697 a_400_62400# 0.32fF
C4157 VN.n3698 a_400_62400# 1.22fF
C4158 VN.n3699 a_400_62400# 0.07fF
C4159 VN.t1318 a_400_62400# 0.03fF
C4160 VN.n3700 a_400_62400# 0.16fF
C4161 VN.n3701 a_400_62400# 0.19fF
C4162 VN.n3703 a_400_62400# 0.33fF
C4163 VN.n3704 a_400_62400# 0.12fF
C4164 VN.n3705 a_400_62400# 0.28fF
C4165 VN.n3706 a_400_62400# 1.72fF
C4166 VN.n3707 a_400_62400# 0.71fF
C4167 VN.n3708 a_400_62400# 2.51fF
C4168 VN.n3709 a_400_62400# 0.16fF
C4169 VN.t1105 a_400_62400# 0.03fF
C4170 VN.n3710 a_400_62400# 0.19fF
C4171 VN.t2254 a_400_62400# 0.03fF
C4172 VN.n3712 a_400_62400# 0.32fF
C4173 VN.n3713 a_400_62400# 0.48fF
C4174 VN.n3714 a_400_62400# 0.81fF
C4175 VN.n3715 a_400_62400# 0.95fF
C4176 VN.n3716 a_400_62400# 2.11fF
C4177 VN.n3717 a_400_62400# 3.28fF
C4178 VN.t563 a_400_62400# 0.03fF
C4179 VN.n3718 a_400_62400# 0.32fF
C4180 VN.n3719 a_400_62400# 1.22fF
C4181 VN.n3720 a_400_62400# 0.07fF
C4182 VN.t1771 a_400_62400# 0.03fF
C4183 VN.n3721 a_400_62400# 0.16fF
C4184 VN.n3722 a_400_62400# 0.19fF
C4185 VN.n3724 a_400_62400# 2.53fF
C4186 VN.n3725 a_400_62400# 0.08fF
C4187 VN.n3726 a_400_62400# 0.04fF
C4188 VN.n3727 a_400_62400# 0.05fF
C4189 VN.n3728 a_400_62400# 1.33fF
C4190 VN.n3729 a_400_62400# 0.03fF
C4191 VN.n3730 a_400_62400# 0.01fF
C4192 VN.n3731 a_400_62400# 0.02fF
C4193 VN.n3732 a_400_62400# 0.11fF
C4194 VN.n3733 a_400_62400# 0.48fF
C4195 VN.n3734 a_400_62400# 2.48fF
C4196 VN.t1390 a_400_62400# 0.03fF
C4197 VN.n3735 a_400_62400# 0.32fF
C4198 VN.n3736 a_400_62400# 0.48fF
C4199 VN.n3737 a_400_62400# 0.81fF
C4200 VN.n3738 a_400_62400# 0.16fF
C4201 VN.t238 a_400_62400# 0.03fF
C4202 VN.n3739 a_400_62400# 0.19fF
C4203 VN.n3741 a_400_62400# 0.93fF
C4204 VN.n3742 a_400_62400# 0.30fF
C4205 VN.n3743 a_400_62400# 0.34fF
C4206 VN.n3744 a_400_62400# 0.12fF
C4207 VN.n3745 a_400_62400# 0.30fF
C4208 VN.n3746 a_400_62400# 0.93fF
C4209 VN.n3747 a_400_62400# 1.55fF
C4210 VN.n3748 a_400_62400# 0.29fF
C4211 VN.n3749 a_400_62400# 0.34fF
C4212 VN.n3750 a_400_62400# 0.12fF
C4213 VN.n3751 a_400_62400# 2.52fF
C4214 VN.t2222 a_400_62400# 0.03fF
C4215 VN.n3752 a_400_62400# 0.32fF
C4216 VN.n3753 a_400_62400# 1.22fF
C4217 VN.n3754 a_400_62400# 0.07fF
C4218 VN.t899 a_400_62400# 0.03fF
C4219 VN.n3755 a_400_62400# 0.16fF
C4220 VN.n3756 a_400_62400# 0.19fF
C4221 VN.n3758 a_400_62400# 27.83fF
C4222 VN.n3759 a_400_62400# 0.09fF
C4223 VN.n3760 a_400_62400# 0.27fF
C4224 VN.n3761 a_400_62400# 0.12fF
C4225 VN.n3762 a_400_62400# 0.28fF
C4226 VN.n3763 a_400_62400# 0.13fF
C4227 VN.n3764 a_400_62400# 0.40fF
C4228 VN.n3765 a_400_62400# 0.93fF
C4229 VN.n3766 a_400_62400# 0.60fF
C4230 VN.n3767 a_400_62400# 3.12fF
C4231 VN.n3768 a_400_62400# 0.16fF
C4232 VN.t1465 a_400_62400# 0.03fF
C4233 VN.n3769 a_400_62400# 0.19fF
C4234 VN.t2583 a_400_62400# 0.03fF
C4235 VN.n3771 a_400_62400# 0.32fF
C4236 VN.n3772 a_400_62400# 0.48fF
C4237 VN.n3773 a_400_62400# 0.81fF
C4238 VN.n3774 a_400_62400# 2.54fF
C4239 VN.n3775 a_400_62400# 0.23fF
C4240 VN.n3776 a_400_62400# 1.02fF
C4241 VN.n3777 a_400_62400# 0.34fF
C4242 VN.n3778 a_400_62400# 0.40fF
C4243 VN.n3779 a_400_62400# 0.42fF
C4244 VN.n3780 a_400_62400# 0.63fF
C4245 VN.n3781 a_400_62400# 0.21fF
C4246 VN.n3782 a_400_62400# 2.58fF
C4247 VN.t2259 a_400_62400# 0.03fF
C4248 VN.n3783 a_400_62400# 0.16fF
C4249 VN.n3784 a_400_62400# 0.19fF
C4250 VN.t888 a_400_62400# 0.03fF
C4251 VN.n3786 a_400_62400# 0.32fF
C4252 VN.n3787 a_400_62400# 1.22fF
C4253 VN.n3788 a_400_62400# 0.07fF
C4254 VN.n3789 a_400_62400# 2.51fF
C4255 VN.n3790 a_400_62400# 0.16fF
C4256 VN.t1888 a_400_62400# 0.03fF
C4257 VN.n3791 a_400_62400# 0.19fF
C4258 VN.t524 a_400_62400# 0.03fF
C4259 VN.n3793 a_400_62400# 0.32fF
C4260 VN.n3794 a_400_62400# 0.48fF
C4261 VN.n3795 a_400_62400# 0.81fF
C4262 VN.n3796 a_400_62400# 1.24fF
C4263 VN.n3797 a_400_62400# 0.43fF
C4264 VN.n3798 a_400_62400# 0.43fF
C4265 VN.n3799 a_400_62400# 1.24fF
C4266 VN.n3800 a_400_62400# 1.46fF
C4267 VN.n3801 a_400_62400# 0.21fF
C4268 VN.n3802 a_400_62400# 6.64fF
C4269 VN.t154 a_400_62400# 0.03fF
C4270 VN.n3803 a_400_62400# 0.16fF
C4271 VN.n3804 a_400_62400# 0.19fF
C4272 VN.t1357 a_400_62400# 0.03fF
C4273 VN.n3806 a_400_62400# 0.32fF
C4274 VN.n3807 a_400_62400# 1.22fF
C4275 VN.n3808 a_400_62400# 0.07fF
C4276 VN.n3809 a_400_62400# 2.51fF
C4277 VN.n3810 a_400_62400# 3.57fF
C4278 VN.t2179 a_400_62400# 0.03fF
C4279 VN.n3811 a_400_62400# 0.32fF
C4280 VN.n3812 a_400_62400# 0.48fF
C4281 VN.n3813 a_400_62400# 0.81fF
C4282 VN.n3814 a_400_62400# 0.16fF
C4283 VN.t1016 a_400_62400# 0.03fF
C4284 VN.n3815 a_400_62400# 0.19fF
C4285 VN.n3817 a_400_62400# 6.91fF
C4286 VN.t1817 a_400_62400# 0.03fF
C4287 VN.n3818 a_400_62400# 0.16fF
C4288 VN.n3819 a_400_62400# 0.19fF
C4289 VN.t490 a_400_62400# 0.03fF
C4290 VN.n3821 a_400_62400# 0.32fF
C4291 VN.n3822 a_400_62400# 1.22fF
C4292 VN.n3823 a_400_62400# 0.07fF
C4293 VN.n3824 a_400_62400# 2.51fF
C4294 VN.n3825 a_400_62400# 3.57fF
C4295 VN.t1311 a_400_62400# 0.03fF
C4296 VN.n3826 a_400_62400# 0.32fF
C4297 VN.n3827 a_400_62400# 0.48fF
C4298 VN.n3828 a_400_62400# 0.81fF
C4299 VN.n3829 a_400_62400# 0.16fF
C4300 VN.t142 a_400_62400# 0.03fF
C4301 VN.n3830 a_400_62400# 0.19fF
C4302 VN.n3832 a_400_62400# 6.92fF
C4303 VN.t944 a_400_62400# 0.03fF
C4304 VN.n3833 a_400_62400# 0.16fF
C4305 VN.n3834 a_400_62400# 0.19fF
C4306 VN.t2145 a_400_62400# 0.03fF
C4307 VN.n3836 a_400_62400# 0.32fF
C4308 VN.n3837 a_400_62400# 1.22fF
C4309 VN.n3838 a_400_62400# 0.07fF
C4310 VN.n3839 a_400_62400# 2.51fF
C4311 VN.n3840 a_400_62400# 3.57fF
C4312 VN.t450 a_400_62400# 0.03fF
C4313 VN.n3841 a_400_62400# 0.32fF
C4314 VN.n3842 a_400_62400# 0.48fF
C4315 VN.n3843 a_400_62400# 0.81fF
C4316 VN.n3844 a_400_62400# 0.16fF
C4317 VN.t1805 a_400_62400# 0.03fF
C4318 VN.n3845 a_400_62400# 0.19fF
C4319 VN.n3847 a_400_62400# 6.92fF
C4320 VN.t19 a_400_62400# 0.03fF
C4321 VN.n3848 a_400_62400# 0.16fF
C4322 VN.n3849 a_400_62400# 0.19fF
C4323 VN.t1275 a_400_62400# 0.03fF
C4324 VN.n3851 a_400_62400# 0.32fF
C4325 VN.n3852 a_400_62400# 1.22fF
C4326 VN.n3853 a_400_62400# 0.07fF
C4327 VN.n3854 a_400_62400# 2.51fF
C4328 VN.n3855 a_400_62400# 3.57fF
C4329 VN.t2096 a_400_62400# 0.03fF
C4330 VN.n3856 a_400_62400# 0.32fF
C4331 VN.n3857 a_400_62400# 0.48fF
C4332 VN.n3858 a_400_62400# 0.81fF
C4333 VN.n3859 a_400_62400# 0.16fF
C4334 VN.t1063 a_400_62400# 0.03fF
C4335 VN.n3860 a_400_62400# 0.19fF
C4336 VN.n3862 a_400_62400# 6.92fF
C4337 VN.t1734 a_400_62400# 0.03fF
C4338 VN.n3863 a_400_62400# 0.16fF
C4339 VN.n3864 a_400_62400# 0.19fF
C4340 VN.t405 a_400_62400# 0.03fF
C4341 VN.n3866 a_400_62400# 0.32fF
C4342 VN.n3867 a_400_62400# 1.22fF
C4343 VN.n3868 a_400_62400# 0.07fF
C4344 VN.n3869 a_400_62400# 2.51fF
C4345 VN.n3870 a_400_62400# 3.57fF
C4346 VN.t1356 a_400_62400# 0.03fF
C4347 VN.n3871 a_400_62400# 0.32fF
C4348 VN.n3872 a_400_62400# 0.48fF
C4349 VN.n3873 a_400_62400# 0.81fF
C4350 VN.n3874 a_400_62400# 0.16fF
C4351 VN.t189 a_400_62400# 0.03fF
C4352 VN.n3875 a_400_62400# 0.19fF
C4353 VN.n3877 a_400_62400# 6.92fF
C4354 VN.t860 a_400_62400# 0.03fF
C4355 VN.n3878 a_400_62400# 0.16fF
C4356 VN.n3879 a_400_62400# 0.19fF
C4357 VN.t2188 a_400_62400# 0.03fF
C4358 VN.n3881 a_400_62400# 0.32fF
C4359 VN.n3882 a_400_62400# 1.22fF
C4360 VN.n3883 a_400_62400# 0.07fF
C4361 VN.n3884 a_400_62400# 2.51fF
C4362 VN.n3885 a_400_62400# 3.57fF
C4363 VN.t2113 a_400_62400# 0.03fF
C4364 VN.n3886 a_400_62400# 0.32fF
C4365 VN.n3887 a_400_62400# 0.48fF
C4366 VN.n3888 a_400_62400# 0.81fF
C4367 VN.n3889 a_400_62400# 0.16fF
C4368 VN.t938 a_400_62400# 0.03fF
C4369 VN.n3890 a_400_62400# 0.19fF
C4370 VN.n3892 a_400_62400# 6.92fF
C4371 VN.t2522 a_400_62400# 0.03fF
C4372 VN.n3893 a_400_62400# 0.16fF
C4373 VN.n3894 a_400_62400# 0.19fF
C4374 VN.t2006 a_400_62400# 0.03fF
C4375 VN.n3896 a_400_62400# 0.32fF
C4376 VN.n3897 a_400_62400# 1.22fF
C4377 VN.n3898 a_400_62400# 0.07fF
C4378 VN.n3899 a_400_62400# 2.51fF
C4379 VN.n3900 a_400_62400# 3.57fF
C4380 VN.t1235 a_400_62400# 0.03fF
C4381 VN.n3901 a_400_62400# 0.32fF
C4382 VN.n3902 a_400_62400# 0.48fF
C4383 VN.n3903 a_400_62400# 0.81fF
C4384 VN.n3904 a_400_62400# 0.16fF
C4385 VN.t15 a_400_62400# 0.03fF
C4386 VN.n3905 a_400_62400# 0.19fF
C4387 VN.n3907 a_400_62400# 6.92fF
C4388 VN.t754 a_400_62400# 0.03fF
C4389 VN.n3908 a_400_62400# 0.16fF
C4390 VN.n3909 a_400_62400# 0.19fF
C4391 VN.t1133 a_400_62400# 0.03fF
C4392 VN.n3911 a_400_62400# 0.32fF
C4393 VN.n3912 a_400_62400# 1.22fF
C4394 VN.n3913 a_400_62400# 0.07fF
C4395 VN.n3914 a_400_62400# 2.51fF
C4396 VN.n3915 a_400_62400# 3.57fF
C4397 VN.t371 a_400_62400# 0.03fF
C4398 VN.n3916 a_400_62400# 0.32fF
C4399 VN.n3917 a_400_62400# 0.48fF
C4400 VN.n3918 a_400_62400# 0.81fF
C4401 VN.n3919 a_400_62400# 0.16fF
C4402 VN.t1731 a_400_62400# 0.03fF
C4403 VN.n3920 a_400_62400# 0.19fF
C4404 VN.n3922 a_400_62400# 2.51fF
C4405 VN.n3923 a_400_62400# 3.59fF
C4406 VN.t2589 a_400_62400# 0.03fF
C4407 VN.n3924 a_400_62400# 0.32fF
C4408 VN.n3925 a_400_62400# 0.48fF
C4409 VN.n3926 a_400_62400# 0.81fF
C4410 VN.t1694 a_400_62400# 0.03fF
C4411 VN.n3927 a_400_62400# 1.63fF
C4412 VN.n3928 a_400_62400# 0.81fF
C4413 VN.n3929 a_400_62400# 1.21fF
C4414 VN.n3930 a_400_62400# 1.54fF
C4415 VN.n3931 a_400_62400# 4.06fF
C4416 VN.t269 a_400_62400# 28.64fF
C4417 VN.n3932 a_400_62400# 28.43fF
C4418 VN.n3934 a_400_62400# 0.50fF
C4419 VN.n3935 a_400_62400# 0.31fF
C4420 VN.n3936 a_400_62400# 3.88fF
C4421 VN.n3937 a_400_62400# 3.29fF
C4422 VN.n3938 a_400_62400# 2.62fF
C4423 VN.n3939 a_400_62400# 5.27fF
C4424 VN.n3940 a_400_62400# 0.34fF
C4425 VN.n3941 a_400_62400# 0.02fF
C4426 VN.t569 a_400_62400# 0.03fF
C4427 VN.n3942 a_400_62400# 0.34fF
C4428 VN.t1154 a_400_62400# 0.03fF
C4429 VN.n3943 a_400_62400# 1.28fF
C4430 VN.n3944 a_400_62400# 0.94fF
C4431 VN.n3945 a_400_62400# 1.04fF
C4432 VN.n3946 a_400_62400# 2.58fF
C4433 VN.n3947 a_400_62400# 2.51fF
C4434 VN.n3948 a_400_62400# 0.16fF
C4435 VN.t2228 a_400_62400# 0.03fF
C4436 VN.n3949 a_400_62400# 0.19fF
C4437 VN.t824 a_400_62400# 0.03fF
C4438 VN.n3951 a_400_62400# 0.32fF
C4439 VN.n3952 a_400_62400# 0.48fF
C4440 VN.n3953 a_400_62400# 0.81fF
C4441 VN.n3954 a_400_62400# 2.03fF
C4442 VN.n3955 a_400_62400# 4.01fF
C4443 VN.t288 a_400_62400# 0.03fF
C4444 VN.n3956 a_400_62400# 0.32fF
C4445 VN.n3957 a_400_62400# 1.22fF
C4446 VN.n3958 a_400_62400# 0.07fF
C4447 VN.t2296 a_400_62400# 0.03fF
C4448 VN.n3959 a_400_62400# 0.16fF
C4449 VN.n3960 a_400_62400# 0.19fF
C4450 VN.n3962 a_400_62400# 2.53fF
C4451 VN.n3963 a_400_62400# 2.51fF
C4452 VN.t2485 a_400_62400# 0.03fF
C4453 VN.n3964 a_400_62400# 0.32fF
C4454 VN.n3965 a_400_62400# 0.48fF
C4455 VN.n3966 a_400_62400# 0.81fF
C4456 VN.n3967 a_400_62400# 0.16fF
C4457 VN.t1362 a_400_62400# 0.03fF
C4458 VN.n3968 a_400_62400# 0.19fF
C4459 VN.n3970 a_400_62400# 1.55fF
C4460 VN.n3971 a_400_62400# 0.29fF
C4461 VN.n3972 a_400_62400# 2.52fF
C4462 VN.t1940 a_400_62400# 0.03fF
C4463 VN.n3973 a_400_62400# 0.32fF
C4464 VN.n3974 a_400_62400# 1.22fF
C4465 VN.n3975 a_400_62400# 0.07fF
C4466 VN.t1549 a_400_62400# 0.03fF
C4467 VN.n3976 a_400_62400# 0.16fF
C4468 VN.n3977 a_400_62400# 0.19fF
C4469 VN.n3979 a_400_62400# 1.04fF
C4470 VN.n3980 a_400_62400# 2.60fF
C4471 VN.n3981 a_400_62400# 2.51fF
C4472 VN.n3982 a_400_62400# 0.16fF
C4473 VN.t495 a_400_62400# 0.03fF
C4474 VN.n3983 a_400_62400# 0.19fF
C4475 VN.t1621 a_400_62400# 0.03fF
C4476 VN.n3985 a_400_62400# 0.32fF
C4477 VN.n3986 a_400_62400# 0.48fF
C4478 VN.n3987 a_400_62400# 0.81fF
C4479 VN.n3988 a_400_62400# 2.46fF
C4480 VN.n3989 a_400_62400# 4.01fF
C4481 VN.t1067 a_400_62400# 0.03fF
C4482 VN.n3990 a_400_62400# 0.32fF
C4483 VN.n3991 a_400_62400# 1.22fF
C4484 VN.n3992 a_400_62400# 0.07fF
C4485 VN.t676 a_400_62400# 0.03fF
C4486 VN.n3993 a_400_62400# 0.16fF
C4487 VN.n3994 a_400_62400# 0.19fF
C4488 VN.n3996 a_400_62400# 2.53fF
C4489 VN.n3997 a_400_62400# 2.34fF
C4490 VN.t750 a_400_62400# 0.03fF
C4491 VN.n3998 a_400_62400# 0.32fF
C4492 VN.n3999 a_400_62400# 0.48fF
C4493 VN.n4000 a_400_62400# 0.81fF
C4494 VN.n4001 a_400_62400# 0.16fF
C4495 VN.t2152 a_400_62400# 0.03fF
C4496 VN.n4002 a_400_62400# 0.19fF
C4497 VN.n4004 a_400_62400# 1.55fF
C4498 VN.n4005 a_400_62400# 0.29fF
C4499 VN.n4006 a_400_62400# 3.27fF
C4500 VN.t193 a_400_62400# 0.03fF
C4501 VN.n4007 a_400_62400# 0.32fF
C4502 VN.n4008 a_400_62400# 1.22fF
C4503 VN.n4009 a_400_62400# 0.07fF
C4504 VN.t2337 a_400_62400# 0.03fF
C4505 VN.n4010 a_400_62400# 0.16fF
C4506 VN.n4011 a_400_62400# 0.19fF
C4507 VN.n4013 a_400_62400# 2.51fF
C4508 VN.n4014 a_400_62400# 0.56fF
C4509 VN.n4015 a_400_62400# 0.64fF
C4510 VN.n4016 a_400_62400# 0.12fF
C4511 VN.n4017 a_400_62400# 0.44fF
C4512 VN.n4018 a_400_62400# 0.40fF
C4513 VN.n4019 a_400_62400# 1.03fF
C4514 VN.n4020 a_400_62400# 0.79fF
C4515 VN.t1236 a_400_62400# 0.03fF
C4516 VN.n4021 a_400_62400# 0.32fF
C4517 VN.n4022 a_400_62400# 0.48fF
C4518 VN.n4023 a_400_62400# 0.81fF
C4519 VN.n4024 a_400_62400# 0.16fF
C4520 VN.t29 a_400_62400# 0.03fF
C4521 VN.n4025 a_400_62400# 0.19fF
C4522 VN.n4027 a_400_62400# 3.50fF
C4523 VN.n4028 a_400_62400# 2.89fF
C4524 VN.t683 a_400_62400# 0.03fF
C4525 VN.n4029 a_400_62400# 0.32fF
C4526 VN.n4030 a_400_62400# 1.22fF
C4527 VN.n4031 a_400_62400# 0.07fF
C4528 VN.t290 a_400_62400# 0.03fF
C4529 VN.n4032 a_400_62400# 0.16fF
C4530 VN.n4033 a_400_62400# 0.19fF
C4531 VN.n4035 a_400_62400# 1.05fF
C4532 VN.n4036 a_400_62400# 3.07fF
C4533 VN.n4037 a_400_62400# 2.51fF
C4534 VN.n4038 a_400_62400# 0.16fF
C4535 VN.t1738 a_400_62400# 0.03fF
C4536 VN.n4039 a_400_62400# 0.19fF
C4537 VN.t372 a_400_62400# 0.03fF
C4538 VN.n4041 a_400_62400# 0.32fF
C4539 VN.n4042 a_400_62400# 0.48fF
C4540 VN.n4043 a_400_62400# 0.81fF
C4541 VN.n4044 a_400_62400# 1.86fF
C4542 VN.n4045 a_400_62400# 1.53fF
C4543 VN.n4046 a_400_62400# 0.47fF
C4544 VN.n4047 a_400_62400# 2.71fF
C4545 VN.t2343 a_400_62400# 0.03fF
C4546 VN.n4048 a_400_62400# 0.32fF
C4547 VN.n4049 a_400_62400# 1.22fF
C4548 VN.n4050 a_400_62400# 0.07fF
C4549 VN.t1942 a_400_62400# 0.03fF
C4550 VN.n4051 a_400_62400# 0.16fF
C4551 VN.n4052 a_400_62400# 0.19fF
C4552 VN.n4054 a_400_62400# 2.53fF
C4553 VN.n4055 a_400_62400# 2.51fF
C4554 VN.t2024 a_400_62400# 0.03fF
C4555 VN.n4056 a_400_62400# 0.32fF
C4556 VN.n4057 a_400_62400# 0.48fF
C4557 VN.n4058 a_400_62400# 0.81fF
C4558 VN.n4059 a_400_62400# 0.16fF
C4559 VN.t998 a_400_62400# 0.03fF
C4560 VN.n4060 a_400_62400# 0.19fF
C4561 VN.n4062 a_400_62400# 1.55fF
C4562 VN.n4063 a_400_62400# 0.29fF
C4563 VN.n4064 a_400_62400# 2.52fF
C4564 VN.t1475 a_400_62400# 0.03fF
C4565 VN.n4065 a_400_62400# 0.32fF
C4566 VN.n4066 a_400_62400# 1.22fF
C4567 VN.n4067 a_400_62400# 0.07fF
C4568 VN.t1071 a_400_62400# 0.03fF
C4569 VN.n4068 a_400_62400# 0.16fF
C4570 VN.n4069 a_400_62400# 0.19fF
C4571 VN.n4071 a_400_62400# 27.83fF
C4572 VN.n4072 a_400_62400# 3.93fF
C4573 VN.n4073 a_400_62400# 2.51fF
C4574 VN.n4074 a_400_62400# 0.16fF
C4575 VN.t117 a_400_62400# 0.03fF
C4576 VN.n4075 a_400_62400# 0.19fF
C4577 VN.t1291 a_400_62400# 0.03fF
C4578 VN.n4077 a_400_62400# 0.32fF
C4579 VN.n4078 a_400_62400# 0.48fF
C4580 VN.n4079 a_400_62400# 0.81fF
C4581 VN.n4080 a_400_62400# 1.46fF
C4582 VN.n4081 a_400_62400# 0.21fF
C4583 VN.n4082 a_400_62400# 2.81fF
C4584 VN.t197 a_400_62400# 0.03fF
C4585 VN.n4083 a_400_62400# 0.16fF
C4586 VN.n4084 a_400_62400# 0.19fF
C4587 VN.t730 a_400_62400# 0.03fF
C4588 VN.n4086 a_400_62400# 0.32fF
C4589 VN.n4087 a_400_62400# 1.22fF
C4590 VN.n4088 a_400_62400# 0.07fF
C4591 VN.n4089 a_400_62400# 2.51fF
C4592 VN.n4090 a_400_62400# 3.57fF
C4593 VN.t424 a_400_62400# 0.03fF
C4594 VN.n4091 a_400_62400# 0.32fF
C4595 VN.n4092 a_400_62400# 0.48fF
C4596 VN.n4093 a_400_62400# 0.81fF
C4597 VN.n4094 a_400_62400# 0.16fF
C4598 VN.t1785 a_400_62400# 0.03fF
C4599 VN.n4095 a_400_62400# 0.19fF
C4600 VN.n4097 a_400_62400# 3.93fF
C4601 VN.n4098 a_400_62400# 3.08fF
C4602 VN.t1854 a_400_62400# 0.03fF
C4603 VN.n4099 a_400_62400# 0.16fF
C4604 VN.n4100 a_400_62400# 0.19fF
C4605 VN.t2384 a_400_62400# 0.03fF
C4606 VN.n4102 a_400_62400# 0.32fF
C4607 VN.n4103 a_400_62400# 1.22fF
C4608 VN.n4104 a_400_62400# 0.07fF
C4609 VN.n4105 a_400_62400# 2.51fF
C4610 VN.n4106 a_400_62400# 3.57fF
C4611 VN.t2069 a_400_62400# 0.03fF
C4612 VN.n4107 a_400_62400# 0.32fF
C4613 VN.n4108 a_400_62400# 0.48fF
C4614 VN.n4109 a_400_62400# 0.81fF
C4615 VN.n4110 a_400_62400# 0.16fF
C4616 VN.t907 a_400_62400# 0.03fF
C4617 VN.n4111 a_400_62400# 0.19fF
C4618 VN.n4113 a_400_62400# 3.75fF
C4619 VN.n4114 a_400_62400# 3.08fF
C4620 VN.t985 a_400_62400# 0.03fF
C4621 VN.n4115 a_400_62400# 0.16fF
C4622 VN.n4116 a_400_62400# 0.19fF
C4623 VN.t1515 a_400_62400# 0.03fF
C4624 VN.n4118 a_400_62400# 0.32fF
C4625 VN.n4119 a_400_62400# 1.22fF
C4626 VN.n4120 a_400_62400# 0.07fF
C4627 VN.n4121 a_400_62400# 2.51fF
C4628 VN.n4122 a_400_62400# 3.57fF
C4629 VN.t1199 a_400_62400# 0.03fF
C4630 VN.n4123 a_400_62400# 0.32fF
C4631 VN.n4124 a_400_62400# 0.48fF
C4632 VN.n4125 a_400_62400# 0.81fF
C4633 VN.n4126 a_400_62400# 0.16fF
C4634 VN.t2570 a_400_62400# 0.03fF
C4635 VN.n4127 a_400_62400# 0.19fF
C4636 VN.n4129 a_400_62400# 3.75fF
C4637 VN.n4130 a_400_62400# 3.08fF
C4638 VN.t96 a_400_62400# 0.03fF
C4639 VN.n4131 a_400_62400# 0.16fF
C4640 VN.n4132 a_400_62400# 0.19fF
C4641 VN.t647 a_400_62400# 0.03fF
C4642 VN.n4134 a_400_62400# 0.32fF
C4643 VN.n4135 a_400_62400# 1.22fF
C4644 VN.n4136 a_400_62400# 0.07fF
C4645 VN.n4137 a_400_62400# 2.51fF
C4646 VN.n4138 a_400_62400# 3.57fF
C4647 VN.t331 a_400_62400# 0.03fF
C4648 VN.n4139 a_400_62400# 0.32fF
C4649 VN.n4140 a_400_62400# 0.48fF
C4650 VN.n4141 a_400_62400# 0.81fF
C4651 VN.n4142 a_400_62400# 0.16fF
C4652 VN.t1699 a_400_62400# 0.03fF
C4653 VN.n4143 a_400_62400# 0.19fF
C4654 VN.n4145 a_400_62400# 3.75fF
C4655 VN.n4146 a_400_62400# 3.08fF
C4656 VN.t1896 a_400_62400# 0.03fF
C4657 VN.n4147 a_400_62400# 0.16fF
C4658 VN.n4148 a_400_62400# 0.19fF
C4659 VN.t2306 a_400_62400# 0.03fF
C4660 VN.n4150 a_400_62400# 0.32fF
C4661 VN.n4151 a_400_62400# 1.22fF
C4662 VN.n4152 a_400_62400# 0.07fF
C4663 VN.n4153 a_400_62400# 2.51fF
C4664 VN.n4154 a_400_62400# 3.57fF
C4665 VN.t1977 a_400_62400# 0.03fF
C4666 VN.n4155 a_400_62400# 0.32fF
C4667 VN.n4156 a_400_62400# 0.48fF
C4668 VN.n4157 a_400_62400# 0.81fF
C4669 VN.n4158 a_400_62400# 0.16fF
C4670 VN.t829 a_400_62400# 0.03fF
C4671 VN.n4159 a_400_62400# 0.19fF
C4672 VN.n4161 a_400_62400# 3.75fF
C4673 VN.n4162 a_400_62400# 3.08fF
C4674 VN.t1021 a_400_62400# 0.03fF
C4675 VN.n4163 a_400_62400# 0.16fF
C4676 VN.n4164 a_400_62400# 0.19fF
C4677 VN.t1435 a_400_62400# 0.03fF
C4678 VN.n4166 a_400_62400# 0.32fF
C4679 VN.n4167 a_400_62400# 1.22fF
C4680 VN.n4168 a_400_62400# 0.07fF
C4681 VN.n4169 a_400_62400# 2.51fF
C4682 VN.n4170 a_400_62400# 3.57fF
C4683 VN.t1803 a_400_62400# 0.03fF
C4684 VN.n4171 a_400_62400# 0.32fF
C4685 VN.n4172 a_400_62400# 0.48fF
C4686 VN.n4173 a_400_62400# 0.81fF
C4687 VN.n4174 a_400_62400# 0.16fF
C4688 VN.t666 a_400_62400# 0.03fF
C4689 VN.n4175 a_400_62400# 0.19fF
C4690 VN.n4177 a_400_62400# 3.75fF
C4691 VN.n4178 a_400_62400# 3.08fF
C4692 VN.t843 a_400_62400# 0.03fF
C4693 VN.n4179 a_400_62400# 0.16fF
C4694 VN.n4180 a_400_62400# 0.19fF
C4695 VN.t221 a_400_62400# 0.03fF
C4696 VN.n4182 a_400_62400# 0.32fF
C4697 VN.n4183 a_400_62400# 1.22fF
C4698 VN.n4184 a_400_62400# 0.07fF
C4699 VN.n4185 a_400_62400# 2.51fF
C4700 VN.n4186 a_400_62400# 3.57fF
C4701 VN.t927 a_400_62400# 0.03fF
C4702 VN.n4187 a_400_62400# 0.32fF
C4703 VN.n4188 a_400_62400# 0.48fF
C4704 VN.n4189 a_400_62400# 0.81fF
C4705 VN.n4190 a_400_62400# 0.16fF
C4706 VN.t2324 a_400_62400# 0.03fF
C4707 VN.n4191 a_400_62400# 0.19fF
C4708 VN.n4193 a_400_62400# 3.75fF
C4709 VN.n4194 a_400_62400# 3.08fF
C4710 VN.t2507 a_400_62400# 0.03fF
C4711 VN.n4195 a_400_62400# 0.16fF
C4712 VN.n4196 a_400_62400# 0.19fF
C4713 VN.t1871 a_400_62400# 0.03fF
C4714 VN.n4198 a_400_62400# 0.32fF
C4715 VN.n4199 a_400_62400# 1.22fF
C4716 VN.n4200 a_400_62400# 0.07fF
C4717 VN.n4201 a_400_62400# 3.65fF
C4718 VN.n4202 a_400_62400# 2.14fF
C4719 VN.n4203 a_400_62400# 0.16fF
C4720 VN.t709 a_400_62400# 0.03fF
C4721 VN.n4204 a_400_62400# 0.19fF
C4722 VN.t1721 a_400_62400# 0.03fF
C4723 VN.n4206 a_400_62400# 0.32fF
C4724 VN.n4207 a_400_62400# 0.48fF
C4725 VN.n4208 a_400_62400# 0.81fF
C4726 VN.n4209 a_400_62400# 0.09fF
C4727 VN.n4210 a_400_62400# 0.01fF
C4728 VN.n4211 a_400_62400# 0.02fF
C4729 VN.n4212 a_400_62400# 0.02fF
C4730 VN.n4213 a_400_62400# 0.32fF
C4731 VN.n4214 a_400_62400# 1.56fF
C4732 VN.n4215 a_400_62400# 1.81fF
C4733 VN.n4216 a_400_62400# 3.08fF
C4734 VN.t773 a_400_62400# 0.03fF
C4735 VN.n4217 a_400_62400# 0.16fF
C4736 VN.n4218 a_400_62400# 0.19fF
C4737 VN.t123 a_400_62400# 0.03fF
C4738 VN.n4220 a_400_62400# 0.32fF
C4739 VN.n4221 a_400_62400# 1.22fF
C4740 VN.n4222 a_400_62400# 0.07fF
C4741 VN.t28 a_400_62400# 64.69fF
C4742 VN.t1001 a_400_62400# 0.03fF
C4743 VN.n4223 a_400_62400# 0.32fF
C4744 VN.n4224 a_400_62400# 1.22fF
C4745 VN.n4225 a_400_62400# 0.07fF
C4746 VN.t1644 a_400_62400# 0.03fF
C4747 VN.n4226 a_400_62400# 0.16fF
C4748 VN.n4227 a_400_62400# 0.19fF
C4749 VN.n4229 a_400_62400# 0.16fF
C4750 VN.t1458 a_400_62400# 0.03fF
C4751 VN.n4230 a_400_62400# 0.19fF
C4752 VN.n4232 a_400_62400# 6.92fF
C4753 VN.n4233 a_400_62400# 6.56fF
C4754 VN.t2411 a_400_62400# 0.03fF
C4755 VN.n4234 a_400_62400# 0.16fF
C4756 VN.n4235 a_400_62400# 0.19fF
C4757 VN.t270 a_400_62400# 0.03fF
C4758 VN.n4237 a_400_62400# 0.32fF
C4759 VN.n4238 a_400_62400# 1.22fF
C4760 VN.n4239 a_400_62400# 0.07fF
C4761 VN.n4240 a_400_62400# 2.51fF
C4762 VN.n4241 a_400_62400# 3.58fF
C4763 VN.t2023 a_400_62400# 0.03fF
C4764 VN.n4242 a_400_62400# 0.32fF
C4765 VN.n4243 a_400_62400# 0.48fF
C4766 VN.n4244 a_400_62400# 0.81fF
C4767 VN.n4245 a_400_62400# 0.16fF
C4768 VN.t855 a_400_62400# 0.03fF
C4769 VN.n4246 a_400_62400# 0.19fF
C4770 VN.n4248 a_400_62400# 7.29fF
C4771 VN.t1548 a_400_62400# 0.03fF
C4772 VN.n4249 a_400_62400# 0.16fF
C4773 VN.n4250 a_400_62400# 0.19fF
C4774 VN.t1920 a_400_62400# 0.03fF
C4775 VN.n4252 a_400_62400# 0.32fF
C4776 VN.n4253 a_400_62400# 1.22fF
C4777 VN.n4254 a_400_62400# 0.07fF
C4778 VN.t14 a_400_62400# 64.17fF
C4779 VN.t1045 a_400_62400# 0.03fF
C4780 VN.n4255 a_400_62400# 1.60fF
C4781 VN.n4256 a_400_62400# 0.07fF
C4782 VN.t800 a_400_62400# 0.03fF
C4783 VN.n4257 a_400_62400# 0.02fF
C4784 VN.n4258 a_400_62400# 0.34fF
C4785 VN.n4260 a_400_62400# 2.01fF
C4786 VN.n4261 a_400_62400# 1.75fF
C4787 VN.n4262 a_400_62400# 0.37fF
C4788 VN.n4263 a_400_62400# 0.33fF
C4789 VN.n4264 a_400_62400# 5.88fF
C4790 VN.n4265 a_400_62400# 0.02fF
C4791 VN.n4266 a_400_62400# 0.02fF
C4792 VN.n4267 a_400_62400# 0.03fF
C4793 VN.n4268 a_400_62400# 0.05fF
C4794 VN.n4269 a_400_62400# 0.23fF
C4795 VN.n4270 a_400_62400# 0.02fF
C4796 VN.n4271 a_400_62400# 0.03fF
C4797 VN.n4272 a_400_62400# 0.01fF
C4798 VN.n4273 a_400_62400# 0.01fF
C4799 VN.n4274 a_400_62400# 0.01fF
C4800 VN.n4275 a_400_62400# 0.02fF
C4801 VN.n4276 a_400_62400# 0.03fF
C4802 VN.n4277 a_400_62400# 0.06fF
C4803 VN.n4278 a_400_62400# 0.05fF
C4804 VN.n4279 a_400_62400# 0.15fF
C4805 VN.n4280 a_400_62400# 0.51fF
C4806 VN.n4281 a_400_62400# 0.27fF
C4807 VN.n4282 a_400_62400# 37.46fF
C4808 VN.n4283 a_400_62400# 37.46fF
C4809 VN.n4284 a_400_62400# 0.79fF
C4810 VN.n4285 a_400_62400# 0.23fF
C4811 VN.n4286 a_400_62400# 1.18fF
C4812 VN.t122 a_400_62400# 28.64fF
C4813 VN.n4287 a_400_62400# 0.79fF
C4814 VN.n4288 a_400_62400# 0.11fF
C4815 VN.n4289 a_400_62400# 4.98fF
C4816 VN.n4290 a_400_62400# 0.80fF
C4817 VN.n4291 a_400_62400# 0.29fF
C4818 VN.n4292 a_400_62400# 1.96fF
C4819 VN.n4294 a_400_62400# 25.18fF
C4820 VN.n4296 a_400_62400# 1.87fF
C4821 VN.n4297 a_400_62400# 5.36fF
C4822 VN.n4298 a_400_62400# 1.81fF
C4823 VN.t1989 a_400_62400# 0.03fF
C4824 VN.n4299 a_400_62400# 0.85fF
C4825 VN.n4300 a_400_62400# 0.81fF
C4826 VN.n4301 a_400_62400# 0.33fF
C4827 VN.n4302 a_400_62400# 0.12fF
C4828 VN.n4303 a_400_62400# 0.28fF
C4829 VN.n4304 a_400_62400# 1.23fF
C4830 VN.n4305 a_400_62400# 0.59fF
C4831 VN.n4306 a_400_62400# 2.51fF
C4832 VN.n4307 a_400_62400# 0.16fF
C4833 VN.t988 a_400_62400# 0.03fF
C4834 VN.n4308 a_400_62400# 0.19fF
C4835 VN.t2013 a_400_62400# 0.03fF
C4836 VN.n4310 a_400_62400# 0.32fF
C4837 VN.n4311 a_400_62400# 0.48fF
C4838 VN.n4312 a_400_62400# 0.81fF
C4839 VN.n4313 a_400_62400# 0.03fF
C4840 VN.n4314 a_400_62400# 0.01fF
C4841 VN.n4315 a_400_62400# 0.02fF
C4842 VN.n4316 a_400_62400# 0.11fF
C4843 VN.n4317 a_400_62400# 0.08fF
C4844 VN.n4318 a_400_62400# 0.04fF
C4845 VN.n4319 a_400_62400# 0.05fF
C4846 VN.n4320 a_400_62400# 1.34fF
C4847 VN.n4321 a_400_62400# 0.48fF
C4848 VN.n4322 a_400_62400# 2.51fF
C4849 VN.n4323 a_400_62400# 2.67fF
C4850 VN.t326 a_400_62400# 0.03fF
C4851 VN.n4324 a_400_62400# 0.32fF
C4852 VN.n4325 a_400_62400# 1.22fF
C4853 VN.n4326 a_400_62400# 0.07fF
C4854 VN.t1665 a_400_62400# 0.03fF
C4855 VN.n4327 a_400_62400# 0.16fF
C4856 VN.n4328 a_400_62400# 0.19fF
C4857 VN.n4330 a_400_62400# 2.53fF
C4858 VN.n4331 a_400_62400# 0.08fF
C4859 VN.n4332 a_400_62400# 0.04fF
C4860 VN.n4333 a_400_62400# 0.05fF
C4861 VN.n4334 a_400_62400# 1.33fF
C4862 VN.n4335 a_400_62400# 0.03fF
C4863 VN.n4336 a_400_62400# 0.01fF
C4864 VN.n4337 a_400_62400# 0.02fF
C4865 VN.n4338 a_400_62400# 0.11fF
C4866 VN.n4339 a_400_62400# 0.48fF
C4867 VN.n4340 a_400_62400# 2.48fF
C4868 VN.t1279 a_400_62400# 0.03fF
C4869 VN.n4341 a_400_62400# 0.32fF
C4870 VN.n4342 a_400_62400# 0.48fF
C4871 VN.n4343 a_400_62400# 0.81fF
C4872 VN.n4344 a_400_62400# 0.16fF
C4873 VN.t100 a_400_62400# 0.03fF
C4874 VN.n4345 a_400_62400# 0.19fF
C4875 VN.n4347 a_400_62400# 0.93fF
C4876 VN.n4348 a_400_62400# 0.30fF
C4877 VN.n4349 a_400_62400# 0.34fF
C4878 VN.n4350 a_400_62400# 0.12fF
C4879 VN.n4351 a_400_62400# 0.30fF
C4880 VN.n4352 a_400_62400# 0.93fF
C4881 VN.n4353 a_400_62400# 1.55fF
C4882 VN.n4354 a_400_62400# 0.29fF
C4883 VN.n4355 a_400_62400# 0.34fF
C4884 VN.n4356 a_400_62400# 0.12fF
C4885 VN.n4357 a_400_62400# 2.52fF
C4886 VN.t2115 a_400_62400# 0.03fF
C4887 VN.n4358 a_400_62400# 0.32fF
C4888 VN.n4359 a_400_62400# 1.22fF
C4889 VN.n4360 a_400_62400# 0.07fF
C4890 VN.t799 a_400_62400# 0.03fF
C4891 VN.n4361 a_400_62400# 0.16fF
C4892 VN.n4362 a_400_62400# 0.19fF
C4893 VN.n4364 a_400_62400# 0.33fF
C4894 VN.n4365 a_400_62400# 0.12fF
C4895 VN.n4366 a_400_62400# 0.28fF
C4896 VN.n4367 a_400_62400# 1.23fF
C4897 VN.n4368 a_400_62400# 0.59fF
C4898 VN.n4369 a_400_62400# 2.51fF
C4899 VN.n4370 a_400_62400# 0.16fF
C4900 VN.t1772 a_400_62400# 0.03fF
C4901 VN.n4371 a_400_62400# 0.19fF
C4902 VN.t412 a_400_62400# 0.03fF
C4903 VN.n4373 a_400_62400# 0.32fF
C4904 VN.n4374 a_400_62400# 0.48fF
C4905 VN.n4375 a_400_62400# 0.81fF
C4906 VN.n4376 a_400_62400# 0.03fF
C4907 VN.n4377 a_400_62400# 0.01fF
C4908 VN.n4378 a_400_62400# 0.02fF
C4909 VN.n4379 a_400_62400# 0.11fF
C4910 VN.n4380 a_400_62400# 0.08fF
C4911 VN.n4381 a_400_62400# 0.04fF
C4912 VN.n4382 a_400_62400# 0.05fF
C4913 VN.n4383 a_400_62400# 1.34fF
C4914 VN.n4384 a_400_62400# 0.48fF
C4915 VN.n4385 a_400_62400# 2.51fF
C4916 VN.n4386 a_400_62400# 2.67fF
C4917 VN.t1237 a_400_62400# 0.03fF
C4918 VN.n4387 a_400_62400# 0.32fF
C4919 VN.n4388 a_400_62400# 1.22fF
C4920 VN.n4389 a_400_62400# 0.07fF
C4921 VN.t2454 a_400_62400# 0.03fF
C4922 VN.n4390 a_400_62400# 0.16fF
C4923 VN.n4391 a_400_62400# 0.19fF
C4924 VN.n4393 a_400_62400# 2.53fF
C4925 VN.n4394 a_400_62400# 0.05fF
C4926 VN.n4395 a_400_62400# 0.09fF
C4927 VN.n4396 a_400_62400# 0.07fF
C4928 VN.n4397 a_400_62400# 1.16fF
C4929 VN.n4398 a_400_62400# 0.01fF
C4930 VN.n4399 a_400_62400# 0.01fF
C4931 VN.n4400 a_400_62400# 0.01fF
C4932 VN.n4401 a_400_62400# 0.09fF
C4933 VN.n4402 a_400_62400# 0.91fF
C4934 VN.n4403 a_400_62400# 0.96fF
C4935 VN.t862 a_400_62400# 0.03fF
C4936 VN.n4404 a_400_62400# 0.32fF
C4937 VN.n4405 a_400_62400# 0.48fF
C4938 VN.n4406 a_400_62400# 0.81fF
C4939 VN.n4407 a_400_62400# 0.16fF
C4940 VN.t2265 a_400_62400# 0.03fF
C4941 VN.n4408 a_400_62400# 0.19fF
C4942 VN.n4410 a_400_62400# 0.93fF
C4943 VN.n4411 a_400_62400# 0.30fF
C4944 VN.n4412 a_400_62400# 0.34fF
C4945 VN.n4413 a_400_62400# 0.12fF
C4946 VN.n4414 a_400_62400# 0.30fF
C4947 VN.n4415 a_400_62400# 0.93fF
C4948 VN.n4416 a_400_62400# 1.55fF
C4949 VN.n4417 a_400_62400# 0.29fF
C4950 VN.n4418 a_400_62400# 0.34fF
C4951 VN.n4419 a_400_62400# 0.12fF
C4952 VN.n4420 a_400_62400# 3.10fF
C4953 VN.t1701 a_400_62400# 0.03fF
C4954 VN.n4421 a_400_62400# 0.32fF
C4955 VN.n4422 a_400_62400# 1.22fF
C4956 VN.n4423 a_400_62400# 0.07fF
C4957 VN.t1590 a_400_62400# 0.03fF
C4958 VN.n4424 a_400_62400# 0.16fF
C4959 VN.n4425 a_400_62400# 0.19fF
C4960 VN.n4427 a_400_62400# 2.51fF
C4961 VN.n4428 a_400_62400# 0.61fF
C4962 VN.n4429 a_400_62400# 0.30fF
C4963 VN.n4430 a_400_62400# 0.51fF
C4964 VN.n4431 a_400_62400# 0.21fF
C4965 VN.n4432 a_400_62400# 0.38fF
C4966 VN.n4433 a_400_62400# 0.29fF
C4967 VN.n4434 a_400_62400# 0.40fF
C4968 VN.n4435 a_400_62400# 0.28fF
C4969 VN.t2524 a_400_62400# 0.03fF
C4970 VN.n4436 a_400_62400# 0.32fF
C4971 VN.n4437 a_400_62400# 0.48fF
C4972 VN.n4438 a_400_62400# 0.81fF
C4973 VN.n4439 a_400_62400# 0.16fF
C4974 VN.t1400 a_400_62400# 0.03fF
C4975 VN.n4440 a_400_62400# 0.19fF
C4976 VN.n4442 a_400_62400# 0.06fF
C4977 VN.n4443 a_400_62400# 0.04fF
C4978 VN.n4444 a_400_62400# 0.04fF
C4979 VN.n4445 a_400_62400# 0.14fF
C4980 VN.n4446 a_400_62400# 0.48fF
C4981 VN.n4447 a_400_62400# 0.50fF
C4982 VN.n4448 a_400_62400# 0.14fF
C4983 VN.n4449 a_400_62400# 0.16fF
C4984 VN.n4450 a_400_62400# 0.09fF
C4985 VN.n4451 a_400_62400# 0.16fF
C4986 VN.n4452 a_400_62400# 0.24fF
C4987 VN.n4453 a_400_62400# 5.35fF
C4988 VN.t830 a_400_62400# 0.03fF
C4989 VN.n4454 a_400_62400# 0.32fF
C4990 VN.n4455 a_400_62400# 1.22fF
C4991 VN.n4456 a_400_62400# 0.07fF
C4992 VN.t2078 a_400_62400# 0.03fF
C4993 VN.n4457 a_400_62400# 0.16fF
C4994 VN.n4458 a_400_62400# 0.19fF
C4995 VN.n4460 a_400_62400# 0.33fF
C4996 VN.n4461 a_400_62400# 0.12fF
C4997 VN.n4462 a_400_62400# 0.28fF
C4998 VN.n4463 a_400_62400# 1.72fF
C4999 VN.n4464 a_400_62400# 0.71fF
C5000 VN.n4465 a_400_62400# 2.51fF
C5001 VN.n4466 a_400_62400# 0.16fF
C5002 VN.t539 a_400_62400# 0.03fF
C5003 VN.n4467 a_400_62400# 0.19fF
C5004 VN.t1661 a_400_62400# 0.03fF
C5005 VN.n4469 a_400_62400# 0.32fF
C5006 VN.n4470 a_400_62400# 0.48fF
C5007 VN.n4471 a_400_62400# 0.81fF
C5008 VN.n4472 a_400_62400# 0.95fF
C5009 VN.n4473 a_400_62400# 2.11fF
C5010 VN.n4474 a_400_62400# 3.28fF
C5011 VN.t2493 a_400_62400# 0.03fF
C5012 VN.n4475 a_400_62400# 0.32fF
C5013 VN.n4476 a_400_62400# 1.22fF
C5014 VN.n4477 a_400_62400# 0.07fF
C5015 VN.t1206 a_400_62400# 0.03fF
C5016 VN.n4478 a_400_62400# 0.16fF
C5017 VN.n4479 a_400_62400# 0.19fF
C5018 VN.n4481 a_400_62400# 2.53fF
C5019 VN.n4482 a_400_62400# 0.08fF
C5020 VN.n4483 a_400_62400# 0.04fF
C5021 VN.n4484 a_400_62400# 0.05fF
C5022 VN.n4485 a_400_62400# 1.33fF
C5023 VN.n4486 a_400_62400# 0.03fF
C5024 VN.n4487 a_400_62400# 0.01fF
C5025 VN.n4488 a_400_62400# 0.02fF
C5026 VN.n4489 a_400_62400# 0.11fF
C5027 VN.n4490 a_400_62400# 0.48fF
C5028 VN.n4491 a_400_62400# 2.48fF
C5029 VN.t793 a_400_62400# 0.03fF
C5030 VN.n4492 a_400_62400# 0.32fF
C5031 VN.n4493 a_400_62400# 0.48fF
C5032 VN.n4494 a_400_62400# 0.81fF
C5033 VN.n4495 a_400_62400# 0.16fF
C5034 VN.t2195 a_400_62400# 0.03fF
C5035 VN.n4496 a_400_62400# 0.19fF
C5036 VN.n4498 a_400_62400# 0.93fF
C5037 VN.n4499 a_400_62400# 0.30fF
C5038 VN.n4500 a_400_62400# 0.34fF
C5039 VN.n4501 a_400_62400# 0.12fF
C5040 VN.n4502 a_400_62400# 0.30fF
C5041 VN.n4503 a_400_62400# 0.93fF
C5042 VN.n4504 a_400_62400# 1.55fF
C5043 VN.n4505 a_400_62400# 0.29fF
C5044 VN.n4506 a_400_62400# 0.34fF
C5045 VN.n4507 a_400_62400# 0.12fF
C5046 VN.n4508 a_400_62400# 2.52fF
C5047 VN.t1629 a_400_62400# 0.03fF
C5048 VN.n4509 a_400_62400# 0.32fF
C5049 VN.n4510 a_400_62400# 1.22fF
C5050 VN.n4511 a_400_62400# 0.07fF
C5051 VN.t477 a_400_62400# 0.03fF
C5052 VN.n4512 a_400_62400# 0.16fF
C5053 VN.n4513 a_400_62400# 0.19fF
C5054 VN.n4515 a_400_62400# 27.83fF
C5055 VN.n4516 a_400_62400# 2.30fF
C5056 VN.n4517 a_400_62400# 4.08fF
C5057 VN.t363 a_400_62400# 0.03fF
C5058 VN.n4518 a_400_62400# 0.32fF
C5059 VN.n4519 a_400_62400# 0.48fF
C5060 VN.n4520 a_400_62400# 0.81fF
C5061 VN.n4521 a_400_62400# 0.16fF
C5062 VN.t1730 a_400_62400# 0.03fF
C5063 VN.n4522 a_400_62400# 0.19fF
C5064 VN.n4524 a_400_62400# 0.42fF
C5065 VN.n4525 a_400_62400# 0.34fF
C5066 VN.n4526 a_400_62400# 0.12fF
C5067 VN.n4527 a_400_62400# 0.30fF
C5068 VN.n4528 a_400_62400# 0.88fF
C5069 VN.n4529 a_400_62400# 1.28fF
C5070 VN.n4530 a_400_62400# 0.30fF
C5071 VN.n4531 a_400_62400# 0.28fF
C5072 VN.n4532 a_400_62400# 0.27fF
C5073 VN.n4533 a_400_62400# 0.09fF
C5074 VN.n4534 a_400_62400# 0.12fF
C5075 VN.n4535 a_400_62400# 0.13fF
C5076 VN.n4536 a_400_62400# 2.66fF
C5077 VN.t2529 a_400_62400# 0.03fF
C5078 VN.n4537 a_400_62400# 0.16fF
C5079 VN.n4538 a_400_62400# 0.19fF
C5080 VN.t1195 a_400_62400# 0.03fF
C5081 VN.n4540 a_400_62400# 0.32fF
C5082 VN.n4541 a_400_62400# 1.22fF
C5083 VN.n4542 a_400_62400# 0.07fF
C5084 VN.n4543 a_400_62400# 2.51fF
C5085 VN.n4544 a_400_62400# 0.16fF
C5086 VN.t1325 a_400_62400# 0.03fF
C5087 VN.n4545 a_400_62400# 0.19fF
C5088 VN.t2448 a_400_62400# 0.03fF
C5089 VN.n4547 a_400_62400# 0.32fF
C5090 VN.n4548 a_400_62400# 0.48fF
C5091 VN.n4549 a_400_62400# 0.81fF
C5092 VN.n4550 a_400_62400# 1.24fF
C5093 VN.n4551 a_400_62400# 0.43fF
C5094 VN.n4552 a_400_62400# 0.43fF
C5095 VN.n4553 a_400_62400# 1.24fF
C5096 VN.n4554 a_400_62400# 1.46fF
C5097 VN.n4555 a_400_62400# 0.21fF
C5098 VN.n4556 a_400_62400# 6.64fF
C5099 VN.t2131 a_400_62400# 0.03fF
C5100 VN.n4557 a_400_62400# 0.16fF
C5101 VN.n4558 a_400_62400# 0.19fF
C5102 VN.t759 a_400_62400# 0.03fF
C5103 VN.n4560 a_400_62400# 0.32fF
C5104 VN.n4561 a_400_62400# 1.22fF
C5105 VN.n4562 a_400_62400# 0.07fF
C5106 VN.n4563 a_400_62400# 2.51fF
C5107 VN.n4564 a_400_62400# 3.57fF
C5108 VN.t1583 a_400_62400# 0.03fF
C5109 VN.n4565 a_400_62400# 0.32fF
C5110 VN.n4566 a_400_62400# 0.48fF
C5111 VN.n4567 a_400_62400# 0.81fF
C5112 VN.n4568 a_400_62400# 0.16fF
C5113 VN.t463 a_400_62400# 0.03fF
C5114 VN.n4569 a_400_62400# 0.19fF
C5115 VN.n4571 a_400_62400# 6.91fF
C5116 VN.t1255 a_400_62400# 0.03fF
C5117 VN.n4572 a_400_62400# 0.16fF
C5118 VN.n4573 a_400_62400# 0.19fF
C5119 VN.t2412 a_400_62400# 0.03fF
C5120 VN.n4575 a_400_62400# 0.32fF
C5121 VN.n4576 a_400_62400# 1.22fF
C5122 VN.n4577 a_400_62400# 0.07fF
C5123 VN.n4578 a_400_62400# 2.51fF
C5124 VN.n4579 a_400_62400# 3.57fF
C5125 VN.t719 a_400_62400# 0.03fF
C5126 VN.n4580 a_400_62400# 0.32fF
C5127 VN.n4581 a_400_62400# 0.48fF
C5128 VN.n4582 a_400_62400# 0.81fF
C5129 VN.n4583 a_400_62400# 0.16fF
C5130 VN.t2112 a_400_62400# 0.03fF
C5131 VN.n4584 a_400_62400# 0.19fF
C5132 VN.n4586 a_400_62400# 6.92fF
C5133 VN.t385 a_400_62400# 0.03fF
C5134 VN.n4587 a_400_62400# 0.16fF
C5135 VN.n4588 a_400_62400# 0.19fF
C5136 VN.t1551 a_400_62400# 0.03fF
C5137 VN.n4590 a_400_62400# 0.32fF
C5138 VN.n4591 a_400_62400# 1.22fF
C5139 VN.n4592 a_400_62400# 0.07fF
C5140 VN.n4593 a_400_62400# 2.51fF
C5141 VN.n4594 a_400_62400# 3.57fF
C5142 VN.t2373 a_400_62400# 0.03fF
C5143 VN.n4595 a_400_62400# 0.32fF
C5144 VN.n4596 a_400_62400# 0.48fF
C5145 VN.n4597 a_400_62400# 0.81fF
C5146 VN.n4598 a_400_62400# 0.16fF
C5147 VN.t1368 a_400_62400# 0.03fF
C5148 VN.n4599 a_400_62400# 0.19fF
C5149 VN.n4601 a_400_62400# 6.92fF
C5150 VN.t2039 a_400_62400# 0.03fF
C5151 VN.n4602 a_400_62400# 0.16fF
C5152 VN.n4603 a_400_62400# 0.19fF
C5153 VN.t678 a_400_62400# 0.03fF
C5154 VN.n4605 a_400_62400# 0.32fF
C5155 VN.n4606 a_400_62400# 1.22fF
C5156 VN.n4607 a_400_62400# 0.07fF
C5157 VN.n4608 a_400_62400# 2.51fF
C5158 VN.n4609 a_400_62400# 3.57fF
C5159 VN.t1626 a_400_62400# 0.03fF
C5160 VN.n4610 a_400_62400# 0.32fF
C5161 VN.n4611 a_400_62400# 0.48fF
C5162 VN.n4612 a_400_62400# 0.81fF
C5163 VN.n4613 a_400_62400# 0.16fF
C5164 VN.t501 a_400_62400# 0.03fF
C5165 VN.n4614 a_400_62400# 0.19fF
C5166 VN.n4616 a_400_62400# 6.92fF
C5167 VN.t1167 a_400_62400# 0.03fF
C5168 VN.n4617 a_400_62400# 0.16fF
C5169 VN.n4618 a_400_62400# 0.19fF
C5170 VN.t2457 a_400_62400# 0.03fF
C5171 VN.n4620 a_400_62400# 0.32fF
C5172 VN.n4621 a_400_62400# 1.22fF
C5173 VN.n4622 a_400_62400# 0.07fF
C5174 VN.n4623 a_400_62400# 2.51fF
C5175 VN.n4624 a_400_62400# 3.57fF
C5176 VN.t438 a_400_62400# 0.03fF
C5177 VN.n4625 a_400_62400# 0.32fF
C5178 VN.n4626 a_400_62400# 0.48fF
C5179 VN.n4627 a_400_62400# 0.81fF
C5180 VN.n4628 a_400_62400# 0.16fF
C5181 VN.t1787 a_400_62400# 0.03fF
C5182 VN.n4629 a_400_62400# 0.19fF
C5183 VN.n4631 a_400_62400# 6.92fF
C5184 VN.t296 a_400_62400# 0.03fF
C5185 VN.n4632 a_400_62400# 0.16fF
C5186 VN.n4633 a_400_62400# 0.19fF
C5187 VN.t329 a_400_62400# 0.03fF
C5188 VN.n4635 a_400_62400# 0.32fF
C5189 VN.n4636 a_400_62400# 1.22fF
C5190 VN.n4637 a_400_62400# 0.07fF
C5191 VN.n4638 a_400_62400# 2.51fF
C5192 VN.n4639 a_400_62400# 3.57fF
C5193 VN.t2083 a_400_62400# 0.03fF
C5194 VN.n4640 a_400_62400# 0.32fF
C5195 VN.n4641 a_400_62400# 0.48fF
C5196 VN.n4642 a_400_62400# 0.81fF
C5197 VN.n4643 a_400_62400# 0.16fF
C5198 VN.t912 a_400_62400# 0.03fF
C5199 VN.n4644 a_400_62400# 0.19fF
C5200 VN.n4646 a_400_62400# 6.92fF
C5201 VN.t1600 a_400_62400# 0.03fF
C5202 VN.n4647 a_400_62400# 0.16fF
C5203 VN.n4648 a_400_62400# 0.19fF
C5204 VN.t1975 a_400_62400# 0.03fF
C5205 VN.n4650 a_400_62400# 0.32fF
C5206 VN.n4651 a_400_62400# 1.22fF
C5207 VN.n4652 a_400_62400# 0.07fF
C5208 VN.n4653 a_400_62400# 2.51fF
C5209 VN.n4654 a_400_62400# 3.57fF
C5210 VN.t1209 a_400_62400# 0.03fF
C5211 VN.n4655 a_400_62400# 0.32fF
C5212 VN.n4656 a_400_62400# 0.48fF
C5213 VN.n4657 a_400_62400# 0.81fF
C5214 VN.n4658 a_400_62400# 0.16fF
C5215 VN.t2574 a_400_62400# 0.03fF
C5216 VN.n4659 a_400_62400# 0.19fF
C5217 VN.n4661 a_400_62400# 2.51fF
C5218 VN.n4662 a_400_62400# 3.59fF
C5219 VN.t901 a_400_62400# 0.03fF
C5220 VN.n4663 a_400_62400# 0.32fF
C5221 VN.n4664 a_400_62400# 0.48fF
C5222 VN.n4665 a_400_62400# 0.81fF
C5223 VN.t1987 a_400_62400# 0.03fF
C5224 VN.n4666 a_400_62400# 1.63fF
C5225 VN.n4667 a_400_62400# 0.49fF
C5226 VN.n4668 a_400_62400# 1.64fF
C5227 VN.n4669 a_400_62400# 0.81fF
C5228 VN.n4670 a_400_62400# 1.21fF
C5229 VN.n4671 a_400_62400# 1.54fF
C5230 VN.n4672 a_400_62400# 4.06fF
C5231 VN.t103 a_400_62400# 28.64fF
C5232 VN.n4673 a_400_62400# 28.43fF
C5233 VN.n4675 a_400_62400# 0.50fF
C5234 VN.n4676 a_400_62400# 0.31fF
C5235 VN.n4677 a_400_62400# 3.74fF
C5236 VN.n4678 a_400_62400# 3.29fF
C5237 VN.n4679 a_400_62400# 5.35fF
C5238 VN.n4680 a_400_62400# 0.34fF
C5239 VN.n4681 a_400_62400# 0.02fF
C5240 VN.t838 a_400_62400# 0.03fF
C5241 VN.n4682 a_400_62400# 0.34fF
C5242 VN.t1446 a_400_62400# 0.03fF
C5243 VN.n4683 a_400_62400# 1.28fF
C5244 VN.n4684 a_400_62400# 0.94fF
C5245 VN.n4685 a_400_62400# 2.53fF
C5246 VN.n4686 a_400_62400# 2.51fF
C5247 VN.t1114 a_400_62400# 0.03fF
C5248 VN.n4687 a_400_62400# 0.32fF
C5249 VN.n4688 a_400_62400# 0.48fF
C5250 VN.n4689 a_400_62400# 0.81fF
C5251 VN.n4690 a_400_62400# 0.16fF
C5252 VN.t2501 a_400_62400# 0.03fF
C5253 VN.n4691 a_400_62400# 0.19fF
C5254 VN.n4693 a_400_62400# 1.55fF
C5255 VN.n4694 a_400_62400# 0.29fF
C5256 VN.n4695 a_400_62400# 2.52fF
C5257 VN.t578 a_400_62400# 0.03fF
C5258 VN.n4696 a_400_62400# 0.32fF
C5259 VN.n4697 a_400_62400# 1.22fF
C5260 VN.n4698 a_400_62400# 0.07fF
C5261 VN.t2565 a_400_62400# 0.03fF
C5262 VN.n4699 a_400_62400# 0.16fF
C5263 VN.n4700 a_400_62400# 0.19fF
C5264 VN.n4702 a_400_62400# 1.04fF
C5265 VN.n4703 a_400_62400# 2.60fF
C5266 VN.n4704 a_400_62400# 2.51fF
C5267 VN.n4705 a_400_62400# 0.16fF
C5268 VN.t1638 a_400_62400# 0.03fF
C5269 VN.n4706 a_400_62400# 0.19fF
C5270 VN.t250 a_400_62400# 0.03fF
C5271 VN.n4708 a_400_62400# 0.32fF
C5272 VN.n4709 a_400_62400# 0.48fF
C5273 VN.n4710 a_400_62400# 0.81fF
C5274 VN.n4711 a_400_62400# 2.46fF
C5275 VN.n4712 a_400_62400# 4.01fF
C5276 VN.t2236 a_400_62400# 0.03fF
C5277 VN.n4713 a_400_62400# 0.32fF
C5278 VN.n4714 a_400_62400# 1.22fF
C5279 VN.n4715 a_400_62400# 0.07fF
C5280 VN.t1826 a_400_62400# 0.03fF
C5281 VN.n4716 a_400_62400# 0.16fF
C5282 VN.n4717 a_400_62400# 0.19fF
C5283 VN.n4719 a_400_62400# 2.53fF
C5284 VN.n4720 a_400_62400# 2.51fF
C5285 VN.t1900 a_400_62400# 0.03fF
C5286 VN.n4721 a_400_62400# 0.32fF
C5287 VN.n4722 a_400_62400# 0.48fF
C5288 VN.n4723 a_400_62400# 0.81fF
C5289 VN.n4724 a_400_62400# 0.16fF
C5290 VN.t767 a_400_62400# 0.03fF
C5291 VN.n4725 a_400_62400# 0.19fF
C5292 VN.n4727 a_400_62400# 1.55fF
C5293 VN.n4728 a_400_62400# 0.29fF
C5294 VN.n4729 a_400_62400# 2.52fF
C5295 VN.t1371 a_400_62400# 0.03fF
C5296 VN.n4730 a_400_62400# 0.32fF
C5297 VN.n4731 a_400_62400# 1.22fF
C5298 VN.n4732 a_400_62400# 0.07fF
C5299 VN.t950 a_400_62400# 0.03fF
C5300 VN.n4733 a_400_62400# 0.16fF
C5301 VN.n4734 a_400_62400# 0.19fF
C5302 VN.n4736 a_400_62400# 1.04fF
C5303 VN.n4737 a_400_62400# 2.60fF
C5304 VN.n4738 a_400_62400# 2.51fF
C5305 VN.n4739 a_400_62400# 0.16fF
C5306 VN.t2421 a_400_62400# 0.03fF
C5307 VN.n4740 a_400_62400# 0.19fF
C5308 VN.t1025 a_400_62400# 0.03fF
C5309 VN.n4742 a_400_62400# 0.32fF
C5310 VN.n4743 a_400_62400# 0.48fF
C5311 VN.n4744 a_400_62400# 0.81fF
C5312 VN.n4745 a_400_62400# 2.46fF
C5313 VN.n4746 a_400_62400# 4.01fF
C5314 VN.t506 a_400_62400# 0.03fF
C5315 VN.n4747 a_400_62400# 0.32fF
C5316 VN.n4748 a_400_62400# 1.22fF
C5317 VN.n4749 a_400_62400# 0.07fF
C5318 VN.t33 a_400_62400# 0.03fF
C5319 VN.n4750 a_400_62400# 0.16fF
C5320 VN.n4751 a_400_62400# 0.19fF
C5321 VN.n4753 a_400_62400# 2.53fF
C5322 VN.n4754 a_400_62400# 2.34fF
C5323 VN.t1520 a_400_62400# 0.03fF
C5324 VN.n4755 a_400_62400# 0.32fF
C5325 VN.n4756 a_400_62400# 0.48fF
C5326 VN.n4757 a_400_62400# 0.81fF
C5327 VN.n4758 a_400_62400# 0.16fF
C5328 VN.t391 a_400_62400# 0.03fF
C5329 VN.n4759 a_400_62400# 0.19fF
C5330 VN.n4761 a_400_62400# 1.55fF
C5331 VN.n4762 a_400_62400# 0.29fF
C5332 VN.n4763 a_400_62400# 3.27fF
C5333 VN.t957 a_400_62400# 0.03fF
C5334 VN.n4764 a_400_62400# 0.32fF
C5335 VN.n4765 a_400_62400# 1.22fF
C5336 VN.n4766 a_400_62400# 0.07fF
C5337 VN.t581 a_400_62400# 0.03fF
C5338 VN.n4767 a_400_62400# 0.16fF
C5339 VN.n4768 a_400_62400# 0.19fF
C5340 VN.n4770 a_400_62400# 2.51fF
C5341 VN.n4771 a_400_62400# 0.56fF
C5342 VN.n4772 a_400_62400# 0.64fF
C5343 VN.n4773 a_400_62400# 0.12fF
C5344 VN.n4774 a_400_62400# 0.44fF
C5345 VN.n4775 a_400_62400# 0.40fF
C5346 VN.n4776 a_400_62400# 1.03fF
C5347 VN.n4777 a_400_62400# 0.79fF
C5348 VN.t652 a_400_62400# 0.03fF
C5349 VN.n4778 a_400_62400# 0.32fF
C5350 VN.n4779 a_400_62400# 0.48fF
C5351 VN.n4780 a_400_62400# 0.81fF
C5352 VN.n4781 a_400_62400# 0.16fF
C5353 VN.t2044 a_400_62400# 0.03fF
C5354 VN.n4782 a_400_62400# 0.19fF
C5355 VN.n4784 a_400_62400# 3.50fF
C5356 VN.n4785 a_400_62400# 2.89fF
C5357 VN.t48 a_400_62400# 0.03fF
C5358 VN.n4786 a_400_62400# 0.32fF
C5359 VN.n4787 a_400_62400# 1.22fF
C5360 VN.n4788 a_400_62400# 0.07fF
C5361 VN.t2238 a_400_62400# 0.03fF
C5362 VN.n4789 a_400_62400# 0.16fF
C5363 VN.n4790 a_400_62400# 0.19fF
C5364 VN.n4792 a_400_62400# 1.05fF
C5365 VN.n4793 a_400_62400# 3.07fF
C5366 VN.n4794 a_400_62400# 2.51fF
C5367 VN.n4795 a_400_62400# 0.16fF
C5368 VN.t1308 a_400_62400# 0.03fF
C5369 VN.n4796 a_400_62400# 0.19fF
C5370 VN.t2311 a_400_62400# 0.03fF
C5371 VN.n4798 a_400_62400# 0.32fF
C5372 VN.n4799 a_400_62400# 0.48fF
C5373 VN.n4800 a_400_62400# 0.81fF
C5374 VN.n4801 a_400_62400# 1.86fF
C5375 VN.n4802 a_400_62400# 1.53fF
C5376 VN.n4803 a_400_62400# 0.47fF
C5377 VN.n4804 a_400_62400# 2.71fF
C5378 VN.t1745 a_400_62400# 0.03fF
C5379 VN.n4805 a_400_62400# 0.32fF
C5380 VN.n4806 a_400_62400# 1.22fF
C5381 VN.n4807 a_400_62400# 0.07fF
C5382 VN.t1373 a_400_62400# 0.03fF
C5383 VN.n4808 a_400_62400# 0.16fF
C5384 VN.n4809 a_400_62400# 0.19fF
C5385 VN.n4811 a_400_62400# 2.53fF
C5386 VN.n4812 a_400_62400# 2.51fF
C5387 VN.t1564 a_400_62400# 0.03fF
C5388 VN.n4813 a_400_62400# 0.32fF
C5389 VN.n4814 a_400_62400# 0.48fF
C5390 VN.n4815 a_400_62400# 0.81fF
C5391 VN.n4816 a_400_62400# 0.16fF
C5392 VN.t447 a_400_62400# 0.03fF
C5393 VN.n4817 a_400_62400# 0.19fF
C5394 VN.n4819 a_400_62400# 1.55fF
C5395 VN.n4820 a_400_62400# 0.29fF
C5396 VN.n4821 a_400_62400# 2.52fF
C5397 VN.t1003 a_400_62400# 0.03fF
C5398 VN.n4822 a_400_62400# 0.32fF
C5399 VN.n4823 a_400_62400# 1.22fF
C5400 VN.n4824 a_400_62400# 0.07fF
C5401 VN.t510 a_400_62400# 0.03fF
C5402 VN.n4825 a_400_62400# 0.16fF
C5403 VN.n4826 a_400_62400# 0.19fF
C5404 VN.n4828 a_400_62400# 27.83fF
C5405 VN.n4829 a_400_62400# 3.93fF
C5406 VN.n4830 a_400_62400# 2.51fF
C5407 VN.n4831 a_400_62400# 0.16fF
C5408 VN.t2093 a_400_62400# 0.03fF
C5409 VN.n4832 a_400_62400# 0.19fF
C5410 VN.t694 a_400_62400# 0.03fF
C5411 VN.n4834 a_400_62400# 0.32fF
C5412 VN.n4835 a_400_62400# 0.48fF
C5413 VN.n4836 a_400_62400# 0.81fF
C5414 VN.n4837 a_400_62400# 1.46fF
C5415 VN.n4838 a_400_62400# 0.21fF
C5416 VN.n4839 a_400_62400# 2.81fF
C5417 VN.t2162 a_400_62400# 0.03fF
C5418 VN.n4840 a_400_62400# 0.16fF
C5419 VN.n4841 a_400_62400# 0.19fF
C5420 VN.t127 a_400_62400# 0.03fF
C5421 VN.n4843 a_400_62400# 0.32fF
C5422 VN.n4844 a_400_62400# 1.22fF
C5423 VN.n4845 a_400_62400# 0.07fF
C5424 VN.n4846 a_400_62400# 2.51fF
C5425 VN.n4847 a_400_62400# 3.57fF
C5426 VN.t2353 a_400_62400# 0.03fF
C5427 VN.n4848 a_400_62400# 0.32fF
C5428 VN.n4849 a_400_62400# 0.48fF
C5429 VN.n4850 a_400_62400# 0.81fF
C5430 VN.n4851 a_400_62400# 0.16fF
C5431 VN.t1216 a_400_62400# 0.03fF
C5432 VN.n4852 a_400_62400# 0.19fF
C5433 VN.n4854 a_400_62400# 3.93fF
C5434 VN.n4855 a_400_62400# 3.08fF
C5435 VN.t1294 a_400_62400# 0.03fF
C5436 VN.n4856 a_400_62400# 0.16fF
C5437 VN.n4857 a_400_62400# 0.19fF
C5438 VN.t1791 a_400_62400# 0.03fF
C5439 VN.n4859 a_400_62400# 0.32fF
C5440 VN.n4860 a_400_62400# 1.22fF
C5441 VN.n4861 a_400_62400# 0.07fF
C5442 VN.n4862 a_400_62400# 2.51fF
C5443 VN.n4863 a_400_62400# 3.57fF
C5444 VN.t1485 a_400_62400# 0.03fF
C5445 VN.n4864 a_400_62400# 0.32fF
C5446 VN.n4865 a_400_62400# 0.48fF
C5447 VN.n4866 a_400_62400# 0.81fF
C5448 VN.n4867 a_400_62400# 0.16fF
C5449 VN.t354 a_400_62400# 0.03fF
C5450 VN.n4868 a_400_62400# 0.19fF
C5451 VN.n4870 a_400_62400# 3.75fF
C5452 VN.n4871 a_400_62400# 3.08fF
C5453 VN.t429 a_400_62400# 0.03fF
C5454 VN.n4872 a_400_62400# 0.16fF
C5455 VN.n4873 a_400_62400# 0.19fF
C5456 VN.t916 a_400_62400# 0.03fF
C5457 VN.n4875 a_400_62400# 0.32fF
C5458 VN.n4876 a_400_62400# 1.22fF
C5459 VN.n4877 a_400_62400# 0.07fF
C5460 VN.n4878 a_400_62400# 2.51fF
C5461 VN.n4879 a_400_62400# 3.57fF
C5462 VN.t618 a_400_62400# 0.03fF
C5463 VN.n4880 a_400_62400# 0.32fF
C5464 VN.n4881 a_400_62400# 0.48fF
C5465 VN.n4882 a_400_62400# 0.81fF
C5466 VN.n4883 a_400_62400# 0.16fF
C5467 VN.t1999 a_400_62400# 0.03fF
C5468 VN.n4884 a_400_62400# 0.19fF
C5469 VN.n4886 a_400_62400# 3.75fF
C5470 VN.n4887 a_400_62400# 3.08fF
C5471 VN.t2203 a_400_62400# 0.03fF
C5472 VN.n4888 a_400_62400# 0.16fF
C5473 VN.n4889 a_400_62400# 0.19fF
C5474 VN.t2579 a_400_62400# 0.03fF
C5475 VN.n4891 a_400_62400# 0.32fF
C5476 VN.n4892 a_400_62400# 1.22fF
C5477 VN.n4893 a_400_62400# 0.07fF
C5478 VN.n4894 a_400_62400# 2.51fF
C5479 VN.n4895 a_400_62400# 3.57fF
C5480 VN.t2270 a_400_62400# 0.03fF
C5481 VN.n4896 a_400_62400# 0.32fF
C5482 VN.n4897 a_400_62400# 0.48fF
C5483 VN.n4898 a_400_62400# 0.81fF
C5484 VN.n4899 a_400_62400# 0.16fF
C5485 VN.t1125 a_400_62400# 0.03fF
C5486 VN.n4900 a_400_62400# 0.19fF
C5487 VN.n4902 a_400_62400# 3.75fF
C5488 VN.n4903 a_400_62400# 3.08fF
C5489 VN.t1335 a_400_62400# 0.03fF
C5490 VN.n4904 a_400_62400# 0.16fF
C5491 VN.n4905 a_400_62400# 0.19fF
C5492 VN.t1709 a_400_62400# 0.03fF
C5493 VN.n4907 a_400_62400# 0.32fF
C5494 VN.n4908 a_400_62400# 1.22fF
C5495 VN.n4909 a_400_62400# 0.07fF
C5496 VN.n4910 a_400_62400# 2.51fF
C5497 VN.n4911 a_400_62400# 3.57fF
C5498 VN.t104 a_400_62400# 0.03fF
C5499 VN.n4912 a_400_62400# 0.32fF
C5500 VN.n4913 a_400_62400# 0.48fF
C5501 VN.n4914 a_400_62400# 0.81fF
C5502 VN.n4915 a_400_62400# 0.16fF
C5503 VN.t1507 a_400_62400# 0.03fF
C5504 VN.n4916 a_400_62400# 0.19fF
C5505 VN.n4918 a_400_62400# 3.75fF
C5506 VN.n4919 a_400_62400# 3.08fF
C5507 VN.t1689 a_400_62400# 0.03fF
C5508 VN.n4920 a_400_62400# 0.16fF
C5509 VN.n4921 a_400_62400# 0.19fF
C5510 VN.t1060 a_400_62400# 0.03fF
C5511 VN.n4923 a_400_62400# 0.32fF
C5512 VN.n4924 a_400_62400# 1.22fF
C5513 VN.n4925 a_400_62400# 0.07fF
C5514 VN.n4926 a_400_62400# 2.51fF
C5515 VN.n4927 a_400_62400# 3.57fF
C5516 VN.t1775 a_400_62400# 0.03fF
C5517 VN.n4928 a_400_62400# 0.32fF
C5518 VN.n4929 a_400_62400# 0.48fF
C5519 VN.n4930 a_400_62400# 0.81fF
C5520 VN.n4931 a_400_62400# 0.16fF
C5521 VN.t640 a_400_62400# 0.03fF
C5522 VN.n4932 a_400_62400# 0.19fF
C5523 VN.n4934 a_400_62400# 3.75fF
C5524 VN.n4935 a_400_62400# 3.08fF
C5525 VN.t821 a_400_62400# 0.03fF
C5526 VN.n4936 a_400_62400# 0.16fF
C5527 VN.n4937 a_400_62400# 0.19fF
C5528 VN.t186 a_400_62400# 0.03fF
C5529 VN.n4939 a_400_62400# 0.32fF
C5530 VN.n4940 a_400_62400# 1.22fF
C5531 VN.n4941 a_400_62400# 0.07fF
C5532 VN.n4942 a_400_62400# 3.65fF
C5533 VN.n4943 a_400_62400# 2.14fF
C5534 VN.n4944 a_400_62400# 0.16fF
C5535 VN.t1550 a_400_62400# 0.03fF
C5536 VN.n4945 a_400_62400# 0.19fF
C5537 VN.t2563 a_400_62400# 0.03fF
C5538 VN.n4947 a_400_62400# 0.32fF
C5539 VN.n4948 a_400_62400# 0.48fF
C5540 VN.n4949 a_400_62400# 0.81fF
C5541 VN.n4950 a_400_62400# 0.09fF
C5542 VN.n4951 a_400_62400# 0.01fF
C5543 VN.n4952 a_400_62400# 0.02fF
C5544 VN.n4953 a_400_62400# 0.02fF
C5545 VN.n4954 a_400_62400# 0.32fF
C5546 VN.n4955 a_400_62400# 1.56fF
C5547 VN.n4956 a_400_62400# 1.81fF
C5548 VN.n4957 a_400_62400# 3.08fF
C5549 VN.t1618 a_400_62400# 0.03fF
C5550 VN.n4958 a_400_62400# 0.16fF
C5551 VN.n4959 a_400_62400# 0.19fF
C5552 VN.t971 a_400_62400# 0.03fF
C5553 VN.n4961 a_400_62400# 0.32fF
C5554 VN.n4962 a_400_62400# 1.22fF
C5555 VN.n4963 a_400_62400# 0.07fF
C5556 VN.t32 a_400_62400# 64.69fF
C5557 VN.t1843 a_400_62400# 0.03fF
C5558 VN.n4964 a_400_62400# 0.32fF
C5559 VN.n4965 a_400_62400# 1.22fF
C5560 VN.n4966 a_400_62400# 0.07fF
C5561 VN.t2481 a_400_62400# 0.03fF
C5562 VN.n4967 a_400_62400# 0.16fF
C5563 VN.n4968 a_400_62400# 0.19fF
C5564 VN.n4970 a_400_62400# 0.16fF
C5565 VN.t2299 a_400_62400# 0.03fF
C5566 VN.n4971 a_400_62400# 0.19fF
C5567 VN.n4973 a_400_62400# 6.92fF
C5568 VN.n4974 a_400_62400# 6.56fF
C5569 VN.t734 a_400_62400# 0.03fF
C5570 VN.n4975 a_400_62400# 0.16fF
C5571 VN.n4976 a_400_62400# 0.19fF
C5572 VN.t1108 a_400_62400# 0.03fF
C5573 VN.n4978 a_400_62400# 0.32fF
C5574 VN.n4979 a_400_62400# 1.22fF
C5575 VN.n4980 a_400_62400# 0.07fF
C5576 VN.n4981 a_400_62400# 2.51fF
C5577 VN.n4982 a_400_62400# 3.58fF
C5578 VN.t346 a_400_62400# 0.03fF
C5579 VN.n4983 a_400_62400# 0.32fF
C5580 VN.n4984 a_400_62400# 0.48fF
C5581 VN.n4985 a_400_62400# 0.81fF
C5582 VN.n4986 a_400_62400# 0.16fF
C5583 VN.t1702 a_400_62400# 0.03fF
C5584 VN.n4987 a_400_62400# 0.19fF
C5585 VN.n4989 a_400_62400# 7.29fF
C5586 VN.t2389 a_400_62400# 0.03fF
C5587 VN.n4990 a_400_62400# 0.16fF
C5588 VN.n4991 a_400_62400# 0.19fF
C5589 VN.t240 a_400_62400# 0.03fF
C5590 VN.n4993 a_400_62400# 0.32fF
C5591 VN.n4994 a_400_62400# 1.22fF
C5592 VN.n4995 a_400_62400# 0.07fF
C5593 VN.t99 a_400_62400# 64.17fF
C5594 VN.t1889 a_400_62400# 0.03fF
C5595 VN.n4996 a_400_62400# 1.60fF
C5596 VN.n4997 a_400_62400# 0.07fF
C5597 VN.t1649 a_400_62400# 0.03fF
C5598 VN.n4998 a_400_62400# 0.02fF
C5599 VN.n4999 a_400_62400# 0.34fF
C5600 VN.n5001 a_400_62400# 2.01fF
C5601 VN.n5002 a_400_62400# 1.75fF
C5602 VN.n5003 a_400_62400# 0.37fF
C5603 VN.n5004 a_400_62400# 0.33fF
C5604 VN.n5005 a_400_62400# 5.88fF
C5605 VN.n5006 a_400_62400# 0.02fF
C5606 VN.n5007 a_400_62400# 0.02fF
C5607 VN.n5008 a_400_62400# 0.03fF
C5608 VN.n5009 a_400_62400# 0.05fF
C5609 VN.n5010 a_400_62400# 0.23fF
C5610 VN.n5011 a_400_62400# 0.02fF
C5611 VN.n5012 a_400_62400# 0.03fF
C5612 VN.n5013 a_400_62400# 0.01fF
C5613 VN.n5014 a_400_62400# 0.01fF
C5614 VN.n5015 a_400_62400# 0.01fF
C5615 VN.n5016 a_400_62400# 0.02fF
C5616 VN.n5017 a_400_62400# 0.03fF
C5617 VN.n5018 a_400_62400# 0.06fF
C5618 VN.n5019 a_400_62400# 0.05fF
C5619 VN.n5020 a_400_62400# 0.15fF
C5620 VN.n5021 a_400_62400# 0.51fF
C5621 VN.n5022 a_400_62400# 0.27fF
C5622 VN.n5023 a_400_62400# 37.46fF
C5623 VN.n5024 a_400_62400# 37.46fF
C5624 VN.n5025 a_400_62400# 0.79fF
C5625 VN.n5026 a_400_62400# 0.23fF
C5626 VN.n5027 a_400_62400# 1.18fF
C5627 VN.t47 a_400_62400# 28.64fF
C5628 VN.n5028 a_400_62400# 0.79fF
C5629 VN.n5029 a_400_62400# 0.11fF
C5630 VN.n5030 a_400_62400# 4.98fF
C5631 VN.n5031 a_400_62400# 0.80fF
C5632 VN.n5032 a_400_62400# 0.29fF
C5633 VN.n5033 a_400_62400# 1.96fF
C5634 VN.n5035 a_400_62400# 25.18fF
C5635 VN.n5037 a_400_62400# 1.87fF
C5636 VN.n5038 a_400_62400# 5.36fF
C5637 VN.n5039 a_400_62400# 1.81fF
C5638 VN.t314 a_400_62400# 0.03fF
C5639 VN.n5040 a_400_62400# 0.85fF
C5640 VN.n5041 a_400_62400# 0.81fF
C5641 VN.n5042 a_400_62400# 2.53fF
C5642 VN.n5043 a_400_62400# 0.08fF
C5643 VN.n5044 a_400_62400# 0.04fF
C5644 VN.n5045 a_400_62400# 0.05fF
C5645 VN.n5046 a_400_62400# 1.33fF
C5646 VN.n5047 a_400_62400# 0.03fF
C5647 VN.n5048 a_400_62400# 0.01fF
C5648 VN.n5049 a_400_62400# 0.02fF
C5649 VN.n5050 a_400_62400# 0.11fF
C5650 VN.n5051 a_400_62400# 0.48fF
C5651 VN.n5052 a_400_62400# 2.48fF
C5652 VN.t2302 a_400_62400# 0.03fF
C5653 VN.n5053 a_400_62400# 0.32fF
C5654 VN.n5054 a_400_62400# 0.48fF
C5655 VN.n5055 a_400_62400# 0.81fF
C5656 VN.n5056 a_400_62400# 0.16fF
C5657 VN.t1298 a_400_62400# 0.03fF
C5658 VN.n5057 a_400_62400# 0.19fF
C5659 VN.n5059 a_400_62400# 0.93fF
C5660 VN.n5060 a_400_62400# 0.30fF
C5661 VN.n5061 a_400_62400# 0.34fF
C5662 VN.n5062 a_400_62400# 0.12fF
C5663 VN.n5063 a_400_62400# 0.30fF
C5664 VN.n5064 a_400_62400# 0.93fF
C5665 VN.n5065 a_400_62400# 1.55fF
C5666 VN.n5066 a_400_62400# 0.29fF
C5667 VN.n5067 a_400_62400# 0.34fF
C5668 VN.n5068 a_400_62400# 0.12fF
C5669 VN.n5069 a_400_62400# 2.52fF
C5670 VN.t612 a_400_62400# 0.03fF
C5671 VN.n5070 a_400_62400# 0.32fF
C5672 VN.n5071 a_400_62400# 1.22fF
C5673 VN.n5072 a_400_62400# 0.07fF
C5674 VN.t1957 a_400_62400# 0.03fF
C5675 VN.n5073 a_400_62400# 0.16fF
C5676 VN.n5074 a_400_62400# 0.19fF
C5677 VN.n5076 a_400_62400# 0.33fF
C5678 VN.n5077 a_400_62400# 0.12fF
C5679 VN.n5078 a_400_62400# 0.28fF
C5680 VN.n5079 a_400_62400# 1.23fF
C5681 VN.n5080 a_400_62400# 0.59fF
C5682 VN.n5081 a_400_62400# 2.51fF
C5683 VN.n5082 a_400_62400# 0.16fF
C5684 VN.t432 a_400_62400# 0.03fF
C5685 VN.n5083 a_400_62400# 0.19fF
C5686 VN.t1555 a_400_62400# 0.03fF
C5687 VN.n5085 a_400_62400# 0.32fF
C5688 VN.n5086 a_400_62400# 0.48fF
C5689 VN.n5087 a_400_62400# 0.81fF
C5690 VN.n5088 a_400_62400# 0.03fF
C5691 VN.n5089 a_400_62400# 0.01fF
C5692 VN.n5090 a_400_62400# 0.02fF
C5693 VN.n5091 a_400_62400# 0.11fF
C5694 VN.n5092 a_400_62400# 0.08fF
C5695 VN.n5093 a_400_62400# 0.04fF
C5696 VN.n5094 a_400_62400# 0.05fF
C5697 VN.n5095 a_400_62400# 1.34fF
C5698 VN.n5096 a_400_62400# 0.48fF
C5699 VN.n5097 a_400_62400# 2.51fF
C5700 VN.n5098 a_400_62400# 2.67fF
C5701 VN.t2391 a_400_62400# 0.03fF
C5702 VN.n5099 a_400_62400# 0.32fF
C5703 VN.n5100 a_400_62400# 1.22fF
C5704 VN.n5101 a_400_62400# 0.07fF
C5705 VN.t1090 a_400_62400# 0.03fF
C5706 VN.n5102 a_400_62400# 0.16fF
C5707 VN.n5103 a_400_62400# 0.19fF
C5708 VN.n5105 a_400_62400# 2.53fF
C5709 VN.n5106 a_400_62400# 0.08fF
C5710 VN.n5107 a_400_62400# 0.04fF
C5711 VN.n5108 a_400_62400# 0.05fF
C5712 VN.n5109 a_400_62400# 1.33fF
C5713 VN.n5110 a_400_62400# 0.03fF
C5714 VN.n5111 a_400_62400# 0.01fF
C5715 VN.n5112 a_400_62400# 0.02fF
C5716 VN.n5113 a_400_62400# 0.11fF
C5717 VN.n5114 a_400_62400# 0.48fF
C5718 VN.n5115 a_400_62400# 2.48fF
C5719 VN.t684 a_400_62400# 0.03fF
C5720 VN.n5116 a_400_62400# 0.32fF
C5721 VN.n5117 a_400_62400# 0.48fF
C5722 VN.n5118 a_400_62400# 0.81fF
C5723 VN.n5119 a_400_62400# 0.16fF
C5724 VN.t2079 a_400_62400# 0.03fF
C5725 VN.n5120 a_400_62400# 0.19fF
C5726 VN.n5122 a_400_62400# 0.93fF
C5727 VN.n5123 a_400_62400# 0.30fF
C5728 VN.n5124 a_400_62400# 0.34fF
C5729 VN.n5125 a_400_62400# 0.12fF
C5730 VN.n5126 a_400_62400# 0.30fF
C5731 VN.n5127 a_400_62400# 0.93fF
C5732 VN.n5128 a_400_62400# 1.55fF
C5733 VN.n5129 a_400_62400# 0.29fF
C5734 VN.n5130 a_400_62400# 0.34fF
C5735 VN.n5131 a_400_62400# 0.12fF
C5736 VN.n5132 a_400_62400# 2.52fF
C5737 VN.t1522 a_400_62400# 0.03fF
C5738 VN.n5133 a_400_62400# 0.32fF
C5739 VN.n5134 a_400_62400# 1.22fF
C5740 VN.n5135 a_400_62400# 0.07fF
C5741 VN.t217 a_400_62400# 0.03fF
C5742 VN.n5136 a_400_62400# 0.16fF
C5743 VN.n5137 a_400_62400# 0.19fF
C5744 VN.n5139 a_400_62400# 0.33fF
C5745 VN.n5140 a_400_62400# 0.12fF
C5746 VN.n5141 a_400_62400# 0.28fF
C5747 VN.n5142 a_400_62400# 1.23fF
C5748 VN.n5143 a_400_62400# 0.59fF
C5749 VN.n5144 a_400_62400# 2.51fF
C5750 VN.n5145 a_400_62400# 0.16fF
C5751 VN.t2540 a_400_62400# 0.03fF
C5752 VN.n5146 a_400_62400# 0.19fF
C5753 VN.t1170 a_400_62400# 0.03fF
C5754 VN.n5148 a_400_62400# 0.32fF
C5755 VN.n5149 a_400_62400# 0.48fF
C5756 VN.n5150 a_400_62400# 0.81fF
C5757 VN.n5151 a_400_62400# 0.03fF
C5758 VN.n5152 a_400_62400# 0.01fF
C5759 VN.n5153 a_400_62400# 0.02fF
C5760 VN.n5154 a_400_62400# 0.11fF
C5761 VN.n5155 a_400_62400# 0.08fF
C5762 VN.n5156 a_400_62400# 0.04fF
C5763 VN.n5157 a_400_62400# 0.05fF
C5764 VN.n5158 a_400_62400# 1.34fF
C5765 VN.n5159 a_400_62400# 0.48fF
C5766 VN.n5160 a_400_62400# 2.51fF
C5767 VN.n5161 a_400_62400# 2.67fF
C5768 VN.t2001 a_400_62400# 0.03fF
C5769 VN.n5162 a_400_62400# 0.32fF
C5770 VN.n5163 a_400_62400# 1.22fF
C5771 VN.n5164 a_400_62400# 0.07fF
C5772 VN.t1868 a_400_62400# 0.03fF
C5773 VN.n5165 a_400_62400# 0.16fF
C5774 VN.n5166 a_400_62400# 0.19fF
C5775 VN.n5168 a_400_62400# 2.53fF
C5776 VN.n5169 a_400_62400# 0.09fF
C5777 VN.n5170 a_400_62400# 0.05fF
C5778 VN.n5171 a_400_62400# 0.07fF
C5779 VN.n5172 a_400_62400# 1.16fF
C5780 VN.n5173 a_400_62400# 0.01fF
C5781 VN.n5174 a_400_62400# 0.01fF
C5782 VN.n5175 a_400_62400# 0.01fF
C5783 VN.n5176 a_400_62400# 0.09fF
C5784 VN.n5177 a_400_62400# 0.91fF
C5785 VN.n5178 a_400_62400# 0.96fF
C5786 VN.t301 a_400_62400# 0.03fF
C5787 VN.n5179 a_400_62400# 0.32fF
C5788 VN.n5180 a_400_62400# 0.48fF
C5789 VN.n5181 a_400_62400# 0.81fF
C5790 VN.n5182 a_400_62400# 0.16fF
C5791 VN.t1675 a_400_62400# 0.03fF
C5792 VN.n5183 a_400_62400# 0.19fF
C5793 VN.n5185 a_400_62400# 0.93fF
C5794 VN.n5186 a_400_62400# 0.30fF
C5795 VN.n5187 a_400_62400# 0.34fF
C5796 VN.n5188 a_400_62400# 0.12fF
C5797 VN.n5189 a_400_62400# 0.30fF
C5798 VN.n5190 a_400_62400# 0.93fF
C5799 VN.n5191 a_400_62400# 1.55fF
C5800 VN.n5192 a_400_62400# 0.29fF
C5801 VN.n5193 a_400_62400# 0.34fF
C5802 VN.n5194 a_400_62400# 0.12fF
C5803 VN.n5195 a_400_62400# 3.10fF
C5804 VN.t1126 a_400_62400# 0.03fF
C5805 VN.n5196 a_400_62400# 0.32fF
C5806 VN.n5197 a_400_62400# 1.22fF
C5807 VN.n5198 a_400_62400# 0.07fF
C5808 VN.t2359 a_400_62400# 0.03fF
C5809 VN.n5199 a_400_62400# 0.16fF
C5810 VN.n5200 a_400_62400# 0.19fF
C5811 VN.n5202 a_400_62400# 2.51fF
C5812 VN.n5203 a_400_62400# 0.61fF
C5813 VN.n5204 a_400_62400# 0.30fF
C5814 VN.n5205 a_400_62400# 0.51fF
C5815 VN.n5206 a_400_62400# 0.21fF
C5816 VN.n5207 a_400_62400# 0.38fF
C5817 VN.n5208 a_400_62400# 0.29fF
C5818 VN.n5209 a_400_62400# 0.40fF
C5819 VN.n5210 a_400_62400# 0.28fF
C5820 VN.t1949 a_400_62400# 0.03fF
C5821 VN.n5211 a_400_62400# 0.32fF
C5822 VN.n5212 a_400_62400# 0.48fF
C5823 VN.n5213 a_400_62400# 0.81fF
C5824 VN.n5214 a_400_62400# 0.16fF
C5825 VN.t809 a_400_62400# 0.03fF
C5826 VN.n5215 a_400_62400# 0.19fF
C5827 VN.n5217 a_400_62400# 0.06fF
C5828 VN.n5218 a_400_62400# 0.04fF
C5829 VN.n5219 a_400_62400# 0.04fF
C5830 VN.n5220 a_400_62400# 0.14fF
C5831 VN.n5221 a_400_62400# 0.48fF
C5832 VN.n5222 a_400_62400# 0.50fF
C5833 VN.n5223 a_400_62400# 0.14fF
C5834 VN.n5224 a_400_62400# 0.16fF
C5835 VN.n5225 a_400_62400# 0.09fF
C5836 VN.n5226 a_400_62400# 0.16fF
C5837 VN.n5227 a_400_62400# 0.24fF
C5838 VN.n5228 a_400_62400# 5.35fF
C5839 VN.t262 a_400_62400# 0.03fF
C5840 VN.n5229 a_400_62400# 0.32fF
C5841 VN.n5230 a_400_62400# 1.22fF
C5842 VN.n5231 a_400_62400# 0.07fF
C5843 VN.t1492 a_400_62400# 0.03fF
C5844 VN.n5232 a_400_62400# 0.16fF
C5845 VN.n5233 a_400_62400# 0.19fF
C5846 VN.n5235 a_400_62400# 0.33fF
C5847 VN.n5236 a_400_62400# 0.12fF
C5848 VN.n5237 a_400_62400# 0.28fF
C5849 VN.n5238 a_400_62400# 1.72fF
C5850 VN.n5239 a_400_62400# 0.71fF
C5851 VN.n5240 a_400_62400# 2.51fF
C5852 VN.n5241 a_400_62400# 0.16fF
C5853 VN.t2464 a_400_62400# 0.03fF
C5854 VN.n5242 a_400_62400# 0.19fF
C5855 VN.t1080 a_400_62400# 0.03fF
C5856 VN.n5244 a_400_62400# 0.32fF
C5857 VN.n5245 a_400_62400# 0.48fF
C5858 VN.n5246 a_400_62400# 0.81fF
C5859 VN.n5247 a_400_62400# 0.95fF
C5860 VN.n5248 a_400_62400# 2.11fF
C5861 VN.n5249 a_400_62400# 3.28fF
C5862 VN.t1912 a_400_62400# 0.03fF
C5863 VN.n5250 a_400_62400# 0.32fF
C5864 VN.n5251 a_400_62400# 1.22fF
C5865 VN.n5252 a_400_62400# 0.07fF
C5866 VN.t746 a_400_62400# 0.03fF
C5867 VN.n5253 a_400_62400# 0.16fF
C5868 VN.n5254 a_400_62400# 0.19fF
C5869 VN.n5256 a_400_62400# 2.53fF
C5870 VN.n5257 a_400_62400# 0.08fF
C5871 VN.n5258 a_400_62400# 0.04fF
C5872 VN.n5259 a_400_62400# 0.05fF
C5873 VN.n5260 a_400_62400# 1.33fF
C5874 VN.n5261 a_400_62400# 0.03fF
C5875 VN.n5262 a_400_62400# 0.01fF
C5876 VN.n5263 a_400_62400# 0.02fF
C5877 VN.n5264 a_400_62400# 0.11fF
C5878 VN.n5265 a_400_62400# 0.48fF
C5879 VN.n5266 a_400_62400# 2.48fF
C5880 VN.t206 a_400_62400# 0.03fF
C5881 VN.n5267 a_400_62400# 0.32fF
C5882 VN.n5268 a_400_62400# 0.48fF
C5883 VN.n5269 a_400_62400# 0.81fF
C5884 VN.n5270 a_400_62400# 0.16fF
C5885 VN.t1598 a_400_62400# 0.03fF
C5886 VN.n5271 a_400_62400# 0.19fF
C5887 VN.n5273 a_400_62400# 0.93fF
C5888 VN.n5274 a_400_62400# 0.30fF
C5889 VN.n5275 a_400_62400# 0.34fF
C5890 VN.n5276 a_400_62400# 0.12fF
C5891 VN.n5277 a_400_62400# 0.30fF
C5892 VN.n5278 a_400_62400# 0.93fF
C5893 VN.n5279 a_400_62400# 1.55fF
C5894 VN.n5280 a_400_62400# 0.29fF
C5895 VN.n5281 a_400_62400# 0.34fF
C5896 VN.n5282 a_400_62400# 0.12fF
C5897 VN.n5283 a_400_62400# 2.52fF
C5898 VN.t1037 a_400_62400# 0.03fF
C5899 VN.n5284 a_400_62400# 0.32fF
C5900 VN.n5285 a_400_62400# 1.22fF
C5901 VN.n5286 a_400_62400# 0.07fF
C5902 VN.t2405 a_400_62400# 0.03fF
C5903 VN.n5287 a_400_62400# 0.16fF
C5904 VN.n5288 a_400_62400# 0.19fF
C5905 VN.n5290 a_400_62400# 27.83fF
C5906 VN.n5291 a_400_62400# 0.09fF
C5907 VN.n5292 a_400_62400# 0.27fF
C5908 VN.n5293 a_400_62400# 0.12fF
C5909 VN.n5294 a_400_62400# 0.28fF
C5910 VN.n5295 a_400_62400# 0.13fF
C5911 VN.n5296 a_400_62400# 0.40fF
C5912 VN.n5297 a_400_62400# 0.93fF
C5913 VN.n5298 a_400_62400# 0.60fF
C5914 VN.n5299 a_400_62400# 3.12fF
C5915 VN.n5300 a_400_62400# 0.16fF
C5916 VN.t2031 a_400_62400# 0.03fF
C5917 VN.n5301 a_400_62400# 0.19fF
C5918 VN.t643 a_400_62400# 0.03fF
C5919 VN.n5303 a_400_62400# 0.32fF
C5920 VN.n5304 a_400_62400# 0.48fF
C5921 VN.n5305 a_400_62400# 0.81fF
C5922 VN.n5306 a_400_62400# 2.54fF
C5923 VN.n5307 a_400_62400# 0.23fF
C5924 VN.n5308 a_400_62400# 1.02fF
C5925 VN.n5309 a_400_62400# 0.34fF
C5926 VN.n5310 a_400_62400# 0.40fF
C5927 VN.n5311 a_400_62400# 0.42fF
C5928 VN.n5312 a_400_62400# 0.63fF
C5929 VN.n5313 a_400_62400# 0.21fF
C5930 VN.n5314 a_400_62400# 2.58fF
C5931 VN.t307 a_400_62400# 0.03fF
C5932 VN.n5315 a_400_62400# 0.16fF
C5933 VN.n5316 a_400_62400# 0.19fF
C5934 VN.t1480 a_400_62400# 0.03fF
C5935 VN.n5318 a_400_62400# 0.32fF
C5936 VN.n5319 a_400_62400# 1.22fF
C5937 VN.n5320 a_400_62400# 0.07fF
C5938 VN.n5321 a_400_62400# 2.51fF
C5939 VN.n5322 a_400_62400# 0.16fF
C5940 VN.t733 a_400_62400# 0.03fF
C5941 VN.n5323 a_400_62400# 0.19fF
C5942 VN.t1859 a_400_62400# 0.03fF
C5943 VN.n5325 a_400_62400# 0.32fF
C5944 VN.n5326 a_400_62400# 0.48fF
C5945 VN.n5327 a_400_62400# 0.81fF
C5946 VN.n5328 a_400_62400# 1.24fF
C5947 VN.n5329 a_400_62400# 0.43fF
C5948 VN.n5330 a_400_62400# 0.43fF
C5949 VN.n5331 a_400_62400# 1.24fF
C5950 VN.n5332 a_400_62400# 1.46fF
C5951 VN.n5333 a_400_62400# 0.21fF
C5952 VN.n5334 a_400_62400# 6.64fF
C5953 VN.t1538 a_400_62400# 0.03fF
C5954 VN.n5335 a_400_62400# 0.16fF
C5955 VN.n5336 a_400_62400# 0.19fF
C5956 VN.t165 a_400_62400# 0.03fF
C5957 VN.n5338 a_400_62400# 0.32fF
C5958 VN.n5339 a_400_62400# 1.22fF
C5959 VN.n5340 a_400_62400# 0.07fF
C5960 VN.n5341 a_400_62400# 2.51fF
C5961 VN.n5342 a_400_62400# 3.57fF
C5962 VN.t990 a_400_62400# 0.03fF
C5963 VN.n5343 a_400_62400# 0.32fF
C5964 VN.n5344 a_400_62400# 0.48fF
C5965 VN.n5345 a_400_62400# 0.81fF
C5966 VN.n5346 a_400_62400# 0.16fF
C5967 VN.t2386 a_400_62400# 0.03fF
C5968 VN.n5347 a_400_62400# 0.19fF
C5969 VN.n5349 a_400_62400# 6.91fF
C5970 VN.t667 a_400_62400# 0.03fF
C5971 VN.n5350 a_400_62400# 0.16fF
C5972 VN.n5351 a_400_62400# 0.19fF
C5973 VN.t1828 a_400_62400# 0.03fF
C5974 VN.n5353 a_400_62400# 0.32fF
C5975 VN.n5354 a_400_62400# 1.22fF
C5976 VN.n5355 a_400_62400# 0.07fF
C5977 VN.n5356 a_400_62400# 2.51fF
C5978 VN.n5357 a_400_62400# 3.57fF
C5979 VN.t105 a_400_62400# 0.03fF
C5980 VN.n5358 a_400_62400# 0.32fF
C5981 VN.n5359 a_400_62400# 0.48fF
C5982 VN.n5360 a_400_62400# 0.81fF
C5983 VN.n5361 a_400_62400# 0.16fF
C5984 VN.t1645 a_400_62400# 0.03fF
C5985 VN.n5362 a_400_62400# 0.19fF
C5986 VN.n5364 a_400_62400# 6.92fF
C5987 VN.t2327 a_400_62400# 0.03fF
C5988 VN.n5365 a_400_62400# 0.16fF
C5989 VN.n5366 a_400_62400# 0.19fF
C5990 VN.t951 a_400_62400# 0.03fF
C5991 VN.n5368 a_400_62400# 0.32fF
C5992 VN.n5369 a_400_62400# 1.22fF
C5993 VN.n5370 a_400_62400# 0.07fF
C5994 VN.n5371 a_400_62400# 2.51fF
C5995 VN.n5372 a_400_62400# 3.57fF
C5996 VN.t1905 a_400_62400# 0.03fF
C5997 VN.n5373 a_400_62400# 0.32fF
C5998 VN.n5374 a_400_62400# 0.48fF
C5999 VN.n5375 a_400_62400# 0.81fF
C6000 VN.n5376 a_400_62400# 0.16fF
C6001 VN.t774 a_400_62400# 0.03fF
C6002 VN.n5377 a_400_62400# 0.19fF
C6003 VN.n5379 a_400_62400# 6.92fF
C6004 VN.t1462 a_400_62400# 0.03fF
C6005 VN.n5380 a_400_62400# 0.16fF
C6006 VN.n5381 a_400_62400# 0.19fF
C6007 VN.t220 a_400_62400# 0.03fF
C6008 VN.n5383 a_400_62400# 0.32fF
C6009 VN.n5384 a_400_62400# 1.22fF
C6010 VN.n5385 a_400_62400# 0.07fF
C6011 VN.n5386 a_400_62400# 2.51fF
C6012 VN.n5387 a_400_62400# 3.57fF
C6013 VN.t1274 a_400_62400# 0.03fF
C6014 VN.n5388 a_400_62400# 0.32fF
C6015 VN.n5389 a_400_62400# 0.48fF
C6016 VN.n5390 a_400_62400# 0.81fF
C6017 VN.n5391 a_400_62400# 0.16fF
C6018 VN.t72 a_400_62400# 0.03fF
C6019 VN.n5392 a_400_62400# 0.19fF
C6020 VN.n5394 a_400_62400# 6.92fF
C6021 VN.t589 a_400_62400# 0.03fF
C6022 VN.n5395 a_400_62400# 0.16fF
C6023 VN.n5396 a_400_62400# 0.19fF
C6024 VN.t1173 a_400_62400# 0.03fF
C6025 VN.n5398 a_400_62400# 0.32fF
C6026 VN.n5399 a_400_62400# 1.22fF
C6027 VN.n5400 a_400_62400# 0.07fF
C6028 VN.n5401 a_400_62400# 2.51fF
C6029 VN.n5402 a_400_62400# 3.57fF
C6030 VN.t404 a_400_62400# 0.03fF
C6031 VN.n5403 a_400_62400# 0.32fF
C6032 VN.n5404 a_400_62400# 0.48fF
C6033 VN.n5405 a_400_62400# 0.81fF
C6034 VN.n5406 a_400_62400# 0.16fF
C6035 VN.t1759 a_400_62400# 0.03fF
C6036 VN.n5407 a_400_62400# 0.19fF
C6037 VN.n5409 a_400_62400# 6.92fF
C6038 VN.t2441 a_400_62400# 0.03fF
C6039 VN.n5410 a_400_62400# 0.16fF
C6040 VN.n5411 a_400_62400# 0.19fF
C6041 VN.t305 a_400_62400# 0.03fF
C6042 VN.n5413 a_400_62400# 0.32fF
C6043 VN.n5414 a_400_62400# 1.22fF
C6044 VN.n5415 a_400_62400# 0.07fF
C6045 VN.n5416 a_400_62400# 2.51fF
C6046 VN.n5417 a_400_62400# 3.57fF
C6047 VN.t2054 a_400_62400# 0.03fF
C6048 VN.n5418 a_400_62400# 0.32fF
C6049 VN.n5419 a_400_62400# 0.48fF
C6050 VN.n5420 a_400_62400# 0.81fF
C6051 VN.n5421 a_400_62400# 0.16fF
C6052 VN.t886 a_400_62400# 0.03fF
C6053 VN.n5422 a_400_62400# 0.19fF
C6054 VN.n5424 a_400_62400# 2.51fF
C6055 VN.n5425 a_400_62400# 3.59fF
C6056 VN.t1748 a_400_62400# 0.03fF
C6057 VN.n5426 a_400_62400# 0.32fF
C6058 VN.n5427 a_400_62400# 0.48fF
C6059 VN.n5428 a_400_62400# 0.81fF
C6060 VN.t2279 a_400_62400# 0.03fF
C6061 VN.n5429 a_400_62400# 1.63fF
C6062 VN.n5430 a_400_62400# 0.81fF
C6063 VN.n5431 a_400_62400# 1.21fF
C6064 VN.n5432 a_400_62400# 1.54fF
C6065 VN.n5433 a_400_62400# 4.06fF
C6066 VN.t55 a_400_62400# 28.64fF
C6067 VN.n5434 a_400_62400# 28.43fF
C6068 VN.n5436 a_400_62400# 0.50fF
C6069 VN.n5437 a_400_62400# 0.31fF
C6070 VN.n5438 a_400_62400# 3.88fF
C6071 VN.n5439 a_400_62400# 3.29fF
C6072 VN.n5440 a_400_62400# 2.62fF
C6073 VN.n5441 a_400_62400# 5.27fF
C6074 VN.n5442 a_400_62400# 0.34fF
C6075 VN.n5443 a_400_62400# 0.02fF
C6076 VN.t1134 a_400_62400# 0.03fF
C6077 VN.n5444 a_400_62400# 0.34fF
C6078 VN.t1719 a_400_62400# 0.03fF
C6079 VN.n5445 a_400_62400# 1.28fF
C6080 VN.n5446 a_400_62400# 0.94fF
C6081 VN.n5447 a_400_62400# 1.04fF
C6082 VN.n5448 a_400_62400# 2.58fF
C6083 VN.n5449 a_400_62400# 2.51fF
C6084 VN.n5450 a_400_62400# 0.16fF
C6085 VN.t271 a_400_62400# 0.03fF
C6086 VN.n5451 a_400_62400# 0.19fF
C6087 VN.t1411 a_400_62400# 0.03fF
C6088 VN.n5453 a_400_62400# 0.32fF
C6089 VN.n5454 a_400_62400# 0.48fF
C6090 VN.n5455 a_400_62400# 0.81fF
C6091 VN.n5456 a_400_62400# 2.03fF
C6092 VN.n5457 a_400_62400# 4.01fF
C6093 VN.t846 a_400_62400# 0.03fF
C6094 VN.n5458 a_400_62400# 0.32fF
C6095 VN.n5459 a_400_62400# 1.22fF
C6096 VN.n5460 a_400_62400# 0.07fF
C6097 VN.t344 a_400_62400# 0.03fF
C6098 VN.n5461 a_400_62400# 0.16fF
C6099 VN.n5462 a_400_62400# 0.19fF
C6100 VN.n5464 a_400_62400# 2.53fF
C6101 VN.n5465 a_400_62400# 2.51fF
C6102 VN.t551 a_400_62400# 0.03fF
C6103 VN.n5466 a_400_62400# 0.32fF
C6104 VN.n5467 a_400_62400# 0.48fF
C6105 VN.n5468 a_400_62400# 0.81fF
C6106 VN.n5469 a_400_62400# 0.16fF
C6107 VN.t1921 a_400_62400# 0.03fF
C6108 VN.n5470 a_400_62400# 0.19fF
C6109 VN.n5472 a_400_62400# 1.55fF
C6110 VN.n5473 a_400_62400# 0.29fF
C6111 VN.n5474 a_400_62400# 2.52fF
C6112 VN.t2510 a_400_62400# 0.03fF
C6113 VN.n5475 a_400_62400# 0.32fF
C6114 VN.n5476 a_400_62400# 1.22fF
C6115 VN.n5477 a_400_62400# 0.07fF
C6116 VN.t2136 a_400_62400# 0.03fF
C6117 VN.n5478 a_400_62400# 0.16fF
C6118 VN.n5479 a_400_62400# 0.19fF
C6119 VN.n5481 a_400_62400# 1.04fF
C6120 VN.n5482 a_400_62400# 2.60fF
C6121 VN.n5483 a_400_62400# 2.51fF
C6122 VN.n5484 a_400_62400# 0.16fF
C6123 VN.t1046 a_400_62400# 0.03fF
C6124 VN.n5485 a_400_62400# 0.19fF
C6125 VN.t2206 a_400_62400# 0.03fF
C6126 VN.n5487 a_400_62400# 0.32fF
C6127 VN.n5488 a_400_62400# 0.48fF
C6128 VN.n5489 a_400_62400# 0.81fF
C6129 VN.n5490 a_400_62400# 2.46fF
C6130 VN.n5491 a_400_62400# 4.01fF
C6131 VN.t1647 a_400_62400# 0.03fF
C6132 VN.n5492 a_400_62400# 0.32fF
C6133 VN.n5493 a_400_62400# 1.22fF
C6134 VN.n5494 a_400_62400# 0.07fF
C6135 VN.t1262 a_400_62400# 0.03fF
C6136 VN.n5495 a_400_62400# 0.16fF
C6137 VN.n5496 a_400_62400# 0.19fF
C6138 VN.n5498 a_400_62400# 2.53fF
C6139 VN.n5499 a_400_62400# 2.51fF
C6140 VN.t1339 a_400_62400# 0.03fF
C6141 VN.n5500 a_400_62400# 0.32fF
C6142 VN.n5501 a_400_62400# 0.48fF
C6143 VN.n5502 a_400_62400# 0.81fF
C6144 VN.n5503 a_400_62400# 0.16fF
C6145 VN.t177 a_400_62400# 0.03fF
C6146 VN.n5504 a_400_62400# 0.19fF
C6147 VN.n5506 a_400_62400# 1.55fF
C6148 VN.n5507 a_400_62400# 0.29fF
C6149 VN.n5508 a_400_62400# 2.52fF
C6150 VN.t777 a_400_62400# 0.03fF
C6151 VN.n5509 a_400_62400# 0.32fF
C6152 VN.n5510 a_400_62400# 1.22fF
C6153 VN.n5511 a_400_62400# 0.07fF
C6154 VN.t394 a_400_62400# 0.03fF
C6155 VN.n5512 a_400_62400# 0.16fF
C6156 VN.n5513 a_400_62400# 0.19fF
C6157 VN.n5515 a_400_62400# 1.04fF
C6158 VN.n5516 a_400_62400# 2.60fF
C6159 VN.n5517 a_400_62400# 2.51fF
C6160 VN.n5518 a_400_62400# 0.16fF
C6161 VN.t670 a_400_62400# 0.03fF
C6162 VN.n5519 a_400_62400# 0.19fF
C6163 VN.t1797 a_400_62400# 0.03fF
C6164 VN.n5521 a_400_62400# 0.32fF
C6165 VN.n5522 a_400_62400# 0.48fF
C6166 VN.n5523 a_400_62400# 0.81fF
C6167 VN.n5524 a_400_62400# 2.46fF
C6168 VN.n5525 a_400_62400# 4.01fF
C6169 VN.t1269 a_400_62400# 0.03fF
C6170 VN.n5526 a_400_62400# 0.32fF
C6171 VN.n5527 a_400_62400# 1.22fF
C6172 VN.n5528 a_400_62400# 0.07fF
C6173 VN.t849 a_400_62400# 0.03fF
C6174 VN.n5529 a_400_62400# 0.16fF
C6175 VN.n5530 a_400_62400# 0.19fF
C6176 VN.n5532 a_400_62400# 2.53fF
C6177 VN.n5533 a_400_62400# 2.34fF
C6178 VN.t922 a_400_62400# 0.03fF
C6179 VN.n5534 a_400_62400# 0.32fF
C6180 VN.n5535 a_400_62400# 0.48fF
C6181 VN.n5536 a_400_62400# 0.81fF
C6182 VN.n5537 a_400_62400# 0.16fF
C6183 VN.t2330 a_400_62400# 0.03fF
C6184 VN.n5538 a_400_62400# 0.19fF
C6185 VN.n5540 a_400_62400# 1.55fF
C6186 VN.n5541 a_400_62400# 0.29fF
C6187 VN.n5542 a_400_62400# 3.27fF
C6188 VN.t401 a_400_62400# 0.03fF
C6189 VN.n5543 a_400_62400# 0.32fF
C6190 VN.n5544 a_400_62400# 1.22fF
C6191 VN.n5545 a_400_62400# 0.07fF
C6192 VN.t2513 a_400_62400# 0.03fF
C6193 VN.n5546 a_400_62400# 0.16fF
C6194 VN.n5547 a_400_62400# 0.19fF
C6195 VN.n5549 a_400_62400# 2.51fF
C6196 VN.n5550 a_400_62400# 0.56fF
C6197 VN.n5551 a_400_62400# 0.64fF
C6198 VN.n5552 a_400_62400# 0.12fF
C6199 VN.n5553 a_400_62400# 0.44fF
C6200 VN.n5554 a_400_62400# 0.40fF
C6201 VN.n5555 a_400_62400# 1.03fF
C6202 VN.n5556 a_400_62400# 0.79fF
C6203 VN.t2584 a_400_62400# 0.03fF
C6204 VN.n5557 a_400_62400# 0.32fF
C6205 VN.n5558 a_400_62400# 0.48fF
C6206 VN.n5559 a_400_62400# 0.81fF
C6207 VN.n5560 a_400_62400# 0.16fF
C6208 VN.t1580 a_400_62400# 0.03fF
C6209 VN.n5561 a_400_62400# 0.19fF
C6210 VN.n5563 a_400_62400# 3.50fF
C6211 VN.n5564 a_400_62400# 2.89fF
C6212 VN.t2049 a_400_62400# 0.03fF
C6213 VN.n5565 a_400_62400# 0.32fF
C6214 VN.n5566 a_400_62400# 1.22fF
C6215 VN.n5567 a_400_62400# 0.07fF
C6216 VN.t1650 a_400_62400# 0.03fF
C6217 VN.n5568 a_400_62400# 0.16fF
C6218 VN.n5569 a_400_62400# 0.19fF
C6219 VN.n5571 a_400_62400# 1.05fF
C6220 VN.n5572 a_400_62400# 3.07fF
C6221 VN.n5573 a_400_62400# 2.51fF
C6222 VN.n5574 a_400_62400# 0.16fF
C6223 VN.t715 a_400_62400# 0.03fF
C6224 VN.n5575 a_400_62400# 0.19fF
C6225 VN.t1840 a_400_62400# 0.03fF
C6226 VN.n5577 a_400_62400# 0.32fF
C6227 VN.n5578 a_400_62400# 0.48fF
C6228 VN.n5579 a_400_62400# 0.81fF
C6229 VN.n5580 a_400_62400# 1.86fF
C6230 VN.n5581 a_400_62400# 1.53fF
C6231 VN.n5582 a_400_62400# 0.47fF
C6232 VN.n5583 a_400_62400# 2.71fF
C6233 VN.t1314 a_400_62400# 0.03fF
C6234 VN.n5584 a_400_62400# 0.32fF
C6235 VN.n5585 a_400_62400# 1.22fF
C6236 VN.n5586 a_400_62400# 0.07fF
C6237 VN.t780 a_400_62400# 0.03fF
C6238 VN.n5587 a_400_62400# 0.16fF
C6239 VN.n5588 a_400_62400# 0.19fF
C6240 VN.n5590 a_400_62400# 2.53fF
C6241 VN.n5591 a_400_62400# 2.51fF
C6242 VN.t969 a_400_62400# 0.03fF
C6243 VN.n5592 a_400_62400# 0.32fF
C6244 VN.n5593 a_400_62400# 0.48fF
C6245 VN.n5594 a_400_62400# 0.81fF
C6246 VN.n5595 a_400_62400# 0.16fF
C6247 VN.t2370 a_400_62400# 0.03fF
C6248 VN.n5596 a_400_62400# 0.19fF
C6249 VN.n5598 a_400_62400# 1.55fF
C6250 VN.n5599 a_400_62400# 0.29fF
C6251 VN.n5600 a_400_62400# 2.52fF
C6252 VN.t453 a_400_62400# 0.03fF
C6253 VN.n5601 a_400_62400# 0.32fF
C6254 VN.n5602 a_400_62400# 1.22fF
C6255 VN.n5603 a_400_62400# 0.07fF
C6256 VN.t2429 a_400_62400# 0.03fF
C6257 VN.n5604 a_400_62400# 0.16fF
C6258 VN.n5605 a_400_62400# 0.19fF
C6259 VN.n5607 a_400_62400# 27.83fF
C6260 VN.n5608 a_400_62400# 3.93fF
C6261 VN.n5609 a_400_62400# 2.51fF
C6262 VN.n5610 a_400_62400# 0.16fF
C6263 VN.t1501 a_400_62400# 0.03fF
C6264 VN.n5611 a_400_62400# 0.19fF
C6265 VN.t70 a_400_62400# 0.03fF
C6266 VN.n5613 a_400_62400# 0.32fF
C6267 VN.n5614 a_400_62400# 0.48fF
C6268 VN.n5615 a_400_62400# 0.81fF
C6269 VN.n5616 a_400_62400# 1.46fF
C6270 VN.n5617 a_400_62400# 0.21fF
C6271 VN.n5618 a_400_62400# 2.81fF
C6272 VN.t1568 a_400_62400# 0.03fF
C6273 VN.n5619 a_400_62400# 0.16fF
C6274 VN.n5620 a_400_62400# 0.19fF
C6275 VN.t2099 a_400_62400# 0.03fF
C6276 VN.n5622 a_400_62400# 0.32fF
C6277 VN.n5623 a_400_62400# 1.22fF
C6278 VN.n5624 a_400_62400# 0.07fF
C6279 VN.n5625 a_400_62400# 2.51fF
C6280 VN.n5626 a_400_62400# 3.57fF
C6281 VN.t1758 a_400_62400# 0.03fF
C6282 VN.n5627 a_400_62400# 0.32fF
C6283 VN.n5628 a_400_62400# 0.48fF
C6284 VN.n5629 a_400_62400# 0.81fF
C6285 VN.n5630 a_400_62400# 0.16fF
C6286 VN.t634 a_400_62400# 0.03fF
C6287 VN.n5631 a_400_62400# 0.19fF
C6288 VN.n5633 a_400_62400# 3.93fF
C6289 VN.n5634 a_400_62400# 3.08fF
C6290 VN.t698 a_400_62400# 0.03fF
C6291 VN.n5635 a_400_62400# 0.16fF
C6292 VN.n5636 a_400_62400# 0.19fF
C6293 VN.t1222 a_400_62400# 0.03fF
C6294 VN.n5638 a_400_62400# 0.32fF
C6295 VN.n5639 a_400_62400# 1.22fF
C6296 VN.n5640 a_400_62400# 0.07fF
C6297 VN.n5641 a_400_62400# 2.51fF
C6298 VN.n5642 a_400_62400# 3.57fF
C6299 VN.t885 a_400_62400# 0.03fF
C6300 VN.n5643 a_400_62400# 0.32fF
C6301 VN.n5644 a_400_62400# 0.48fF
C6302 VN.n5645 a_400_62400# 0.81fF
C6303 VN.n5646 a_400_62400# 0.16fF
C6304 VN.t2291 a_400_62400# 0.03fF
C6305 VN.n5647 a_400_62400# 0.19fF
C6306 VN.n5649 a_400_62400# 3.75fF
C6307 VN.n5650 a_400_62400# 3.08fF
C6308 VN.t2475 a_400_62400# 0.03fF
C6309 VN.n5651 a_400_62400# 0.16fF
C6310 VN.n5652 a_400_62400# 0.19fF
C6311 VN.t358 a_400_62400# 0.03fF
C6312 VN.n5654 a_400_62400# 0.32fF
C6313 VN.n5655 a_400_62400# 1.22fF
C6314 VN.n5656 a_400_62400# 0.07fF
C6315 VN.n5657 a_400_62400# 2.51fF
C6316 VN.n5658 a_400_62400# 3.57fF
C6317 VN.t2546 a_400_62400# 0.03fF
C6318 VN.n5659 a_400_62400# 0.32fF
C6319 VN.n5660 a_400_62400# 0.48fF
C6320 VN.n5661 a_400_62400# 0.81fF
C6321 VN.n5662 a_400_62400# 0.16fF
C6322 VN.t1422 a_400_62400# 0.03fF
C6323 VN.n5663 a_400_62400# 0.19fF
C6324 VN.n5665 a_400_62400# 3.75fF
C6325 VN.n5666 a_400_62400# 3.08fF
C6326 VN.t1614 a_400_62400# 0.03fF
C6327 VN.n5667 a_400_62400# 0.16fF
C6328 VN.n5668 a_400_62400# 0.19fF
C6329 VN.t2007 a_400_62400# 0.03fF
C6330 VN.n5670 a_400_62400# 0.32fF
C6331 VN.n5671 a_400_62400# 1.22fF
C6332 VN.n5672 a_400_62400# 0.07fF
C6333 VN.n5673 a_400_62400# 2.51fF
C6334 VN.n5674 a_400_62400# 3.57fF
C6335 VN.t963 a_400_62400# 0.03fF
C6336 VN.n5675 a_400_62400# 0.32fF
C6337 VN.n5676 a_400_62400# 0.48fF
C6338 VN.n5677 a_400_62400# 0.81fF
C6339 VN.n5678 a_400_62400# 0.16fF
C6340 VN.t2351 a_400_62400# 0.03fF
C6341 VN.n5679 a_400_62400# 0.19fF
C6342 VN.n5681 a_400_62400# 3.75fF
C6343 VN.n5682 a_400_62400# 3.08fF
C6344 VN.t2531 a_400_62400# 0.03fF
C6345 VN.n5683 a_400_62400# 0.16fF
C6346 VN.n5684 a_400_62400# 0.19fF
C6347 VN.t1903 a_400_62400# 0.03fF
C6348 VN.n5686 a_400_62400# 0.32fF
C6349 VN.n5687 a_400_62400# 1.22fF
C6350 VN.n5688 a_400_62400# 0.07fF
C6351 VN.n5689 a_400_62400# 2.51fF
C6352 VN.n5690 a_400_62400# 3.57fF
C6353 VN.t56 a_400_62400# 0.03fF
C6354 VN.n5691 a_400_62400# 0.32fF
C6355 VN.n5692 a_400_62400# 0.48fF
C6356 VN.n5693 a_400_62400# 0.81fF
C6357 VN.n5694 a_400_62400# 0.16fF
C6358 VN.t1482 a_400_62400# 0.03fF
C6359 VN.n5695 a_400_62400# 0.19fF
C6360 VN.n5697 a_400_62400# 3.75fF
C6361 VN.n5698 a_400_62400# 3.08fF
C6362 VN.t1667 a_400_62400# 0.03fF
C6363 VN.n5699 a_400_62400# 0.16fF
C6364 VN.n5700 a_400_62400# 0.19fF
C6365 VN.t1029 a_400_62400# 0.03fF
C6366 VN.n5702 a_400_62400# 0.32fF
C6367 VN.n5703 a_400_62400# 1.22fF
C6368 VN.n5704 a_400_62400# 0.07fF
C6369 VN.n5705 a_400_62400# 3.65fF
C6370 VN.n5706 a_400_62400# 2.14fF
C6371 VN.n5707 a_400_62400# 0.16fF
C6372 VN.t2394 a_400_62400# 0.03fF
C6373 VN.n5708 a_400_62400# 0.19fF
C6374 VN.t875 a_400_62400# 0.03fF
C6375 VN.n5710 a_400_62400# 0.32fF
C6376 VN.n5711 a_400_62400# 0.48fF
C6377 VN.n5712 a_400_62400# 0.81fF
C6378 VN.n5713 a_400_62400# 0.09fF
C6379 VN.n5714 a_400_62400# 0.01fF
C6380 VN.n5715 a_400_62400# 0.02fF
C6381 VN.n5716 a_400_62400# 0.02fF
C6382 VN.n5717 a_400_62400# 0.32fF
C6383 VN.n5718 a_400_62400# 1.56fF
C6384 VN.n5719 a_400_62400# 1.81fF
C6385 VN.n5720 a_400_62400# 3.08fF
C6386 VN.t2455 a_400_62400# 0.03fF
C6387 VN.n5721 a_400_62400# 0.16fF
C6388 VN.n5722 a_400_62400# 0.19fF
C6389 VN.t1821 a_400_62400# 0.03fF
C6390 VN.n5724 a_400_62400# 0.32fF
C6391 VN.n5725 a_400_62400# 1.22fF
C6392 VN.n5726 a_400_62400# 0.07fF
C6393 VN.t176 a_400_62400# 64.69fF
C6394 VN.t159 a_400_62400# 0.03fF
C6395 VN.n5727 a_400_62400# 0.32fF
C6396 VN.n5728 a_400_62400# 1.22fF
C6397 VN.n5729 a_400_62400# 0.07fF
C6398 VN.t802 a_400_62400# 0.03fF
C6399 VN.n5730 a_400_62400# 0.16fF
C6400 VN.n5731 a_400_62400# 0.19fF
C6401 VN.n5733 a_400_62400# 0.16fF
C6402 VN.t616 a_400_62400# 0.03fF
C6403 VN.n5734 a_400_62400# 0.19fF
C6404 VN.n5736 a_400_62400# 6.92fF
C6405 VN.n5737 a_400_62400# 6.56fF
C6406 VN.t1577 a_400_62400# 0.03fF
C6407 VN.n5738 a_400_62400# 0.16fF
C6408 VN.n5739 a_400_62400# 0.19fF
C6409 VN.t1953 a_400_62400# 0.03fF
C6410 VN.n5741 a_400_62400# 0.32fF
C6411 VN.n5742 a_400_62400# 1.22fF
C6412 VN.n5743 a_400_62400# 0.07fF
C6413 VN.n5744 a_400_62400# 2.51fF
C6414 VN.n5745 a_400_62400# 3.58fF
C6415 VN.t1185 a_400_62400# 0.03fF
C6416 VN.n5746 a_400_62400# 0.32fF
C6417 VN.n5747 a_400_62400# 0.48fF
C6418 VN.n5748 a_400_62400# 0.81fF
C6419 VN.n5749 a_400_62400# 0.16fF
C6420 VN.t2547 a_400_62400# 0.03fF
C6421 VN.n5750 a_400_62400# 0.19fF
C6422 VN.n5752 a_400_62400# 7.29fF
C6423 VN.t710 a_400_62400# 0.03fF
C6424 VN.n5753 a_400_62400# 0.16fF
C6425 VN.n5754 a_400_62400# 0.19fF
C6426 VN.t1085 a_400_62400# 0.03fF
C6427 VN.n5756 a_400_62400# 0.32fF
C6428 VN.n5757 a_400_62400# 1.22fF
C6429 VN.n5758 a_400_62400# 0.07fF
C6430 VN.t71 a_400_62400# 64.17fF
C6431 VN.t212 a_400_62400# 0.03fF
C6432 VN.n5759 a_400_62400# 1.60fF
C6433 VN.n5760 a_400_62400# 0.07fF
C6434 VN.t2484 a_400_62400# 0.03fF
C6435 VN.n5761 a_400_62400# 0.02fF
C6436 VN.n5762 a_400_62400# 0.34fF
C6437 VN.n5764 a_400_62400# 2.01fF
C6438 VN.n5765 a_400_62400# 1.75fF
C6439 VN.n5766 a_400_62400# 0.37fF
C6440 VN.n5767 a_400_62400# 0.33fF
C6441 VN.n5768 a_400_62400# 5.88fF
C6442 VN.n5769 a_400_62400# 0.02fF
C6443 VN.n5770 a_400_62400# 0.02fF
C6444 VN.n5771 a_400_62400# 0.03fF
C6445 VN.n5772 a_400_62400# 0.05fF
C6446 VN.n5773 a_400_62400# 0.23fF
C6447 VN.n5774 a_400_62400# 0.02fF
C6448 VN.n5775 a_400_62400# 0.03fF
C6449 VN.n5776 a_400_62400# 0.01fF
C6450 VN.n5777 a_400_62400# 0.01fF
C6451 VN.n5778 a_400_62400# 0.01fF
C6452 VN.n5779 a_400_62400# 0.02fF
C6453 VN.n5780 a_400_62400# 0.03fF
C6454 VN.n5781 a_400_62400# 0.06fF
C6455 VN.n5782 a_400_62400# 0.05fF
C6456 VN.n5783 a_400_62400# 0.15fF
C6457 VN.n5784 a_400_62400# 0.51fF
C6458 VN.n5785 a_400_62400# 0.27fF
C6459 VN.n5786 a_400_62400# 37.46fF
C6460 VN.n5787 a_400_62400# 37.46fF
C6461 VN.n5788 a_400_62400# 0.79fF
C6462 VN.n5789 a_400_62400# 0.23fF
C6463 VN.n5790 a_400_62400# 1.18fF
C6464 VN.t158 a_400_62400# 28.64fF
C6465 VN.n5791 a_400_62400# 0.79fF
C6466 VN.n5792 a_400_62400# 0.11fF
C6467 VN.n5793 a_400_62400# 4.98fF
C6468 VN.n5794 a_400_62400# 0.80fF
C6469 VN.n5795 a_400_62400# 0.29fF
C6470 VN.n5796 a_400_62400# 1.96fF
C6471 VN.n5798 a_400_62400# 25.18fF
C6472 VN.n5800 a_400_62400# 1.87fF
C6473 VN.n5801 a_400_62400# 5.36fF
C6474 VN.n5802 a_400_62400# 1.81fF
C6475 VN.t1156 a_400_62400# 0.03fF
C6476 VN.n5803 a_400_62400# 0.85fF
C6477 VN.n5804 a_400_62400# 0.81fF
C6478 VN.n5805 a_400_62400# 0.33fF
C6479 VN.n5806 a_400_62400# 0.12fF
C6480 VN.n5807 a_400_62400# 0.28fF
C6481 VN.n5808 a_400_62400# 1.23fF
C6482 VN.n5809 a_400_62400# 0.59fF
C6483 VN.n5810 a_400_62400# 2.51fF
C6484 VN.n5811 a_400_62400# 0.16fF
C6485 VN.t1571 a_400_62400# 0.03fF
C6486 VN.n5812 a_400_62400# 0.19fF
C6487 VN.t2573 a_400_62400# 0.03fF
C6488 VN.n5814 a_400_62400# 0.32fF
C6489 VN.n5815 a_400_62400# 0.48fF
C6490 VN.n5816 a_400_62400# 0.81fF
C6491 VN.n5817 a_400_62400# 0.03fF
C6492 VN.n5818 a_400_62400# 0.01fF
C6493 VN.n5819 a_400_62400# 0.02fF
C6494 VN.n5820 a_400_62400# 0.11fF
C6495 VN.n5821 a_400_62400# 0.08fF
C6496 VN.n5822 a_400_62400# 0.04fF
C6497 VN.n5823 a_400_62400# 0.05fF
C6498 VN.n5824 a_400_62400# 1.34fF
C6499 VN.n5825 a_400_62400# 0.48fF
C6500 VN.n5826 a_400_62400# 2.51fF
C6501 VN.n5827 a_400_62400# 2.67fF
C6502 VN.t879 a_400_62400# 0.03fF
C6503 VN.n5828 a_400_62400# 0.32fF
C6504 VN.n5829 a_400_62400# 1.22fF
C6505 VN.n5830 a_400_62400# 0.07fF
C6506 VN.t2249 a_400_62400# 0.03fF
C6507 VN.n5831 a_400_62400# 0.16fF
C6508 VN.n5832 a_400_62400# 0.19fF
C6509 VN.n5834 a_400_62400# 2.53fF
C6510 VN.n5835 a_400_62400# 0.08fF
C6511 VN.n5836 a_400_62400# 0.04fF
C6512 VN.n5837 a_400_62400# 0.05fF
C6513 VN.n5838 a_400_62400# 1.33fF
C6514 VN.n5839 a_400_62400# 0.03fF
C6515 VN.n5840 a_400_62400# 0.01fF
C6516 VN.n5841 a_400_62400# 0.02fF
C6517 VN.n5842 a_400_62400# 0.11fF
C6518 VN.n5843 a_400_62400# 0.48fF
C6519 VN.n5844 a_400_62400# 2.48fF
C6520 VN.t1835 a_400_62400# 0.03fF
C6521 VN.n5845 a_400_62400# 0.32fF
C6522 VN.n5846 a_400_62400# 0.48fF
C6523 VN.n5847 a_400_62400# 0.81fF
C6524 VN.n5848 a_400_62400# 0.16fF
C6525 VN.t701 a_400_62400# 0.03fF
C6526 VN.n5849 a_400_62400# 0.19fF
C6527 VN.n5851 a_400_62400# 0.93fF
C6528 VN.n5852 a_400_62400# 0.30fF
C6529 VN.n5853 a_400_62400# 0.34fF
C6530 VN.n5854 a_400_62400# 0.12fF
C6531 VN.n5855 a_400_62400# 0.30fF
C6532 VN.n5856 a_400_62400# 0.93fF
C6533 VN.n5857 a_400_62400# 1.55fF
C6534 VN.n5858 a_400_62400# 0.29fF
C6535 VN.n5859 a_400_62400# 0.34fF
C6536 VN.n5860 a_400_62400# 0.12fF
C6537 VN.n5861 a_400_62400# 2.52fF
C6538 VN.t137 a_400_62400# 0.03fF
C6539 VN.n5862 a_400_62400# 0.32fF
C6540 VN.n5863 a_400_62400# 1.22fF
C6541 VN.n5864 a_400_62400# 0.07fF
C6542 VN.t1388 a_400_62400# 0.03fF
C6543 VN.n5865 a_400_62400# 0.16fF
C6544 VN.n5866 a_400_62400# 0.19fF
C6545 VN.n5868 a_400_62400# 0.33fF
C6546 VN.n5869 a_400_62400# 0.12fF
C6547 VN.n5870 a_400_62400# 0.28fF
C6548 VN.n5871 a_400_62400# 1.23fF
C6549 VN.n5872 a_400_62400# 0.59fF
C6550 VN.n5873 a_400_62400# 2.51fF
C6551 VN.n5874 a_400_62400# 0.16fF
C6552 VN.t2360 a_400_62400# 0.03fF
C6553 VN.n5875 a_400_62400# 0.19fF
C6554 VN.t959 a_400_62400# 0.03fF
C6555 VN.n5877 a_400_62400# 0.32fF
C6556 VN.n5878 a_400_62400# 0.48fF
C6557 VN.n5879 a_400_62400# 0.81fF
C6558 VN.n5880 a_400_62400# 0.03fF
C6559 VN.n5881 a_400_62400# 0.01fF
C6560 VN.n5882 a_400_62400# 0.02fF
C6561 VN.n5883 a_400_62400# 0.11fF
C6562 VN.n5884 a_400_62400# 0.08fF
C6563 VN.n5885 a_400_62400# 0.04fF
C6564 VN.n5886 a_400_62400# 0.05fF
C6565 VN.n5887 a_400_62400# 1.34fF
C6566 VN.n5888 a_400_62400# 0.48fF
C6567 VN.n5889 a_400_62400# 2.51fF
C6568 VN.n5890 a_400_62400# 2.67fF
C6569 VN.t1798 a_400_62400# 0.03fF
C6570 VN.n5891 a_400_62400# 0.32fF
C6571 VN.n5892 a_400_62400# 1.22fF
C6572 VN.n5893 a_400_62400# 0.07fF
C6573 VN.t522 a_400_62400# 0.03fF
C6574 VN.n5894 a_400_62400# 0.16fF
C6575 VN.n5895 a_400_62400# 0.19fF
C6576 VN.n5897 a_400_62400# 2.53fF
C6577 VN.n5898 a_400_62400# 0.08fF
C6578 VN.n5899 a_400_62400# 0.04fF
C6579 VN.n5900 a_400_62400# 0.05fF
C6580 VN.n5901 a_400_62400# 1.33fF
C6581 VN.n5902 a_400_62400# 0.03fF
C6582 VN.n5903 a_400_62400# 0.01fF
C6583 VN.n5904 a_400_62400# 0.02fF
C6584 VN.n5905 a_400_62400# 0.11fF
C6585 VN.n5906 a_400_62400# 0.48fF
C6586 VN.n5907 a_400_62400# 2.48fF
C6587 VN.t1464 a_400_62400# 0.03fF
C6588 VN.n5908 a_400_62400# 0.32fF
C6589 VN.n5909 a_400_62400# 0.48fF
C6590 VN.n5910 a_400_62400# 0.81fF
C6591 VN.n5911 a_400_62400# 0.16fF
C6592 VN.t313 a_400_62400# 0.03fF
C6593 VN.n5912 a_400_62400# 0.19fF
C6594 VN.n5914 a_400_62400# 0.93fF
C6595 VN.n5915 a_400_62400# 0.30fF
C6596 VN.n5916 a_400_62400# 0.34fF
C6597 VN.n5917 a_400_62400# 0.12fF
C6598 VN.n5918 a_400_62400# 0.30fF
C6599 VN.n5919 a_400_62400# 0.93fF
C6600 VN.n5920 a_400_62400# 1.55fF
C6601 VN.n5921 a_400_62400# 0.29fF
C6602 VN.n5922 a_400_62400# 0.34fF
C6603 VN.n5923 a_400_62400# 0.12fF
C6604 VN.n5924 a_400_62400# 2.52fF
C6605 VN.t2292 a_400_62400# 0.03fF
C6606 VN.n5925 a_400_62400# 0.32fF
C6607 VN.n5926 a_400_62400# 1.22fF
C6608 VN.n5927 a_400_62400# 0.07fF
C6609 VN.t2175 a_400_62400# 0.03fF
C6610 VN.n5928 a_400_62400# 0.16fF
C6611 VN.n5929 a_400_62400# 0.19fF
C6612 VN.n5931 a_400_62400# 0.33fF
C6613 VN.n5932 a_400_62400# 0.12fF
C6614 VN.n5933 a_400_62400# 0.28fF
C6615 VN.n5934 a_400_62400# 1.23fF
C6616 VN.n5935 a_400_62400# 0.59fF
C6617 VN.n5936 a_400_62400# 2.51fF
C6618 VN.n5937 a_400_62400# 0.16fF
C6619 VN.t1962 a_400_62400# 0.03fF
C6620 VN.n5938 a_400_62400# 0.19fF
C6621 VN.t592 a_400_62400# 0.03fF
C6622 VN.n5940 a_400_62400# 0.32fF
C6623 VN.n5941 a_400_62400# 0.48fF
C6624 VN.n5942 a_400_62400# 0.81fF
C6625 VN.n5943 a_400_62400# 0.03fF
C6626 VN.n5944 a_400_62400# 0.01fF
C6627 VN.n5945 a_400_62400# 0.02fF
C6628 VN.n5946 a_400_62400# 0.11fF
C6629 VN.n5947 a_400_62400# 0.08fF
C6630 VN.n5948 a_400_62400# 0.04fF
C6631 VN.n5949 a_400_62400# 0.05fF
C6632 VN.n5950 a_400_62400# 1.34fF
C6633 VN.n5951 a_400_62400# 0.48fF
C6634 VN.n5952 a_400_62400# 2.51fF
C6635 VN.n5953 a_400_62400# 2.67fF
C6636 VN.t1423 a_400_62400# 0.03fF
C6637 VN.n5954 a_400_62400# 0.32fF
C6638 VN.n5955 a_400_62400# 1.22fF
C6639 VN.n5956 a_400_62400# 0.07fF
C6640 VN.t75 a_400_62400# 0.03fF
C6641 VN.n5957 a_400_62400# 0.16fF
C6642 VN.n5958 a_400_62400# 0.19fF
C6643 VN.n5960 a_400_62400# 2.53fF
C6644 VN.n5961 a_400_62400# 0.05fF
C6645 VN.n5962 a_400_62400# 0.09fF
C6646 VN.n5963 a_400_62400# 0.07fF
C6647 VN.n5964 a_400_62400# 1.16fF
C6648 VN.n5965 a_400_62400# 0.01fF
C6649 VN.n5966 a_400_62400# 0.01fF
C6650 VN.n5967 a_400_62400# 0.01fF
C6651 VN.n5968 a_400_62400# 0.09fF
C6652 VN.n5969 a_400_62400# 0.91fF
C6653 VN.n5970 a_400_62400# 0.96fF
C6654 VN.t2245 a_400_62400# 0.03fF
C6655 VN.n5971 a_400_62400# 0.32fF
C6656 VN.n5972 a_400_62400# 0.48fF
C6657 VN.n5973 a_400_62400# 0.81fF
C6658 VN.n5974 a_400_62400# 0.16fF
C6659 VN.t1097 a_400_62400# 0.03fF
C6660 VN.n5975 a_400_62400# 0.19fF
C6661 VN.n5977 a_400_62400# 0.93fF
C6662 VN.n5978 a_400_62400# 0.30fF
C6663 VN.n5979 a_400_62400# 0.34fF
C6664 VN.n5980 a_400_62400# 0.12fF
C6665 VN.n5981 a_400_62400# 0.30fF
C6666 VN.n5982 a_400_62400# 0.93fF
C6667 VN.n5983 a_400_62400# 1.55fF
C6668 VN.n5984 a_400_62400# 0.29fF
C6669 VN.n5985 a_400_62400# 0.34fF
C6670 VN.n5986 a_400_62400# 0.12fF
C6671 VN.n5987 a_400_62400# 3.10fF
C6672 VN.t558 a_400_62400# 0.03fF
C6673 VN.n5988 a_400_62400# 0.32fF
C6674 VN.n5989 a_400_62400# 1.22fF
C6675 VN.n5990 a_400_62400# 0.07fF
C6676 VN.t1762 a_400_62400# 0.03fF
C6677 VN.n5991 a_400_62400# 0.16fF
C6678 VN.n5992 a_400_62400# 0.19fF
C6679 VN.n5994 a_400_62400# 2.51fF
C6680 VN.n5995 a_400_62400# 0.61fF
C6681 VN.n5996 a_400_62400# 0.30fF
C6682 VN.n5997 a_400_62400# 0.51fF
C6683 VN.n5998 a_400_62400# 0.21fF
C6684 VN.n5999 a_400_62400# 0.38fF
C6685 VN.n6000 a_400_62400# 0.29fF
C6686 VN.n6001 a_400_62400# 0.40fF
C6687 VN.n6002 a_400_62400# 0.28fF
C6688 VN.t1383 a_400_62400# 0.03fF
C6689 VN.n6003 a_400_62400# 0.32fF
C6690 VN.n6004 a_400_62400# 0.48fF
C6691 VN.n6005 a_400_62400# 0.81fF
C6692 VN.n6006 a_400_62400# 0.16fF
C6693 VN.t230 a_400_62400# 0.03fF
C6694 VN.n6007 a_400_62400# 0.19fF
C6695 VN.n6009 a_400_62400# 0.06fF
C6696 VN.n6010 a_400_62400# 0.04fF
C6697 VN.n6011 a_400_62400# 0.04fF
C6698 VN.n6012 a_400_62400# 0.14fF
C6699 VN.n6013 a_400_62400# 0.48fF
C6700 VN.n6014 a_400_62400# 0.50fF
C6701 VN.n6015 a_400_62400# 0.14fF
C6702 VN.n6016 a_400_62400# 0.16fF
C6703 VN.n6017 a_400_62400# 0.09fF
C6704 VN.n6018 a_400_62400# 0.16fF
C6705 VN.n6019 a_400_62400# 0.24fF
C6706 VN.n6020 a_400_62400# 5.35fF
C6707 VN.t2215 a_400_62400# 0.03fF
C6708 VN.n6021 a_400_62400# 0.32fF
C6709 VN.n6022 a_400_62400# 1.22fF
C6710 VN.n6023 a_400_62400# 0.07fF
C6711 VN.t1017 a_400_62400# 0.03fF
C6712 VN.n6024 a_400_62400# 0.16fF
C6713 VN.n6025 a_400_62400# 0.19fF
C6714 VN.n6027 a_400_62400# 0.33fF
C6715 VN.n6028 a_400_62400# 0.12fF
C6716 VN.n6029 a_400_62400# 0.28fF
C6717 VN.n6030 a_400_62400# 1.72fF
C6718 VN.n6031 a_400_62400# 0.71fF
C6719 VN.n6032 a_400_62400# 2.51fF
C6720 VN.n6033 a_400_62400# 0.16fF
C6721 VN.t1877 a_400_62400# 0.03fF
C6722 VN.n6034 a_400_62400# 0.19fF
C6723 VN.t518 a_400_62400# 0.03fF
C6724 VN.n6036 a_400_62400# 0.32fF
C6725 VN.n6037 a_400_62400# 0.48fF
C6726 VN.n6038 a_400_62400# 0.81fF
C6727 VN.n6039 a_400_62400# 0.95fF
C6728 VN.n6040 a_400_62400# 2.11fF
C6729 VN.n6041 a_400_62400# 3.28fF
C6730 VN.t1348 a_400_62400# 0.03fF
C6731 VN.n6042 a_400_62400# 0.32fF
C6732 VN.n6043 a_400_62400# 1.22fF
C6733 VN.n6044 a_400_62400# 0.07fF
C6734 VN.t144 a_400_62400# 0.03fF
C6735 VN.n6045 a_400_62400# 0.16fF
C6736 VN.n6046 a_400_62400# 0.19fF
C6737 VN.n6048 a_400_62400# 2.53fF
C6738 VN.n6049 a_400_62400# 0.08fF
C6739 VN.n6050 a_400_62400# 0.04fF
C6740 VN.n6051 a_400_62400# 0.05fF
C6741 VN.n6052 a_400_62400# 1.33fF
C6742 VN.n6053 a_400_62400# 0.03fF
C6743 VN.n6054 a_400_62400# 0.01fF
C6744 VN.n6055 a_400_62400# 0.02fF
C6745 VN.n6056 a_400_62400# 0.11fF
C6746 VN.n6057 a_400_62400# 0.48fF
C6747 VN.n6058 a_400_62400# 2.48fF
C6748 VN.t2169 a_400_62400# 0.03fF
C6749 VN.n6059 a_400_62400# 0.32fF
C6750 VN.n6060 a_400_62400# 0.48fF
C6751 VN.n6061 a_400_62400# 0.81fF
C6752 VN.n6062 a_400_62400# 0.16fF
C6753 VN.t1008 a_400_62400# 0.03fF
C6754 VN.n6063 a_400_62400# 0.19fF
C6755 VN.n6065 a_400_62400# 0.93fF
C6756 VN.n6066 a_400_62400# 0.30fF
C6757 VN.n6067 a_400_62400# 0.34fF
C6758 VN.n6068 a_400_62400# 0.12fF
C6759 VN.n6069 a_400_62400# 0.30fF
C6760 VN.n6070 a_400_62400# 0.93fF
C6761 VN.n6071 a_400_62400# 1.55fF
C6762 VN.n6072 a_400_62400# 0.29fF
C6763 VN.n6073 a_400_62400# 0.34fF
C6764 VN.n6074 a_400_62400# 0.12fF
C6765 VN.n6075 a_400_62400# 2.52fF
C6766 VN.t483 a_400_62400# 0.03fF
C6767 VN.n6076 a_400_62400# 0.32fF
C6768 VN.n6077 a_400_62400# 1.22fF
C6769 VN.n6078 a_400_62400# 0.07fF
C6770 VN.t1809 a_400_62400# 0.03fF
C6771 VN.n6079 a_400_62400# 0.16fF
C6772 VN.n6080 a_400_62400# 0.19fF
C6773 VN.n6082 a_400_62400# 27.83fF
C6774 VN.n6083 a_400_62400# 2.30fF
C6775 VN.n6084 a_400_62400# 4.08fF
C6776 VN.t911 a_400_62400# 0.03fF
C6777 VN.n6085 a_400_62400# 0.32fF
C6778 VN.n6086 a_400_62400# 0.48fF
C6779 VN.n6087 a_400_62400# 0.81fF
C6780 VN.n6088 a_400_62400# 0.16fF
C6781 VN.t2318 a_400_62400# 0.03fF
C6782 VN.n6089 a_400_62400# 0.19fF
C6783 VN.n6091 a_400_62400# 0.42fF
C6784 VN.n6092 a_400_62400# 0.34fF
C6785 VN.n6093 a_400_62400# 0.12fF
C6786 VN.n6094 a_400_62400# 0.30fF
C6787 VN.n6095 a_400_62400# 0.88fF
C6788 VN.n6096 a_400_62400# 1.28fF
C6789 VN.n6097 a_400_62400# 0.30fF
C6790 VN.n6098 a_400_62400# 0.28fF
C6791 VN.n6099 a_400_62400# 0.27fF
C6792 VN.n6100 a_400_62400# 0.09fF
C6793 VN.n6101 a_400_62400# 0.12fF
C6794 VN.n6102 a_400_62400# 0.13fF
C6795 VN.n6103 a_400_62400# 2.66fF
C6796 VN.t594 a_400_62400# 0.03fF
C6797 VN.n6104 a_400_62400# 0.16fF
C6798 VN.n6105 a_400_62400# 0.19fF
C6799 VN.t1753 a_400_62400# 0.03fF
C6800 VN.n6107 a_400_62400# 0.32fF
C6801 VN.n6108 a_400_62400# 1.22fF
C6802 VN.n6109 a_400_62400# 0.07fF
C6803 VN.n6110 a_400_62400# 2.51fF
C6804 VN.n6111 a_400_62400# 0.16fF
C6805 VN.t133 a_400_62400# 0.03fF
C6806 VN.n6112 a_400_62400# 0.19fF
C6807 VN.t1302 a_400_62400# 0.03fF
C6808 VN.n6114 a_400_62400# 0.32fF
C6809 VN.n6115 a_400_62400# 0.48fF
C6810 VN.n6116 a_400_62400# 0.81fF
C6811 VN.n6117 a_400_62400# 1.24fF
C6812 VN.n6118 a_400_62400# 0.43fF
C6813 VN.n6119 a_400_62400# 0.43fF
C6814 VN.n6120 a_400_62400# 1.24fF
C6815 VN.n6121 a_400_62400# 1.46fF
C6816 VN.n6122 a_400_62400# 0.21fF
C6817 VN.n6123 a_400_62400# 6.64fF
C6818 VN.t934 a_400_62400# 0.03fF
C6819 VN.n6124 a_400_62400# 0.16fF
C6820 VN.n6125 a_400_62400# 0.19fF
C6821 VN.t2137 a_400_62400# 0.03fF
C6822 VN.n6127 a_400_62400# 0.32fF
C6823 VN.n6128 a_400_62400# 1.22fF
C6824 VN.n6129 a_400_62400# 0.07fF
C6825 VN.n6130 a_400_62400# 2.51fF
C6826 VN.n6131 a_400_62400# 3.57fF
C6827 VN.t436 a_400_62400# 0.03fF
C6828 VN.n6132 a_400_62400# 0.32fF
C6829 VN.n6133 a_400_62400# 0.48fF
C6830 VN.n6134 a_400_62400# 0.81fF
C6831 VN.n6135 a_400_62400# 0.16fF
C6832 VN.t1929 a_400_62400# 0.03fF
C6833 VN.n6136 a_400_62400# 0.19fF
C6834 VN.n6138 a_400_62400# 6.91fF
C6835 VN.t11 a_400_62400# 0.03fF
C6836 VN.n6139 a_400_62400# 0.16fF
C6837 VN.n6140 a_400_62400# 0.19fF
C6838 VN.t1263 a_400_62400# 0.03fF
C6839 VN.n6142 a_400_62400# 0.32fF
C6840 VN.n6143 a_400_62400# 1.22fF
C6841 VN.n6144 a_400_62400# 0.07fF
C6842 VN.n6145 a_400_62400# 2.51fF
C6843 VN.n6146 a_400_62400# 3.57fF
C6844 VN.t2211 a_400_62400# 0.03fF
C6845 VN.n6147 a_400_62400# 0.32fF
C6846 VN.n6148 a_400_62400# 0.48fF
C6847 VN.n6149 a_400_62400# 0.81fF
C6848 VN.n6150 a_400_62400# 0.16fF
C6849 VN.t1054 a_400_62400# 0.03fF
C6850 VN.n6151 a_400_62400# 0.19fF
C6851 VN.n6153 a_400_62400# 6.92fF
C6852 VN.t1728 a_400_62400# 0.03fF
C6853 VN.n6154 a_400_62400# 0.16fF
C6854 VN.n6155 a_400_62400# 0.19fF
C6855 VN.t525 a_400_62400# 0.03fF
C6856 VN.n6157 a_400_62400# 0.32fF
C6857 VN.n6158 a_400_62400# 1.22fF
C6858 VN.n6159 a_400_62400# 0.07fF
C6859 VN.n6160 a_400_62400# 2.51fF
C6860 VN.n6161 a_400_62400# 3.57fF
C6861 VN.t2118 a_400_62400# 0.03fF
C6862 VN.n6162 a_400_62400# 0.32fF
C6863 VN.n6163 a_400_62400# 0.48fF
C6864 VN.n6164 a_400_62400# 0.81fF
C6865 VN.n6165 a_400_62400# 0.16fF
C6866 VN.t943 a_400_62400# 0.03fF
C6867 VN.n6166 a_400_62400# 0.19fF
C6868 VN.n6168 a_400_62400# 6.92fF
C6869 VN.t852 a_400_62400# 0.03fF
C6870 VN.n6169 a_400_62400# 0.16fF
C6871 VN.n6170 a_400_62400# 0.19fF
C6872 VN.t2014 a_400_62400# 0.03fF
C6873 VN.n6172 a_400_62400# 0.32fF
C6874 VN.n6173 a_400_62400# 1.22fF
C6875 VN.n6174 a_400_62400# 0.07fF
C6876 VN.n6175 a_400_62400# 2.51fF
C6877 VN.n6176 a_400_62400# 3.57fF
C6878 VN.t1241 a_400_62400# 0.03fF
C6879 VN.n6177 a_400_62400# 0.32fF
C6880 VN.n6178 a_400_62400# 0.48fF
C6881 VN.n6179 a_400_62400# 0.81fF
C6882 VN.n6180 a_400_62400# 0.16fF
C6883 VN.t18 a_400_62400# 0.03fF
C6884 VN.n6181 a_400_62400# 0.19fF
C6885 VN.n6183 a_400_62400# 6.92fF
C6886 VN.t758 a_400_62400# 0.03fF
C6887 VN.n6184 a_400_62400# 0.16fF
C6888 VN.n6185 a_400_62400# 0.19fF
C6889 VN.t1141 a_400_62400# 0.03fF
C6890 VN.n6187 a_400_62400# 0.32fF
C6891 VN.n6188 a_400_62400# 1.22fF
C6892 VN.n6189 a_400_62400# 0.07fF
C6893 VN.n6190 a_400_62400# 2.51fF
C6894 VN.n6191 a_400_62400# 3.57fF
C6895 VN.t376 a_400_62400# 0.03fF
C6896 VN.n6192 a_400_62400# 0.32fF
C6897 VN.n6193 a_400_62400# 0.48fF
C6898 VN.n6194 a_400_62400# 0.81fF
C6899 VN.n6195 a_400_62400# 0.16fF
C6900 VN.t1732 a_400_62400# 0.03fF
C6901 VN.n6196 a_400_62400# 0.19fF
C6902 VN.n6198 a_400_62400# 2.51fF
C6903 VN.n6199 a_400_62400# 3.59fF
C6904 VN.t7 a_400_62400# 0.03fF
C6905 VN.n6200 a_400_62400# 0.32fF
C6906 VN.n6201 a_400_62400# 0.48fF
C6907 VN.n6202 a_400_62400# 0.81fF
C6908 VN.t2554 a_400_62400# 0.03fF
C6909 VN.n6203 a_400_62400# 1.63fF
C6910 VN.n6204 a_400_62400# 0.81fF
C6911 VN.n6205 a_400_62400# 1.21fF
C6912 VN.n6206 a_400_62400# 1.54fF
C6913 VN.n6207 a_400_62400# 4.06fF
C6914 VN.t6 a_400_62400# 28.64fF
C6915 VN.n6208 a_400_62400# 28.43fF
C6916 VN.n6210 a_400_62400# 0.50fF
C6917 VN.n6211 a_400_62400# 0.31fF
C6918 VN.n6212 a_400_62400# 3.74fF
C6919 VN.n6213 a_400_62400# 3.29fF
C6920 VN.n6214 a_400_62400# 1.64fF
C6921 VN.n6215 a_400_62400# 0.49fF
C6922 VN.n6216 a_400_62400# 5.34fF
C6923 VN.n6217 a_400_62400# 0.34fF
C6924 VN.n6218 a_400_62400# 0.02fF
C6925 VN.t1695 a_400_62400# 0.03fF
C6926 VN.n6219 a_400_62400# 0.34fF
C6927 VN.t2017 a_400_62400# 0.03fF
C6928 VN.n6220 a_400_62400# 1.28fF
C6929 VN.n6221 a_400_62400# 0.94fF
C6930 VN.n6222 a_400_62400# 2.53fF
C6931 VN.n6223 a_400_62400# 2.51fF
C6932 VN.t1685 a_400_62400# 0.03fF
C6933 VN.n6224 a_400_62400# 0.32fF
C6934 VN.n6225 a_400_62400# 0.48fF
C6935 VN.n6226 a_400_62400# 0.81fF
C6936 VN.n6227 a_400_62400# 0.16fF
C6937 VN.t825 a_400_62400# 0.03fF
C6938 VN.n6228 a_400_62400# 0.19fF
C6939 VN.n6230 a_400_62400# 1.55fF
C6940 VN.n6231 a_400_62400# 0.29fF
C6941 VN.n6232 a_400_62400# 2.52fF
C6942 VN.t1144 a_400_62400# 0.03fF
C6943 VN.n6233 a_400_62400# 0.32fF
C6944 VN.n6234 a_400_62400# 1.22fF
C6945 VN.n6235 a_400_62400# 0.07fF
C6946 VN.t892 a_400_62400# 0.03fF
C6947 VN.n6236 a_400_62400# 0.16fF
C6948 VN.n6237 a_400_62400# 0.19fF
C6949 VN.n6239 a_400_62400# 1.04fF
C6950 VN.n6240 a_400_62400# 2.60fF
C6951 VN.n6241 a_400_62400# 2.51fF
C6952 VN.n6242 a_400_62400# 0.16fF
C6953 VN.t2489 a_400_62400# 0.03fF
C6954 VN.n6243 a_400_62400# 0.19fF
C6955 VN.t819 a_400_62400# 0.03fF
C6956 VN.n6245 a_400_62400# 0.32fF
C6957 VN.n6246 a_400_62400# 0.48fF
C6958 VN.n6247 a_400_62400# 0.81fF
C6959 VN.n6248 a_400_62400# 2.46fF
C6960 VN.n6249 a_400_62400# 4.01fF
C6961 VN.t280 a_400_62400# 0.03fF
C6962 VN.n6250 a_400_62400# 0.32fF
C6963 VN.n6251 a_400_62400# 1.22fF
C6964 VN.n6252 a_400_62400# 0.07fF
C6965 VN.t147 a_400_62400# 0.03fF
C6966 VN.n6253 a_400_62400# 0.16fF
C6967 VN.n6254 a_400_62400# 0.19fF
C6968 VN.n6256 a_400_62400# 2.53fF
C6969 VN.n6257 a_400_62400# 2.51fF
C6970 VN.t2476 a_400_62400# 0.03fF
C6971 VN.n6258 a_400_62400# 0.32fF
C6972 VN.n6259 a_400_62400# 0.48fF
C6973 VN.n6260 a_400_62400# 0.81fF
C6974 VN.n6261 a_400_62400# 0.16fF
C6975 VN.t1624 a_400_62400# 0.03fF
C6976 VN.n6262 a_400_62400# 0.19fF
C6977 VN.n6264 a_400_62400# 1.55fF
C6978 VN.n6265 a_400_62400# 0.29fF
C6979 VN.n6266 a_400_62400# 2.52fF
C6980 VN.t1931 a_400_62400# 0.03fF
C6981 VN.n6267 a_400_62400# 0.32fF
C6982 VN.n6268 a_400_62400# 1.22fF
C6983 VN.n6269 a_400_62400# 0.07fF
C6984 VN.t1811 a_400_62400# 0.03fF
C6985 VN.n6270 a_400_62400# 0.16fF
C6986 VN.n6271 a_400_62400# 0.19fF
C6987 VN.n6273 a_400_62400# 1.04fF
C6988 VN.n6274 a_400_62400# 2.60fF
C6989 VN.n6275 a_400_62400# 2.51fF
C6990 VN.n6276 a_400_62400# 0.16fF
C6991 VN.t753 a_400_62400# 0.03fF
C6992 VN.n6277 a_400_62400# 0.19fF
C6993 VN.t1615 a_400_62400# 0.03fF
C6994 VN.n6279 a_400_62400# 0.32fF
C6995 VN.n6280 a_400_62400# 0.48fF
C6996 VN.n6281 a_400_62400# 0.81fF
C6997 VN.n6282 a_400_62400# 2.46fF
C6998 VN.n6283 a_400_62400# 4.01fF
C6999 VN.t1056 a_400_62400# 0.03fF
C7000 VN.n6284 a_400_62400# 0.32fF
C7001 VN.n6285 a_400_62400# 1.22fF
C7002 VN.n6286 a_400_62400# 0.07fF
C7003 VN.t936 a_400_62400# 0.03fF
C7004 VN.n6287 a_400_62400# 0.16fF
C7005 VN.n6288 a_400_62400# 0.19fF
C7006 VN.n6290 a_400_62400# 2.53fF
C7007 VN.n6291 a_400_62400# 2.51fF
C7008 VN.t2106 a_400_62400# 0.03fF
C7009 VN.n6292 a_400_62400# 0.32fF
C7010 VN.n6293 a_400_62400# 0.48fF
C7011 VN.n6294 a_400_62400# 0.81fF
C7012 VN.n6295 a_400_62400# 0.16fF
C7013 VN.t1242 a_400_62400# 0.03fF
C7014 VN.n6296 a_400_62400# 0.19fF
C7015 VN.n6298 a_400_62400# 1.55fF
C7016 VN.n6299 a_400_62400# 0.29fF
C7017 VN.n6300 a_400_62400# 2.52fF
C7018 VN.t1543 a_400_62400# 0.03fF
C7019 VN.n6301 a_400_62400# 0.32fF
C7020 VN.n6302 a_400_62400# 1.22fF
C7021 VN.n6303 a_400_62400# 0.07fF
C7022 VN.t1434 a_400_62400# 0.03fF
C7023 VN.n6304 a_400_62400# 0.16fF
C7024 VN.n6305 a_400_62400# 0.19fF
C7025 VN.n6307 a_400_62400# 1.04fF
C7026 VN.n6308 a_400_62400# 2.60fF
C7027 VN.n6309 a_400_62400# 2.51fF
C7028 VN.n6310 a_400_62400# 0.16fF
C7029 VN.t377 a_400_62400# 0.03fF
C7030 VN.n6311 a_400_62400# 0.19fF
C7031 VN.t1229 a_400_62400# 0.03fF
C7032 VN.n6313 a_400_62400# 0.32fF
C7033 VN.n6314 a_400_62400# 0.48fF
C7034 VN.n6315 a_400_62400# 0.81fF
C7035 VN.n6316 a_400_62400# 2.46fF
C7036 VN.n6317 a_400_62400# 4.01fF
C7037 VN.t674 a_400_62400# 0.03fF
C7038 VN.n6318 a_400_62400# 0.32fF
C7039 VN.n6319 a_400_62400# 1.22fF
C7040 VN.n6320 a_400_62400# 0.07fF
C7041 VN.t568 a_400_62400# 0.03fF
C7042 VN.n6321 a_400_62400# 0.16fF
C7043 VN.n6322 a_400_62400# 0.19fF
C7044 VN.n6324 a_400_62400# 2.53fF
C7045 VN.n6325 a_400_62400# 2.34fF
C7046 VN.t364 a_400_62400# 0.03fF
C7047 VN.n6326 a_400_62400# 0.32fF
C7048 VN.n6327 a_400_62400# 0.48fF
C7049 VN.n6328 a_400_62400# 0.81fF
C7050 VN.n6329 a_400_62400# 0.16fF
C7051 VN.t2164 a_400_62400# 0.03fF
C7052 VN.n6330 a_400_62400# 0.19fF
C7053 VN.n6332 a_400_62400# 1.55fF
C7054 VN.n6333 a_400_62400# 0.29fF
C7055 VN.n6334 a_400_62400# 3.27fF
C7056 VN.t2333 a_400_62400# 0.03fF
C7057 VN.n6335 a_400_62400# 0.32fF
C7058 VN.n6336 a_400_62400# 1.22fF
C7059 VN.n6337 a_400_62400# 0.07fF
C7060 VN.t2227 a_400_62400# 0.03fF
C7061 VN.n6338 a_400_62400# 0.16fF
C7062 VN.n6339 a_400_62400# 0.19fF
C7063 VN.n6341 a_400_62400# 2.51fF
C7064 VN.n6342 a_400_62400# 0.56fF
C7065 VN.n6343 a_400_62400# 0.64fF
C7066 VN.n6344 a_400_62400# 0.12fF
C7067 VN.n6345 a_400_62400# 0.44fF
C7068 VN.n6346 a_400_62400# 0.40fF
C7069 VN.n6347 a_400_62400# 1.03fF
C7070 VN.n6348 a_400_62400# 0.79fF
C7071 VN.t2149 a_400_62400# 0.03fF
C7072 VN.n6349 a_400_62400# 0.32fF
C7073 VN.n6350 a_400_62400# 0.48fF
C7074 VN.n6351 a_400_62400# 0.81fF
C7075 VN.n6352 a_400_62400# 0.16fF
C7076 VN.t1297 a_400_62400# 0.03fF
C7077 VN.n6353 a_400_62400# 0.19fF
C7078 VN.n6355 a_400_62400# 3.50fF
C7079 VN.n6356 a_400_62400# 2.89fF
C7080 VN.t1586 a_400_62400# 0.03fF
C7081 VN.n6357 a_400_62400# 0.32fF
C7082 VN.n6358 a_400_62400# 1.22fF
C7083 VN.n6359 a_400_62400# 0.07fF
C7084 VN.t1361 a_400_62400# 0.03fF
C7085 VN.n6360 a_400_62400# 0.16fF
C7086 VN.n6361 a_400_62400# 0.19fF
C7087 VN.n6363 a_400_62400# 1.05fF
C7088 VN.n6364 a_400_62400# 3.07fF
C7089 VN.n6365 a_400_62400# 2.51fF
C7090 VN.n6366 a_400_62400# 0.16fF
C7091 VN.t431 a_400_62400# 0.03fF
C7092 VN.n6367 a_400_62400# 0.19fF
C7093 VN.t1280 a_400_62400# 0.03fF
C7094 VN.n6369 a_400_62400# 0.32fF
C7095 VN.n6370 a_400_62400# 0.48fF
C7096 VN.n6371 a_400_62400# 0.81fF
C7097 VN.n6372 a_400_62400# 1.86fF
C7098 VN.n6373 a_400_62400# 1.53fF
C7099 VN.n6374 a_400_62400# 0.47fF
C7100 VN.n6375 a_400_62400# 2.71fF
C7101 VN.t721 a_400_62400# 0.03fF
C7102 VN.n6376 a_400_62400# 0.32fF
C7103 VN.n6377 a_400_62400# 1.22fF
C7104 VN.n6378 a_400_62400# 0.07fF
C7105 VN.t494 a_400_62400# 0.03fF
C7106 VN.n6379 a_400_62400# 0.16fF
C7107 VN.n6380 a_400_62400# 0.19fF
C7108 VN.n6382 a_400_62400# 2.53fF
C7109 VN.n6383 a_400_62400# 2.51fF
C7110 VN.t413 a_400_62400# 0.03fF
C7111 VN.n6384 a_400_62400# 0.32fF
C7112 VN.n6385 a_400_62400# 0.48fF
C7113 VN.n6386 a_400_62400# 0.81fF
C7114 VN.n6387 a_400_62400# 0.16fF
C7115 VN.t2076 a_400_62400# 0.03fF
C7116 VN.n6388 a_400_62400# 0.19fF
C7117 VN.n6390 a_400_62400# 1.55fF
C7118 VN.n6391 a_400_62400# 0.29fF
C7119 VN.n6392 a_400_62400# 2.52fF
C7120 VN.t2374 a_400_62400# 0.03fF
C7121 VN.n6393 a_400_62400# 0.32fF
C7122 VN.n6394 a_400_62400# 1.22fF
C7123 VN.n6395 a_400_62400# 0.07fF
C7124 VN.t2151 a_400_62400# 0.03fF
C7125 VN.n6396 a_400_62400# 0.16fF
C7126 VN.n6397 a_400_62400# 0.19fF
C7127 VN.n6399 a_400_62400# 27.83fF
C7128 VN.n6400 a_400_62400# 3.93fF
C7129 VN.n6401 a_400_62400# 2.51fF
C7130 VN.n6402 a_400_62400# 0.16fF
C7131 VN.t1204 a_400_62400# 0.03fF
C7132 VN.n6403 a_400_62400# 0.19fF
C7133 VN.t2061 a_400_62400# 0.03fF
C7134 VN.n6405 a_400_62400# 0.32fF
C7135 VN.n6406 a_400_62400# 0.48fF
C7136 VN.n6407 a_400_62400# 0.81fF
C7137 VN.n6408 a_400_62400# 1.46fF
C7138 VN.n6409 a_400_62400# 0.21fF
C7139 VN.n6410 a_400_62400# 2.81fF
C7140 VN.t1283 a_400_62400# 0.03fF
C7141 VN.n6411 a_400_62400# 0.16fF
C7142 VN.n6412 a_400_62400# 0.19fF
C7143 VN.t1506 a_400_62400# 0.03fF
C7144 VN.n6414 a_400_62400# 0.32fF
C7145 VN.n6415 a_400_62400# 1.22fF
C7146 VN.n6416 a_400_62400# 0.07fF
C7147 VN.n6417 a_400_62400# 2.51fF
C7148 VN.n6418 a_400_62400# 3.57fF
C7149 VN.t1190 a_400_62400# 0.03fF
C7150 VN.n6419 a_400_62400# 0.32fF
C7151 VN.n6420 a_400_62400# 0.48fF
C7152 VN.n6421 a_400_62400# 0.81fF
C7153 VN.n6422 a_400_62400# 0.16fF
C7154 VN.t339 a_400_62400# 0.03fF
C7155 VN.n6423 a_400_62400# 0.19fF
C7156 VN.n6425 a_400_62400# 3.93fF
C7157 VN.n6426 a_400_62400# 3.08fF
C7158 VN.t538 a_400_62400# 0.03fF
C7159 VN.n6427 a_400_62400# 0.16fF
C7160 VN.n6428 a_400_62400# 0.19fF
C7161 VN.t639 a_400_62400# 0.03fF
C7162 VN.n6430 a_400_62400# 0.32fF
C7163 VN.n6431 a_400_62400# 1.22fF
C7164 VN.n6432 a_400_62400# 0.07fF
C7165 VN.n6433 a_400_62400# 2.51fF
C7166 VN.n6434 a_400_62400# 3.57fF
C7167 VN.t320 a_400_62400# 0.03fF
C7168 VN.n6435 a_400_62400# 0.32fF
C7169 VN.n6436 a_400_62400# 0.48fF
C7170 VN.n6437 a_400_62400# 0.81fF
C7171 VN.n6438 a_400_62400# 0.16fF
C7172 VN.t1982 a_400_62400# 0.03fF
C7173 VN.n6439 a_400_62400# 0.19fF
C7174 VN.n6441 a_400_62400# 3.75fF
C7175 VN.n6442 a_400_62400# 3.08fF
C7176 VN.t2193 a_400_62400# 0.03fF
C7177 VN.n6443 a_400_62400# 0.16fF
C7178 VN.n6444 a_400_62400# 0.19fF
C7179 VN.t2298 a_400_62400# 0.03fF
C7180 VN.n6446 a_400_62400# 0.32fF
C7181 VN.n6447 a_400_62400# 1.22fF
C7182 VN.n6448 a_400_62400# 0.07fF
C7183 VN.n6449 a_400_62400# 2.51fF
C7184 VN.n6450 a_400_62400# 3.57fF
C7185 VN.t1807 a_400_62400# 0.03fF
C7186 VN.n6451 a_400_62400# 0.32fF
C7187 VN.n6452 a_400_62400# 0.48fF
C7188 VN.n6453 a_400_62400# 0.81fF
C7189 VN.n6454 a_400_62400# 0.16fF
C7190 VN.t2339 a_400_62400# 0.03fF
C7191 VN.n6455 a_400_62400# 0.19fF
C7192 VN.n6457 a_400_62400# 3.75fF
C7193 VN.n6458 a_400_62400# 3.08fF
C7194 VN.t2519 a_400_62400# 0.03fF
C7195 VN.n6459 a_400_62400# 0.16fF
C7196 VN.n6460 a_400_62400# 0.19fF
C7197 VN.t229 a_400_62400# 0.03fF
C7198 VN.n6462 a_400_62400# 0.32fF
C7199 VN.n6463 a_400_62400# 1.22fF
C7200 VN.n6464 a_400_62400# 0.07fF
C7201 VN.n6465 a_400_62400# 2.51fF
C7202 VN.n6466 a_400_62400# 3.57fF
C7203 VN.t931 a_400_62400# 0.03fF
C7204 VN.n6467 a_400_62400# 0.32fF
C7205 VN.n6468 a_400_62400# 0.48fF
C7206 VN.n6469 a_400_62400# 0.81fF
C7207 VN.n6470 a_400_62400# 0.16fF
C7208 VN.t1472 a_400_62400# 0.03fF
C7209 VN.n6471 a_400_62400# 0.19fF
C7210 VN.n6473 a_400_62400# 3.75fF
C7211 VN.n6474 a_400_62400# 3.08fF
C7212 VN.t1659 a_400_62400# 0.03fF
C7213 VN.n6475 a_400_62400# 0.16fF
C7214 VN.n6476 a_400_62400# 0.19fF
C7215 VN.t1876 a_400_62400# 0.03fF
C7216 VN.n6478 a_400_62400# 0.32fF
C7217 VN.n6479 a_400_62400# 1.22fF
C7218 VN.n6480 a_400_62400# 0.07fF
C7219 VN.n6481 a_400_62400# 3.65fF
C7220 VN.n6482 a_400_62400# 2.14fF
C7221 VN.n6483 a_400_62400# 0.16fF
C7222 VN.t2382 a_400_62400# 0.03fF
C7223 VN.n6484 a_400_62400# 0.19fF
C7224 VN.t1724 a_400_62400# 0.03fF
C7225 VN.n6486 a_400_62400# 0.32fF
C7226 VN.n6487 a_400_62400# 0.48fF
C7227 VN.n6488 a_400_62400# 0.81fF
C7228 VN.n6489 a_400_62400# 0.09fF
C7229 VN.n6490 a_400_62400# 0.01fF
C7230 VN.n6491 a_400_62400# 0.02fF
C7231 VN.n6492 a_400_62400# 0.02fF
C7232 VN.n6493 a_400_62400# 0.32fF
C7233 VN.n6494 a_400_62400# 1.56fF
C7234 VN.n6495 a_400_62400# 1.81fF
C7235 VN.n6496 a_400_62400# 3.08fF
C7236 VN.t2444 a_400_62400# 0.03fF
C7237 VN.n6497 a_400_62400# 0.16fF
C7238 VN.n6498 a_400_62400# 0.19fF
C7239 VN.t132 a_400_62400# 0.03fF
C7240 VN.n6500 a_400_62400# 0.32fF
C7241 VN.n6501 a_400_62400# 1.22fF
C7242 VN.n6502 a_400_62400# 0.07fF
C7243 VN.t146 a_400_62400# 64.69fF
C7244 VN.t1007 a_400_62400# 0.03fF
C7245 VN.n6503 a_400_62400# 0.32fF
C7246 VN.n6504 a_400_62400# 1.22fF
C7247 VN.n6505 a_400_62400# 0.07fF
C7248 VN.t791 a_400_62400# 0.03fF
C7249 VN.n6506 a_400_62400# 0.16fF
C7250 VN.n6507 a_400_62400# 0.19fF
C7251 VN.n6509 a_400_62400# 0.16fF
C7252 VN.t605 a_400_62400# 0.03fF
C7253 VN.n6510 a_400_62400# 0.19fF
C7254 VN.n6512 a_400_62400# 6.92fF
C7255 VN.n6513 a_400_62400# 6.56fF
C7256 VN.t2414 a_400_62400# 0.03fF
C7257 VN.n6514 a_400_62400# 0.16fF
C7258 VN.n6515 a_400_62400# 0.19fF
C7259 VN.t276 a_400_62400# 0.03fF
C7260 VN.n6517 a_400_62400# 0.32fF
C7261 VN.n6518 a_400_62400# 1.22fF
C7262 VN.n6519 a_400_62400# 0.07fF
C7263 VN.n6520 a_400_62400# 2.51fF
C7264 VN.n6521 a_400_62400# 3.58fF
C7265 VN.t2030 a_400_62400# 0.03fF
C7266 VN.n6522 a_400_62400# 0.32fF
C7267 VN.n6523 a_400_62400# 0.48fF
C7268 VN.n6524 a_400_62400# 0.81fF
C7269 VN.n6525 a_400_62400# 0.16fF
C7270 VN.t857 a_400_62400# 0.03fF
C7271 VN.n6526 a_400_62400# 0.19fF
C7272 VN.n6528 a_400_62400# 7.29fF
C7273 VN.t1552 a_400_62400# 0.03fF
C7274 VN.n6529 a_400_62400# 0.16fF
C7275 VN.n6530 a_400_62400# 0.19fF
C7276 VN.t1926 a_400_62400# 0.03fF
C7277 VN.n6532 a_400_62400# 0.32fF
C7278 VN.n6533 a_400_62400# 1.22fF
C7279 VN.n6534 a_400_62400# 0.07fF
C7280 VN.t10 a_400_62400# 64.17fF
C7281 VN.t1050 a_400_62400# 0.03fF
C7282 VN.n6535 a_400_62400# 1.60fF
C7283 VN.n6536 a_400_62400# 0.07fF
C7284 VN.t804 a_400_62400# 0.03fF
C7285 VN.n6537 a_400_62400# 0.02fF
C7286 VN.n6538 a_400_62400# 0.34fF
C7287 VN.n6540 a_400_62400# 2.01fF
C7288 VN.n6541 a_400_62400# 1.75fF
C7289 VN.n6542 a_400_62400# 0.37fF
C7290 VN.n6543 a_400_62400# 0.33fF
C7291 VN.n6544 a_400_62400# 5.88fF
C7292 VN.n6545 a_400_62400# 0.02fF
C7293 VN.n6546 a_400_62400# 0.02fF
C7294 VN.n6547 a_400_62400# 0.03fF
C7295 VN.n6548 a_400_62400# 0.05fF
C7296 VN.n6549 a_400_62400# 0.23fF
C7297 VN.n6550 a_400_62400# 0.02fF
C7298 VN.n6551 a_400_62400# 0.03fF
C7299 VN.n6552 a_400_62400# 0.01fF
C7300 VN.n6553 a_400_62400# 0.01fF
C7301 VN.n6554 a_400_62400# 0.01fF
C7302 VN.n6555 a_400_62400# 0.02fF
C7303 VN.n6556 a_400_62400# 0.03fF
C7304 VN.n6557 a_400_62400# 0.06fF
C7305 VN.n6558 a_400_62400# 0.05fF
C7306 VN.n6559 a_400_62400# 0.15fF
C7307 VN.n6560 a_400_62400# 0.51fF
C7308 VN.n6561 a_400_62400# 0.27fF
C7309 VN.n6562 a_400_62400# 37.46fF
C7310 VN.n6563 a_400_62400# 37.46fF
C7311 VN.n6564 a_400_62400# 0.79fF
C7312 VN.n6565 a_400_62400# 0.23fF
C7313 VN.n6566 a_400_62400# 1.18fF
C7314 VN.t131 a_400_62400# 28.64fF
C7315 VN.n6567 a_400_62400# 0.79fF
C7316 VN.n6568 a_400_62400# 0.11fF
C7317 VN.n6569 a_400_62400# 4.98fF
C7318 VN.n6570 a_400_62400# 0.80fF
C7319 VN.n6571 a_400_62400# 0.29fF
C7320 VN.n6572 a_400_62400# 1.96fF
C7321 VN.n6574 a_400_62400# 25.18fF
C7322 VN.n6576 a_400_62400# 1.87fF
C7323 VN.n6577 a_400_62400# 5.36fF
C7324 VN.n6578 a_400_62400# 1.81fF
C7325 VN.t1998 a_400_62400# 0.03fF
C7326 VN.n6579 a_400_62400# 0.85fF
C7327 VN.n6580 a_400_62400# 0.81fF
C7328 VN.n6581 a_400_62400# 0.16fF
C7329 VN.t2590 a_400_62400# 0.03fF
C7330 VN.n6582 a_400_62400# 0.19fF
C7331 VN.t2336 a_400_62400# 0.03fF
C7332 VN.n6583 a_400_62400# 0.32fF
C7333 VN.n6584 a_400_62400# 1.24fF
C7334 VN.n6585 a_400_62400# 0.27fF
C7335 VN.n6586 a_400_62400# 0.09fF
C7336 VN.n6587 a_400_62400# 0.12fF
C7337 VN.n6588 a_400_62400# 0.28fF
C7338 VN.n6589 a_400_62400# 0.13fF
C7339 VN.n6590 a_400_62400# 0.41fF
C7340 VN.n6591 a_400_62400# 1.45fF
C7341 VN.n6592 a_400_62400# 0.72fF
C7342 VN.n6593 a_400_62400# 3.13fF
C7343 VN.n6594 a_400_62400# 2.54fF
C7344 VN.n6595 a_400_62400# 0.23fF
C7345 VN.n6596 a_400_62400# 1.02fF
C7346 VN.n6597 a_400_62400# 0.34fF
C7347 VN.n6598 a_400_62400# 0.40fF
C7348 VN.n6599 a_400_62400# 0.42fF
C7349 VN.n6600 a_400_62400# 0.63fF
C7350 VN.n6601 a_400_62400# 0.21fF
C7351 VN.t856 a_400_62400# 0.03fF
C7352 VN.n6602 a_400_62400# 0.16fF
C7353 VN.n6603 a_400_62400# 0.19fF
C7354 VN.n6604 a_400_62400# 2.51fF
C7355 VN.n6605 a_400_62400# 3.58fF
C7356 VN.t353 a_400_62400# 0.03fF
C7357 VN.n6606 a_400_62400# 0.32fF
C7358 VN.n6607 a_400_62400# 0.48fF
C7359 VN.n6608 a_400_62400# 0.81fF
C7360 VN.n6609 a_400_62400# 0.16fF
C7361 VN.t1708 a_400_62400# 0.03fF
C7362 VN.n6610 a_400_62400# 0.19fF
C7363 VN.n6612 a_400_62400# 7.29fF
C7364 VN.t1908 a_400_62400# 0.03fF
C7365 VN.n6613 a_400_62400# 0.32fF
C7366 VN.n6614 a_400_62400# 1.22fF
C7367 VN.n6615 a_400_62400# 0.07fF
C7368 VN.t2396 a_400_62400# 0.03fF
C7369 VN.n6616 a_400_62400# 0.16fF
C7370 VN.n6617 a_400_62400# 0.19fF
C7371 VN.n6619 a_400_62400# 2.51fF
C7372 VN.n6620 a_400_62400# 3.57fF
C7373 VN.t1215 a_400_62400# 0.03fF
C7374 VN.n6621 a_400_62400# 0.32fF
C7375 VN.n6622 a_400_62400# 0.48fF
C7376 VN.n6623 a_400_62400# 0.81fF
C7377 VN.n6624 a_400_62400# 0.16fF
C7378 VN.t2578 a_400_62400# 0.03fF
C7379 VN.n6625 a_400_62400# 0.19fF
C7380 VN.n6627 a_400_62400# 2.51fF
C7381 VN.n6628 a_400_62400# 3.59fF
C7382 VN.t2581 a_400_62400# 0.03fF
C7383 VN.n6629 a_400_62400# 0.32fF
C7384 VN.n6630 a_400_62400# 0.48fF
C7385 VN.n6631 a_400_62400# 0.81fF
C7386 VN.t614 a_400_62400# 0.03fF
C7387 VN.n6632 a_400_62400# 1.63fF
C7388 VN.n6633 a_400_62400# 0.81fF
C7389 VN.n6634 a_400_62400# 1.21fF
C7390 VN.n6635 a_400_62400# 1.54fF
C7391 VN.n6636 a_400_62400# 4.06fF
C7392 VN.t37 a_400_62400# 28.64fF
C7393 VN.n6637 a_400_62400# 28.43fF
C7394 VN.n6639 a_400_62400# 0.50fF
C7395 VN.n6640 a_400_62400# 0.31fF
C7396 VN.n6641 a_400_62400# 3.88fF
C7397 VN.n6642 a_400_62400# 3.29fF
C7398 VN.n6643 a_400_62400# 2.62fF
C7399 VN.n6644 a_400_62400# 5.27fF
C7400 VN.n6645 a_400_62400# 0.34fF
C7401 VN.n6646 a_400_62400# 0.02fF
C7402 VN.t1991 a_400_62400# 0.03fF
C7403 VN.n6647 a_400_62400# 0.34fF
C7404 VN.t2304 a_400_62400# 0.03fF
C7405 VN.n6648 a_400_62400# 1.28fF
C7406 VN.n6649 a_400_62400# 0.94fF
C7407 VN.n6650 a_400_62400# 1.05fF
C7408 VN.n6651 a_400_62400# 3.03fF
C7409 VN.n6652 a_400_62400# 2.51fF
C7410 VN.n6653 a_400_62400# 0.16fF
C7411 VN.t1117 a_400_62400# 0.03fF
C7412 VN.n6654 a_400_62400# 0.19fF
C7413 VN.t2266 a_400_62400# 0.03fF
C7414 VN.n6656 a_400_62400# 0.32fF
C7415 VN.n6657 a_400_62400# 0.48fF
C7416 VN.n6658 a_400_62400# 0.81fF
C7417 VN.n6659 a_400_62400# 2.03fF
C7418 VN.n6660 a_400_62400# 2.91fF
C7419 VN.t1432 a_400_62400# 0.03fF
C7420 VN.n6661 a_400_62400# 0.32fF
C7421 VN.n6662 a_400_62400# 1.22fF
C7422 VN.n6663 a_400_62400# 0.07fF
C7423 VN.t1197 a_400_62400# 0.03fF
C7424 VN.n6664 a_400_62400# 0.16fF
C7425 VN.n6665 a_400_62400# 0.19fF
C7426 VN.n6667 a_400_62400# 2.53fF
C7427 VN.n6668 a_400_62400# 2.51fF
C7428 VN.t1401 a_400_62400# 0.03fF
C7429 VN.n6669 a_400_62400# 0.32fF
C7430 VN.n6670 a_400_62400# 0.48fF
C7431 VN.n6671 a_400_62400# 0.81fF
C7432 VN.n6672 a_400_62400# 0.16fF
C7433 VN.t254 a_400_62400# 0.03fF
C7434 VN.n6673 a_400_62400# 0.19fF
C7435 VN.n6675 a_400_62400# 1.55fF
C7436 VN.n6676 a_400_62400# 0.29fF
C7437 VN.n6677 a_400_62400# 2.52fF
C7438 VN.t565 a_400_62400# 0.03fF
C7439 VN.n6678 a_400_62400# 0.32fF
C7440 VN.n6679 a_400_62400# 1.22fF
C7441 VN.n6680 a_400_62400# 0.07fF
C7442 VN.t468 a_400_62400# 0.03fF
C7443 VN.n6681 a_400_62400# 0.16fF
C7444 VN.n6682 a_400_62400# 0.19fF
C7445 VN.n6684 a_400_62400# 1.04fF
C7446 VN.n6685 a_400_62400# 2.60fF
C7447 VN.n6686 a_400_62400# 2.51fF
C7448 VN.n6687 a_400_62400# 0.16fF
C7449 VN.t1904 a_400_62400# 0.03fF
C7450 VN.n6688 a_400_62400# 0.19fF
C7451 VN.t540 a_400_62400# 0.03fF
C7452 VN.n6690 a_400_62400# 0.32fF
C7453 VN.n6691 a_400_62400# 0.48fF
C7454 VN.n6692 a_400_62400# 0.81fF
C7455 VN.n6693 a_400_62400# 2.46fF
C7456 VN.n6694 a_400_62400# 4.01fF
C7457 VN.t2225 a_400_62400# 0.03fF
C7458 VN.n6695 a_400_62400# 0.32fF
C7459 VN.n6696 a_400_62400# 1.22fF
C7460 VN.n6697 a_400_62400# 0.07fF
C7461 VN.t2119 a_400_62400# 0.03fF
C7462 VN.n6698 a_400_62400# 0.16fF
C7463 VN.n6699 a_400_62400# 0.19fF
C7464 VN.n6701 a_400_62400# 2.53fF
C7465 VN.n6702 a_400_62400# 2.51fF
C7466 VN.t2196 a_400_62400# 0.03fF
C7467 VN.n6703 a_400_62400# 0.32fF
C7468 VN.n6704 a_400_62400# 0.48fF
C7469 VN.n6705 a_400_62400# 0.81fF
C7470 VN.n6706 a_400_62400# 0.16fF
C7471 VN.t1030 a_400_62400# 0.03fF
C7472 VN.n6707 a_400_62400# 0.19fF
C7473 VN.n6709 a_400_62400# 1.55fF
C7474 VN.n6710 a_400_62400# 0.29fF
C7475 VN.n6711 a_400_62400# 2.52fF
C7476 VN.t1360 a_400_62400# 0.03fF
C7477 VN.n6712 a_400_62400# 0.32fF
C7478 VN.n6713 a_400_62400# 1.22fF
C7479 VN.n6714 a_400_62400# 0.07fF
C7480 VN.t1243 a_400_62400# 0.03fF
C7481 VN.n6715 a_400_62400# 0.16fF
C7482 VN.n6716 a_400_62400# 0.19fF
C7483 VN.n6718 a_400_62400# 1.04fF
C7484 VN.n6719 a_400_62400# 2.60fF
C7485 VN.n6720 a_400_62400# 2.51fF
C7486 VN.n6721 a_400_62400# 0.16fF
C7487 VN.t1526 a_400_62400# 0.03fF
C7488 VN.n6722 a_400_62400# 0.19fF
C7489 VN.t116 a_400_62400# 0.03fF
C7490 VN.n6724 a_400_62400# 0.32fF
C7491 VN.n6725 a_400_62400# 0.48fF
C7492 VN.n6726 a_400_62400# 0.81fF
C7493 VN.n6727 a_400_62400# 2.46fF
C7494 VN.n6728 a_400_62400# 4.01fF
C7495 VN.t1818 a_400_62400# 0.03fF
C7496 VN.n6729 a_400_62400# 0.32fF
C7497 VN.n6730 a_400_62400# 1.22fF
C7498 VN.n6731 a_400_62400# 0.07fF
C7499 VN.t1707 a_400_62400# 0.03fF
C7500 VN.n6732 a_400_62400# 0.16fF
C7501 VN.n6733 a_400_62400# 0.19fF
C7502 VN.n6735 a_400_62400# 2.53fF
C7503 VN.n6736 a_400_62400# 2.51fF
C7504 VN.t1784 a_400_62400# 0.03fF
C7505 VN.n6737 a_400_62400# 0.32fF
C7506 VN.n6738 a_400_62400# 0.48fF
C7507 VN.n6739 a_400_62400# 0.81fF
C7508 VN.n6740 a_400_62400# 0.16fF
C7509 VN.t658 a_400_62400# 0.03fF
C7510 VN.n6741 a_400_62400# 0.19fF
C7511 VN.n6743 a_400_62400# 1.55fF
C7512 VN.n6744 a_400_62400# 0.29fF
C7513 VN.n6745 a_400_62400# 2.52fF
C7514 VN.t946 a_400_62400# 0.03fF
C7515 VN.n6746 a_400_62400# 0.32fF
C7516 VN.n6747 a_400_62400# 1.22fF
C7517 VN.n6748 a_400_62400# 0.07fF
C7518 VN.t837 a_400_62400# 0.03fF
C7519 VN.n6749 a_400_62400# 0.16fF
C7520 VN.n6750 a_400_62400# 0.19fF
C7521 VN.n6752 a_400_62400# 1.04fF
C7522 VN.n6753 a_400_62400# 2.60fF
C7523 VN.n6754 a_400_62400# 2.51fF
C7524 VN.n6755 a_400_62400# 0.16fF
C7525 VN.t2431 a_400_62400# 0.03fF
C7526 VN.n6756 a_400_62400# 0.19fF
C7527 VN.t908 a_400_62400# 0.03fF
C7528 VN.n6758 a_400_62400# 0.32fF
C7529 VN.n6759 a_400_62400# 0.48fF
C7530 VN.n6760 a_400_62400# 0.81fF
C7531 VN.n6761 a_400_62400# 2.46fF
C7532 VN.n6762 a_400_62400# 4.01fF
C7533 VN.t23 a_400_62400# 0.03fF
C7534 VN.n6763 a_400_62400# 0.32fF
C7535 VN.n6764 a_400_62400# 1.22fF
C7536 VN.n6765 a_400_62400# 0.07fF
C7537 VN.t2500 a_400_62400# 0.03fF
C7538 VN.n6766 a_400_62400# 0.16fF
C7539 VN.n6767 a_400_62400# 0.19fF
C7540 VN.n6769 a_400_62400# 2.53fF
C7541 VN.n6770 a_400_62400# 2.34fF
C7542 VN.t170 a_400_62400# 0.03fF
C7543 VN.n6771 a_400_62400# 0.32fF
C7544 VN.n6772 a_400_62400# 0.48fF
C7545 VN.n6773 a_400_62400# 0.81fF
C7546 VN.n6774 a_400_62400# 0.16fF
C7547 VN.t1570 a_400_62400# 0.03fF
C7548 VN.n6775 a_400_62400# 0.19fF
C7549 VN.n6777 a_400_62400# 1.55fF
C7550 VN.n6778 a_400_62400# 0.29fF
C7551 VN.n6779 a_400_62400# 3.27fF
C7552 VN.t1864 a_400_62400# 0.03fF
C7553 VN.n6780 a_400_62400# 0.32fF
C7554 VN.n6781 a_400_62400# 1.22fF
C7555 VN.n6782 a_400_62400# 0.07fF
C7556 VN.t1637 a_400_62400# 0.03fF
C7557 VN.n6783 a_400_62400# 0.16fF
C7558 VN.n6784 a_400_62400# 0.19fF
C7559 VN.n6786 a_400_62400# 2.51fF
C7560 VN.n6787 a_400_62400# 0.56fF
C7561 VN.n6788 a_400_62400# 0.64fF
C7562 VN.n6789 a_400_62400# 0.12fF
C7563 VN.n6790 a_400_62400# 0.44fF
C7564 VN.n6791 a_400_62400# 0.40fF
C7565 VN.n6792 a_400_62400# 1.03fF
C7566 VN.n6793 a_400_62400# 0.79fF
C7567 VN.t1831 a_400_62400# 0.03fF
C7568 VN.n6794 a_400_62400# 0.32fF
C7569 VN.n6795 a_400_62400# 0.48fF
C7570 VN.n6796 a_400_62400# 0.81fF
C7571 VN.n6797 a_400_62400# 0.16fF
C7572 VN.t700 a_400_62400# 0.03fF
C7573 VN.n6798 a_400_62400# 0.19fF
C7574 VN.n6800 a_400_62400# 3.50fF
C7575 VN.n6801 a_400_62400# 2.89fF
C7576 VN.t994 a_400_62400# 0.03fF
C7577 VN.n6802 a_400_62400# 0.32fF
C7578 VN.n6803 a_400_62400# 1.22fF
C7579 VN.n6804 a_400_62400# 0.07fF
C7580 VN.t765 a_400_62400# 0.03fF
C7581 VN.n6805 a_400_62400# 0.16fF
C7582 VN.n6806 a_400_62400# 0.19fF
C7583 VN.n6808 a_400_62400# 1.05fF
C7584 VN.n6809 a_400_62400# 3.07fF
C7585 VN.n6810 a_400_62400# 2.51fF
C7586 VN.n6811 a_400_62400# 0.16fF
C7587 VN.t2357 a_400_62400# 0.03fF
C7588 VN.n6812 a_400_62400# 0.19fF
C7589 VN.t954 a_400_62400# 0.03fF
C7590 VN.n6814 a_400_62400# 0.32fF
C7591 VN.n6815 a_400_62400# 0.48fF
C7592 VN.n6816 a_400_62400# 0.81fF
C7593 VN.n6817 a_400_62400# 1.86fF
C7594 VN.n6818 a_400_62400# 1.53fF
C7595 VN.n6819 a_400_62400# 0.47fF
C7596 VN.n6820 a_400_62400# 2.71fF
C7597 VN.t112 a_400_62400# 0.03fF
C7598 VN.n6821 a_400_62400# 0.32fF
C7599 VN.n6822 a_400_62400# 1.22fF
C7600 VN.n6823 a_400_62400# 0.07fF
C7601 VN.t2419 a_400_62400# 0.03fF
C7602 VN.n6824 a_400_62400# 0.16fF
C7603 VN.n6825 a_400_62400# 0.19fF
C7604 VN.n6827 a_400_62400# 2.53fF
C7605 VN.n6828 a_400_62400# 2.51fF
C7606 VN.t38 a_400_62400# 0.03fF
C7607 VN.n6829 a_400_62400# 0.32fF
C7608 VN.n6830 a_400_62400# 0.48fF
C7609 VN.n6831 a_400_62400# 0.81fF
C7610 VN.n6832 a_400_62400# 0.16fF
C7611 VN.t1489 a_400_62400# 0.03fF
C7612 VN.n6833 a_400_62400# 0.19fF
C7613 VN.n6835 a_400_62400# 1.55fF
C7614 VN.n6836 a_400_62400# 0.29fF
C7615 VN.n6837 a_400_62400# 2.52fF
C7616 VN.t1780 a_400_62400# 0.03fF
C7617 VN.n6838 a_400_62400# 0.32fF
C7618 VN.n6839 a_400_62400# 1.22fF
C7619 VN.n6840 a_400_62400# 0.07fF
C7620 VN.t1557 a_400_62400# 0.03fF
C7621 VN.n6841 a_400_62400# 0.16fF
C7622 VN.n6842 a_400_62400# 0.19fF
C7623 VN.n6844 a_400_62400# 27.83fF
C7624 VN.n6845 a_400_62400# 3.93fF
C7625 VN.n6846 a_400_62400# 2.51fF
C7626 VN.n6847 a_400_62400# 0.16fF
C7627 VN.t623 a_400_62400# 0.03fF
C7628 VN.n6848 a_400_62400# 0.19fF
C7629 VN.t1741 a_400_62400# 0.03fF
C7630 VN.n6850 a_400_62400# 0.32fF
C7631 VN.n6851 a_400_62400# 0.48fF
C7632 VN.n6852 a_400_62400# 0.81fF
C7633 VN.n6853 a_400_62400# 1.46fF
C7634 VN.n6854 a_400_62400# 0.21fF
C7635 VN.n6855 a_400_62400# 2.81fF
C7636 VN.t807 a_400_62400# 0.03fF
C7637 VN.n6856 a_400_62400# 0.16fF
C7638 VN.n6857 a_400_62400# 0.19fF
C7639 VN.t905 a_400_62400# 0.03fF
C7640 VN.n6859 a_400_62400# 0.32fF
C7641 VN.n6860 a_400_62400# 1.22fF
C7642 VN.n6861 a_400_62400# 0.07fF
C7643 VN.n6862 a_400_62400# 2.51fF
C7644 VN.n6863 a_400_62400# 3.57fF
C7645 VN.t869 a_400_62400# 0.03fF
C7646 VN.n6864 a_400_62400# 0.32fF
C7647 VN.n6865 a_400_62400# 0.48fF
C7648 VN.n6866 a_400_62400# 0.81fF
C7649 VN.n6867 a_400_62400# 0.16fF
C7650 VN.t2274 a_400_62400# 0.03fF
C7651 VN.n6868 a_400_62400# 0.19fF
C7652 VN.n6870 a_400_62400# 3.93fF
C7653 VN.n6871 a_400_62400# 3.08fF
C7654 VN.t2461 a_400_62400# 0.03fF
C7655 VN.n6872 a_400_62400# 0.16fF
C7656 VN.n6873 a_400_62400# 0.19fF
C7657 VN.t2567 a_400_62400# 0.03fF
C7658 VN.n6875 a_400_62400# 0.32fF
C7659 VN.n6876 a_400_62400# 1.22fF
C7660 VN.n6877 a_400_62400# 0.07fF
C7661 VN.n6878 a_400_62400# 2.51fF
C7662 VN.n6879 a_400_62400# 3.57fF
C7663 VN.t1794 a_400_62400# 0.03fF
C7664 VN.n6880 a_400_62400# 0.32fF
C7665 VN.n6881 a_400_62400# 0.48fF
C7666 VN.n6882 a_400_62400# 0.81fF
C7667 VN.n6883 a_400_62400# 0.16fF
C7668 VN.t657 a_400_62400# 0.03fF
C7669 VN.n6884 a_400_62400# 0.19fF
C7670 VN.n6886 a_400_62400# 3.75fF
C7671 VN.n6887 a_400_62400# 3.08fF
C7672 VN.t836 a_400_62400# 0.03fF
C7673 VN.n6888 a_400_62400# 0.16fF
C7674 VN.n6889 a_400_62400# 0.19fF
C7675 VN.t1069 a_400_62400# 0.03fF
C7676 VN.n6891 a_400_62400# 0.32fF
C7677 VN.n6892 a_400_62400# 1.22fF
C7678 VN.n6893 a_400_62400# 0.07fF
C7679 VN.n6894 a_400_62400# 2.51fF
C7680 VN.n6895 a_400_62400# 3.57fF
C7681 VN.t919 a_400_62400# 0.03fF
C7682 VN.n6896 a_400_62400# 0.32fF
C7683 VN.n6897 a_400_62400# 0.48fF
C7684 VN.n6898 a_400_62400# 0.81fF
C7685 VN.n6899 a_400_62400# 0.16fF
C7686 VN.t2317 a_400_62400# 0.03fF
C7687 VN.n6900 a_400_62400# 0.19fF
C7688 VN.n6902 a_400_62400# 3.75fF
C7689 VN.n6903 a_400_62400# 3.08fF
C7690 VN.t2499 a_400_62400# 0.03fF
C7691 VN.n6904 a_400_62400# 0.16fF
C7692 VN.n6905 a_400_62400# 0.19fF
C7693 VN.t196 a_400_62400# 0.03fF
C7694 VN.n6907 a_400_62400# 0.32fF
C7695 VN.n6908 a_400_62400# 1.22fF
C7696 VN.n6909 a_400_62400# 0.07fF
C7697 VN.n6910 a_400_62400# 3.65fF
C7698 VN.n6911 a_400_62400# 2.14fF
C7699 VN.n6912 a_400_62400# 0.16fF
C7700 VN.t699 a_400_62400# 0.03fF
C7701 VN.n6913 a_400_62400# 0.19fF
C7702 VN.t1712 a_400_62400# 0.03fF
C7703 VN.n6915 a_400_62400# 0.32fF
C7704 VN.n6916 a_400_62400# 0.48fF
C7705 VN.n6917 a_400_62400# 0.81fF
C7706 VN.n6918 a_400_62400# 0.09fF
C7707 VN.n6919 a_400_62400# 0.01fF
C7708 VN.n6920 a_400_62400# 0.02fF
C7709 VN.n6921 a_400_62400# 0.02fF
C7710 VN.n6922 a_400_62400# 0.32fF
C7711 VN.n6923 a_400_62400# 1.56fF
C7712 VN.n6924 a_400_62400# 1.81fF
C7713 VN.n6925 a_400_62400# 3.08fF
C7714 VN.t764 a_400_62400# 0.03fF
C7715 VN.n6926 a_400_62400# 0.16fF
C7716 VN.n6927 a_400_62400# 0.19fF
C7717 VN.t981 a_400_62400# 0.03fF
C7718 VN.n6929 a_400_62400# 0.32fF
C7719 VN.n6930 a_400_62400# 1.22fF
C7720 VN.n6931 a_400_62400# 0.07fF
C7721 VN.t253 a_400_62400# 64.69fF
C7722 VN.t1852 a_400_62400# 0.03fF
C7723 VN.n6932 a_400_62400# 0.32fF
C7724 VN.n6933 a_400_62400# 1.22fF
C7725 VN.n6934 a_400_62400# 0.07fF
C7726 VN.t1636 a_400_62400# 0.03fF
C7727 VN.n6935 a_400_62400# 0.16fF
C7728 VN.n6936 a_400_62400# 0.19fF
C7729 VN.n6938 a_400_62400# 0.16fF
C7730 VN.t1449 a_400_62400# 0.03fF
C7731 VN.n6939 a_400_62400# 0.19fF
C7732 VN.n6941 a_400_62400# 6.92fF
C7733 VN.n6942 a_400_62400# 6.56fF
C7734 VN.t259 a_400_62400# 0.03fF
C7735 VN.n6943 a_400_62400# 0.32fF
C7736 VN.n6944 a_400_62400# 1.22fF
C7737 VN.n6945 a_400_62400# 0.07fF
C7738 VN.t739 a_400_62400# 0.03fF
C7739 VN.n6946 a_400_62400# 0.16fF
C7740 VN.n6947 a_400_62400# 0.19fF
C7741 VN.n6949 a_400_62400# 2.51fF
C7742 VN.n6950 a_400_62400# 3.57fF
C7743 VN.t2092 a_400_62400# 0.03fF
C7744 VN.n6951 a_400_62400# 0.32fF
C7745 VN.n6952 a_400_62400# 0.48fF
C7746 VN.n6953 a_400_62400# 0.81fF
C7747 VN.n6954 a_400_62400# 0.16fF
C7748 VN.t914 a_400_62400# 0.03fF
C7749 VN.n6955 a_400_62400# 0.19fF
C7750 VN.n6957 a_400_62400# 6.92fF
C7751 VN.t1122 a_400_62400# 0.03fF
C7752 VN.n6958 a_400_62400# 0.32fF
C7753 VN.n6959 a_400_62400# 1.22fF
C7754 VN.n6960 a_400_62400# 0.07fF
C7755 VN.t1606 a_400_62400# 0.03fF
C7756 VN.n6961 a_400_62400# 0.16fF
C7757 VN.n6962 a_400_62400# 0.19fF
C7758 VN.n6964 a_400_62400# 2.51fF
C7759 VN.n6965 a_400_62400# 3.57fF
C7760 VN.t445 a_400_62400# 0.03fF
C7761 VN.n6966 a_400_62400# 0.32fF
C7762 VN.n6967 a_400_62400# 0.48fF
C7763 VN.n6968 a_400_62400# 0.81fF
C7764 VN.n6969 a_400_62400# 0.16fF
C7765 VN.t1789 a_400_62400# 0.03fF
C7766 VN.n6970 a_400_62400# 0.19fF
C7767 VN.n6972 a_400_62400# 6.92fF
C7768 VN.t1995 a_400_62400# 0.03fF
C7769 VN.n6973 a_400_62400# 0.32fF
C7770 VN.n6974 a_400_62400# 1.22fF
C7771 VN.n6975 a_400_62400# 0.07fF
C7772 VN.t1152 a_400_62400# 0.03fF
C7773 VN.n6976 a_400_62400# 0.16fF
C7774 VN.n6977 a_400_62400# 0.19fF
C7775 VN.n6979 a_400_62400# 2.51fF
C7776 VN.n6980 a_400_62400# 3.57fF
C7777 VN.t2480 a_400_62400# 0.03fF
C7778 VN.n6981 a_400_62400# 0.32fF
C7779 VN.n6982 a_400_62400# 0.48fF
C7780 VN.n6983 a_400_62400# 0.81fF
C7781 VN.n6984 a_400_62400# 0.16fF
C7782 VN.t1359 a_400_62400# 0.03fF
C7783 VN.n6985 a_400_62400# 0.19fF
C7784 VN.n6987 a_400_62400# 6.91fF
C7785 VN.t1077 a_400_62400# 0.03fF
C7786 VN.n6988 a_400_62400# 0.32fF
C7787 VN.n6989 a_400_62400# 1.22fF
C7788 VN.n6990 a_400_62400# 0.07fF
C7789 VN.t2027 a_400_62400# 0.03fF
C7790 VN.n6991 a_400_62400# 0.16fF
C7791 VN.n6992 a_400_62400# 0.19fF
C7792 VN.n6994 a_400_62400# 2.51fF
C7793 VN.n6995 a_400_62400# 0.16fF
C7794 VN.t2224 a_400_62400# 0.03fF
C7795 VN.n6996 a_400_62400# 0.19fF
C7796 VN.t707 a_400_62400# 0.03fF
C7797 VN.n6998 a_400_62400# 0.32fF
C7798 VN.n6999 a_400_62400# 0.48fF
C7799 VN.n7000 a_400_62400# 0.81fF
C7800 VN.n7001 a_400_62400# 1.24fF
C7801 VN.n7002 a_400_62400# 0.43fF
C7802 VN.n7003 a_400_62400# 0.43fF
C7803 VN.n7004 a_400_62400# 1.24fF
C7804 VN.n7005 a_400_62400# 1.46fF
C7805 VN.n7006 a_400_62400# 0.21fF
C7806 VN.n7007 a_400_62400# 6.64fF
C7807 VN.t1813 a_400_62400# 0.03fF
C7808 VN.n7008 a_400_62400# 0.32fF
C7809 VN.n7009 a_400_62400# 1.22fF
C7810 VN.n7010 a_400_62400# 0.07fF
C7811 VN.t374 a_400_62400# 0.03fF
C7812 VN.n7011 a_400_62400# 0.16fF
C7813 VN.n7012 a_400_62400# 0.19fF
C7814 VN.n7014 a_400_62400# 2.53fF
C7815 VN.n7015 a_400_62400# 0.08fF
C7816 VN.n7016 a_400_62400# 0.04fF
C7817 VN.n7017 a_400_62400# 0.05fF
C7818 VN.n7018 a_400_62400# 1.33fF
C7819 VN.n7019 a_400_62400# 0.03fF
C7820 VN.n7020 a_400_62400# 0.01fF
C7821 VN.n7021 a_400_62400# 0.02fF
C7822 VN.n7022 a_400_62400# 0.11fF
C7823 VN.n7023 a_400_62400# 0.48fF
C7824 VN.n7024 a_400_62400# 2.48fF
C7825 VN.t356 a_400_62400# 0.03fF
C7826 VN.n7025 a_400_62400# 0.32fF
C7827 VN.n7026 a_400_62400# 0.48fF
C7828 VN.n7027 a_400_62400# 0.81fF
C7829 VN.n7028 a_400_62400# 0.16fF
C7830 VN.t1844 a_400_62400# 0.03fF
C7831 VN.n7029 a_400_62400# 0.19fF
C7832 VN.n7031 a_400_62400# 0.93fF
C7833 VN.n7032 a_400_62400# 0.30fF
C7834 VN.n7033 a_400_62400# 0.34fF
C7835 VN.n7034 a_400_62400# 0.12fF
C7836 VN.n7035 a_400_62400# 0.30fF
C7837 VN.n7036 a_400_62400# 0.93fF
C7838 VN.n7037 a_400_62400# 1.55fF
C7839 VN.n7038 a_400_62400# 0.29fF
C7840 VN.n7039 a_400_62400# 0.34fF
C7841 VN.n7040 a_400_62400# 0.12fF
C7842 VN.n7041 a_400_62400# 2.52fF
C7843 VN.t1471 a_400_62400# 0.03fF
C7844 VN.n7042 a_400_62400# 0.32fF
C7845 VN.n7043 a_400_62400# 1.22fF
C7846 VN.n7044 a_400_62400# 0.07fF
C7847 VN.t2518 a_400_62400# 0.03fF
C7848 VN.n7045 a_400_62400# 0.16fF
C7849 VN.n7046 a_400_62400# 0.19fF
C7850 VN.n7048 a_400_62400# 0.33fF
C7851 VN.n7049 a_400_62400# 0.12fF
C7852 VN.n7050 a_400_62400# 0.28fF
C7853 VN.n7051 a_400_62400# 1.23fF
C7854 VN.n7052 a_400_62400# 0.59fF
C7855 VN.n7053 a_400_62400# 2.51fF
C7856 VN.n7054 a_400_62400# 0.16fF
C7857 VN.t972 a_400_62400# 0.03fF
C7858 VN.n7055 a_400_62400# 0.19fF
C7859 VN.t2144 a_400_62400# 0.03fF
C7860 VN.n7057 a_400_62400# 0.32fF
C7861 VN.n7058 a_400_62400# 0.48fF
C7862 VN.n7059 a_400_62400# 0.81fF
C7863 VN.n7060 a_400_62400# 0.03fF
C7864 VN.n7061 a_400_62400# 0.01fF
C7865 VN.n7062 a_400_62400# 0.02fF
C7866 VN.n7063 a_400_62400# 0.11fF
C7867 VN.n7064 a_400_62400# 0.08fF
C7868 VN.n7065 a_400_62400# 0.04fF
C7869 VN.n7066 a_400_62400# 0.05fF
C7870 VN.n7067 a_400_62400# 1.34fF
C7871 VN.n7068 a_400_62400# 0.48fF
C7872 VN.n7069 a_400_62400# 2.51fF
C7873 VN.n7070 a_400_62400# 2.67fF
C7874 VN.t727 a_400_62400# 0.03fF
C7875 VN.n7071 a_400_62400# 0.32fF
C7876 VN.n7072 a_400_62400# 1.22fF
C7877 VN.n7073 a_400_62400# 0.07fF
C7878 VN.t1658 a_400_62400# 0.03fF
C7879 VN.n7074 a_400_62400# 0.16fF
C7880 VN.n7075 a_400_62400# 0.19fF
C7881 VN.n7077 a_400_62400# 2.53fF
C7882 VN.n7078 a_400_62400# 0.08fF
C7883 VN.n7079 a_400_62400# 0.04fF
C7884 VN.n7080 a_400_62400# 0.05fF
C7885 VN.n7081 a_400_62400# 1.33fF
C7886 VN.n7082 a_400_62400# 0.03fF
C7887 VN.n7083 a_400_62400# 0.01fF
C7888 VN.n7084 a_400_62400# 0.02fF
C7889 VN.n7085 a_400_62400# 0.11fF
C7890 VN.n7086 a_400_62400# 0.48fF
C7891 VN.n7087 a_400_62400# 2.48fF
C7892 VN.t1270 a_400_62400# 0.03fF
C7893 VN.n7088 a_400_62400# 0.32fF
C7894 VN.n7089 a_400_62400# 0.48fF
C7895 VN.n7090 a_400_62400# 0.81fF
C7896 VN.n7091 a_400_62400# 0.16fF
C7897 VN.t77 a_400_62400# 0.03fF
C7898 VN.n7092 a_400_62400# 0.19fF
C7899 VN.n7094 a_400_62400# 0.93fF
C7900 VN.n7095 a_400_62400# 0.30fF
C7901 VN.n7096 a_400_62400# 0.34fF
C7902 VN.n7097 a_400_62400# 0.12fF
C7903 VN.n7098 a_400_62400# 0.30fF
C7904 VN.n7099 a_400_62400# 0.93fF
C7905 VN.n7100 a_400_62400# 1.55fF
C7906 VN.n7101 a_400_62400# 0.29fF
C7907 VN.n7102 a_400_62400# 0.34fF
C7908 VN.n7103 a_400_62400# 0.12fF
C7909 VN.n7104 a_400_62400# 2.52fF
C7910 VN.t2378 a_400_62400# 0.03fF
C7911 VN.n7105 a_400_62400# 0.32fF
C7912 VN.n7106 a_400_62400# 1.22fF
C7913 VN.n7107 a_400_62400# 0.07fF
C7914 VN.t790 a_400_62400# 0.03fF
C7915 VN.n7108 a_400_62400# 0.16fF
C7916 VN.n7109 a_400_62400# 0.19fF
C7917 VN.n7111 a_400_62400# 0.33fF
C7918 VN.n7112 a_400_62400# 0.12fF
C7919 VN.n7113 a_400_62400# 0.28fF
C7920 VN.n7114 a_400_62400# 1.23fF
C7921 VN.n7115 a_400_62400# 0.59fF
C7922 VN.n7116 a_400_62400# 2.51fF
C7923 VN.n7117 a_400_62400# 0.16fF
C7924 VN.t604 a_400_62400# 0.03fF
C7925 VN.n7118 a_400_62400# 0.19fF
C7926 VN.t1729 a_400_62400# 0.03fF
C7927 VN.n7120 a_400_62400# 0.32fF
C7928 VN.n7121 a_400_62400# 0.48fF
C7929 VN.n7122 a_400_62400# 0.81fF
C7930 VN.n7123 a_400_62400# 0.03fF
C7931 VN.n7124 a_400_62400# 0.01fF
C7932 VN.n7125 a_400_62400# 0.02fF
C7933 VN.n7126 a_400_62400# 0.11fF
C7934 VN.n7127 a_400_62400# 0.08fF
C7935 VN.n7128 a_400_62400# 0.04fF
C7936 VN.n7129 a_400_62400# 0.05fF
C7937 VN.n7130 a_400_62400# 1.34fF
C7938 VN.n7131 a_400_62400# 0.48fF
C7939 VN.n7132 a_400_62400# 2.51fF
C7940 VN.n7133 a_400_62400# 2.67fF
C7941 VN.t342 a_400_62400# 0.03fF
C7942 VN.n7134 a_400_62400# 0.32fF
C7943 VN.n7135 a_400_62400# 1.22fF
C7944 VN.n7136 a_400_62400# 0.07fF
C7945 VN.t2443 a_400_62400# 0.03fF
C7946 VN.n7137 a_400_62400# 0.16fF
C7947 VN.n7138 a_400_62400# 0.19fF
C7948 VN.n7140 a_400_62400# 2.53fF
C7949 VN.n7141 a_400_62400# 0.08fF
C7950 VN.n7142 a_400_62400# 0.04fF
C7951 VN.n7143 a_400_62400# 0.05fF
C7952 VN.n7144 a_400_62400# 1.33fF
C7953 VN.n7145 a_400_62400# 0.03fF
C7954 VN.n7146 a_400_62400# 0.01fF
C7955 VN.n7147 a_400_62400# 0.02fF
C7956 VN.n7148 a_400_62400# 0.11fF
C7957 VN.n7149 a_400_62400# 0.48fF
C7958 VN.n7150 a_400_62400# 2.48fF
C7959 VN.t854 a_400_62400# 0.03fF
C7960 VN.n7151 a_400_62400# 0.32fF
C7961 VN.n7152 a_400_62400# 0.48fF
C7962 VN.n7153 a_400_62400# 0.81fF
C7963 VN.n7154 a_400_62400# 0.16fF
C7964 VN.t2257 a_400_62400# 0.03fF
C7965 VN.n7155 a_400_62400# 0.19fF
C7966 VN.n7157 a_400_62400# 0.93fF
C7967 VN.n7158 a_400_62400# 0.30fF
C7968 VN.n7159 a_400_62400# 0.34fF
C7969 VN.n7160 a_400_62400# 0.12fF
C7970 VN.n7161 a_400_62400# 0.30fF
C7971 VN.n7162 a_400_62400# 0.93fF
C7972 VN.n7163 a_400_62400# 1.55fF
C7973 VN.n7164 a_400_62400# 0.29fF
C7974 VN.n7165 a_400_62400# 0.34fF
C7975 VN.n7166 a_400_62400# 0.12fF
C7976 VN.n7167 a_400_62400# 2.52fF
C7977 VN.t1986 a_400_62400# 0.03fF
C7978 VN.n7168 a_400_62400# 0.32fF
C7979 VN.n7169 a_400_62400# 1.22fF
C7980 VN.n7170 a_400_62400# 0.07fF
C7981 VN.t418 a_400_62400# 0.03fF
C7982 VN.n7171 a_400_62400# 0.16fF
C7983 VN.n7172 a_400_62400# 0.19fF
C7984 VN.n7174 a_400_62400# 0.33fF
C7985 VN.n7175 a_400_62400# 0.12fF
C7986 VN.n7176 a_400_62400# 0.28fF
C7987 VN.n7177 a_400_62400# 1.23fF
C7988 VN.n7178 a_400_62400# 0.59fF
C7989 VN.n7179 a_400_62400# 2.51fF
C7990 VN.n7180 a_400_62400# 0.16fF
C7991 VN.t1394 a_400_62400# 0.03fF
C7992 VN.n7181 a_400_62400# 0.19fF
C7993 VN.t2516 a_400_62400# 0.03fF
C7994 VN.n7183 a_400_62400# 0.32fF
C7995 VN.n7184 a_400_62400# 0.48fF
C7996 VN.n7185 a_400_62400# 0.81fF
C7997 VN.n7186 a_400_62400# 0.03fF
C7998 VN.n7187 a_400_62400# 0.01fF
C7999 VN.n7188 a_400_62400# 0.02fF
C8000 VN.n7189 a_400_62400# 0.11fF
C8001 VN.n7190 a_400_62400# 0.08fF
C8002 VN.n7191 a_400_62400# 0.04fF
C8003 VN.n7192 a_400_62400# 0.05fF
C8004 VN.n7193 a_400_62400# 1.34fF
C8005 VN.n7194 a_400_62400# 0.48fF
C8006 VN.n7195 a_400_62400# 2.51fF
C8007 VN.n7196 a_400_62400# 2.67fF
C8008 VN.t1112 a_400_62400# 0.03fF
C8009 VN.n7197 a_400_62400# 0.32fF
C8010 VN.n7198 a_400_62400# 1.22fF
C8011 VN.n7199 a_400_62400# 0.07fF
C8012 VN.t2067 a_400_62400# 0.03fF
C8013 VN.n7200 a_400_62400# 0.16fF
C8014 VN.n7201 a_400_62400# 0.19fF
C8015 VN.n7203 a_400_62400# 2.53fF
C8016 VN.n7204 a_400_62400# 0.09fF
C8017 VN.n7205 a_400_62400# 0.05fF
C8018 VN.n7206 a_400_62400# 0.07fF
C8019 VN.n7207 a_400_62400# 1.16fF
C8020 VN.n7208 a_400_62400# 0.01fF
C8021 VN.n7209 a_400_62400# 0.01fF
C8022 VN.n7210 a_400_62400# 0.01fF
C8023 VN.n7211 a_400_62400# 0.09fF
C8024 VN.n7212 a_400_62400# 0.91fF
C8025 VN.n7213 a_400_62400# 0.96fF
C8026 VN.t1654 a_400_62400# 0.03fF
C8027 VN.n7214 a_400_62400# 0.32fF
C8028 VN.n7215 a_400_62400# 0.48fF
C8029 VN.n7216 a_400_62400# 0.81fF
C8030 VN.n7217 a_400_62400# 0.16fF
C8031 VN.t529 a_400_62400# 0.03fF
C8032 VN.n7218 a_400_62400# 0.19fF
C8033 VN.n7220 a_400_62400# 0.93fF
C8034 VN.n7221 a_400_62400# 0.30fF
C8035 VN.n7222 a_400_62400# 0.34fF
C8036 VN.n7223 a_400_62400# 0.12fF
C8037 VN.n7224 a_400_62400# 0.30fF
C8038 VN.n7225 a_400_62400# 0.93fF
C8039 VN.n7226 a_400_62400# 1.55fF
C8040 VN.n7227 a_400_62400# 0.29fF
C8041 VN.n7228 a_400_62400# 0.34fF
C8042 VN.n7229 a_400_62400# 0.12fF
C8043 VN.n7230 a_400_62400# 3.10fF
C8044 VN.t248 a_400_62400# 0.03fF
C8045 VN.n7231 a_400_62400# 0.32fF
C8046 VN.n7232 a_400_62400# 1.22fF
C8047 VN.n7233 a_400_62400# 0.07fF
C8048 VN.t1328 a_400_62400# 0.03fF
C8049 VN.n7234 a_400_62400# 0.16fF
C8050 VN.n7235 a_400_62400# 0.19fF
C8051 VN.n7237 a_400_62400# 2.51fF
C8052 VN.n7238 a_400_62400# 0.61fF
C8053 VN.n7239 a_400_62400# 0.30fF
C8054 VN.n7240 a_400_62400# 0.51fF
C8055 VN.n7241 a_400_62400# 0.21fF
C8056 VN.n7242 a_400_62400# 0.38fF
C8057 VN.n7243 a_400_62400# 0.29fF
C8058 VN.n7244 a_400_62400# 0.40fF
C8059 VN.n7245 a_400_62400# 0.28fF
C8060 VN.t785 a_400_62400# 0.03fF
C8061 VN.n7246 a_400_62400# 0.32fF
C8062 VN.n7247 a_400_62400# 0.48fF
C8063 VN.n7248 a_400_62400# 0.81fF
C8064 VN.n7249 a_400_62400# 0.16fF
C8065 VN.t2184 a_400_62400# 0.03fF
C8066 VN.n7250 a_400_62400# 0.19fF
C8067 VN.n7252 a_400_62400# 0.06fF
C8068 VN.n7253 a_400_62400# 0.04fF
C8069 VN.n7254 a_400_62400# 0.04fF
C8070 VN.n7255 a_400_62400# 0.14fF
C8071 VN.n7256 a_400_62400# 0.48fF
C8072 VN.n7257 a_400_62400# 0.50fF
C8073 VN.n7258 a_400_62400# 0.14fF
C8074 VN.n7259 a_400_62400# 0.16fF
C8075 VN.n7260 a_400_62400# 0.09fF
C8076 VN.n7261 a_400_62400# 0.16fF
C8077 VN.n7262 a_400_62400# 0.24fF
C8078 VN.n7263 a_400_62400# 5.35fF
C8079 VN.t1897 a_400_62400# 0.03fF
C8080 VN.n7264 a_400_62400# 0.32fF
C8081 VN.n7265 a_400_62400# 1.22fF
C8082 VN.n7266 a_400_62400# 0.07fF
C8083 VN.t466 a_400_62400# 0.03fF
C8084 VN.n7267 a_400_62400# 0.16fF
C8085 VN.n7268 a_400_62400# 0.19fF
C8086 VN.n7270 a_400_62400# 0.33fF
C8087 VN.n7271 a_400_62400# 0.12fF
C8088 VN.n7272 a_400_62400# 0.28fF
C8089 VN.n7273 a_400_62400# 1.72fF
C8090 VN.n7274 a_400_62400# 0.71fF
C8091 VN.n7275 a_400_62400# 2.51fF
C8092 VN.n7276 a_400_62400# 0.16fF
C8093 VN.t1319 a_400_62400# 0.03fF
C8094 VN.n7277 a_400_62400# 0.19fF
C8095 VN.t2439 a_400_62400# 0.03fF
C8096 VN.n7279 a_400_62400# 0.32fF
C8097 VN.n7280 a_400_62400# 0.48fF
C8098 VN.n7281 a_400_62400# 0.81fF
C8099 VN.n7282 a_400_62400# 0.95fF
C8100 VN.n7283 a_400_62400# 2.11fF
C8101 VN.n7284 a_400_62400# 3.28fF
C8102 VN.t1022 a_400_62400# 0.03fF
C8103 VN.n7285 a_400_62400# 0.32fF
C8104 VN.n7286 a_400_62400# 1.22fF
C8105 VN.n7287 a_400_62400# 0.07fF
C8106 VN.t2116 a_400_62400# 0.03fF
C8107 VN.n7288 a_400_62400# 0.16fF
C8108 VN.n7289 a_400_62400# 0.19fF
C8109 VN.n7291 a_400_62400# 2.53fF
C8110 VN.n7292 a_400_62400# 0.08fF
C8111 VN.n7293 a_400_62400# 0.04fF
C8112 VN.n7294 a_400_62400# 0.05fF
C8113 VN.n7295 a_400_62400# 1.33fF
C8114 VN.n7296 a_400_62400# 0.03fF
C8115 VN.n7297 a_400_62400# 0.01fF
C8116 VN.n7298 a_400_62400# 0.02fF
C8117 VN.n7299 a_400_62400# 0.11fF
C8118 VN.n7300 a_400_62400# 0.48fF
C8119 VN.n7301 a_400_62400# 2.48fF
C8120 VN.t1576 a_400_62400# 0.03fF
C8121 VN.n7302 a_400_62400# 0.32fF
C8122 VN.n7303 a_400_62400# 0.48fF
C8123 VN.n7304 a_400_62400# 0.81fF
C8124 VN.n7305 a_400_62400# 0.16fF
C8125 VN.t456 a_400_62400# 0.03fF
C8126 VN.n7306 a_400_62400# 0.19fF
C8127 VN.n7308 a_400_62400# 0.93fF
C8128 VN.n7309 a_400_62400# 0.30fF
C8129 VN.n7310 a_400_62400# 0.34fF
C8130 VN.n7311 a_400_62400# 0.12fF
C8131 VN.n7312 a_400_62400# 0.30fF
C8132 VN.n7313 a_400_62400# 0.93fF
C8133 VN.n7314 a_400_62400# 1.55fF
C8134 VN.n7315 a_400_62400# 0.29fF
C8135 VN.n7316 a_400_62400# 0.34fF
C8136 VN.n7317 a_400_62400# 0.12fF
C8137 VN.n7318 a_400_62400# 2.52fF
C8138 VN.t150 a_400_62400# 0.03fF
C8139 VN.n7319 a_400_62400# 0.32fF
C8140 VN.n7320 a_400_62400# 1.22fF
C8141 VN.n7321 a_400_62400# 0.07fF
C8142 VN.t1239 a_400_62400# 0.03fF
C8143 VN.n7322 a_400_62400# 0.16fF
C8144 VN.n7323 a_400_62400# 0.19fF
C8145 VN.n7325 a_400_62400# 27.83fF
C8146 VN.t1219 a_400_62400# 0.03fF
C8147 VN.n7326 a_400_62400# 0.32fF
C8148 VN.n7327 a_400_62400# 1.22fF
C8149 VN.t76 a_400_62400# 66.88fF
C8150 VN.t1033 a_400_62400# 0.03fF
C8151 VN.n7328 a_400_62400# 1.60fF
C8152 VN.n7329 a_400_62400# 0.07fF
C8153 VN.t1652 a_400_62400# 0.03fF
C8154 VN.n7330 a_400_62400# 0.02fF
C8155 VN.n7331 a_400_62400# 0.34fF
C8156 VN.n7333 a_400_62400# 2.01fF
C8157 VN.n7334 a_400_62400# 1.75fF
C8158 VN.n7335 a_400_62400# 0.37fF
C8159 VN.n7336 a_400_62400# 0.33fF
C8160 VN.n7337 a_400_62400# 5.88fF
C8161 VN.n7338 a_400_62400# 0.02fF
C8162 VN.n7339 a_400_62400# 0.02fF
C8163 VN.n7340 a_400_62400# 0.03fF
C8164 VN.n7341 a_400_62400# 0.05fF
C8165 VN.n7342 a_400_62400# 0.23fF
C8166 VN.n7343 a_400_62400# 0.02fF
C8167 VN.n7344 a_400_62400# 0.03fF
C8168 VN.n7345 a_400_62400# 0.01fF
C8169 VN.n7346 a_400_62400# 0.01fF
C8170 VN.n7347 a_400_62400# 0.01fF
C8171 VN.n7348 a_400_62400# 0.02fF
C8172 VN.n7349 a_400_62400# 0.03fF
C8173 VN.n7350 a_400_62400# 0.06fF
C8174 VN.n7351 a_400_62400# 0.05fF
C8175 VN.n7352 a_400_62400# 0.15fF
C8176 VN.n7353 a_400_62400# 0.51fF
C8177 VN.n7354 a_400_62400# 0.27fF
C8178 VN.n7355 a_400_62400# 37.46fF
C8179 VN.n7356 a_400_62400# 37.46fF
C8180 VN.n7357 a_400_62400# 0.79fF
C8181 VN.n7358 a_400_62400# 0.23fF
C8182 VN.n7359 a_400_62400# 1.18fF
C8183 VN.t22 a_400_62400# 28.64fF
C8184 VN.n7360 a_400_62400# 0.79fF
C8185 VN.n7361 a_400_62400# 0.11fF
C8186 VN.n7362 a_400_62400# 4.98fF
C8187 VN.n7363 a_400_62400# 0.80fF
C8188 VN.n7364 a_400_62400# 0.29fF
C8189 VN.n7365 a_400_62400# 1.96fF
C8190 VN.n7367 a_400_62400# 25.18fF
C8191 VN.n7369 a_400_62400# 1.87fF
C8192 VN.n7370 a_400_62400# 5.36fF
C8193 VN.n7371 a_400_62400# 1.81fF
C8194 VN.t321 a_400_62400# 0.03fF
C8195 VN.n7372 a_400_62400# 0.85fF
C8196 VN.n7373 a_400_62400# 0.81fF
C8197 VN.n7374 a_400_62400# 0.33fF
C8198 VN.n7375 a_400_62400# 0.12fF
C8199 VN.n7376 a_400_62400# 0.28fF
C8200 VN.n7377 a_400_62400# 1.72fF
C8201 VN.n7378 a_400_62400# 0.71fF
C8202 VN.n7379 a_400_62400# 2.51fF
C8203 VN.n7380 a_400_62400# 0.16fF
C8204 VN.t2155 a_400_62400# 0.03fF
C8205 VN.n7381 a_400_62400# 0.19fF
C8206 VN.t636 a_400_62400# 0.03fF
C8207 VN.n7383 a_400_62400# 0.32fF
C8208 VN.n7384 a_400_62400# 0.48fF
C8209 VN.n7385 a_400_62400# 0.81fF
C8210 VN.n7386 a_400_62400# 0.03fF
C8211 VN.n7387 a_400_62400# 0.01fF
C8212 VN.n7388 a_400_62400# 0.02fF
C8213 VN.n7389 a_400_62400# 0.11fF
C8214 VN.n7390 a_400_62400# 0.08fF
C8215 VN.n7391 a_400_62400# 0.04fF
C8216 VN.n7392 a_400_62400# 0.05fF
C8217 VN.n7393 a_400_62400# 1.34fF
C8218 VN.n7394 a_400_62400# 0.48fF
C8219 VN.n7395 a_400_62400# 2.51fF
C8220 VN.n7396 a_400_62400# 2.67fF
C8221 VN.t1739 a_400_62400# 0.03fF
C8222 VN.n7397 a_400_62400# 0.32fF
C8223 VN.n7398 a_400_62400# 1.22fF
C8224 VN.n7399 a_400_62400# 0.07fF
C8225 VN.t293 a_400_62400# 0.03fF
C8226 VN.n7400 a_400_62400# 0.16fF
C8227 VN.n7401 a_400_62400# 0.19fF
C8228 VN.n7403 a_400_62400# 2.53fF
C8229 VN.n7404 a_400_62400# 0.08fF
C8230 VN.n7405 a_400_62400# 0.04fF
C8231 VN.n7406 a_400_62400# 0.05fF
C8232 VN.n7407 a_400_62400# 1.33fF
C8233 VN.n7408 a_400_62400# 0.03fF
C8234 VN.n7409 a_400_62400# 0.01fF
C8235 VN.n7410 a_400_62400# 0.02fF
C8236 VN.n7411 a_400_62400# 0.11fF
C8237 VN.n7412 a_400_62400# 0.48fF
C8238 VN.n7413 a_400_62400# 2.48fF
C8239 VN.t2409 a_400_62400# 0.03fF
C8240 VN.n7414 a_400_62400# 0.32fF
C8241 VN.n7415 a_400_62400# 0.48fF
C8242 VN.n7416 a_400_62400# 0.81fF
C8243 VN.n7417 a_400_62400# 0.16fF
C8244 VN.t1287 a_400_62400# 0.03fF
C8245 VN.n7418 a_400_62400# 0.19fF
C8246 VN.n7420 a_400_62400# 0.93fF
C8247 VN.n7421 a_400_62400# 0.30fF
C8248 VN.n7422 a_400_62400# 0.34fF
C8249 VN.n7423 a_400_62400# 0.12fF
C8250 VN.n7424 a_400_62400# 0.30fF
C8251 VN.n7425 a_400_62400# 0.93fF
C8252 VN.n7426 a_400_62400# 1.55fF
C8253 VN.n7427 a_400_62400# 0.29fF
C8254 VN.n7428 a_400_62400# 0.34fF
C8255 VN.n7429 a_400_62400# 0.12fF
C8256 VN.n7430 a_400_62400# 2.52fF
C8257 VN.t999 a_400_62400# 0.03fF
C8258 VN.n7431 a_400_62400# 0.32fF
C8259 VN.n7432 a_400_62400# 1.22fF
C8260 VN.n7433 a_400_62400# 0.07fF
C8261 VN.t1944 a_400_62400# 0.03fF
C8262 VN.n7434 a_400_62400# 0.16fF
C8263 VN.n7435 a_400_62400# 0.19fF
C8264 VN.n7437 a_400_62400# 0.33fF
C8265 VN.n7438 a_400_62400# 0.12fF
C8266 VN.n7439 a_400_62400# 0.28fF
C8267 VN.n7440 a_400_62400# 1.23fF
C8268 VN.n7441 a_400_62400# 0.59fF
C8269 VN.n7442 a_400_62400# 2.51fF
C8270 VN.n7443 a_400_62400# 0.16fF
C8271 VN.t420 a_400_62400# 0.03fF
C8272 VN.n7444 a_400_62400# 0.19fF
C8273 VN.t1544 a_400_62400# 0.03fF
C8274 VN.n7446 a_400_62400# 0.32fF
C8275 VN.n7447 a_400_62400# 0.48fF
C8276 VN.n7448 a_400_62400# 0.81fF
C8277 VN.n7449 a_400_62400# 0.03fF
C8278 VN.n7450 a_400_62400# 0.01fF
C8279 VN.n7451 a_400_62400# 0.02fF
C8280 VN.n7452 a_400_62400# 0.11fF
C8281 VN.n7453 a_400_62400# 0.08fF
C8282 VN.n7454 a_400_62400# 0.04fF
C8283 VN.n7455 a_400_62400# 0.05fF
C8284 VN.n7456 a_400_62400# 1.34fF
C8285 VN.n7457 a_400_62400# 0.48fF
C8286 VN.n7458 a_400_62400# 2.51fF
C8287 VN.n7459 a_400_62400# 2.67fF
C8288 VN.t118 a_400_62400# 0.03fF
C8289 VN.n7460 a_400_62400# 0.32fF
C8290 VN.n7461 a_400_62400# 1.22fF
C8291 VN.n7462 a_400_62400# 0.07fF
C8292 VN.t1074 a_400_62400# 0.03fF
C8293 VN.n7463 a_400_62400# 0.16fF
C8294 VN.n7464 a_400_62400# 0.19fF
C8295 VN.n7466 a_400_62400# 2.53fF
C8296 VN.n7467 a_400_62400# 0.08fF
C8297 VN.n7468 a_400_62400# 0.04fF
C8298 VN.n7469 a_400_62400# 0.05fF
C8299 VN.n7470 a_400_62400# 1.33fF
C8300 VN.n7471 a_400_62400# 0.03fF
C8301 VN.n7472 a_400_62400# 0.01fF
C8302 VN.n7473 a_400_62400# 0.02fF
C8303 VN.n7474 a_400_62400# 0.11fF
C8304 VN.n7475 a_400_62400# 0.48fF
C8305 VN.n7476 a_400_62400# 2.48fF
C8306 VN.t2029 a_400_62400# 0.03fF
C8307 VN.n7477 a_400_62400# 0.32fF
C8308 VN.n7478 a_400_62400# 0.48fF
C8309 VN.n7479 a_400_62400# 0.81fF
C8310 VN.n7480 a_400_62400# 0.16fF
C8311 VN.t866 a_400_62400# 0.03fF
C8312 VN.n7481 a_400_62400# 0.19fF
C8313 VN.n7483 a_400_62400# 0.93fF
C8314 VN.n7484 a_400_62400# 0.30fF
C8315 VN.n7485 a_400_62400# 0.34fF
C8316 VN.n7486 a_400_62400# 0.12fF
C8317 VN.n7487 a_400_62400# 0.30fF
C8318 VN.n7488 a_400_62400# 0.93fF
C8319 VN.n7489 a_400_62400# 1.55fF
C8320 VN.n7490 a_400_62400# 0.29fF
C8321 VN.n7491 a_400_62400# 0.34fF
C8322 VN.n7492 a_400_62400# 0.12fF
C8323 VN.n7493 a_400_62400# 2.52fF
C8324 VN.t626 a_400_62400# 0.03fF
C8325 VN.n7494 a_400_62400# 0.32fF
C8326 VN.n7495 a_400_62400# 1.22fF
C8327 VN.n7496 a_400_62400# 0.07fF
C8328 VN.t199 a_400_62400# 0.03fF
C8329 VN.n7497 a_400_62400# 0.16fF
C8330 VN.n7498 a_400_62400# 0.19fF
C8331 VN.n7500 a_400_62400# 0.33fF
C8332 VN.n7501 a_400_62400# 0.12fF
C8333 VN.n7502 a_400_62400# 0.28fF
C8334 VN.n7503 a_400_62400# 1.23fF
C8335 VN.n7504 a_400_62400# 0.59fF
C8336 VN.n7505 a_400_62400# 2.51fF
C8337 VN.n7506 a_400_62400# 0.16fF
C8338 VN.t2530 a_400_62400# 0.03fF
C8339 VN.n7507 a_400_62400# 0.19fF
C8340 VN.t1155 a_400_62400# 0.03fF
C8341 VN.n7509 a_400_62400# 0.32fF
C8342 VN.n7510 a_400_62400# 0.48fF
C8343 VN.n7511 a_400_62400# 0.81fF
C8344 VN.n7512 a_400_62400# 0.03fF
C8345 VN.n7513 a_400_62400# 0.01fF
C8346 VN.n7514 a_400_62400# 0.02fF
C8347 VN.n7515 a_400_62400# 0.11fF
C8348 VN.n7516 a_400_62400# 0.08fF
C8349 VN.n7517 a_400_62400# 0.04fF
C8350 VN.n7518 a_400_62400# 0.05fF
C8351 VN.n7519 a_400_62400# 1.34fF
C8352 VN.n7520 a_400_62400# 0.48fF
C8353 VN.n7521 a_400_62400# 2.51fF
C8354 VN.n7522 a_400_62400# 2.67fF
C8355 VN.t2278 a_400_62400# 0.03fF
C8356 VN.n7523 a_400_62400# 0.32fF
C8357 VN.n7524 a_400_62400# 1.22fF
C8358 VN.n7525 a_400_62400# 0.07fF
C8359 VN.t689 a_400_62400# 0.03fF
C8360 VN.n7526 a_400_62400# 0.16fF
C8361 VN.n7527 a_400_62400# 0.19fF
C8362 VN.n7529 a_400_62400# 2.53fF
C8363 VN.n7530 a_400_62400# 0.08fF
C8364 VN.n7531 a_400_62400# 0.04fF
C8365 VN.n7532 a_400_62400# 0.05fF
C8366 VN.n7533 a_400_62400# 1.33fF
C8367 VN.n7534 a_400_62400# 0.03fF
C8368 VN.n7535 a_400_62400# 0.01fF
C8369 VN.n7536 a_400_62400# 0.02fF
C8370 VN.n7537 a_400_62400# 0.11fF
C8371 VN.n7538 a_400_62400# 0.48fF
C8372 VN.n7539 a_400_62400# 2.48fF
C8373 VN.t287 a_400_62400# 0.03fF
C8374 VN.n7540 a_400_62400# 0.32fF
C8375 VN.n7541 a_400_62400# 0.48fF
C8376 VN.n7542 a_400_62400# 0.81fF
C8377 VN.n7543 a_400_62400# 0.16fF
C8378 VN.t1666 a_400_62400# 0.03fF
C8379 VN.n7544 a_400_62400# 0.19fF
C8380 VN.n7546 a_400_62400# 0.93fF
C8381 VN.n7547 a_400_62400# 0.30fF
C8382 VN.n7548 a_400_62400# 0.34fF
C8383 VN.n7549 a_400_62400# 0.12fF
C8384 VN.n7550 a_400_62400# 0.30fF
C8385 VN.n7551 a_400_62400# 0.93fF
C8386 VN.n7552 a_400_62400# 1.55fF
C8387 VN.n7553 a_400_62400# 0.29fF
C8388 VN.n7554 a_400_62400# 0.34fF
C8389 VN.n7555 a_400_62400# 0.12fF
C8390 VN.n7556 a_400_62400# 2.52fF
C8391 VN.t1409 a_400_62400# 0.03fF
C8392 VN.n7557 a_400_62400# 0.32fF
C8393 VN.n7558 a_400_62400# 1.22fF
C8394 VN.n7559 a_400_62400# 0.07fF
C8395 VN.t2349 a_400_62400# 0.03fF
C8396 VN.n7560 a_400_62400# 0.16fF
C8397 VN.n7561 a_400_62400# 0.19fF
C8398 VN.n7563 a_400_62400# 0.33fF
C8399 VN.n7564 a_400_62400# 0.12fF
C8400 VN.n7565 a_400_62400# 0.28fF
C8401 VN.n7566 a_400_62400# 1.23fF
C8402 VN.n7567 a_400_62400# 0.59fF
C8403 VN.n7568 a_400_62400# 2.51fF
C8404 VN.n7569 a_400_62400# 0.16fF
C8405 VN.t798 a_400_62400# 0.03fF
C8406 VN.n7570 a_400_62400# 0.19fF
C8407 VN.t1939 a_400_62400# 0.03fF
C8408 VN.n7572 a_400_62400# 0.32fF
C8409 VN.n7573 a_400_62400# 0.48fF
C8410 VN.n7574 a_400_62400# 0.81fF
C8411 VN.n7575 a_400_62400# 0.03fF
C8412 VN.n7576 a_400_62400# 0.01fF
C8413 VN.n7577 a_400_62400# 0.02fF
C8414 VN.n7578 a_400_62400# 0.11fF
C8415 VN.n7579 a_400_62400# 0.08fF
C8416 VN.n7580 a_400_62400# 0.04fF
C8417 VN.n7581 a_400_62400# 0.05fF
C8418 VN.n7582 a_400_62400# 1.34fF
C8419 VN.n7583 a_400_62400# 0.48fF
C8420 VN.n7584 a_400_62400# 2.51fF
C8421 VN.n7585 a_400_62400# 2.67fF
C8422 VN.t549 a_400_62400# 0.03fF
C8423 VN.n7586 a_400_62400# 0.32fF
C8424 VN.n7587 a_400_62400# 1.22fF
C8425 VN.n7588 a_400_62400# 0.07fF
C8426 VN.t1601 a_400_62400# 0.03fF
C8427 VN.n7589 a_400_62400# 0.16fF
C8428 VN.n7590 a_400_62400# 0.19fF
C8429 VN.n7592 a_400_62400# 2.53fF
C8430 VN.n7593 a_400_62400# 0.09fF
C8431 VN.n7594 a_400_62400# 0.05fF
C8432 VN.n7595 a_400_62400# 0.07fF
C8433 VN.n7596 a_400_62400# 1.16fF
C8434 VN.n7597 a_400_62400# 0.01fF
C8435 VN.n7598 a_400_62400# 0.01fF
C8436 VN.n7599 a_400_62400# 0.01fF
C8437 VN.n7600 a_400_62400# 0.09fF
C8438 VN.n7601 a_400_62400# 0.91fF
C8439 VN.n7602 a_400_62400# 0.96fF
C8440 VN.t1068 a_400_62400# 0.03fF
C8441 VN.n7603 a_400_62400# 0.32fF
C8442 VN.n7604 a_400_62400# 0.48fF
C8443 VN.n7605 a_400_62400# 0.81fF
C8444 VN.n7606 a_400_62400# 0.16fF
C8445 VN.t2453 a_400_62400# 0.03fF
C8446 VN.n7607 a_400_62400# 0.19fF
C8447 VN.n7609 a_400_62400# 0.93fF
C8448 VN.n7610 a_400_62400# 0.30fF
C8449 VN.n7611 a_400_62400# 0.34fF
C8450 VN.n7612 a_400_62400# 0.12fF
C8451 VN.n7613 a_400_62400# 0.30fF
C8452 VN.n7614 a_400_62400# 0.93fF
C8453 VN.n7615 a_400_62400# 1.55fF
C8454 VN.n7616 a_400_62400# 0.29fF
C8455 VN.n7617 a_400_62400# 0.34fF
C8456 VN.n7618 a_400_62400# 0.12fF
C8457 VN.n7619 a_400_62400# 3.10fF
C8458 VN.t2204 a_400_62400# 0.03fF
C8459 VN.n7620 a_400_62400# 0.32fF
C8460 VN.n7621 a_400_62400# 1.22fF
C8461 VN.n7622 a_400_62400# 0.07fF
C8462 VN.t736 a_400_62400# 0.03fF
C8463 VN.n7623 a_400_62400# 0.16fF
C8464 VN.n7624 a_400_62400# 0.19fF
C8465 VN.n7626 a_400_62400# 2.51fF
C8466 VN.n7627 a_400_62400# 0.61fF
C8467 VN.n7628 a_400_62400# 0.30fF
C8468 VN.n7629 a_400_62400# 0.51fF
C8469 VN.n7630 a_400_62400# 0.21fF
C8470 VN.n7631 a_400_62400# 0.38fF
C8471 VN.n7632 a_400_62400# 0.29fF
C8472 VN.n7633 a_400_62400# 0.40fF
C8473 VN.n7634 a_400_62400# 0.28fF
C8474 VN.t194 a_400_62400# 0.03fF
C8475 VN.n7635 a_400_62400# 0.32fF
C8476 VN.n7636 a_400_62400# 0.48fF
C8477 VN.n7637 a_400_62400# 0.81fF
C8478 VN.n7638 a_400_62400# 0.16fF
C8479 VN.t1591 a_400_62400# 0.03fF
C8480 VN.n7639 a_400_62400# 0.19fF
C8481 VN.n7641 a_400_62400# 0.06fF
C8482 VN.n7642 a_400_62400# 0.04fF
C8483 VN.n7643 a_400_62400# 0.04fF
C8484 VN.n7644 a_400_62400# 0.14fF
C8485 VN.n7645 a_400_62400# 0.48fF
C8486 VN.n7646 a_400_62400# 0.50fF
C8487 VN.n7647 a_400_62400# 0.14fF
C8488 VN.n7648 a_400_62400# 0.16fF
C8489 VN.n7649 a_400_62400# 0.09fF
C8490 VN.n7650 a_400_62400# 0.16fF
C8491 VN.n7651 a_400_62400# 0.24fF
C8492 VN.n7652 a_400_62400# 5.35fF
C8493 VN.t1336 a_400_62400# 0.03fF
C8494 VN.n7653 a_400_62400# 0.32fF
C8495 VN.n7654 a_400_62400# 1.22fF
C8496 VN.n7655 a_400_62400# 0.07fF
C8497 VN.t2392 a_400_62400# 0.03fF
C8498 VN.n7656 a_400_62400# 0.16fF
C8499 VN.n7657 a_400_62400# 0.19fF
C8500 VN.n7659 a_400_62400# 0.33fF
C8501 VN.n7660 a_400_62400# 0.12fF
C8502 VN.n7661 a_400_62400# 0.28fF
C8503 VN.n7662 a_400_62400# 1.72fF
C8504 VN.n7663 a_400_62400# 0.71fF
C8505 VN.n7664 a_400_62400# 2.51fF
C8506 VN.n7665 a_400_62400# 0.16fF
C8507 VN.t724 a_400_62400# 0.03fF
C8508 VN.n7666 a_400_62400# 0.19fF
C8509 VN.t1850 a_400_62400# 0.03fF
C8510 VN.n7668 a_400_62400# 0.32fF
C8511 VN.n7669 a_400_62400# 0.48fF
C8512 VN.n7670 a_400_62400# 0.81fF
C8513 VN.n7671 a_400_62400# 0.95fF
C8514 VN.n7672 a_400_62400# 2.11fF
C8515 VN.n7673 a_400_62400# 3.28fF
C8516 VN.t472 a_400_62400# 0.03fF
C8517 VN.n7674 a_400_62400# 0.32fF
C8518 VN.n7675 a_400_62400# 1.22fF
C8519 VN.n7676 a_400_62400# 0.07fF
C8520 VN.t1524 a_400_62400# 0.03fF
C8521 VN.n7677 a_400_62400# 0.16fF
C8522 VN.n7678 a_400_62400# 0.19fF
C8523 VN.n7680 a_400_62400# 2.53fF
C8524 VN.n7681 a_400_62400# 0.08fF
C8525 VN.n7682 a_400_62400# 0.04fF
C8526 VN.n7683 a_400_62400# 0.05fF
C8527 VN.n7684 a_400_62400# 1.33fF
C8528 VN.n7685 a_400_62400# 0.03fF
C8529 VN.n7686 a_400_62400# 0.01fF
C8530 VN.n7687 a_400_62400# 0.02fF
C8531 VN.n7688 a_400_62400# 0.11fF
C8532 VN.n7689 a_400_62400# 0.48fF
C8533 VN.n7690 a_400_62400# 2.48fF
C8534 VN.t978 a_400_62400# 0.03fF
C8535 VN.n7691 a_400_62400# 0.32fF
C8536 VN.n7692 a_400_62400# 0.48fF
C8537 VN.n7693 a_400_62400# 0.81fF
C8538 VN.n7694 a_400_62400# 0.16fF
C8539 VN.t2496 a_400_62400# 0.03fF
C8540 VN.n7695 a_400_62400# 0.19fF
C8541 VN.n7697 a_400_62400# 0.93fF
C8542 VN.n7698 a_400_62400# 0.30fF
C8543 VN.n7699 a_400_62400# 0.34fF
C8544 VN.n7700 a_400_62400# 0.12fF
C8545 VN.n7701 a_400_62400# 0.30fF
C8546 VN.n7702 a_400_62400# 0.93fF
C8547 VN.n7703 a_400_62400# 1.55fF
C8548 VN.n7704 a_400_62400# 0.29fF
C8549 VN.n7705 a_400_62400# 0.34fF
C8550 VN.n7706 a_400_62400# 0.12fF
C8551 VN.n7707 a_400_62400# 2.52fF
C8552 VN.t2125 a_400_62400# 0.03fF
C8553 VN.n7708 a_400_62400# 0.32fF
C8554 VN.n7709 a_400_62400# 1.22fF
C8555 VN.n7710 a_400_62400# 0.07fF
C8556 VN.t654 a_400_62400# 0.03fF
C8557 VN.n7711 a_400_62400# 0.16fF
C8558 VN.n7712 a_400_62400# 0.19fF
C8559 VN.n7714 a_400_62400# 27.83fF
C8560 VN.n7715 a_400_62400# 2.30fF
C8561 VN.n7716 a_400_62400# 4.08fF
C8562 VN.t1503 a_400_62400# 0.03fF
C8563 VN.n7717 a_400_62400# 0.32fF
C8564 VN.n7718 a_400_62400# 0.48fF
C8565 VN.n7719 a_400_62400# 0.81fF
C8566 VN.n7720 a_400_62400# 0.16fF
C8567 VN.t368 a_400_62400# 0.03fF
C8568 VN.n7721 a_400_62400# 0.19fF
C8569 VN.n7723 a_400_62400# 0.42fF
C8570 VN.n7724 a_400_62400# 0.34fF
C8571 VN.n7725 a_400_62400# 0.12fF
C8572 VN.n7726 a_400_62400# 0.30fF
C8573 VN.n7727 a_400_62400# 0.88fF
C8574 VN.n7728 a_400_62400# 1.28fF
C8575 VN.n7729 a_400_62400# 0.30fF
C8576 VN.n7730 a_400_62400# 0.28fF
C8577 VN.n7731 a_400_62400# 0.27fF
C8578 VN.n7732 a_400_62400# 0.09fF
C8579 VN.n7733 a_400_62400# 0.12fF
C8580 VN.n7734 a_400_62400# 0.13fF
C8581 VN.n7735 a_400_62400# 2.66fF
C8582 VN.t1161 a_400_62400# 0.03fF
C8583 VN.n7736 a_400_62400# 0.16fF
C8584 VN.n7737 a_400_62400# 0.19fF
C8585 VN.t31 a_400_62400# 0.03fF
C8586 VN.n7739 a_400_62400# 0.32fF
C8587 VN.n7740 a_400_62400# 1.22fF
C8588 VN.n7741 a_400_62400# 0.07fF
C8589 VN.n7742 a_400_62400# 2.51fF
C8590 VN.n7743 a_400_62400# 0.16fF
C8591 VN.t1633 a_400_62400# 0.03fF
C8592 VN.n7744 a_400_62400# 0.19fF
C8593 VN.t245 a_400_62400# 0.03fF
C8594 VN.n7746 a_400_62400# 0.32fF
C8595 VN.n7747 a_400_62400# 0.48fF
C8596 VN.n7748 a_400_62400# 0.81fF
C8597 VN.n7749 a_400_62400# 1.24fF
C8598 VN.n7750 a_400_62400# 0.43fF
C8599 VN.n7751 a_400_62400# 0.43fF
C8600 VN.n7752 a_400_62400# 1.24fF
C8601 VN.n7753 a_400_62400# 1.46fF
C8602 VN.n7754 a_400_62400# 0.21fF
C8603 VN.n7755 a_400_62400# 6.64fF
C8604 VN.t2313 a_400_62400# 0.03fF
C8605 VN.n7756 a_400_62400# 0.16fF
C8606 VN.n7757 a_400_62400# 0.19fF
C8607 VN.t1381 a_400_62400# 0.03fF
C8608 VN.n7759 a_400_62400# 0.32fF
C8609 VN.n7760 a_400_62400# 1.22fF
C8610 VN.n7761 a_400_62400# 0.07fF
C8611 VN.n7762 a_400_62400# 2.51fF
C8612 VN.n7763 a_400_62400# 3.57fF
C8613 VN.t1281 a_400_62400# 0.03fF
C8614 VN.n7764 a_400_62400# 0.32fF
C8615 VN.n7765 a_400_62400# 0.48fF
C8616 VN.n7766 a_400_62400# 0.81fF
C8617 VN.n7767 a_400_62400# 0.16fF
C8618 VN.t81 a_400_62400# 0.03fF
C8619 VN.n7768 a_400_62400# 0.19fF
C8620 VN.n7770 a_400_62400# 6.91fF
C8621 VN.t1443 a_400_62400# 0.03fF
C8622 VN.n7771 a_400_62400# 0.16fF
C8623 VN.n7772 a_400_62400# 0.19fF
C8624 VN.t318 a_400_62400# 0.03fF
C8625 VN.n7774 a_400_62400# 0.32fF
C8626 VN.n7775 a_400_62400# 1.22fF
C8627 VN.n7776 a_400_62400# 0.07fF
C8628 VN.n7777 a_400_62400# 2.51fF
C8629 VN.n7778 a_400_62400# 3.57fF
C8630 VN.t415 a_400_62400# 0.03fF
C8631 VN.n7779 a_400_62400# 0.32fF
C8632 VN.n7780 a_400_62400# 0.48fF
C8633 VN.n7781 a_400_62400# 0.81fF
C8634 VN.n7782 a_400_62400# 0.16fF
C8635 VN.t1763 a_400_62400# 0.03fF
C8636 VN.n7783 a_400_62400# 0.19fF
C8637 VN.n7785 a_400_62400# 6.92fF
C8638 VN.t2445 a_400_62400# 0.03fF
C8639 VN.n7786 a_400_62400# 0.16fF
C8640 VN.n7787 a_400_62400# 0.19fF
C8641 VN.t1967 a_400_62400# 0.03fF
C8642 VN.n7789 a_400_62400# 0.32fF
C8643 VN.n7790 a_400_62400# 1.22fF
C8644 VN.n7791 a_400_62400# 0.07fF
C8645 VN.n7792 a_400_62400# 2.51fF
C8646 VN.n7793 a_400_62400# 3.57fF
C8647 VN.t2063 a_400_62400# 0.03fF
C8648 VN.n7794 a_400_62400# 0.32fF
C8649 VN.n7795 a_400_62400# 0.48fF
C8650 VN.n7796 a_400_62400# 0.81fF
C8651 VN.n7797 a_400_62400# 0.16fF
C8652 VN.t891 a_400_62400# 0.03fF
C8653 VN.n7798 a_400_62400# 0.19fF
C8654 VN.n7800 a_400_62400# 2.51fF
C8655 VN.n7801 a_400_62400# 3.59fF
C8656 VN.t893 a_400_62400# 0.03fF
C8657 VN.n7802 a_400_62400# 0.32fF
C8658 VN.n7803 a_400_62400# 0.48fF
C8659 VN.n7804 a_400_62400# 0.81fF
C8660 VN.t881 a_400_62400# 0.03fF
C8661 VN.n7805 a_400_62400# 1.63fF
C8662 VN.n7806 a_400_62400# 0.49fF
C8663 VN.n7807 a_400_62400# 1.64fF
C8664 VN.n7808 a_400_62400# 0.81fF
C8665 VN.n7809 a_400_62400# 1.21fF
C8666 VN.n7810 a_400_62400# 1.54fF
C8667 VN.n7811 a_400_62400# 4.06fF
C8668 VN.t30 a_400_62400# 28.64fF
C8669 VN.n7812 a_400_62400# 28.43fF
C8670 VN.n7814 a_400_62400# 0.50fF
C8671 VN.n7815 a_400_62400# 0.31fF
C8672 VN.n7816 a_400_62400# 3.74fF
C8673 VN.n7817 a_400_62400# 3.29fF
C8674 VN.n7818 a_400_62400# 5.35fF
C8675 VN.n7819 a_400_62400# 0.34fF
C8676 VN.n7820 a_400_62400# 0.02fF
C8677 VN.t2283 a_400_62400# 0.03fF
C8678 VN.n7821 a_400_62400# 0.34fF
C8679 VN.t2576 a_400_62400# 0.03fF
C8680 VN.n7822 a_400_62400# 1.28fF
C8681 VN.n7823 a_400_62400# 0.94fF
C8682 VN.n7824 a_400_62400# 2.53fF
C8683 VN.n7825 a_400_62400# 2.51fF
C8684 VN.t2541 a_400_62400# 0.03fF
C8685 VN.n7826 a_400_62400# 0.32fF
C8686 VN.n7827 a_400_62400# 0.48fF
C8687 VN.n7828 a_400_62400# 0.81fF
C8688 VN.n7829 a_400_62400# 0.16fF
C8689 VN.t1414 a_400_62400# 0.03fF
C8690 VN.n7830 a_400_62400# 0.19fF
C8691 VN.n7832 a_400_62400# 1.55fF
C8692 VN.n7833 a_400_62400# 0.29fF
C8693 VN.n7834 a_400_62400# 2.52fF
C8694 VN.t1705 a_400_62400# 0.03fF
C8695 VN.n7835 a_400_62400# 0.32fF
C8696 VN.n7836 a_400_62400# 1.22fF
C8697 VN.n7837 a_400_62400# 0.07fF
C8698 VN.t1483 a_400_62400# 0.03fF
C8699 VN.n7838 a_400_62400# 0.16fF
C8700 VN.n7839 a_400_62400# 0.19fF
C8701 VN.n7841 a_400_62400# 1.05fF
C8702 VN.n7842 a_400_62400# 3.07fF
C8703 VN.n7843 a_400_62400# 2.51fF
C8704 VN.n7844 a_400_62400# 0.16fF
C8705 VN.t552 a_400_62400# 0.03fF
C8706 VN.n7845 a_400_62400# 0.19fF
C8707 VN.t1676 a_400_62400# 0.03fF
C8708 VN.n7847 a_400_62400# 0.32fF
C8709 VN.n7848 a_400_62400# 0.48fF
C8710 VN.n7849 a_400_62400# 0.81fF
C8711 VN.n7850 a_400_62400# 2.46fF
C8712 VN.n7851 a_400_62400# 2.91fF
C8713 VN.t833 a_400_62400# 0.03fF
C8714 VN.n7852 a_400_62400# 0.32fF
C8715 VN.n7853 a_400_62400# 1.22fF
C8716 VN.n7854 a_400_62400# 0.07fF
C8717 VN.t738 a_400_62400# 0.03fF
C8718 VN.n7855 a_400_62400# 0.16fF
C8719 VN.n7856 a_400_62400# 0.19fF
C8720 VN.n7858 a_400_62400# 2.53fF
C8721 VN.n7859 a_400_62400# 2.51fF
C8722 VN.t810 a_400_62400# 0.03fF
C8723 VN.n7860 a_400_62400# 0.32fF
C8724 VN.n7861 a_400_62400# 0.48fF
C8725 VN.n7862 a_400_62400# 0.81fF
C8726 VN.n7863 a_400_62400# 0.16fF
C8727 VN.t2208 a_400_62400# 0.03fF
C8728 VN.n7864 a_400_62400# 0.19fF
C8729 VN.n7866 a_400_62400# 1.55fF
C8730 VN.n7867 a_400_62400# 0.29fF
C8731 VN.n7868 a_400_62400# 2.52fF
C8732 VN.t2498 a_400_62400# 0.03fF
C8733 VN.n7869 a_400_62400# 0.32fF
C8734 VN.n7870 a_400_62400# 1.22fF
C8735 VN.n7871 a_400_62400# 0.07fF
C8736 VN.t2395 a_400_62400# 0.03fF
C8737 VN.n7872 a_400_62400# 0.16fF
C8738 VN.n7873 a_400_62400# 0.19fF
C8739 VN.n7875 a_400_62400# 1.04fF
C8740 VN.n7876 a_400_62400# 2.60fF
C8741 VN.n7877 a_400_62400# 2.51fF
C8742 VN.n7878 a_400_62400# 0.16fF
C8743 VN.t1343 a_400_62400# 0.03fF
C8744 VN.n7879 a_400_62400# 0.19fF
C8745 VN.t2465 a_400_62400# 0.03fF
C8746 VN.n7881 a_400_62400# 0.32fF
C8747 VN.n7882 a_400_62400# 0.48fF
C8748 VN.n7883 a_400_62400# 0.81fF
C8749 VN.n7884 a_400_62400# 2.46fF
C8750 VN.n7885 a_400_62400# 4.01fF
C8751 VN.t1635 a_400_62400# 0.03fF
C8752 VN.n7886 a_400_62400# 0.32fF
C8753 VN.n7887 a_400_62400# 1.22fF
C8754 VN.n7888 a_400_62400# 0.07fF
C8755 VN.t1527 a_400_62400# 0.03fF
C8756 VN.n7889 a_400_62400# 0.16fF
C8757 VN.n7890 a_400_62400# 0.19fF
C8758 VN.n7892 a_400_62400# 2.53fF
C8759 VN.n7893 a_400_62400# 2.51fF
C8760 VN.t444 a_400_62400# 0.03fF
C8761 VN.n7894 a_400_62400# 0.32fF
C8762 VN.n7895 a_400_62400# 0.48fF
C8763 VN.n7896 a_400_62400# 0.81fF
C8764 VN.n7897 a_400_62400# 0.16fF
C8765 VN.t1802 a_400_62400# 0.03fF
C8766 VN.n7898 a_400_62400# 0.19fF
C8767 VN.n7900 a_400_62400# 1.55fF
C8768 VN.n7901 a_400_62400# 0.29fF
C8769 VN.n7902 a_400_62400# 2.52fF
C8770 VN.t2132 a_400_62400# 0.03fF
C8771 VN.n7903 a_400_62400# 0.32fF
C8772 VN.n7904 a_400_62400# 1.22fF
C8773 VN.n7905 a_400_62400# 0.07fF
C8774 VN.t2005 a_400_62400# 0.03fF
C8775 VN.n7906 a_400_62400# 0.16fF
C8776 VN.n7907 a_400_62400# 0.19fF
C8777 VN.n7909 a_400_62400# 1.04fF
C8778 VN.n7910 a_400_62400# 2.60fF
C8779 VN.n7911 a_400_62400# 2.51fF
C8780 VN.n7912 a_400_62400# 0.16fF
C8781 VN.t926 a_400_62400# 0.03fF
C8782 VN.n7913 a_400_62400# 0.19fF
C8783 VN.t2091 a_400_62400# 0.03fF
C8784 VN.n7915 a_400_62400# 0.32fF
C8785 VN.n7916 a_400_62400# 0.48fF
C8786 VN.n7917 a_400_62400# 0.81fF
C8787 VN.n7918 a_400_62400# 2.46fF
C8788 VN.n7919 a_400_62400# 4.01fF
C8789 VN.t1257 a_400_62400# 0.03fF
C8790 VN.n7920 a_400_62400# 0.32fF
C8791 VN.n7921 a_400_62400# 1.22fF
C8792 VN.n7922 a_400_62400# 0.07fF
C8793 VN.t1132 a_400_62400# 0.03fF
C8794 VN.n7923 a_400_62400# 0.16fF
C8795 VN.n7924 a_400_62400# 0.19fF
C8796 VN.n7926 a_400_62400# 2.53fF
C8797 VN.n7927 a_400_62400# 2.51fF
C8798 VN.t1217 a_400_62400# 0.03fF
C8799 VN.n7928 a_400_62400# 0.32fF
C8800 VN.n7929 a_400_62400# 0.48fF
C8801 VN.n7930 a_400_62400# 0.81fF
C8802 VN.n7931 a_400_62400# 0.16fF
C8803 VN.t185 a_400_62400# 0.03fF
C8804 VN.n7932 a_400_62400# 0.19fF
C8805 VN.n7934 a_400_62400# 1.55fF
C8806 VN.n7935 a_400_62400# 0.29fF
C8807 VN.n7936 a_400_62400# 2.52fF
C8808 VN.t388 a_400_62400# 0.03fF
C8809 VN.n7937 a_400_62400# 0.32fF
C8810 VN.n7938 a_400_62400# 1.22fF
C8811 VN.n7939 a_400_62400# 0.07fF
C8812 VN.t268 a_400_62400# 0.03fF
C8813 VN.n7940 a_400_62400# 0.16fF
C8814 VN.n7941 a_400_62400# 0.19fF
C8815 VN.n7943 a_400_62400# 1.04fF
C8816 VN.n7944 a_400_62400# 2.60fF
C8817 VN.n7945 a_400_62400# 2.51fF
C8818 VN.n7946 a_400_62400# 0.16fF
C8819 VN.t1842 a_400_62400# 0.03fF
C8820 VN.n7947 a_400_62400# 0.19fF
C8821 VN.t487 a_400_62400# 0.03fF
C8822 VN.n7949 a_400_62400# 0.32fF
C8823 VN.n7950 a_400_62400# 0.48fF
C8824 VN.n7951 a_400_62400# 0.81fF
C8825 VN.n7952 a_400_62400# 2.46fF
C8826 VN.n7953 a_400_62400# 4.01fF
C8827 VN.t2173 a_400_62400# 0.03fF
C8828 VN.n7954 a_400_62400# 0.32fF
C8829 VN.n7955 a_400_62400# 1.22fF
C8830 VN.n7956 a_400_62400# 0.07fF
C8831 VN.t1919 a_400_62400# 0.03fF
C8832 VN.n7957 a_400_62400# 0.16fF
C8833 VN.n7958 a_400_62400# 0.19fF
C8834 VN.n7960 a_400_62400# 2.53fF
C8835 VN.n7961 a_400_62400# 2.34fF
C8836 VN.t2141 a_400_62400# 0.03fF
C8837 VN.n7962 a_400_62400# 0.32fF
C8838 VN.n7963 a_400_62400# 0.48fF
C8839 VN.n7964 a_400_62400# 0.81fF
C8840 VN.n7965 a_400_62400# 0.16fF
C8841 VN.t970 a_400_62400# 0.03fF
C8842 VN.n7966 a_400_62400# 0.19fF
C8843 VN.n7968 a_400_62400# 1.55fF
C8844 VN.n7969 a_400_62400# 0.29fF
C8845 VN.n7970 a_400_62400# 3.27fF
C8846 VN.t1306 a_400_62400# 0.03fF
C8847 VN.n7971 a_400_62400# 0.32fF
C8848 VN.n7972 a_400_62400# 1.22fF
C8849 VN.n7973 a_400_62400# 0.07fF
C8850 VN.t1044 a_400_62400# 0.03fF
C8851 VN.n7974 a_400_62400# 0.16fF
C8852 VN.n7975 a_400_62400# 0.19fF
C8853 VN.n7977 a_400_62400# 2.51fF
C8854 VN.n7978 a_400_62400# 0.56fF
C8855 VN.n7979 a_400_62400# 0.64fF
C8856 VN.n7980 a_400_62400# 0.12fF
C8857 VN.n7981 a_400_62400# 0.44fF
C8858 VN.n7982 a_400_62400# 0.40fF
C8859 VN.n7983 a_400_62400# 1.03fF
C8860 VN.n7984 a_400_62400# 0.79fF
C8861 VN.t1267 a_400_62400# 0.03fF
C8862 VN.n7985 a_400_62400# 0.32fF
C8863 VN.n7986 a_400_62400# 0.48fF
C8864 VN.n7987 a_400_62400# 0.81fF
C8865 VN.n7988 a_400_62400# 0.16fF
C8866 VN.t74 a_400_62400# 0.03fF
C8867 VN.n7989 a_400_62400# 0.19fF
C8868 VN.n7991 a_400_62400# 3.50fF
C8869 VN.n7992 a_400_62400# 2.89fF
C8870 VN.t442 a_400_62400# 0.03fF
C8871 VN.n7993 a_400_62400# 0.32fF
C8872 VN.n7994 a_400_62400# 1.22fF
C8873 VN.n7995 a_400_62400# 0.07fF
C8874 VN.t175 a_400_62400# 0.03fF
C8875 VN.n7996 a_400_62400# 0.16fF
C8876 VN.n7997 a_400_62400# 0.19fF
C8877 VN.n7999 a_400_62400# 1.05fF
C8878 VN.n8000 a_400_62400# 3.07fF
C8879 VN.n8001 a_400_62400# 2.51fF
C8880 VN.n8002 a_400_62400# 0.16fF
C8881 VN.t1760 a_400_62400# 0.03fF
C8882 VN.n8003 a_400_62400# 0.19fF
C8883 VN.t398 a_400_62400# 0.03fF
C8884 VN.n8005 a_400_62400# 0.32fF
C8885 VN.n8006 a_400_62400# 0.48fF
C8886 VN.n8007 a_400_62400# 0.81fF
C8887 VN.n8008 a_400_62400# 1.86fF
C8888 VN.n8009 a_400_62400# 1.53fF
C8889 VN.n8010 a_400_62400# 0.47fF
C8890 VN.n8011 a_400_62400# 2.71fF
C8891 VN.t2087 a_400_62400# 0.03fF
C8892 VN.n8012 a_400_62400# 0.32fF
C8893 VN.n8013 a_400_62400# 1.22fF
C8894 VN.n8014 a_400_62400# 0.07fF
C8895 VN.t1837 a_400_62400# 0.03fF
C8896 VN.n8015 a_400_62400# 0.16fF
C8897 VN.n8016 a_400_62400# 0.19fF
C8898 VN.n8018 a_400_62400# 2.53fF
C8899 VN.n8019 a_400_62400# 2.51fF
C8900 VN.t2047 a_400_62400# 0.03fF
C8901 VN.n8020 a_400_62400# 0.32fF
C8902 VN.n8021 a_400_62400# 0.48fF
C8903 VN.n8022 a_400_62400# 0.81fF
C8904 VN.n8023 a_400_62400# 0.16fF
C8905 VN.t889 a_400_62400# 0.03fF
C8906 VN.n8024 a_400_62400# 0.19fF
C8907 VN.n8026 a_400_62400# 1.55fF
C8908 VN.n8027 a_400_62400# 0.29fF
C8909 VN.n8028 a_400_62400# 2.52fF
C8910 VN.t1211 a_400_62400# 0.03fF
C8911 VN.n8029 a_400_62400# 0.32fF
C8912 VN.n8030 a_400_62400# 1.22fF
C8913 VN.n8031 a_400_62400# 0.07fF
C8914 VN.t1095 a_400_62400# 0.03fF
C8915 VN.n8032 a_400_62400# 0.16fF
C8916 VN.n8033 a_400_62400# 0.19fF
C8917 VN.n8035 a_400_62400# 27.83fF
C8918 VN.n8036 a_400_62400# 3.93fF
C8919 VN.n8037 a_400_62400# 2.51fF
C8920 VN.n8038 a_400_62400# 0.16fF
C8921 VN.t2550 a_400_62400# 0.03fF
C8922 VN.n8039 a_400_62400# 0.19fF
C8923 VN.t1179 a_400_62400# 0.03fF
C8924 VN.n8041 a_400_62400# 0.32fF
C8925 VN.n8042 a_400_62400# 0.48fF
C8926 VN.n8043 a_400_62400# 0.81fF
C8927 VN.n8044 a_400_62400# 1.46fF
C8928 VN.n8045 a_400_62400# 0.21fF
C8929 VN.n8046 a_400_62400# 2.81fF
C8930 VN.t226 a_400_62400# 0.03fF
C8931 VN.n8047 a_400_62400# 0.16fF
C8932 VN.n8048 a_400_62400# 0.19fF
C8933 VN.t348 a_400_62400# 0.03fF
C8934 VN.n8050 a_400_62400# 0.32fF
C8935 VN.n8051 a_400_62400# 1.22fF
C8936 VN.n8052 a_400_62400# 0.07fF
C8937 VN.n8053 a_400_62400# 2.51fF
C8938 VN.n8054 a_400_62400# 3.57fF
C8939 VN.t85 a_400_62400# 0.03fF
C8940 VN.n8055 a_400_62400# 0.32fF
C8941 VN.n8056 a_400_62400# 0.48fF
C8942 VN.n8057 a_400_62400# 0.81fF
C8943 VN.n8058 a_400_62400# 0.16fF
C8944 VN.t1499 a_400_62400# 0.03fF
C8945 VN.n8059 a_400_62400# 0.19fF
C8946 VN.n8061 a_400_62400# 3.93fF
C8947 VN.n8062 a_400_62400# 3.08fF
C8948 VN.t1683 a_400_62400# 0.03fF
C8949 VN.n8063 a_400_62400# 0.16fF
C8950 VN.n8064 a_400_62400# 0.19fF
C8951 VN.t1910 a_400_62400# 0.03fF
C8952 VN.n8066 a_400_62400# 0.32fF
C8953 VN.n8067 a_400_62400# 1.22fF
C8954 VN.n8068 a_400_62400# 0.07fF
C8955 VN.n8069 a_400_62400# 2.51fF
C8956 VN.n8070 a_400_62400# 3.57fF
C8957 VN.t1764 a_400_62400# 0.03fF
C8958 VN.n8071 a_400_62400# 0.32fF
C8959 VN.n8072 a_400_62400# 0.48fF
C8960 VN.n8073 a_400_62400# 0.81fF
C8961 VN.n8074 a_400_62400# 0.16fF
C8962 VN.t633 a_400_62400# 0.03fF
C8963 VN.n8075 a_400_62400# 0.19fF
C8964 VN.n8077 a_400_62400# 3.75fF
C8965 VN.n8078 a_400_62400# 3.08fF
C8966 VN.t817 a_400_62400# 0.03fF
C8967 VN.n8079 a_400_62400# 0.16fF
C8968 VN.n8080 a_400_62400# 0.19fF
C8969 VN.t1035 a_400_62400# 0.03fF
C8970 VN.n8082 a_400_62400# 0.32fF
C8971 VN.n8083 a_400_62400# 1.22fF
C8972 VN.n8084 a_400_62400# 0.07fF
C8973 VN.n8085 a_400_62400# 3.65fF
C8974 VN.n8086 a_400_62400# 2.14fF
C8975 VN.n8087 a_400_62400# 0.16fF
C8976 VN.t1542 a_400_62400# 0.03fF
C8977 VN.n8088 a_400_62400# 0.19fF
C8978 VN.t2555 a_400_62400# 0.03fF
C8979 VN.n8090 a_400_62400# 0.32fF
C8980 VN.n8091 a_400_62400# 0.48fF
C8981 VN.n8092 a_400_62400# 0.81fF
C8982 VN.n8093 a_400_62400# 0.09fF
C8983 VN.n8094 a_400_62400# 0.01fF
C8984 VN.n8095 a_400_62400# 0.02fF
C8985 VN.n8096 a_400_62400# 0.02fF
C8986 VN.n8097 a_400_62400# 0.32fF
C8987 VN.n8098 a_400_62400# 1.56fF
C8988 VN.n8099 a_400_62400# 1.81fF
C8989 VN.n8100 a_400_62400# 3.08fF
C8990 VN.t1613 a_400_62400# 0.03fF
C8991 VN.n8101 a_400_62400# 0.16fF
C8992 VN.n8102 a_400_62400# 0.19fF
C8993 VN.t1827 a_400_62400# 0.03fF
C8994 VN.n8104 a_400_62400# 0.32fF
C8995 VN.n8105 a_400_62400# 1.22fF
C8996 VN.n8106 a_400_62400# 0.07fF
C8997 VN.t73 a_400_62400# 64.69fF
C8998 VN.t163 a_400_62400# 0.03fF
C8999 VN.n8107 a_400_62400# 0.32fF
C9000 VN.n8108 a_400_62400# 1.22fF
C9001 VN.n8109 a_400_62400# 0.07fF
C9002 VN.t2474 a_400_62400# 0.03fF
C9003 VN.n8110 a_400_62400# 0.16fF
C9004 VN.n8111 a_400_62400# 0.19fF
C9005 VN.n8113 a_400_62400# 0.16fF
C9006 VN.t2290 a_400_62400# 0.03fF
C9007 VN.n8114 a_400_62400# 0.19fF
C9008 VN.n8116 a_400_62400# 6.92fF
C9009 VN.n8117 a_400_62400# 6.56fF
C9010 VN.t1582 a_400_62400# 0.03fF
C9011 VN.n8118 a_400_62400# 0.16fF
C9012 VN.n8119 a_400_62400# 0.19fF
C9013 VN.t1100 a_400_62400# 0.03fF
C9014 VN.n8121 a_400_62400# 0.32fF
C9015 VN.n8122 a_400_62400# 1.22fF
C9016 VN.n8123 a_400_62400# 0.07fF
C9017 VN.n8124 a_400_62400# 2.51fF
C9018 VN.n8125 a_400_62400# 3.58fF
C9019 VN.t1191 a_400_62400# 0.03fF
C9020 VN.n8126 a_400_62400# 0.32fF
C9021 VN.n8127 a_400_62400# 0.48fF
C9022 VN.n8128 a_400_62400# 0.81fF
C9023 VN.n8129 a_400_62400# 0.16fF
C9024 VN.t2553 a_400_62400# 0.03fF
C9025 VN.n8130 a_400_62400# 0.19fF
C9026 VN.n8132 a_400_62400# 7.29fF
C9027 VN.t717 a_400_62400# 0.03fF
C9028 VN.n8133 a_400_62400# 0.16fF
C9029 VN.n8134 a_400_62400# 0.19fF
C9030 VN.t233 a_400_62400# 0.03fF
C9031 VN.n8136 a_400_62400# 0.32fF
C9032 VN.n8137 a_400_62400# 1.22fF
C9033 VN.n8138 a_400_62400# 0.07fF
C9034 VN.t80 a_400_62400# 64.17fF
C9035 VN.t1880 a_400_62400# 0.03fF
C9036 VN.n8139 a_400_62400# 1.60fF
C9037 VN.n8140 a_400_62400# 0.07fF
C9038 VN.t2488 a_400_62400# 0.03fF
C9039 VN.n8141 a_400_62400# 0.02fF
C9040 VN.n8142 a_400_62400# 0.34fF
C9041 VN.n8144 a_400_62400# 2.01fF
C9042 VN.n8145 a_400_62400# 1.75fF
C9043 VN.n8146 a_400_62400# 0.37fF
C9044 VN.n8147 a_400_62400# 0.33fF
C9045 VN.n8148 a_400_62400# 5.88fF
C9046 VN.n8149 a_400_62400# 0.02fF
C9047 VN.n8150 a_400_62400# 0.02fF
C9048 VN.n8151 a_400_62400# 0.03fF
C9049 VN.n8152 a_400_62400# 0.05fF
C9050 VN.n8153 a_400_62400# 0.23fF
C9051 VN.n8154 a_400_62400# 0.02fF
C9052 VN.n8155 a_400_62400# 0.03fF
C9053 VN.n8156 a_400_62400# 0.01fF
C9054 VN.n8157 a_400_62400# 0.01fF
C9055 VN.n8158 a_400_62400# 0.01fF
C9056 VN.n8159 a_400_62400# 0.02fF
C9057 VN.n8160 a_400_62400# 0.03fF
C9058 VN.n8161 a_400_62400# 0.06fF
C9059 VN.n8162 a_400_62400# 0.05fF
C9060 VN.n8163 a_400_62400# 0.15fF
C9061 VN.n8164 a_400_62400# 0.51fF
C9062 VN.n8165 a_400_62400# 0.27fF
C9063 VN.n8166 a_400_62400# 37.46fF
C9064 VN.n8167 a_400_62400# 37.46fF
C9065 VN.n8168 a_400_62400# 0.79fF
C9066 VN.n8169 a_400_62400# 0.23fF
C9067 VN.n8170 a_400_62400# 1.18fF
C9068 VN.t155 a_400_62400# 28.64fF
C9069 VN.n8171 a_400_62400# 0.79fF
C9070 VN.n8172 a_400_62400# 0.11fF
C9071 VN.n8173 a_400_62400# 4.98fF
C9072 VN.n8174 a_400_62400# 0.80fF
C9073 VN.n8175 a_400_62400# 0.29fF
C9074 VN.n8176 a_400_62400# 1.96fF
C9075 VN.n8178 a_400_62400# 25.18fF
C9076 VN.n8180 a_400_62400# 1.87fF
C9077 VN.n8181 a_400_62400# 5.36fF
C9078 VN.n8182 a_400_62400# 1.81fF
C9079 VN.t1160 a_400_62400# 0.03fF
C9080 VN.n8183 a_400_62400# 0.85fF
C9081 VN.n8184 a_400_62400# 0.81fF
C9082 VN.n8185 a_400_62400# 2.53fF
C9083 VN.n8186 a_400_62400# 0.08fF
C9084 VN.n8187 a_400_62400# 0.04fF
C9085 VN.n8188 a_400_62400# 0.05fF
C9086 VN.n8189 a_400_62400# 1.33fF
C9087 VN.n8190 a_400_62400# 0.03fF
C9088 VN.n8191 a_400_62400# 0.01fF
C9089 VN.n8192 a_400_62400# 0.02fF
C9090 VN.n8193 a_400_62400# 0.11fF
C9091 VN.n8194 a_400_62400# 0.48fF
C9092 VN.n8195 a_400_62400# 2.48fF
C9093 VN.t902 a_400_62400# 0.03fF
C9094 VN.n8196 a_400_62400# 0.32fF
C9095 VN.n8197 a_400_62400# 0.48fF
C9096 VN.n8198 a_400_62400# 0.81fF
C9097 VN.n8199 a_400_62400# 0.16fF
C9098 VN.t2423 a_400_62400# 0.03fF
C9099 VN.n8200 a_400_62400# 0.19fF
C9100 VN.n8202 a_400_62400# 0.93fF
C9101 VN.n8203 a_400_62400# 0.30fF
C9102 VN.n8204 a_400_62400# 0.34fF
C9103 VN.n8205 a_400_62400# 0.12fF
C9104 VN.n8206 a_400_62400# 0.30fF
C9105 VN.n8207 a_400_62400# 0.93fF
C9106 VN.n8208 a_400_62400# 1.55fF
C9107 VN.n8209 a_400_62400# 0.29fF
C9108 VN.n8210 a_400_62400# 0.34fF
C9109 VN.n8211 a_400_62400# 0.12fF
C9110 VN.n8212 a_400_62400# 2.52fF
C9111 VN.t940 a_400_62400# 0.03fF
C9112 VN.n8213 a_400_62400# 0.32fF
C9113 VN.n8214 a_400_62400# 1.22fF
C9114 VN.n8215 a_400_62400# 0.07fF
C9115 VN.t585 a_400_62400# 0.03fF
C9116 VN.n8216 a_400_62400# 0.16fF
C9117 VN.n8217 a_400_62400# 0.19fF
C9118 VN.n8219 a_400_62400# 0.33fF
C9119 VN.n8220 a_400_62400# 0.12fF
C9120 VN.n8221 a_400_62400# 0.28fF
C9121 VN.n8222 a_400_62400# 1.72fF
C9122 VN.n8223 a_400_62400# 0.71fF
C9123 VN.n8224 a_400_62400# 2.51fF
C9124 VN.n8225 a_400_62400# 0.16fF
C9125 VN.t1561 a_400_62400# 0.03fF
C9126 VN.n8226 a_400_62400# 0.19fF
C9127 VN.t156 a_400_62400# 0.03fF
C9128 VN.n8228 a_400_62400# 0.32fF
C9129 VN.n8229 a_400_62400# 0.48fF
C9130 VN.n8230 a_400_62400# 0.81fF
C9131 VN.n8231 a_400_62400# 0.03fF
C9132 VN.n8232 a_400_62400# 0.01fF
C9133 VN.n8233 a_400_62400# 0.02fF
C9134 VN.n8234 a_400_62400# 0.11fF
C9135 VN.n8235 a_400_62400# 0.08fF
C9136 VN.n8236 a_400_62400# 0.04fF
C9137 VN.n8237 a_400_62400# 0.05fF
C9138 VN.n8238 a_400_62400# 1.34fF
C9139 VN.n8239 a_400_62400# 0.48fF
C9140 VN.n8240 a_400_62400# 2.51fF
C9141 VN.n8241 a_400_62400# 2.67fF
C9142 VN.t205 a_400_62400# 0.03fF
C9143 VN.n8242 a_400_62400# 0.32fF
C9144 VN.n8243 a_400_62400# 1.22fF
C9145 VN.n8244 a_400_62400# 0.07fF
C9146 VN.t2241 a_400_62400# 0.03fF
C9147 VN.n8245 a_400_62400# 0.16fF
C9148 VN.n8246 a_400_62400# 0.19fF
C9149 VN.n8248 a_400_62400# 2.53fF
C9150 VN.n8249 a_400_62400# 0.08fF
C9151 VN.n8250 a_400_62400# 0.04fF
C9152 VN.n8251 a_400_62400# 0.05fF
C9153 VN.n8252 a_400_62400# 1.33fF
C9154 VN.n8253 a_400_62400# 0.03fF
C9155 VN.n8254 a_400_62400# 0.01fF
C9156 VN.n8255 a_400_62400# 0.02fF
C9157 VN.n8256 a_400_62400# 0.11fF
C9158 VN.n8257 a_400_62400# 0.48fF
C9159 VN.n8258 a_400_62400# 2.48fF
C9160 VN.t1819 a_400_62400# 0.03fF
C9161 VN.n8259 a_400_62400# 0.32fF
C9162 VN.n8260 a_400_62400# 0.48fF
C9163 VN.n8261 a_400_62400# 0.81fF
C9164 VN.n8262 a_400_62400# 0.16fF
C9165 VN.t691 a_400_62400# 0.03fF
C9166 VN.n8263 a_400_62400# 0.19fF
C9167 VN.n8265 a_400_62400# 0.93fF
C9168 VN.n8266 a_400_62400# 0.30fF
C9169 VN.n8267 a_400_62400# 0.34fF
C9170 VN.n8268 a_400_62400# 0.12fF
C9171 VN.n8269 a_400_62400# 0.30fF
C9172 VN.n8270 a_400_62400# 0.93fF
C9173 VN.n8271 a_400_62400# 1.55fF
C9174 VN.n8272 a_400_62400# 0.29fF
C9175 VN.n8273 a_400_62400# 0.34fF
C9176 VN.n8274 a_400_62400# 0.12fF
C9177 VN.n8275 a_400_62400# 2.52fF
C9178 VN.t1857 a_400_62400# 0.03fF
C9179 VN.n8276 a_400_62400# 0.32fF
C9180 VN.n8277 a_400_62400# 1.22fF
C9181 VN.n8278 a_400_62400# 0.07fF
C9182 VN.t1377 a_400_62400# 0.03fF
C9183 VN.n8279 a_400_62400# 0.16fF
C9184 VN.n8280 a_400_62400# 0.19fF
C9185 VN.n8282 a_400_62400# 0.33fF
C9186 VN.n8283 a_400_62400# 0.12fF
C9187 VN.n8284 a_400_62400# 0.28fF
C9188 VN.n8285 a_400_62400# 1.23fF
C9189 VN.n8286 a_400_62400# 0.59fF
C9190 VN.n8287 a_400_62400# 2.51fF
C9191 VN.n8288 a_400_62400# 0.16fF
C9192 VN.t1176 a_400_62400# 0.03fF
C9193 VN.n8289 a_400_62400# 0.19fF
C9194 VN.t2316 a_400_62400# 0.03fF
C9195 VN.n8291 a_400_62400# 0.32fF
C9196 VN.n8292 a_400_62400# 0.48fF
C9197 VN.n8293 a_400_62400# 0.81fF
C9198 VN.n8294 a_400_62400# 0.03fF
C9199 VN.n8295 a_400_62400# 0.01fF
C9200 VN.n8296 a_400_62400# 0.02fF
C9201 VN.n8297 a_400_62400# 0.11fF
C9202 VN.n8298 a_400_62400# 0.08fF
C9203 VN.n8299 a_400_62400# 0.04fF
C9204 VN.n8300 a_400_62400# 0.05fF
C9205 VN.n8301 a_400_62400# 1.34fF
C9206 VN.n8302 a_400_62400# 0.48fF
C9207 VN.n8303 a_400_62400# 2.51fF
C9208 VN.n8304 a_400_62400# 2.67fF
C9209 VN.t2352 a_400_62400# 0.03fF
C9210 VN.n8305 a_400_62400# 0.32fF
C9211 VN.n8306 a_400_62400# 1.22fF
C9212 VN.n8307 a_400_62400# 0.07fF
C9213 VN.t512 a_400_62400# 0.03fF
C9214 VN.n8308 a_400_62400# 0.16fF
C9215 VN.n8309 a_400_62400# 0.19fF
C9216 VN.n8311 a_400_62400# 2.53fF
C9217 VN.n8312 a_400_62400# 0.08fF
C9218 VN.n8313 a_400_62400# 0.04fF
C9219 VN.n8314 a_400_62400# 0.05fF
C9220 VN.n8315 a_400_62400# 1.33fF
C9221 VN.n8316 a_400_62400# 0.03fF
C9222 VN.n8317 a_400_62400# 0.01fF
C9223 VN.n8318 a_400_62400# 0.02fF
C9224 VN.n8319 a_400_62400# 0.11fF
C9225 VN.n8320 a_400_62400# 0.48fF
C9226 VN.n8321 a_400_62400# 2.48fF
C9227 VN.t1447 a_400_62400# 0.03fF
C9228 VN.n8322 a_400_62400# 0.32fF
C9229 VN.n8323 a_400_62400# 0.48fF
C9230 VN.n8324 a_400_62400# 0.81fF
C9231 VN.n8325 a_400_62400# 0.16fF
C9232 VN.t308 a_400_62400# 0.03fF
C9233 VN.n8326 a_400_62400# 0.19fF
C9234 VN.n8328 a_400_62400# 0.93fF
C9235 VN.n8329 a_400_62400# 0.30fF
C9236 VN.n8330 a_400_62400# 0.34fF
C9237 VN.n8331 a_400_62400# 0.12fF
C9238 VN.n8332 a_400_62400# 0.30fF
C9239 VN.n8333 a_400_62400# 0.93fF
C9240 VN.n8334 a_400_62400# 1.55fF
C9241 VN.n8335 a_400_62400# 0.29fF
C9242 VN.n8336 a_400_62400# 0.34fF
C9243 VN.n8337 a_400_62400# 0.12fF
C9244 VN.n8338 a_400_62400# 2.52fF
C9245 VN.t1484 a_400_62400# 0.03fF
C9246 VN.n8339 a_400_62400# 0.32fF
C9247 VN.n8340 a_400_62400# 1.22fF
C9248 VN.n8341 a_400_62400# 0.07fF
C9249 VN.t965 a_400_62400# 0.03fF
C9250 VN.n8342 a_400_62400# 0.16fF
C9251 VN.n8343 a_400_62400# 0.19fF
C9252 VN.n8345 a_400_62400# 0.33fF
C9253 VN.n8346 a_400_62400# 0.12fF
C9254 VN.n8347 a_400_62400# 0.28fF
C9255 VN.n8348 a_400_62400# 1.23fF
C9256 VN.n8349 a_400_62400# 0.59fF
C9257 VN.n8350 a_400_62400# 2.51fF
C9258 VN.n8351 a_400_62400# 0.16fF
C9259 VN.t1956 a_400_62400# 0.03fF
C9260 VN.n8352 a_400_62400# 0.19fF
C9261 VN.t577 a_400_62400# 0.03fF
C9262 VN.n8354 a_400_62400# 0.32fF
C9263 VN.n8355 a_400_62400# 0.48fF
C9264 VN.n8356 a_400_62400# 0.81fF
C9265 VN.n8357 a_400_62400# 0.03fF
C9266 VN.n8358 a_400_62400# 0.01fF
C9267 VN.n8359 a_400_62400# 0.02fF
C9268 VN.n8360 a_400_62400# 0.11fF
C9269 VN.n8361 a_400_62400# 0.08fF
C9270 VN.n8362 a_400_62400# 0.04fF
C9271 VN.n8363 a_400_62400# 0.05fF
C9272 VN.n8364 a_400_62400# 1.34fF
C9273 VN.n8365 a_400_62400# 0.48fF
C9274 VN.n8366 a_400_62400# 2.51fF
C9275 VN.n8367 a_400_62400# 2.67fF
C9276 VN.t617 a_400_62400# 0.03fF
C9277 VN.n8368 a_400_62400# 0.32fF
C9278 VN.n8369 a_400_62400# 1.22fF
C9279 VN.n8370 a_400_62400# 0.07fF
C9280 VN.t61 a_400_62400# 0.03fF
C9281 VN.n8371 a_400_62400# 0.16fF
C9282 VN.n8372 a_400_62400# 0.19fF
C9283 VN.n8374 a_400_62400# 2.53fF
C9284 VN.n8375 a_400_62400# 0.08fF
C9285 VN.n8376 a_400_62400# 0.04fF
C9286 VN.n8377 a_400_62400# 0.05fF
C9287 VN.n8378 a_400_62400# 1.33fF
C9288 VN.n8379 a_400_62400# 0.03fF
C9289 VN.n8380 a_400_62400# 0.01fF
C9290 VN.n8381 a_400_62400# 0.02fF
C9291 VN.n8382 a_400_62400# 0.11fF
C9292 VN.n8383 a_400_62400# 0.48fF
C9293 VN.n8384 a_400_62400# 2.48fF
C9294 VN.t2235 a_400_62400# 0.03fF
C9295 VN.n8385 a_400_62400# 0.32fF
C9296 VN.n8386 a_400_62400# 0.48fF
C9297 VN.n8387 a_400_62400# 0.81fF
C9298 VN.n8388 a_400_62400# 0.16fF
C9299 VN.t1089 a_400_62400# 0.03fF
C9300 VN.n8389 a_400_62400# 0.19fF
C9301 VN.n8391 a_400_62400# 0.93fF
C9302 VN.n8392 a_400_62400# 0.30fF
C9303 VN.n8393 a_400_62400# 0.34fF
C9304 VN.n8394 a_400_62400# 0.12fF
C9305 VN.n8395 a_400_62400# 0.30fF
C9306 VN.n8396 a_400_62400# 0.93fF
C9307 VN.n8397 a_400_62400# 1.55fF
C9308 VN.n8398 a_400_62400# 0.29fF
C9309 VN.n8399 a_400_62400# 0.34fF
C9310 VN.n8400 a_400_62400# 0.12fF
C9311 VN.n8401 a_400_62400# 2.52fF
C9312 VN.t2269 a_400_62400# 0.03fF
C9313 VN.n8402 a_400_62400# 0.32fF
C9314 VN.n8403 a_400_62400# 1.22fF
C9315 VN.n8404 a_400_62400# 0.07fF
C9316 VN.t1879 a_400_62400# 0.03fF
C9317 VN.n8405 a_400_62400# 0.16fF
C9318 VN.n8406 a_400_62400# 0.19fF
C9319 VN.n8408 a_400_62400# 0.33fF
C9320 VN.n8409 a_400_62400# 0.12fF
C9321 VN.n8410 a_400_62400# 0.28fF
C9322 VN.n8411 a_400_62400# 1.23fF
C9323 VN.n8412 a_400_62400# 0.59fF
C9324 VN.n8413 a_400_62400# 2.51fF
C9325 VN.n8414 a_400_62400# 0.16fF
C9326 VN.t219 a_400_62400# 0.03fF
C9327 VN.n8415 a_400_62400# 0.19fF
C9328 VN.t1372 a_400_62400# 0.03fF
C9329 VN.n8417 a_400_62400# 0.32fF
C9330 VN.n8418 a_400_62400# 0.48fF
C9331 VN.n8419 a_400_62400# 0.81fF
C9332 VN.n8420 a_400_62400# 0.03fF
C9333 VN.n8421 a_400_62400# 0.01fF
C9334 VN.n8422 a_400_62400# 0.02fF
C9335 VN.n8423 a_400_62400# 0.11fF
C9336 VN.n8424 a_400_62400# 0.08fF
C9337 VN.n8425 a_400_62400# 0.04fF
C9338 VN.n8426 a_400_62400# 0.05fF
C9339 VN.n8427 a_400_62400# 1.34fF
C9340 VN.n8428 a_400_62400# 0.48fF
C9341 VN.n8429 a_400_62400# 2.51fF
C9342 VN.n8430 a_400_62400# 2.67fF
C9343 VN.t1405 a_400_62400# 0.03fF
C9344 VN.n8431 a_400_62400# 0.32fF
C9345 VN.n8432 a_400_62400# 1.22fF
C9346 VN.n8433 a_400_62400# 0.07fF
C9347 VN.t1011 a_400_62400# 0.03fF
C9348 VN.n8434 a_400_62400# 0.16fF
C9349 VN.n8435 a_400_62400# 0.19fF
C9350 VN.n8437 a_400_62400# 2.53fF
C9351 VN.n8438 a_400_62400# 0.09fF
C9352 VN.n8439 a_400_62400# 0.05fF
C9353 VN.n8440 a_400_62400# 0.07fF
C9354 VN.n8441 a_400_62400# 1.16fF
C9355 VN.n8442 a_400_62400# 0.01fF
C9356 VN.n8443 a_400_62400# 0.01fF
C9357 VN.n8444 a_400_62400# 0.01fF
C9358 VN.n8445 a_400_62400# 0.09fF
C9359 VN.n8446 a_400_62400# 0.91fF
C9360 VN.n8447 a_400_62400# 0.96fF
C9361 VN.t505 a_400_62400# 0.03fF
C9362 VN.n8448 a_400_62400# 0.32fF
C9363 VN.n8449 a_400_62400# 0.48fF
C9364 VN.n8450 a_400_62400# 0.81fF
C9365 VN.n8451 a_400_62400# 0.16fF
C9366 VN.t1869 a_400_62400# 0.03fF
C9367 VN.n8452 a_400_62400# 0.19fF
C9368 VN.n8454 a_400_62400# 0.93fF
C9369 VN.n8455 a_400_62400# 0.30fF
C9370 VN.n8456 a_400_62400# 0.34fF
C9371 VN.n8457 a_400_62400# 0.12fF
C9372 VN.n8458 a_400_62400# 0.30fF
C9373 VN.n8459 a_400_62400# 0.93fF
C9374 VN.n8460 a_400_62400# 1.55fF
C9375 VN.n8461 a_400_62400# 0.29fF
C9376 VN.n8462 a_400_62400# 0.34fF
C9377 VN.n8463 a_400_62400# 0.12fF
C9378 VN.n8464 a_400_62400# 3.10fF
C9379 VN.t543 a_400_62400# 0.03fF
C9380 VN.n8465 a_400_62400# 0.32fF
C9381 VN.n8466 a_400_62400# 1.22fF
C9382 VN.n8467 a_400_62400# 0.07fF
C9383 VN.t138 a_400_62400# 0.03fF
C9384 VN.n8468 a_400_62400# 0.16fF
C9385 VN.n8469 a_400_62400# 0.19fF
C9386 VN.n8471 a_400_62400# 2.51fF
C9387 VN.n8472 a_400_62400# 0.61fF
C9388 VN.n8473 a_400_62400# 0.30fF
C9389 VN.n8474 a_400_62400# 0.51fF
C9390 VN.n8475 a_400_62400# 0.21fF
C9391 VN.n8476 a_400_62400# 0.38fF
C9392 VN.n8477 a_400_62400# 0.29fF
C9393 VN.n8478 a_400_62400# 0.40fF
C9394 VN.n8479 a_400_62400# 0.28fF
C9395 VN.t2159 a_400_62400# 0.03fF
C9396 VN.n8480 a_400_62400# 0.32fF
C9397 VN.n8481 a_400_62400# 0.48fF
C9398 VN.n8482 a_400_62400# 0.81fF
C9399 VN.n8483 a_400_62400# 0.16fF
C9400 VN.t997 a_400_62400# 0.03fF
C9401 VN.n8484 a_400_62400# 0.19fF
C9402 VN.n8486 a_400_62400# 0.06fF
C9403 VN.n8487 a_400_62400# 0.04fF
C9404 VN.n8488 a_400_62400# 0.04fF
C9405 VN.n8489 a_400_62400# 0.14fF
C9406 VN.n8490 a_400_62400# 0.48fF
C9407 VN.n8491 a_400_62400# 0.50fF
C9408 VN.n8492 a_400_62400# 0.14fF
C9409 VN.n8493 a_400_62400# 0.16fF
C9410 VN.n8494 a_400_62400# 0.09fF
C9411 VN.n8495 a_400_62400# 0.16fF
C9412 VN.n8496 a_400_62400# 0.24fF
C9413 VN.n8497 a_400_62400# 5.35fF
C9414 VN.t2199 a_400_62400# 0.03fF
C9415 VN.n8498 a_400_62400# 0.32fF
C9416 VN.n8499 a_400_62400# 1.22fF
C9417 VN.n8500 a_400_62400# 0.07fF
C9418 VN.t1801 a_400_62400# 0.03fF
C9419 VN.n8501 a_400_62400# 0.16fF
C9420 VN.n8502 a_400_62400# 0.19fF
C9421 VN.n8504 a_400_62400# 0.33fF
C9422 VN.n8505 a_400_62400# 0.12fF
C9423 VN.n8506 a_400_62400# 0.28fF
C9424 VN.n8507 a_400_62400# 1.72fF
C9425 VN.n8508 a_400_62400# 0.71fF
C9426 VN.n8509 a_400_62400# 2.51fF
C9427 VN.n8510 a_400_62400# 0.16fF
C9428 VN.t266 a_400_62400# 0.03fF
C9429 VN.n8511 a_400_62400# 0.19fF
C9430 VN.t1290 a_400_62400# 0.03fF
C9431 VN.n8513 a_400_62400# 0.32fF
C9432 VN.n8514 a_400_62400# 0.48fF
C9433 VN.n8515 a_400_62400# 0.81fF
C9434 VN.n8516 a_400_62400# 0.95fF
C9435 VN.n8517 a_400_62400# 2.11fF
C9436 VN.n8518 a_400_62400# 3.28fF
C9437 VN.t1327 a_400_62400# 0.03fF
C9438 VN.n8519 a_400_62400# 0.32fF
C9439 VN.n8520 a_400_62400# 1.22fF
C9440 VN.n8521 a_400_62400# 0.07fF
C9441 VN.t924 a_400_62400# 0.03fF
C9442 VN.n8522 a_400_62400# 0.16fF
C9443 VN.n8523 a_400_62400# 0.19fF
C9444 VN.n8525 a_400_62400# 2.53fF
C9445 VN.n8526 a_400_62400# 0.08fF
C9446 VN.n8527 a_400_62400# 0.04fF
C9447 VN.n8528 a_400_62400# 0.05fF
C9448 VN.n8529 a_400_62400# 1.33fF
C9449 VN.n8530 a_400_62400# 0.03fF
C9450 VN.n8531 a_400_62400# 0.01fF
C9451 VN.n8532 a_400_62400# 0.02fF
C9452 VN.n8533 a_400_62400# 0.11fF
C9453 VN.n8534 a_400_62400# 0.48fF
C9454 VN.n8535 a_400_62400# 2.48fF
C9455 VN.t545 a_400_62400# 0.03fF
C9456 VN.n8536 a_400_62400# 0.32fF
C9457 VN.n8537 a_400_62400# 0.48fF
C9458 VN.n8538 a_400_62400# 0.81fF
C9459 VN.n8539 a_400_62400# 0.16fF
C9460 VN.t1917 a_400_62400# 0.03fF
C9461 VN.n8540 a_400_62400# 0.19fF
C9462 VN.n8542 a_400_62400# 0.93fF
C9463 VN.n8543 a_400_62400# 0.30fF
C9464 VN.n8544 a_400_62400# 0.34fF
C9465 VN.n8545 a_400_62400# 0.12fF
C9466 VN.n8546 a_400_62400# 0.30fF
C9467 VN.n8547 a_400_62400# 0.93fF
C9468 VN.n8548 a_400_62400# 1.55fF
C9469 VN.n8549 a_400_62400# 0.29fF
C9470 VN.n8550 a_400_62400# 0.34fF
C9471 VN.n8551 a_400_62400# 0.12fF
C9472 VN.n8552 a_400_62400# 2.52fF
C9473 VN.t580 a_400_62400# 0.03fF
C9474 VN.n8553 a_400_62400# 0.32fF
C9475 VN.n8554 a_400_62400# 1.22fF
C9476 VN.n8555 a_400_62400# 0.07fF
C9477 VN.t2586 a_400_62400# 0.03fF
C9478 VN.n8556 a_400_62400# 0.16fF
C9479 VN.n8557 a_400_62400# 0.19fF
C9480 VN.n8559 a_400_62400# 27.83fF
C9481 VN.n8560 a_400_62400# 0.09fF
C9482 VN.n8561 a_400_62400# 0.27fF
C9483 VN.n8562 a_400_62400# 0.12fF
C9484 VN.n8563 a_400_62400# 0.28fF
C9485 VN.n8564 a_400_62400# 0.13fF
C9486 VN.n8565 a_400_62400# 0.40fF
C9487 VN.n8566 a_400_62400# 0.93fF
C9488 VN.n8567 a_400_62400# 0.60fF
C9489 VN.n8568 a_400_62400# 3.12fF
C9490 VN.n8569 a_400_62400# 0.16fF
C9491 VN.t646 a_400_62400# 0.03fF
C9492 VN.n8570 a_400_62400# 0.19fF
C9493 VN.t1774 a_400_62400# 0.03fF
C9494 VN.n8572 a_400_62400# 0.32fF
C9495 VN.n8573 a_400_62400# 0.48fF
C9496 VN.n8574 a_400_62400# 0.81fF
C9497 VN.n8575 a_400_62400# 2.54fF
C9498 VN.n8576 a_400_62400# 0.23fF
C9499 VN.n8577 a_400_62400# 1.02fF
C9500 VN.n8578 a_400_62400# 0.42fF
C9501 VN.n8579 a_400_62400# 0.34fF
C9502 VN.n8580 a_400_62400# 0.40fF
C9503 VN.n8581 a_400_62400# 0.63fF
C9504 VN.n8582 a_400_62400# 0.21fF
C9505 VN.n8583 a_400_62400# 2.58fF
C9506 VN.t1454 a_400_62400# 0.03fF
C9507 VN.n8584 a_400_62400# 0.16fF
C9508 VN.n8585 a_400_62400# 0.19fF
C9509 VN.t1815 a_400_62400# 0.03fF
C9510 VN.n8587 a_400_62400# 0.32fF
C9511 VN.n8588 a_400_62400# 1.22fF
C9512 VN.n8589 a_400_62400# 0.07fF
C9513 VN.n8590 a_400_62400# 2.51fF
C9514 VN.n8591 a_400_62400# 0.16fF
C9515 VN.t948 a_400_62400# 0.03fF
C9516 VN.n8592 a_400_62400# 0.19fF
C9517 VN.t2124 a_400_62400# 0.03fF
C9518 VN.n8594 a_400_62400# 0.32fF
C9519 VN.n8595 a_400_62400# 0.48fF
C9520 VN.n8596 a_400_62400# 0.81fF
C9521 VN.n8597 a_400_62400# 1.24fF
C9522 VN.n8598 a_400_62400# 0.43fF
C9523 VN.n8599 a_400_62400# 0.43fF
C9524 VN.n8600 a_400_62400# 1.24fF
C9525 VN.n8601 a_400_62400# 1.46fF
C9526 VN.n8602 a_400_62400# 0.21fF
C9527 VN.n8603 a_400_62400# 6.64fF
C9528 VN.t1716 a_400_62400# 0.03fF
C9529 VN.n8604 a_400_62400# 0.16fF
C9530 VN.n8605 a_400_62400# 0.19fF
C9531 VN.t1450 a_400_62400# 0.03fF
C9532 VN.n8607 a_400_62400# 0.32fF
C9533 VN.n8608 a_400_62400# 1.22fF
C9534 VN.n8609 a_400_62400# 0.07fF
C9535 VN.n8610 a_400_62400# 2.51fF
C9536 VN.n8611 a_400_62400# 3.57fF
C9537 VN.t1249 a_400_62400# 0.03fF
C9538 VN.n8612 a_400_62400# 0.32fF
C9539 VN.n8613 a_400_62400# 0.48fF
C9540 VN.n8614 a_400_62400# 0.81fF
C9541 VN.n8615 a_400_62400# 0.16fF
C9542 VN.t27 a_400_62400# 0.03fF
C9543 VN.n8616 a_400_62400# 0.19fF
C9544 VN.n8618 a_400_62400# 6.91fF
C9545 VN.t766 a_400_62400# 0.03fF
C9546 VN.n8619 a_400_62400# 0.16fF
C9547 VN.n8620 a_400_62400# 0.19fF
C9548 VN.t582 a_400_62400# 0.03fF
C9549 VN.n8622 a_400_62400# 0.32fF
C9550 VN.n8623 a_400_62400# 1.22fF
C9551 VN.n8624 a_400_62400# 0.07fF
C9552 VN.n8625 a_400_62400# 2.51fF
C9553 VN.n8626 a_400_62400# 3.57fF
C9554 VN.t381 a_400_62400# 0.03fF
C9555 VN.n8627 a_400_62400# 0.32fF
C9556 VN.n8628 a_400_62400# 0.48fF
C9557 VN.n8629 a_400_62400# 0.81fF
C9558 VN.n8630 a_400_62400# 0.16fF
C9559 VN.t1737 a_400_62400# 0.03fF
C9560 VN.n8631 a_400_62400# 0.19fF
C9561 VN.n8633 a_400_62400# 2.51fF
C9562 VN.n8634 a_400_62400# 3.59fF
C9563 VN.t2045 a_400_62400# 0.03fF
C9564 VN.n8635 a_400_62400# 0.32fF
C9565 VN.n8636 a_400_62400# 0.48fF
C9566 VN.n8637 a_400_62400# 0.81fF
C9567 VN.t46 a_400_62400# 0.03fF
C9568 VN.n8638 a_400_62400# 1.63fF
C9569 VN.n8639 a_400_62400# 0.81fF
C9570 VN.n8640 a_400_62400# 1.21fF
C9571 VN.n8641 a_400_62400# 1.54fF
C9572 VN.n8642 a_400_62400# 4.06fF
C9573 VN.t45 a_400_62400# 28.64fF
C9574 VN.n8643 a_400_62400# 28.43fF
C9575 VN.n8645 a_400_62400# 0.50fF
C9576 VN.n8646 a_400_62400# 0.31fF
C9577 VN.n8647 a_400_62400# 3.88fF
C9578 VN.n8648 a_400_62400# 3.29fF
C9579 VN.n8649 a_400_62400# 2.62fF
C9580 VN.n8650 a_400_62400# 5.27fF
C9581 VN.n8651 a_400_62400# 0.34fF
C9582 VN.n8652 a_400_62400# 0.02fF
C9583 VN.t1491 a_400_62400# 0.03fF
C9584 VN.n8653 a_400_62400# 0.34fF
C9585 VN.t1782 a_400_62400# 0.03fF
C9586 VN.n8654 a_400_62400# 1.28fF
C9587 VN.n8655 a_400_62400# 0.94fF
C9588 VN.n8656 a_400_62400# 1.04fF
C9589 VN.n8657 a_400_62400# 2.58fF
C9590 VN.n8658 a_400_62400# 2.51fF
C9591 VN.n8659 a_400_62400# 0.16fF
C9592 VN.t624 a_400_62400# 0.03fF
C9593 VN.n8660 a_400_62400# 0.19fF
C9594 VN.t1743 a_400_62400# 0.03fF
C9595 VN.n8662 a_400_62400# 0.32fF
C9596 VN.n8663 a_400_62400# 0.48fF
C9597 VN.n8664 a_400_62400# 0.81fF
C9598 VN.n8665 a_400_62400# 2.03fF
C9599 VN.n8666 a_400_62400# 4.01fF
C9600 VN.t906 a_400_62400# 0.03fF
C9601 VN.n8667 a_400_62400# 0.32fF
C9602 VN.n8668 a_400_62400# 1.22fF
C9603 VN.n8669 a_400_62400# 0.07fF
C9604 VN.t686 a_400_62400# 0.03fF
C9605 VN.n8670 a_400_62400# 0.16fF
C9606 VN.n8671 a_400_62400# 0.19fF
C9607 VN.n8673 a_400_62400# 2.53fF
C9608 VN.n8674 a_400_62400# 2.51fF
C9609 VN.t871 a_400_62400# 0.03fF
C9610 VN.n8675 a_400_62400# 0.32fF
C9611 VN.n8676 a_400_62400# 0.48fF
C9612 VN.n8677 a_400_62400# 0.81fF
C9613 VN.n8678 a_400_62400# 0.16fF
C9614 VN.t2276 a_400_62400# 0.03fF
C9615 VN.n8679 a_400_62400# 0.19fF
C9616 VN.n8681 a_400_62400# 1.55fF
C9617 VN.n8682 a_400_62400# 0.29fF
C9618 VN.n8683 a_400_62400# 2.52fF
C9619 VN.t2569 a_400_62400# 0.03fF
C9620 VN.n8684 a_400_62400# 0.32fF
C9621 VN.n8685 a_400_62400# 1.22fF
C9622 VN.n8686 a_400_62400# 0.07fF
C9623 VN.t2463 a_400_62400# 0.03fF
C9624 VN.n8687 a_400_62400# 0.16fF
C9625 VN.n8688 a_400_62400# 0.19fF
C9626 VN.n8690 a_400_62400# 1.05fF
C9627 VN.n8691 a_400_62400# 3.07fF
C9628 VN.n8692 a_400_62400# 2.51fF
C9629 VN.n8693 a_400_62400# 0.16fF
C9630 VN.t1408 a_400_62400# 0.03fF
C9631 VN.n8694 a_400_62400# 0.19fF
C9632 VN.t2533 a_400_62400# 0.03fF
C9633 VN.n8696 a_400_62400# 0.32fF
C9634 VN.n8697 a_400_62400# 0.48fF
C9635 VN.n8698 a_400_62400# 0.81fF
C9636 VN.n8699 a_400_62400# 2.46fF
C9637 VN.n8700 a_400_62400# 2.91fF
C9638 VN.t1698 a_400_62400# 0.03fF
C9639 VN.n8701 a_400_62400# 0.32fF
C9640 VN.n8702 a_400_62400# 1.22fF
C9641 VN.n8703 a_400_62400# 0.07fF
C9642 VN.t1597 a_400_62400# 0.03fF
C9643 VN.n8704 a_400_62400# 0.16fF
C9644 VN.n8705 a_400_62400# 0.19fF
C9645 VN.n8707 a_400_62400# 2.53fF
C9646 VN.n8708 a_400_62400# 2.51fF
C9647 VN.t1669 a_400_62400# 0.03fF
C9648 VN.n8709 a_400_62400# 0.32fF
C9649 VN.n8710 a_400_62400# 0.48fF
C9650 VN.n8711 a_400_62400# 0.81fF
C9651 VN.n8712 a_400_62400# 0.16fF
C9652 VN.t548 a_400_62400# 0.03fF
C9653 VN.n8713 a_400_62400# 0.19fF
C9654 VN.n8715 a_400_62400# 1.55fF
C9655 VN.n8716 a_400_62400# 0.29fF
C9656 VN.n8717 a_400_62400# 2.52fF
C9657 VN.t828 a_400_62400# 0.03fF
C9658 VN.n8718 a_400_62400# 0.32fF
C9659 VN.n8719 a_400_62400# 1.22fF
C9660 VN.n8720 a_400_62400# 0.07fF
C9661 VN.t732 a_400_62400# 0.03fF
C9662 VN.n8721 a_400_62400# 0.16fF
C9663 VN.n8722 a_400_62400# 0.19fF
C9664 VN.n8724 a_400_62400# 1.04fF
C9665 VN.n8725 a_400_62400# 2.60fF
C9666 VN.n8726 a_400_62400# 2.51fF
C9667 VN.n8727 a_400_62400# 0.16fF
C9668 VN.t1005 a_400_62400# 0.03fF
C9669 VN.n8728 a_400_62400# 0.19fF
C9670 VN.t2167 a_400_62400# 0.03fF
C9671 VN.n8730 a_400_62400# 0.32fF
C9672 VN.n8731 a_400_62400# 0.48fF
C9673 VN.n8732 a_400_62400# 0.81fF
C9674 VN.n8733 a_400_62400# 2.46fF
C9675 VN.n8734 a_400_62400# 4.01fF
C9676 VN.t1332 a_400_62400# 0.03fF
C9677 VN.n8735 a_400_62400# 0.32fF
C9678 VN.n8736 a_400_62400# 1.22fF
C9679 VN.n8737 a_400_62400# 0.07fF
C9680 VN.t1213 a_400_62400# 0.03fF
C9681 VN.n8738 a_400_62400# 0.16fF
C9682 VN.n8739 a_400_62400# 0.19fF
C9683 VN.n8741 a_400_62400# 2.53fF
C9684 VN.n8742 a_400_62400# 2.51fF
C9685 VN.t1301 a_400_62400# 0.03fF
C9686 VN.n8743 a_400_62400# 0.32fF
C9687 VN.n8744 a_400_62400# 0.48fF
C9688 VN.n8745 a_400_62400# 0.81fF
C9689 VN.n8746 a_400_62400# 0.16fF
C9690 VN.t128 a_400_62400# 0.03fF
C9691 VN.n8747 a_400_62400# 0.19fF
C9692 VN.n8749 a_400_62400# 1.55fF
C9693 VN.n8750 a_400_62400# 0.29fF
C9694 VN.n8751 a_400_62400# 2.52fF
C9695 VN.t470 a_400_62400# 0.03fF
C9696 VN.n8752 a_400_62400# 0.32fF
C9697 VN.n8753 a_400_62400# 1.22fF
C9698 VN.n8754 a_400_62400# 0.07fF
C9699 VN.t352 a_400_62400# 0.03fF
C9700 VN.n8755 a_400_62400# 0.16fF
C9701 VN.n8756 a_400_62400# 0.19fF
C9702 VN.n8758 a_400_62400# 1.04fF
C9703 VN.n8759 a_400_62400# 2.60fF
C9704 VN.n8760 a_400_62400# 2.51fF
C9705 VN.n8761 a_400_62400# 0.16fF
C9706 VN.t1927 a_400_62400# 0.03fF
C9707 VN.n8762 a_400_62400# 0.19fF
C9708 VN.t435 a_400_62400# 0.03fF
C9709 VN.n8764 a_400_62400# 0.32fF
C9710 VN.n8765 a_400_62400# 0.48fF
C9711 VN.n8766 a_400_62400# 0.81fF
C9712 VN.n8767 a_400_62400# 2.46fF
C9713 VN.n8768 a_400_62400# 4.01fF
C9714 VN.t2122 a_400_62400# 0.03fF
C9715 VN.n8769 a_400_62400# 0.32fF
C9716 VN.n8770 a_400_62400# 1.22fF
C9717 VN.n8771 a_400_62400# 0.07fF
C9718 VN.t1997 a_400_62400# 0.03fF
C9719 VN.n8772 a_400_62400# 0.16fF
C9720 VN.n8773 a_400_62400# 0.19fF
C9721 VN.n8775 a_400_62400# 2.53fF
C9722 VN.n8776 a_400_62400# 2.51fF
C9723 VN.t2210 a_400_62400# 0.03fF
C9724 VN.n8777 a_400_62400# 0.32fF
C9725 VN.n8778 a_400_62400# 0.48fF
C9726 VN.n8779 a_400_62400# 0.81fF
C9727 VN.n8780 a_400_62400# 0.16fF
C9728 VN.t1052 a_400_62400# 0.03fF
C9729 VN.n8781 a_400_62400# 0.19fF
C9730 VN.n8783 a_400_62400# 1.55fF
C9731 VN.n8784 a_400_62400# 0.29fF
C9732 VN.n8785 a_400_62400# 2.52fF
C9733 VN.t1378 a_400_62400# 0.03fF
C9734 VN.n8786 a_400_62400# 0.32fF
C9735 VN.n8787 a_400_62400# 1.22fF
C9736 VN.n8788 a_400_62400# 0.07fF
C9737 VN.t1123 a_400_62400# 0.03fF
C9738 VN.n8789 a_400_62400# 0.16fF
C9739 VN.n8790 a_400_62400# 0.19fF
C9740 VN.n8792 a_400_62400# 1.04fF
C9741 VN.n8793 a_400_62400# 2.60fF
C9742 VN.n8794 a_400_62400# 2.51fF
C9743 VN.n8795 a_400_62400# 0.16fF
C9744 VN.t181 a_400_62400# 0.03fF
C9745 VN.n8796 a_400_62400# 0.19fF
C9746 VN.t1344 a_400_62400# 0.03fF
C9747 VN.n8798 a_400_62400# 0.32fF
C9748 VN.n8799 a_400_62400# 0.48fF
C9749 VN.n8800 a_400_62400# 0.81fF
C9750 VN.n8801 a_400_62400# 2.46fF
C9751 VN.n8802 a_400_62400# 4.01fF
C9752 VN.t513 a_400_62400# 0.03fF
C9753 VN.n8803 a_400_62400# 0.32fF
C9754 VN.n8804 a_400_62400# 1.22fF
C9755 VN.n8805 a_400_62400# 0.07fF
C9756 VN.t260 a_400_62400# 0.03fF
C9757 VN.n8806 a_400_62400# 0.16fF
C9758 VN.n8807 a_400_62400# 0.19fF
C9759 VN.n8809 a_400_62400# 2.53fF
C9760 VN.n8810 a_400_62400# 2.34fF
C9761 VN.t480 a_400_62400# 0.03fF
C9762 VN.n8811 a_400_62400# 0.32fF
C9763 VN.n8812 a_400_62400# 0.48fF
C9764 VN.n8813 a_400_62400# 0.81fF
C9765 VN.n8814 a_400_62400# 0.16fF
C9766 VN.t1839 a_400_62400# 0.03fF
C9767 VN.n8815 a_400_62400# 0.19fF
C9768 VN.n8817 a_400_62400# 1.55fF
C9769 VN.n8818 a_400_62400# 0.29fF
C9770 VN.n8819 a_400_62400# 3.27fF
C9771 VN.t2166 a_400_62400# 0.03fF
C9772 VN.n8820 a_400_62400# 0.32fF
C9773 VN.n8821 a_400_62400# 1.22fF
C9774 VN.n8822 a_400_62400# 0.07fF
C9775 VN.t1909 a_400_62400# 0.03fF
C9776 VN.n8823 a_400_62400# 0.16fF
C9777 VN.n8824 a_400_62400# 0.19fF
C9778 VN.n8826 a_400_62400# 2.51fF
C9779 VN.n8827 a_400_62400# 0.56fF
C9780 VN.n8828 a_400_62400# 0.64fF
C9781 VN.n8829 a_400_62400# 0.12fF
C9782 VN.n8830 a_400_62400# 0.44fF
C9783 VN.n8831 a_400_62400# 0.40fF
C9784 VN.n8832 a_400_62400# 1.03fF
C9785 VN.n8833 a_400_62400# 0.79fF
C9786 VN.t2135 a_400_62400# 0.03fF
C9787 VN.n8834 a_400_62400# 0.32fF
C9788 VN.n8835 a_400_62400# 0.48fF
C9789 VN.n8836 a_400_62400# 0.81fF
C9790 VN.n8837 a_400_62400# 0.16fF
C9791 VN.t967 a_400_62400# 0.03fF
C9792 VN.n8838 a_400_62400# 0.19fF
C9793 VN.n8840 a_400_62400# 3.50fF
C9794 VN.n8841 a_400_62400# 2.89fF
C9795 VN.t1300 a_400_62400# 0.03fF
C9796 VN.n8842 a_400_62400# 0.32fF
C9797 VN.n8843 a_400_62400# 1.22fF
C9798 VN.n8844 a_400_62400# 0.07fF
C9799 VN.t1034 a_400_62400# 0.03fF
C9800 VN.n8845 a_400_62400# 0.16fF
C9801 VN.n8846 a_400_62400# 0.19fF
C9802 VN.n8848 a_400_62400# 1.05fF
C9803 VN.n8849 a_400_62400# 3.07fF
C9804 VN.n8850 a_400_62400# 2.51fF
C9805 VN.n8851 a_400_62400# 0.16fF
C9806 VN.t65 a_400_62400# 0.03fF
C9807 VN.n8852 a_400_62400# 0.19fF
C9808 VN.t1260 a_400_62400# 0.03fF
C9809 VN.n8854 a_400_62400# 0.32fF
C9810 VN.n8855 a_400_62400# 0.48fF
C9811 VN.n8856 a_400_62400# 0.81fF
C9812 VN.n8857 a_400_62400# 1.86fF
C9813 VN.n8858 a_400_62400# 1.53fF
C9814 VN.n8859 a_400_62400# 0.47fF
C9815 VN.n8860 a_400_62400# 2.71fF
C9816 VN.t434 a_400_62400# 0.03fF
C9817 VN.n8861 a_400_62400# 0.32fF
C9818 VN.n8862 a_400_62400# 1.22fF
C9819 VN.n8863 a_400_62400# 0.07fF
C9820 VN.t309 a_400_62400# 0.03fF
C9821 VN.n8864 a_400_62400# 0.16fF
C9822 VN.n8865 a_400_62400# 0.19fF
C9823 VN.n8867 a_400_62400# 2.53fF
C9824 VN.n8868 a_400_62400# 2.51fF
C9825 VN.t392 a_400_62400# 0.03fF
C9826 VN.n8869 a_400_62400# 0.32fF
C9827 VN.n8870 a_400_62400# 0.48fF
C9828 VN.n8871 a_400_62400# 0.81fF
C9829 VN.n8872 a_400_62400# 0.16fF
C9830 VN.t1756 a_400_62400# 0.03fF
C9831 VN.n8873 a_400_62400# 0.19fF
C9832 VN.n8875 a_400_62400# 1.55fF
C9833 VN.n8876 a_400_62400# 0.29fF
C9834 VN.n8877 a_400_62400# 2.52fF
C9835 VN.t2081 a_400_62400# 0.03fF
C9836 VN.n8878 a_400_62400# 0.32fF
C9837 VN.n8879 a_400_62400# 1.22fF
C9838 VN.n8880 a_400_62400# 0.07fF
C9839 VN.t1958 a_400_62400# 0.03fF
C9840 VN.n8881 a_400_62400# 0.16fF
C9841 VN.n8882 a_400_62400# 0.19fF
C9842 VN.n8884 a_400_62400# 27.83fF
C9843 VN.n8885 a_400_62400# 3.93fF
C9844 VN.n8886 a_400_62400# 2.51fF
C9845 VN.n8887 a_400_62400# 0.16fF
C9846 VN.t40 a_400_62400# 0.03fF
C9847 VN.n8888 a_400_62400# 0.19fF
C9848 VN.t1261 a_400_62400# 0.03fF
C9849 VN.n8890 a_400_62400# 0.32fF
C9850 VN.n8891 a_400_62400# 0.48fF
C9851 VN.n8892 a_400_62400# 0.81fF
C9852 VN.n8893 a_400_62400# 1.46fF
C9853 VN.n8894 a_400_62400# 0.21fF
C9854 VN.n8895 a_400_62400# 2.81fF
C9855 VN.t298 a_400_62400# 0.03fF
C9856 VN.n8896 a_400_62400# 0.16fF
C9857 VN.n8897 a_400_62400# 0.19fF
C9858 VN.t532 a_400_62400# 0.03fF
C9859 VN.n8899 a_400_62400# 0.32fF
C9860 VN.n8900 a_400_62400# 1.22fF
C9861 VN.n8901 a_400_62400# 0.07fF
C9862 VN.n8902 a_400_62400# 2.51fF
C9863 VN.n8903 a_400_62400# 3.57fF
C9864 VN.t393 a_400_62400# 0.03fF
C9865 VN.n8904 a_400_62400# 0.32fF
C9866 VN.n8905 a_400_62400# 0.48fF
C9867 VN.n8906 a_400_62400# 0.81fF
C9868 VN.n8907 a_400_62400# 0.16fF
C9869 VN.t1742 a_400_62400# 0.03fF
C9870 VN.n8908 a_400_62400# 0.19fF
C9871 VN.n8910 a_400_62400# 3.93fF
C9872 VN.n8911 a_400_62400# 3.08fF
C9873 VN.t1947 a_400_62400# 0.03fF
C9874 VN.n8912 a_400_62400# 0.16fF
C9875 VN.n8913 a_400_62400# 0.19fF
C9876 VN.t2186 a_400_62400# 0.03fF
C9877 VN.n8915 a_400_62400# 0.32fF
C9878 VN.n8916 a_400_62400# 1.22fF
C9879 VN.n8917 a_400_62400# 0.07fF
C9880 VN.n8918 a_400_62400# 3.65fF
C9881 VN.n8919 a_400_62400# 2.14fF
C9882 VN.n8920 a_400_62400# 0.16fF
C9883 VN.t124 a_400_62400# 0.03fF
C9884 VN.n8921 a_400_62400# 0.19fF
C9885 VN.t1175 a_400_62400# 0.03fF
C9886 VN.n8923 a_400_62400# 0.32fF
C9887 VN.n8924 a_400_62400# 0.48fF
C9888 VN.n8925 a_400_62400# 0.81fF
C9889 VN.n8926 a_400_62400# 0.09fF
C9890 VN.n8927 a_400_62400# 0.01fF
C9891 VN.n8928 a_400_62400# 0.02fF
C9892 VN.n8929 a_400_62400# 0.02fF
C9893 VN.n8930 a_400_62400# 0.32fF
C9894 VN.n8931 a_400_62400# 1.56fF
C9895 VN.n8932 a_400_62400# 1.81fF
C9896 VN.n8933 a_400_62400# 3.08fF
C9897 VN.t203 a_400_62400# 0.03fF
C9898 VN.n8934 a_400_62400# 0.16fF
C9899 VN.n8935 a_400_62400# 0.19fF
C9900 VN.t459 a_400_62400# 0.03fF
C9901 VN.n8937 a_400_62400# 0.32fF
C9902 VN.n8938 a_400_62400# 1.22fF
C9903 VN.n8939 a_400_62400# 0.07fF
C9904 VN.t39 a_400_62400# 64.69fF
C9905 VN.t1321 a_400_62400# 0.03fF
C9906 VN.n8940 a_400_62400# 0.32fF
C9907 VN.n8941 a_400_62400# 1.22fF
C9908 VN.n8942 a_400_62400# 0.07fF
C9909 VN.t1078 a_400_62400# 0.03fF
C9910 VN.n8943 a_400_62400# 0.16fF
C9911 VN.n8944 a_400_62400# 0.19fF
C9912 VN.n8946 a_400_62400# 0.16fF
C9913 VN.t870 a_400_62400# 0.03fF
C9914 VN.n8947 a_400_62400# 0.19fF
C9915 VN.n8949 a_400_62400# 6.92fF
C9916 VN.n8950 a_400_62400# 6.56fF
C9917 VN.t2420 a_400_62400# 0.03fF
C9918 VN.n8951 a_400_62400# 0.16fF
C9919 VN.n8952 a_400_62400# 0.19fF
C9920 VN.t2240 a_400_62400# 0.03fF
C9921 VN.n8954 a_400_62400# 0.32fF
C9922 VN.n8955 a_400_62400# 1.22fF
C9923 VN.n8956 a_400_62400# 0.07fF
C9924 VN.n8957 a_400_62400# 2.51fF
C9925 VN.n8958 a_400_62400# 3.58fF
C9926 VN.t2035 a_400_62400# 0.03fF
C9927 VN.n8959 a_400_62400# 0.32fF
C9928 VN.n8960 a_400_62400# 0.48fF
C9929 VN.n8961 a_400_62400# 0.81fF
C9930 VN.n8962 a_400_62400# 0.16fF
C9931 VN.t865 a_400_62400# 0.03fF
C9932 VN.n8963 a_400_62400# 0.19fF
C9933 VN.n8965 a_400_62400# 7.29fF
C9934 VN.t1558 a_400_62400# 0.03fF
C9935 VN.n8966 a_400_62400# 0.16fF
C9936 VN.n8967 a_400_62400# 0.19fF
C9937 VN.t1375 a_400_62400# 0.03fF
C9938 VN.n8969 a_400_62400# 0.32fF
C9939 VN.n8970 a_400_62400# 1.22fF
C9940 VN.n8971 a_400_62400# 0.07fF
C9941 VN.t26 a_400_62400# 64.17fF
C9942 VN.t509 a_400_62400# 0.03fF
C9943 VN.n8972 a_400_62400# 1.60fF
C9944 VN.n8973 a_400_62400# 0.07fF
C9945 VN.t808 a_400_62400# 0.03fF
C9946 VN.n8974 a_400_62400# 0.02fF
C9947 VN.n8975 a_400_62400# 0.34fF
C9948 VN.n8977 a_400_62400# 2.01fF
C9949 VN.n8978 a_400_62400# 1.75fF
C9950 VN.n8979 a_400_62400# 0.37fF
C9951 VN.n8980 a_400_62400# 0.33fF
C9952 VN.n8981 a_400_62400# 5.88fF
C9953 VN.n8982 a_400_62400# 0.02fF
C9954 VN.n8983 a_400_62400# 0.02fF
C9955 VN.n8984 a_400_62400# 0.03fF
C9956 VN.n8985 a_400_62400# 0.05fF
C9957 VN.n8986 a_400_62400# 0.23fF
C9958 VN.n8987 a_400_62400# 0.02fF
C9959 VN.n8988 a_400_62400# 0.03fF
C9960 VN.n8989 a_400_62400# 0.01fF
C9961 VN.n8990 a_400_62400# 0.01fF
C9962 VN.n8991 a_400_62400# 0.01fF
C9963 VN.n8992 a_400_62400# 0.02fF
C9964 VN.n8993 a_400_62400# 0.03fF
C9965 VN.n8994 a_400_62400# 0.06fF
C9966 VN.n8995 a_400_62400# 0.05fF
C9967 VN.n8996 a_400_62400# 0.15fF
C9968 VN.n8997 a_400_62400# 0.51fF
C9969 VN.n8998 a_400_62400# 0.27fF
C9970 VN.n8999 a_400_62400# 37.46fF
C9971 VN.n9000 a_400_62400# 37.46fF
C9972 VN.n9001 a_400_62400# 0.79fF
C9973 VN.n9002 a_400_62400# 0.23fF
C9974 VN.n9003 a_400_62400# 1.18fF
C9975 VN.t90 a_400_62400# 28.64fF
C9976 VN.n9004 a_400_62400# 0.79fF
C9977 VN.n9005 a_400_62400# 0.11fF
C9978 VN.n9006 a_400_62400# 4.98fF
C9979 VN.n9007 a_400_62400# 0.80fF
C9980 VN.n9008 a_400_62400# 0.29fF
C9981 VN.n9009 a_400_62400# 1.96fF
C9982 VN.n9011 a_400_62400# 25.18fF
C9983 VN.n9013 a_400_62400# 1.87fF
C9984 VN.n9014 a_400_62400# 5.36fF
C9985 VN.n9015 a_400_62400# 1.81fF
C9986 VN.t2295 a_400_62400# 0.03fF
C9987 VN.n9016 a_400_62400# 0.85fF
C9988 VN.n9017 a_400_62400# 0.81fF
C9989 VN.n9018 a_400_62400# 0.33fF
C9990 VN.n9019 a_400_62400# 0.12fF
C9991 VN.n9020 a_400_62400# 0.28fF
C9992 VN.n9021 a_400_62400# 1.23fF
C9993 VN.n9022 a_400_62400# 0.59fF
C9994 VN.n9023 a_400_62400# 2.51fF
C9995 VN.n9024 a_400_62400# 0.16fF
C9996 VN.t1634 a_400_62400# 0.03fF
C9997 VN.n9025 a_400_62400# 0.19fF
C9998 VN.t91 a_400_62400# 0.03fF
C9999 VN.n9027 a_400_62400# 0.32fF
C10000 VN.n9028 a_400_62400# 0.48fF
C10001 VN.n9029 a_400_62400# 0.81fF
C10002 VN.n9030 a_400_62400# 0.03fF
C10003 VN.n9031 a_400_62400# 0.01fF
C10004 VN.n9032 a_400_62400# 0.02fF
C10005 VN.n9033 a_400_62400# 0.11fF
C10006 VN.n9034 a_400_62400# 0.08fF
C10007 VN.n9035 a_400_62400# 0.04fF
C10008 VN.n9036 a_400_62400# 0.05fF
C10009 VN.n9037 a_400_62400# 1.34fF
C10010 VN.n9038 a_400_62400# 0.48fF
C10011 VN.n9039 a_400_62400# 2.51fF
C10012 VN.n9040 a_400_62400# 2.67fF
C10013 VN.t1251 a_400_62400# 0.03fF
C10014 VN.n9041 a_400_62400# 0.32fF
C10015 VN.n9042 a_400_62400# 1.22fF
C10016 VN.n9043 a_400_62400# 0.07fF
C10017 VN.t2315 a_400_62400# 0.03fF
C10018 VN.n9044 a_400_62400# 0.16fF
C10019 VN.n9045 a_400_62400# 0.19fF
C10020 VN.n9047 a_400_62400# 2.53fF
C10021 VN.n9048 a_400_62400# 0.08fF
C10022 VN.n9049 a_400_62400# 0.04fF
C10023 VN.n9050 a_400_62400# 0.05fF
C10024 VN.n9051 a_400_62400# 1.33fF
C10025 VN.n9052 a_400_62400# 0.03fF
C10026 VN.n9053 a_400_62400# 0.01fF
C10027 VN.n9054 a_400_62400# 0.02fF
C10028 VN.n9055 a_400_62400# 0.11fF
C10029 VN.n9056 a_400_62400# 0.48fF
C10030 VN.n9057 a_400_62400# 2.48fF
C10031 VN.t1893 a_400_62400# 0.03fF
C10032 VN.n9058 a_400_62400# 0.32fF
C10033 VN.n9059 a_400_62400# 0.48fF
C10034 VN.n9060 a_400_62400# 0.81fF
C10035 VN.n9061 a_400_62400# 0.16fF
C10036 VN.t762 a_400_62400# 0.03fF
C10037 VN.n9062 a_400_62400# 0.19fF
C10038 VN.n9064 a_400_62400# 0.93fF
C10039 VN.n9065 a_400_62400# 0.30fF
C10040 VN.n9066 a_400_62400# 0.34fF
C10041 VN.n9067 a_400_62400# 0.12fF
C10042 VN.n9068 a_400_62400# 0.30fF
C10043 VN.n9069 a_400_62400# 0.93fF
C10044 VN.n9070 a_400_62400# 1.55fF
C10045 VN.n9071 a_400_62400# 0.29fF
C10046 VN.n9072 a_400_62400# 0.34fF
C10047 VN.n9073 a_400_62400# 0.12fF
C10048 VN.n9074 a_400_62400# 2.52fF
C10049 VN.t517 a_400_62400# 0.03fF
C10050 VN.n9075 a_400_62400# 0.32fF
C10051 VN.n9076 a_400_62400# 1.22fF
C10052 VN.n9077 a_400_62400# 0.07fF
C10053 VN.t1445 a_400_62400# 0.03fF
C10054 VN.n9078 a_400_62400# 0.16fF
C10055 VN.n9079 a_400_62400# 0.19fF
C10056 VN.n9081 a_400_62400# 0.33fF
C10057 VN.n9082 a_400_62400# 0.12fF
C10058 VN.n9083 a_400_62400# 0.28fF
C10059 VN.n9084 a_400_62400# 1.72fF
C10060 VN.n9085 a_400_62400# 0.71fF
C10061 VN.n9086 a_400_62400# 2.51fF
C10062 VN.n9087 a_400_62400# 0.16fF
C10063 VN.t2417 a_400_62400# 0.03fF
C10064 VN.n9088 a_400_62400# 0.19fF
C10065 VN.t1020 a_400_62400# 0.03fF
C10066 VN.n9090 a_400_62400# 0.32fF
C10067 VN.n9091 a_400_62400# 0.48fF
C10068 VN.n9092 a_400_62400# 0.81fF
C10069 VN.n9093 a_400_62400# 0.03fF
C10070 VN.n9094 a_400_62400# 0.01fF
C10071 VN.n9095 a_400_62400# 0.02fF
C10072 VN.n9096 a_400_62400# 0.11fF
C10073 VN.n9097 a_400_62400# 0.08fF
C10074 VN.n9098 a_400_62400# 0.04fF
C10075 VN.n9099 a_400_62400# 0.05fF
C10076 VN.n9100 a_400_62400# 1.34fF
C10077 VN.n9101 a_400_62400# 0.48fF
C10078 VN.n9102 a_400_62400# 2.51fF
C10079 VN.n9103 a_400_62400# 2.67fF
C10080 VN.t2168 a_400_62400# 0.03fF
C10081 VN.n9104 a_400_62400# 0.32fF
C10082 VN.n9105 a_400_62400# 1.22fF
C10083 VN.n9106 a_400_62400# 0.07fF
C10084 VN.t576 a_400_62400# 0.03fF
C10085 VN.n9107 a_400_62400# 0.16fF
C10086 VN.n9108 a_400_62400# 0.19fF
C10087 VN.n9110 a_400_62400# 2.53fF
C10088 VN.n9111 a_400_62400# 0.08fF
C10089 VN.n9112 a_400_62400# 0.04fF
C10090 VN.n9113 a_400_62400# 0.05fF
C10091 VN.n9114 a_400_62400# 1.33fF
C10092 VN.n9115 a_400_62400# 0.03fF
C10093 VN.n9116 a_400_62400# 0.01fF
C10094 VN.n9117 a_400_62400# 0.02fF
C10095 VN.n9118 a_400_62400# 0.11fF
C10096 VN.n9119 a_400_62400# 0.48fF
C10097 VN.n9120 a_400_62400# 2.48fF
C10098 VN.t1516 a_400_62400# 0.03fF
C10099 VN.n9121 a_400_62400# 0.32fF
C10100 VN.n9122 a_400_62400# 0.48fF
C10101 VN.n9123 a_400_62400# 0.81fF
C10102 VN.n9124 a_400_62400# 0.16fF
C10103 VN.t386 a_400_62400# 0.03fF
C10104 VN.n9125 a_400_62400# 0.19fF
C10105 VN.n9127 a_400_62400# 0.93fF
C10106 VN.n9128 a_400_62400# 0.30fF
C10107 VN.n9129 a_400_62400# 0.34fF
C10108 VN.n9130 a_400_62400# 0.12fF
C10109 VN.n9131 a_400_62400# 0.30fF
C10110 VN.n9132 a_400_62400# 0.93fF
C10111 VN.n9133 a_400_62400# 1.55fF
C10112 VN.n9134 a_400_62400# 0.29fF
C10113 VN.n9135 a_400_62400# 0.34fF
C10114 VN.n9136 a_400_62400# 0.12fF
C10115 VN.n9137 a_400_62400# 2.52fF
C10116 VN.t67 a_400_62400# 0.03fF
C10117 VN.n9138 a_400_62400# 0.32fF
C10118 VN.n9139 a_400_62400# 1.22fF
C10119 VN.n9140 a_400_62400# 0.07fF
C10120 VN.t2234 a_400_62400# 0.03fF
C10121 VN.n9141 a_400_62400# 0.16fF
C10122 VN.n9142 a_400_62400# 0.19fF
C10123 VN.n9144 a_400_62400# 0.33fF
C10124 VN.n9145 a_400_62400# 0.12fF
C10125 VN.n9146 a_400_62400# 0.28fF
C10126 VN.n9147 a_400_62400# 1.23fF
C10127 VN.n9148 a_400_62400# 0.59fF
C10128 VN.n9149 a_400_62400# 2.51fF
C10129 VN.n9150 a_400_62400# 0.16fF
C10130 VN.t2040 a_400_62400# 0.03fF
C10131 VN.n9151 a_400_62400# 0.19fF
C10132 VN.t648 a_400_62400# 0.03fF
C10133 VN.n9153 a_400_62400# 0.32fF
C10134 VN.n9154 a_400_62400# 0.48fF
C10135 VN.n9155 a_400_62400# 0.81fF
C10136 VN.n9156 a_400_62400# 0.03fF
C10137 VN.n9157 a_400_62400# 0.01fF
C10138 VN.n9158 a_400_62400# 0.02fF
C10139 VN.n9159 a_400_62400# 0.11fF
C10140 VN.n9160 a_400_62400# 0.08fF
C10141 VN.n9161 a_400_62400# 0.04fF
C10142 VN.n9162 a_400_62400# 0.05fF
C10143 VN.n9163 a_400_62400# 1.34fF
C10144 VN.n9164 a_400_62400# 0.48fF
C10145 VN.n9165 a_400_62400# 2.51fF
C10146 VN.n9166 a_400_62400# 2.67fF
C10147 VN.t1757 a_400_62400# 0.03fF
C10148 VN.n9167 a_400_62400# 0.32fF
C10149 VN.n9168 a_400_62400# 1.22fF
C10150 VN.n9169 a_400_62400# 0.07fF
C10151 VN.t171 a_400_62400# 0.03fF
C10152 VN.n9170 a_400_62400# 0.16fF
C10153 VN.n9171 a_400_62400# 0.19fF
C10154 VN.n9173 a_400_62400# 2.53fF
C10155 VN.n9174 a_400_62400# 0.08fF
C10156 VN.n9175 a_400_62400# 0.04fF
C10157 VN.n9176 a_400_62400# 0.05fF
C10158 VN.n9177 a_400_62400# 1.33fF
C10159 VN.n9178 a_400_62400# 0.03fF
C10160 VN.n9179 a_400_62400# 0.01fF
C10161 VN.n9180 a_400_62400# 0.02fF
C10162 VN.n9181 a_400_62400# 0.11fF
C10163 VN.n9182 a_400_62400# 0.48fF
C10164 VN.n9183 a_400_62400# 2.48fF
C10165 VN.t2307 a_400_62400# 0.03fF
C10166 VN.n9184 a_400_62400# 0.32fF
C10167 VN.n9185 a_400_62400# 0.48fF
C10168 VN.n9186 a_400_62400# 0.81fF
C10169 VN.n9187 a_400_62400# 0.16fF
C10170 VN.t1168 a_400_62400# 0.03fF
C10171 VN.n9188 a_400_62400# 0.19fF
C10172 VN.n9190 a_400_62400# 0.93fF
C10173 VN.n9191 a_400_62400# 0.30fF
C10174 VN.n9192 a_400_62400# 0.34fF
C10175 VN.n9193 a_400_62400# 0.12fF
C10176 VN.n9194 a_400_62400# 0.30fF
C10177 VN.n9195 a_400_62400# 0.93fF
C10178 VN.n9196 a_400_62400# 1.55fF
C10179 VN.n9197 a_400_62400# 0.29fF
C10180 VN.n9198 a_400_62400# 0.34fF
C10181 VN.n9199 a_400_62400# 0.12fF
C10182 VN.n9200 a_400_62400# 2.52fF
C10183 VN.t884 a_400_62400# 0.03fF
C10184 VN.n9201 a_400_62400# 0.32fF
C10185 VN.n9202 a_400_62400# 1.22fF
C10186 VN.n9203 a_400_62400# 0.07fF
C10187 VN.t1832 a_400_62400# 0.03fF
C10188 VN.n9204 a_400_62400# 0.16fF
C10189 VN.n9205 a_400_62400# 0.19fF
C10190 VN.n9207 a_400_62400# 0.33fF
C10191 VN.n9208 a_400_62400# 0.12fF
C10192 VN.n9209 a_400_62400# 0.28fF
C10193 VN.n9210 a_400_62400# 1.23fF
C10194 VN.n9211 a_400_62400# 0.59fF
C10195 VN.n9212 a_400_62400# 2.51fF
C10196 VN.n9213 a_400_62400# 0.16fF
C10197 VN.t299 a_400_62400# 0.03fF
C10198 VN.n9214 a_400_62400# 0.19fF
C10199 VN.t1437 a_400_62400# 0.03fF
C10200 VN.n9216 a_400_62400# 0.32fF
C10201 VN.n9217 a_400_62400# 0.48fF
C10202 VN.n9218 a_400_62400# 0.81fF
C10203 VN.n9219 a_400_62400# 0.03fF
C10204 VN.n9220 a_400_62400# 0.01fF
C10205 VN.n9221 a_400_62400# 0.02fF
C10206 VN.n9222 a_400_62400# 0.11fF
C10207 VN.n9223 a_400_62400# 0.08fF
C10208 VN.n9224 a_400_62400# 0.04fF
C10209 VN.n9225 a_400_62400# 0.05fF
C10210 VN.n9226 a_400_62400# 1.34fF
C10211 VN.n9227 a_400_62400# 0.48fF
C10212 VN.n9228 a_400_62400# 2.51fF
C10213 VN.n9229 a_400_62400# 2.67fF
C10214 VN.t2545 a_400_62400# 0.03fF
C10215 VN.n9230 a_400_62400# 0.32fF
C10216 VN.n9231 a_400_62400# 1.22fF
C10217 VN.n9232 a_400_62400# 0.07fF
C10218 VN.t1093 a_400_62400# 0.03fF
C10219 VN.n9233 a_400_62400# 0.16fF
C10220 VN.n9234 a_400_62400# 0.19fF
C10221 VN.n9236 a_400_62400# 2.53fF
C10222 VN.n9237 a_400_62400# 0.08fF
C10223 VN.n9238 a_400_62400# 0.04fF
C10224 VN.n9239 a_400_62400# 0.05fF
C10225 VN.n9240 a_400_62400# 1.33fF
C10226 VN.n9241 a_400_62400# 0.03fF
C10227 VN.n9242 a_400_62400# 0.01fF
C10228 VN.n9243 a_400_62400# 0.02fF
C10229 VN.n9244 a_400_62400# 0.11fF
C10230 VN.n9245 a_400_62400# 0.48fF
C10231 VN.n9246 a_400_62400# 2.48fF
C10232 VN.t570 a_400_62400# 0.03fF
C10233 VN.n9247 a_400_62400# 0.32fF
C10234 VN.n9248 a_400_62400# 0.48fF
C10235 VN.n9249 a_400_62400# 0.81fF
C10236 VN.n9250 a_400_62400# 0.16fF
C10237 VN.t1948 a_400_62400# 0.03fF
C10238 VN.n9251 a_400_62400# 0.19fF
C10239 VN.n9253 a_400_62400# 0.93fF
C10240 VN.n9254 a_400_62400# 0.30fF
C10241 VN.n9255 a_400_62400# 0.34fF
C10242 VN.n9256 a_400_62400# 0.12fF
C10243 VN.n9257 a_400_62400# 0.30fF
C10244 VN.n9258 a_400_62400# 0.93fF
C10245 VN.n9259 a_400_62400# 1.55fF
C10246 VN.n9260 a_400_62400# 0.29fF
C10247 VN.n9261 a_400_62400# 0.34fF
C10248 VN.n9262 a_400_62400# 0.12fF
C10249 VN.n9263 a_400_62400# 2.52fF
C10250 VN.t1679 a_400_62400# 0.03fF
C10251 VN.n9264 a_400_62400# 0.32fF
C10252 VN.n9265 a_400_62400# 1.22fF
C10253 VN.n9266 a_400_62400# 0.07fF
C10254 VN.t223 a_400_62400# 0.03fF
C10255 VN.n9267 a_400_62400# 0.16fF
C10256 VN.n9268 a_400_62400# 0.19fF
C10257 VN.n9270 a_400_62400# 0.33fF
C10258 VN.n9271 a_400_62400# 0.12fF
C10259 VN.n9272 a_400_62400# 0.28fF
C10260 VN.n9273 a_400_62400# 1.23fF
C10261 VN.n9274 a_400_62400# 0.59fF
C10262 VN.n9275 a_400_62400# 2.51fF
C10263 VN.n9276 a_400_62400# 0.16fF
C10264 VN.t1079 a_400_62400# 0.03fF
C10265 VN.n9277 a_400_62400# 0.19fF
C10266 VN.t2229 a_400_62400# 0.03fF
C10267 VN.n9279 a_400_62400# 0.32fF
C10268 VN.n9280 a_400_62400# 0.48fF
C10269 VN.n9281 a_400_62400# 0.81fF
C10270 VN.n9282 a_400_62400# 0.03fF
C10271 VN.n9283 a_400_62400# 0.01fF
C10272 VN.n9284 a_400_62400# 0.02fF
C10273 VN.n9285 a_400_62400# 0.11fF
C10274 VN.n9286 a_400_62400# 0.08fF
C10275 VN.n9287 a_400_62400# 0.04fF
C10276 VN.n9288 a_400_62400# 0.05fF
C10277 VN.n9289 a_400_62400# 1.34fF
C10278 VN.n9290 a_400_62400# 0.48fF
C10279 VN.n9291 a_400_62400# 2.51fF
C10280 VN.n9292 a_400_62400# 2.67fF
C10281 VN.t812 a_400_62400# 0.03fF
C10282 VN.n9293 a_400_62400# 0.32fF
C10283 VN.n9294 a_400_62400# 1.22fF
C10284 VN.n9295 a_400_62400# 0.07fF
C10285 VN.t1872 a_400_62400# 0.03fF
C10286 VN.n9296 a_400_62400# 0.16fF
C10287 VN.n9297 a_400_62400# 0.19fF
C10288 VN.n9299 a_400_62400# 2.53fF
C10289 VN.n9300 a_400_62400# 0.09fF
C10290 VN.n9301 a_400_62400# 0.05fF
C10291 VN.n9302 a_400_62400# 0.07fF
C10292 VN.n9303 a_400_62400# 1.16fF
C10293 VN.n9304 a_400_62400# 0.01fF
C10294 VN.n9305 a_400_62400# 0.01fF
C10295 VN.n9306 a_400_62400# 0.01fF
C10296 VN.n9307 a_400_62400# 0.09fF
C10297 VN.n9308 a_400_62400# 0.91fF
C10298 VN.n9309 a_400_62400# 0.96fF
C10299 VN.t1364 a_400_62400# 0.03fF
C10300 VN.n9310 a_400_62400# 0.32fF
C10301 VN.n9311 a_400_62400# 0.48fF
C10302 VN.n9312 a_400_62400# 0.81fF
C10303 VN.n9313 a_400_62400# 0.16fF
C10304 VN.t204 a_400_62400# 0.03fF
C10305 VN.n9314 a_400_62400# 0.19fF
C10306 VN.n9316 a_400_62400# 0.93fF
C10307 VN.n9317 a_400_62400# 0.30fF
C10308 VN.n9318 a_400_62400# 0.34fF
C10309 VN.n9319 a_400_62400# 0.12fF
C10310 VN.n9320 a_400_62400# 0.30fF
C10311 VN.n9321 a_400_62400# 0.93fF
C10312 VN.n9322 a_400_62400# 1.55fF
C10313 VN.n9323 a_400_62400# 0.29fF
C10314 VN.n9324 a_400_62400# 0.34fF
C10315 VN.n9325 a_400_62400# 0.12fF
C10316 VN.n9326 a_400_62400# 3.10fF
C10317 VN.t2468 a_400_62400# 0.03fF
C10318 VN.n9327 a_400_62400# 0.32fF
C10319 VN.n9328 a_400_62400# 1.22fF
C10320 VN.n9329 a_400_62400# 0.07fF
C10321 VN.t1002 a_400_62400# 0.03fF
C10322 VN.n9330 a_400_62400# 0.16fF
C10323 VN.n9331 a_400_62400# 0.19fF
C10324 VN.n9333 a_400_62400# 2.51fF
C10325 VN.n9334 a_400_62400# 0.61fF
C10326 VN.n9335 a_400_62400# 0.30fF
C10327 VN.n9336 a_400_62400# 0.51fF
C10328 VN.n9337 a_400_62400# 0.21fF
C10329 VN.n9338 a_400_62400# 0.38fF
C10330 VN.n9339 a_400_62400# 0.29fF
C10331 VN.n9340 a_400_62400# 0.40fF
C10332 VN.n9341 a_400_62400# 0.28fF
C10333 VN.t497 a_400_62400# 0.03fF
C10334 VN.n9342 a_400_62400# 0.32fF
C10335 VN.n9343 a_400_62400# 0.48fF
C10336 VN.n9344 a_400_62400# 0.81fF
C10337 VN.n9345 a_400_62400# 0.16fF
C10338 VN.t1992 a_400_62400# 0.03fF
C10339 VN.n9346 a_400_62400# 0.19fF
C10340 VN.n9348 a_400_62400# 0.06fF
C10341 VN.n9349 a_400_62400# 0.04fF
C10342 VN.n9350 a_400_62400# 0.04fF
C10343 VN.n9351 a_400_62400# 0.14fF
C10344 VN.n9352 a_400_62400# 0.48fF
C10345 VN.n9353 a_400_62400# 0.50fF
C10346 VN.n9354 a_400_62400# 0.14fF
C10347 VN.n9355 a_400_62400# 0.16fF
C10348 VN.n9356 a_400_62400# 0.09fF
C10349 VN.n9357 a_400_62400# 0.16fF
C10350 VN.n9358 a_400_62400# 0.24fF
C10351 VN.n9359 a_400_62400# 5.35fF
C10352 VN.t1602 a_400_62400# 0.03fF
C10353 VN.n9360 a_400_62400# 0.32fF
C10354 VN.n9361 a_400_62400# 1.22fF
C10355 VN.n9362 a_400_62400# 0.07fF
C10356 VN.t126 a_400_62400# 0.03fF
C10357 VN.n9363 a_400_62400# 0.16fF
C10358 VN.n9364 a_400_62400# 0.19fF
C10359 VN.n9366 a_400_62400# 0.33fF
C10360 VN.n9367 a_400_62400# 0.12fF
C10361 VN.n9368 a_400_62400# 0.28fF
C10362 VN.n9369 a_400_62400# 1.72fF
C10363 VN.n9370 a_400_62400# 0.71fF
C10364 VN.n9371 a_400_62400# 2.51fF
C10365 VN.n9372 a_400_62400# 0.16fF
C10366 VN.t1118 a_400_62400# 0.03fF
C10367 VN.n9373 a_400_62400# 0.19fF
C10368 VN.t2268 a_400_62400# 0.03fF
C10369 VN.n9375 a_400_62400# 0.32fF
C10370 VN.n9376 a_400_62400# 0.48fF
C10371 VN.n9377 a_400_62400# 0.81fF
C10372 VN.n9378 a_400_62400# 0.95fF
C10373 VN.n9379 a_400_62400# 2.11fF
C10374 VN.n9380 a_400_62400# 3.28fF
C10375 VN.t848 a_400_62400# 0.03fF
C10376 VN.n9381 a_400_62400# 0.32fF
C10377 VN.n9382 a_400_62400# 1.22fF
C10378 VN.n9383 a_400_62400# 0.07fF
C10379 VN.t1790 a_400_62400# 0.03fF
C10380 VN.n9384 a_400_62400# 0.16fF
C10381 VN.n9385 a_400_62400# 0.19fF
C10382 VN.n9387 a_400_62400# 2.53fF
C10383 VN.n9388 a_400_62400# 0.08fF
C10384 VN.n9389 a_400_62400# 0.04fF
C10385 VN.n9390 a_400_62400# 0.05fF
C10386 VN.n9391 a_400_62400# 1.33fF
C10387 VN.n9392 a_400_62400# 0.03fF
C10388 VN.n9393 a_400_62400# 0.01fF
C10389 VN.n9394 a_400_62400# 0.02fF
C10390 VN.n9395 a_400_62400# 0.11fF
C10391 VN.n9396 a_400_62400# 0.48fF
C10392 VN.n9397 a_400_62400# 2.48fF
C10393 VN.t718 a_400_62400# 0.03fF
C10394 VN.n9398 a_400_62400# 0.32fF
C10395 VN.n9399 a_400_62400# 0.48fF
C10396 VN.n9400 a_400_62400# 0.81fF
C10397 VN.n9401 a_400_62400# 0.16fF
C10398 VN.t2103 a_400_62400# 0.03fF
C10399 VN.n9402 a_400_62400# 0.19fF
C10400 VN.n9404 a_400_62400# 0.93fF
C10401 VN.n9405 a_400_62400# 0.30fF
C10402 VN.n9406 a_400_62400# 0.34fF
C10403 VN.n9407 a_400_62400# 0.12fF
C10404 VN.n9408 a_400_62400# 0.30fF
C10405 VN.n9409 a_400_62400# 0.93fF
C10406 VN.n9410 a_400_62400# 1.55fF
C10407 VN.n9411 a_400_62400# 0.29fF
C10408 VN.n9412 a_400_62400# 0.34fF
C10409 VN.n9413 a_400_62400# 0.12fF
C10410 VN.n9414 a_400_62400# 2.52fF
C10411 VN.t2293 a_400_62400# 0.03fF
C10412 VN.n9415 a_400_62400# 0.32fF
C10413 VN.n9416 a_400_62400# 1.22fF
C10414 VN.n9417 a_400_62400# 0.07fF
C10415 VN.t915 a_400_62400# 0.03fF
C10416 VN.n9418 a_400_62400# 0.16fF
C10417 VN.n9419 a_400_62400# 0.19fF
C10418 VN.n9421 a_400_62400# 27.83fF
C10419 VN.n9422 a_400_62400# 2.30fF
C10420 VN.n9423 a_400_62400# 4.08fF
C10421 VN.t982 a_400_62400# 0.03fF
C10422 VN.n9424 a_400_62400# 0.32fF
C10423 VN.n9425 a_400_62400# 0.48fF
C10424 VN.n9426 a_400_62400# 0.81fF
C10425 VN.n9427 a_400_62400# 0.16fF
C10426 VN.t2380 a_400_62400# 0.03fF
C10427 VN.n9428 a_400_62400# 0.19fF
C10428 VN.n9430 a_400_62400# 0.42fF
C10429 VN.n9431 a_400_62400# 0.34fF
C10430 VN.n9432 a_400_62400# 0.12fF
C10431 VN.n9433 a_400_62400# 0.30fF
C10432 VN.n9434 a_400_62400# 0.88fF
C10433 VN.n9435 a_400_62400# 1.28fF
C10434 VN.n9436 a_400_62400# 0.30fF
C10435 VN.n9437 a_400_62400# 0.28fF
C10436 VN.n9438 a_400_62400# 0.27fF
C10437 VN.n9439 a_400_62400# 0.09fF
C10438 VN.n9440 a_400_62400# 0.12fF
C10439 VN.n9441 a_400_62400# 0.13fF
C10440 VN.n9442 a_400_62400# 2.66fF
C10441 VN.t655 a_400_62400# 0.03fF
C10442 VN.n9443 a_400_62400# 0.16fF
C10443 VN.n9444 a_400_62400# 0.19fF
C10444 VN.t2128 a_400_62400# 0.03fF
C10445 VN.n9446 a_400_62400# 0.32fF
C10446 VN.n9447 a_400_62400# 1.22fF
C10447 VN.n9448 a_400_62400# 0.07fF
C10448 VN.n9449 a_400_62400# 2.51fF
C10449 VN.n9450 a_400_62400# 0.16fF
C10450 VN.t1226 a_400_62400# 0.03fF
C10451 VN.n9451 a_400_62400# 0.19fF
C10452 VN.t2372 a_400_62400# 0.03fF
C10453 VN.n9453 a_400_62400# 0.32fF
C10454 VN.n9454 a_400_62400# 0.48fF
C10455 VN.n9455 a_400_62400# 0.81fF
C10456 VN.n9456 a_400_62400# 1.24fF
C10457 VN.n9457 a_400_62400# 0.43fF
C10458 VN.n9458 a_400_62400# 0.43fF
C10459 VN.n9459 a_400_62400# 1.24fF
C10460 VN.n9460 a_400_62400# 1.46fF
C10461 VN.n9461 a_400_62400# 0.21fF
C10462 VN.n9462 a_400_62400# 6.64fF
C10463 VN.t1887 a_400_62400# 0.03fF
C10464 VN.n9463 a_400_62400# 0.16fF
C10465 VN.n9464 a_400_62400# 0.19fF
C10466 VN.t1425 a_400_62400# 0.03fF
C10467 VN.n9466 a_400_62400# 0.32fF
C10468 VN.n9467 a_400_62400# 1.22fF
C10469 VN.n9468 a_400_62400# 0.07fF
C10470 VN.n9469 a_400_62400# 2.51fF
C10471 VN.n9470 a_400_62400# 3.57fF
C10472 VN.t1504 a_400_62400# 0.03fF
C10473 VN.n9471 a_400_62400# 0.32fF
C10474 VN.n9472 a_400_62400# 0.48fF
C10475 VN.n9473 a_400_62400# 0.81fF
C10476 VN.n9474 a_400_62400# 0.16fF
C10477 VN.t360 a_400_62400# 0.03fF
C10478 VN.n9475 a_400_62400# 0.19fF
C10479 VN.n9477 a_400_62400# 2.51fF
C10480 VN.n9478 a_400_62400# 3.59fF
C10481 VN.t365 a_400_62400# 0.03fF
C10482 VN.n9479 a_400_62400# 0.32fF
C10483 VN.n9480 a_400_62400# 0.48fF
C10484 VN.n9481 a_400_62400# 0.81fF
C10485 VN.t400 a_400_62400# 0.03fF
C10486 VN.n9482 a_400_62400# 1.63fF
C10487 VN.n9483 a_400_62400# 0.49fF
C10488 VN.n9484 a_400_62400# 1.64fF
C10489 VN.n9485 a_400_62400# 0.81fF
C10490 VN.n9486 a_400_62400# 1.21fF
C10491 VN.n9487 a_400_62400# 1.54fF
C10492 VN.n9488 a_400_62400# 4.06fF
C10493 VN.t66 a_400_62400# 28.64fF
C10494 VN.n9489 a_400_62400# 28.43fF
C10495 VN.n9491 a_400_62400# 0.50fF
C10496 VN.n9492 a_400_62400# 0.31fF
C10497 VN.n9493 a_400_62400# 3.74fF
C10498 VN.n9494 a_400_62400# 3.29fF
C10499 VN.n9495 a_400_62400# 5.35fF
C10500 VN.n9496 a_400_62400# 0.34fF
C10501 VN.n9497 a_400_62400# 0.02fF
C10502 VN.t1761 a_400_62400# 0.03fF
C10503 VN.n9498 a_400_62400# 0.34fF
C10504 VN.t2089 a_400_62400# 0.03fF
C10505 VN.n9499 a_400_62400# 1.28fF
C10506 VN.n9500 a_400_62400# 0.94fF
C10507 VN.n9501 a_400_62400# 2.53fF
C10508 VN.n9502 a_400_62400# 2.51fF
C10509 VN.t2048 a_400_62400# 0.03fF
C10510 VN.n9503 a_400_62400# 0.32fF
C10511 VN.n9504 a_400_62400# 0.48fF
C10512 VN.n9505 a_400_62400# 0.81fF
C10513 VN.n9506 a_400_62400# 0.16fF
C10514 VN.t890 a_400_62400# 0.03fF
C10515 VN.n9507 a_400_62400# 0.19fF
C10516 VN.n9509 a_400_62400# 1.55fF
C10517 VN.n9510 a_400_62400# 0.29fF
C10518 VN.n9511 a_400_62400# 2.52fF
C10519 VN.t1212 a_400_62400# 0.03fF
C10520 VN.n9512 a_400_62400# 0.32fF
C10521 VN.n9513 a_400_62400# 1.22fF
C10522 VN.n9514 a_400_62400# 0.07fF
C10523 VN.t962 a_400_62400# 0.03fF
C10524 VN.n9515 a_400_62400# 0.16fF
C10525 VN.n9516 a_400_62400# 0.19fF
C10526 VN.n9518 a_400_62400# 1.04fF
C10527 VN.n9519 a_400_62400# 2.60fF
C10528 VN.n9520 a_400_62400# 2.51fF
C10529 VN.n9521 a_400_62400# 0.16fF
C10530 VN.t2551 a_400_62400# 0.03fF
C10531 VN.n9522 a_400_62400# 0.19fF
C10532 VN.t1180 a_400_62400# 0.03fF
C10533 VN.n9524 a_400_62400# 0.32fF
C10534 VN.n9525 a_400_62400# 0.48fF
C10535 VN.n9526 a_400_62400# 0.81fF
C10536 VN.n9527 a_400_62400# 2.46fF
C10537 VN.n9528 a_400_62400# 4.01fF
C10538 VN.t351 a_400_62400# 0.03fF
C10539 VN.n9529 a_400_62400# 0.32fF
C10540 VN.n9530 a_400_62400# 1.22fF
C10541 VN.n9531 a_400_62400# 0.07fF
C10542 VN.t227 a_400_62400# 0.03fF
C10543 VN.n9532 a_400_62400# 0.16fF
C10544 VN.n9533 a_400_62400# 0.19fF
C10545 VN.n9535 a_400_62400# 2.53fF
C10546 VN.n9536 a_400_62400# 2.51fF
C10547 VN.t310 a_400_62400# 0.03fF
C10548 VN.n9537 a_400_62400# 0.32fF
C10549 VN.n9538 a_400_62400# 0.48fF
C10550 VN.n9539 a_400_62400# 0.81fF
C10551 VN.n9540 a_400_62400# 0.16fF
C10552 VN.t1681 a_400_62400# 0.03fF
C10553 VN.n9541 a_400_62400# 0.19fF
C10554 VN.n9543 a_400_62400# 1.55fF
C10555 VN.n9544 a_400_62400# 0.29fF
C10556 VN.n9545 a_400_62400# 2.52fF
C10557 VN.t1994 a_400_62400# 0.03fF
C10558 VN.n9546 a_400_62400# 0.32fF
C10559 VN.n9547 a_400_62400# 1.22fF
C10560 VN.n9548 a_400_62400# 0.07fF
C10561 VN.t1875 a_400_62400# 0.03fF
C10562 VN.n9549 a_400_62400# 0.16fF
C10563 VN.n9550 a_400_62400# 0.19fF
C10564 VN.n9552 a_400_62400# 1.05fF
C10565 VN.n9553 a_400_62400# 3.07fF
C10566 VN.n9554 a_400_62400# 2.51fF
C10567 VN.n9555 a_400_62400# 0.16fF
C10568 VN.t815 a_400_62400# 0.03fF
C10569 VN.n9556 a_400_62400# 0.19fF
C10570 VN.t1959 a_400_62400# 0.03fF
C10571 VN.n9558 a_400_62400# 0.32fF
C10572 VN.n9559 a_400_62400# 0.48fF
C10573 VN.n9560 a_400_62400# 0.81fF
C10574 VN.n9561 a_400_62400# 2.46fF
C10575 VN.n9562 a_400_62400# 2.91fF
C10576 VN.t1121 a_400_62400# 0.03fF
C10577 VN.n9563 a_400_62400# 0.32fF
C10578 VN.n9564 a_400_62400# 1.22fF
C10579 VN.n9565 a_400_62400# 0.07fF
C10580 VN.t1006 a_400_62400# 0.03fF
C10581 VN.n9566 a_400_62400# 0.16fF
C10582 VN.n9567 a_400_62400# 0.19fF
C10583 VN.n9569 a_400_62400# 2.53fF
C10584 VN.n9570 a_400_62400# 2.51fF
C10585 VN.t2436 a_400_62400# 0.03fF
C10586 VN.n9571 a_400_62400# 0.32fF
C10587 VN.n9572 a_400_62400# 0.48fF
C10588 VN.n9573 a_400_62400# 0.81fF
C10589 VN.n9574 a_400_62400# 0.16fF
C10590 VN.t1315 a_400_62400# 0.03fF
C10591 VN.n9575 a_400_62400# 0.19fF
C10592 VN.n9577 a_400_62400# 1.55fF
C10593 VN.n9578 a_400_62400# 0.29fF
C10594 VN.n9579 a_400_62400# 2.52fF
C10595 VN.t1609 a_400_62400# 0.03fF
C10596 VN.n9580 a_400_62400# 0.32fF
C10597 VN.n9581 a_400_62400# 1.22fF
C10598 VN.n9582 a_400_62400# 0.07fF
C10599 VN.t1497 a_400_62400# 0.03fF
C10600 VN.n9583 a_400_62400# 0.16fF
C10601 VN.n9584 a_400_62400# 0.19fF
C10602 VN.n9586 a_400_62400# 1.04fF
C10603 VN.n9587 a_400_62400# 2.60fF
C10604 VN.n9588 a_400_62400# 2.51fF
C10605 VN.n9589 a_400_62400# 0.16fF
C10606 VN.t455 a_400_62400# 0.03fF
C10607 VN.n9590 a_400_62400# 0.19fF
C10608 VN.t1575 a_400_62400# 0.03fF
C10609 VN.n9592 a_400_62400# 0.32fF
C10610 VN.n9593 a_400_62400# 0.48fF
C10611 VN.n9594 a_400_62400# 0.81fF
C10612 VN.n9595 a_400_62400# 2.46fF
C10613 VN.n9596 a_400_62400# 4.01fF
C10614 VN.t743 a_400_62400# 0.03fF
C10615 VN.n9597 a_400_62400# 0.32fF
C10616 VN.n9598 a_400_62400# 1.22fF
C10617 VN.n9599 a_400_62400# 0.07fF
C10618 VN.t631 a_400_62400# 0.03fF
C10619 VN.n9600 a_400_62400# 0.16fF
C10620 VN.n9601 a_400_62400# 0.19fF
C10621 VN.n9603 a_400_62400# 2.53fF
C10622 VN.n9604 a_400_62400# 2.51fF
C10623 VN.t706 a_400_62400# 0.03fF
C10624 VN.n9605 a_400_62400# 0.32fF
C10625 VN.n9606 a_400_62400# 0.48fF
C10626 VN.n9607 a_400_62400# 0.81fF
C10627 VN.n9608 a_400_62400# 0.16fF
C10628 VN.t2223 a_400_62400# 0.03fF
C10629 VN.n9609 a_400_62400# 0.19fF
C10630 VN.n9611 a_400_62400# 1.55fF
C10631 VN.n9612 a_400_62400# 0.29fF
C10632 VN.n9613 a_400_62400# 2.52fF
C10633 VN.t2399 a_400_62400# 0.03fF
C10634 VN.n9614 a_400_62400# 0.32fF
C10635 VN.n9615 a_400_62400# 1.22fF
C10636 VN.n9616 a_400_62400# 0.07fF
C10637 VN.t2288 a_400_62400# 0.03fF
C10638 VN.n9617 a_400_62400# 0.16fF
C10639 VN.n9618 a_400_62400# 0.19fF
C10640 VN.n9620 a_400_62400# 1.04fF
C10641 VN.n9621 a_400_62400# 2.60fF
C10642 VN.n9622 a_400_62400# 2.51fF
C10643 VN.n9623 a_400_62400# 0.16fF
C10644 VN.t1358 a_400_62400# 0.03fF
C10645 VN.n9624 a_400_62400# 0.19fF
C10646 VN.t2479 a_400_62400# 0.03fF
C10647 VN.n9626 a_400_62400# 0.32fF
C10648 VN.n9627 a_400_62400# 0.48fF
C10649 VN.n9628 a_400_62400# 0.81fF
C10650 VN.n9629 a_400_62400# 2.46fF
C10651 VN.n9630 a_400_62400# 4.01fF
C10652 VN.t1653 a_400_62400# 0.03fF
C10653 VN.n9631 a_400_62400# 0.32fF
C10654 VN.n9632 a_400_62400# 1.22fF
C10655 VN.n9633 a_400_62400# 0.07fF
C10656 VN.t1421 a_400_62400# 0.03fF
C10657 VN.n9634 a_400_62400# 0.16fF
C10658 VN.n9635 a_400_62400# 0.19fF
C10659 VN.n9637 a_400_62400# 2.53fF
C10660 VN.n9638 a_400_62400# 2.51fF
C10661 VN.t1617 a_400_62400# 0.03fF
C10662 VN.n9639 a_400_62400# 0.32fF
C10663 VN.n9640 a_400_62400# 0.48fF
C10664 VN.n9641 a_400_62400# 0.81fF
C10665 VN.n9642 a_400_62400# 0.16fF
C10666 VN.t491 a_400_62400# 0.03fF
C10667 VN.n9643 a_400_62400# 0.19fF
C10668 VN.n9645 a_400_62400# 1.55fF
C10669 VN.n9646 a_400_62400# 0.29fF
C10670 VN.n9647 a_400_62400# 2.52fF
C10671 VN.t782 a_400_62400# 0.03fF
C10672 VN.n9648 a_400_62400# 0.32fF
C10673 VN.n9649 a_400_62400# 1.22fF
C10674 VN.n9650 a_400_62400# 0.07fF
C10675 VN.t556 a_400_62400# 0.03fF
C10676 VN.n9651 a_400_62400# 0.16fF
C10677 VN.n9652 a_400_62400# 0.19fF
C10678 VN.n9654 a_400_62400# 1.04fF
C10679 VN.n9655 a_400_62400# 2.60fF
C10680 VN.n9656 a_400_62400# 2.51fF
C10681 VN.n9657 a_400_62400# 0.16fF
C10682 VN.t2146 a_400_62400# 0.03fF
C10683 VN.n9658 a_400_62400# 0.19fF
C10684 VN.t748 a_400_62400# 0.03fF
C10685 VN.n9660 a_400_62400# 0.32fF
C10686 VN.n9661 a_400_62400# 0.48fF
C10687 VN.n9662 a_400_62400# 0.81fF
C10688 VN.n9663 a_400_62400# 2.46fF
C10689 VN.n9664 a_400_62400# 4.01fF
C10690 VN.t2433 a_400_62400# 0.03fF
C10691 VN.n9665 a_400_62400# 0.32fF
C10692 VN.n9666 a_400_62400# 1.22fF
C10693 VN.n9667 a_400_62400# 0.07fF
C10694 VN.t2214 a_400_62400# 0.03fF
C10695 VN.n9668 a_400_62400# 0.16fF
C10696 VN.n9669 a_400_62400# 0.19fF
C10697 VN.n9671 a_400_62400# 2.53fF
C10698 VN.n9672 a_400_62400# 2.34fF
C10699 VN.t2407 a_400_62400# 0.03fF
C10700 VN.n9673 a_400_62400# 0.32fF
C10701 VN.n9674 a_400_62400# 0.48fF
C10702 VN.n9675 a_400_62400# 0.81fF
C10703 VN.n9676 a_400_62400# 0.16fF
C10704 VN.t1276 a_400_62400# 0.03fF
C10705 VN.n9677 a_400_62400# 0.19fF
C10706 VN.n9679 a_400_62400# 1.55fF
C10707 VN.n9680 a_400_62400# 0.29fF
C10708 VN.n9681 a_400_62400# 3.27fF
C10709 VN.t1573 a_400_62400# 0.03fF
C10710 VN.n9682 a_400_62400# 0.32fF
C10711 VN.n9683 a_400_62400# 1.22fF
C10712 VN.n9684 a_400_62400# 0.07fF
C10713 VN.t1346 a_400_62400# 0.03fF
C10714 VN.n9685 a_400_62400# 0.16fF
C10715 VN.n9686 a_400_62400# 0.19fF
C10716 VN.n9688 a_400_62400# 2.51fF
C10717 VN.n9689 a_400_62400# 0.56fF
C10718 VN.n9690 a_400_62400# 0.64fF
C10719 VN.n9691 a_400_62400# 0.12fF
C10720 VN.n9692 a_400_62400# 0.44fF
C10721 VN.n9693 a_400_62400# 0.40fF
C10722 VN.n9694 a_400_62400# 1.03fF
C10723 VN.n9695 a_400_62400# 0.79fF
C10724 VN.t1540 a_400_62400# 0.03fF
C10725 VN.n9696 a_400_62400# 0.32fF
C10726 VN.n9697 a_400_62400# 0.48fF
C10727 VN.n9698 a_400_62400# 0.81fF
C10728 VN.n9699 a_400_62400# 0.16fF
C10729 VN.t407 a_400_62400# 0.03fF
C10730 VN.n9700 a_400_62400# 0.19fF
C10731 VN.n9702 a_400_62400# 3.50fF
C10732 VN.n9703 a_400_62400# 2.89fF
C10733 VN.t703 a_400_62400# 0.03fF
C10734 VN.n9704 a_400_62400# 0.32fF
C10735 VN.n9705 a_400_62400# 1.22fF
C10736 VN.n9706 a_400_62400# 0.07fF
C10737 VN.t596 a_400_62400# 0.03fF
C10738 VN.n9707 a_400_62400# 0.16fF
C10739 VN.n9708 a_400_62400# 0.19fF
C10740 VN.n9710 a_400_62400# 1.05fF
C10741 VN.n9711 a_400_62400# 3.07fF
C10742 VN.n9712 a_400_62400# 2.51fF
C10743 VN.n9713 a_400_62400# 0.16fF
C10744 VN.t2057 a_400_62400# 0.03fF
C10745 VN.n9714 a_400_62400# 0.19fF
C10746 VN.t671 a_400_62400# 0.03fF
C10747 VN.n9716 a_400_62400# 0.32fF
C10748 VN.n9717 a_400_62400# 0.48fF
C10749 VN.n9718 a_400_62400# 0.81fF
C10750 VN.n9719 a_400_62400# 1.86fF
C10751 VN.n9720 a_400_62400# 1.53fF
C10752 VN.n9721 a_400_62400# 0.47fF
C10753 VN.n9722 a_400_62400# 2.71fF
C10754 VN.t2362 a_400_62400# 0.03fF
C10755 VN.n9723 a_400_62400# 0.32fF
C10756 VN.n9724 a_400_62400# 1.22fF
C10757 VN.n9725 a_400_62400# 0.07fF
C10758 VN.t2251 a_400_62400# 0.03fF
C10759 VN.n9726 a_400_62400# 0.16fF
C10760 VN.n9727 a_400_62400# 0.19fF
C10761 VN.n9729 a_400_62400# 2.53fF
C10762 VN.n9730 a_400_62400# 2.51fF
C10763 VN.t2107 a_400_62400# 0.03fF
C10764 VN.n9731 a_400_62400# 0.32fF
C10765 VN.n9732 a_400_62400# 0.48fF
C10766 VN.n9733 a_400_62400# 0.81fF
C10767 VN.n9734 a_400_62400# 0.16fF
C10768 VN.t928 a_400_62400# 0.03fF
C10769 VN.n9735 a_400_62400# 0.19fF
C10770 VN.n9737 a_400_62400# 1.55fF
C10771 VN.n9738 a_400_62400# 0.29fF
C10772 VN.n9739 a_400_62400# 2.52fF
C10773 VN.t1376 a_400_62400# 0.03fF
C10774 VN.n9740 a_400_62400# 0.32fF
C10775 VN.n9741 a_400_62400# 1.22fF
C10776 VN.n9742 a_400_62400# 0.07fF
C10777 VN.t1136 a_400_62400# 0.03fF
C10778 VN.n9743 a_400_62400# 0.16fF
C10779 VN.n9744 a_400_62400# 0.19fF
C10780 VN.n9746 a_400_62400# 27.83fF
C10781 VN.n9747 a_400_62400# 3.93fF
C10782 VN.n9748 a_400_62400# 2.51fF
C10783 VN.n9749 a_400_62400# 0.16fF
C10784 VN.t1 a_400_62400# 0.03fF
C10785 VN.n9750 a_400_62400# 0.19fF
C10786 VN.t1230 a_400_62400# 0.03fF
C10787 VN.n9752 a_400_62400# 0.32fF
C10788 VN.n9753 a_400_62400# 0.48fF
C10789 VN.n9754 a_400_62400# 0.81fF
C10790 VN.n9755 a_400_62400# 1.46fF
C10791 VN.n9756 a_400_62400# 0.21fF
C10792 VN.n9757 a_400_62400# 2.81fF
C10793 VN.t273 a_400_62400# 0.03fF
C10794 VN.n9758 a_400_62400# 0.16fF
C10795 VN.n9759 a_400_62400# 0.19fF
C10796 VN.t511 a_400_62400# 0.03fF
C10797 VN.n9761 a_400_62400# 0.32fF
C10798 VN.n9762 a_400_62400# 1.22fF
C10799 VN.n9763 a_400_62400# 0.07fF
C10800 VN.n9764 a_400_62400# 3.65fF
C10801 VN.n9765 a_400_62400# 2.14fF
C10802 VN.n9766 a_400_62400# 0.16fF
C10803 VN.t974 a_400_62400# 0.03fF
C10804 VN.n9767 a_400_62400# 0.19fF
C10805 VN.t2015 a_400_62400# 0.03fF
C10806 VN.n9769 a_400_62400# 0.32fF
C10807 VN.n9770 a_400_62400# 0.48fF
C10808 VN.n9771 a_400_62400# 0.81fF
C10809 VN.n9772 a_400_62400# 0.09fF
C10810 VN.n9773 a_400_62400# 0.01fF
C10811 VN.n9774 a_400_62400# 0.02fF
C10812 VN.n9775 a_400_62400# 0.02fF
C10813 VN.n9776 a_400_62400# 0.32fF
C10814 VN.n9777 a_400_62400# 1.56fF
C10815 VN.n9778 a_400_62400# 1.81fF
C10816 VN.n9779 a_400_62400# 3.08fF
C10817 VN.t1048 a_400_62400# 0.03fF
C10818 VN.n9780 a_400_62400# 0.16fF
C10819 VN.n9781 a_400_62400# 0.19fF
C10820 VN.t1296 a_400_62400# 0.03fF
C10821 VN.n9783 a_400_62400# 0.32fF
C10822 VN.n9784 a_400_62400# 1.22fF
C10823 VN.n9785 a_400_62400# 0.07fF
C10824 VN.t0 a_400_62400# 64.69fF
C10825 VN.t2163 a_400_62400# 0.03fF
C10826 VN.n9786 a_400_62400# 0.32fF
C10827 VN.n9787 a_400_62400# 1.22fF
C10828 VN.n9788 a_400_62400# 0.07fF
C10829 VN.t1923 a_400_62400# 0.03fF
C10830 VN.n9789 a_400_62400# 0.16fF
C10831 VN.n9790 a_400_62400# 0.19fF
C10832 VN.n9792 a_400_62400# 0.16fF
C10833 VN.t1722 a_400_62400# 0.03fF
C10834 VN.n9793 a_400_62400# 0.19fF
C10835 VN.n9795 a_400_62400# 6.93fF
C10836 VN.n9796 a_400_62400# 6.54fF
C10837 VN.t1015 a_400_62400# 0.03fF
C10838 VN.n9797 a_400_62400# 0.16fF
C10839 VN.n9798 a_400_62400# 0.19fF
C10840 VN.t559 a_400_62400# 0.03fF
C10841 VN.n9800 a_400_62400# 0.32fF
C10842 VN.n9801 a_400_62400# 1.22fF
C10843 VN.n9802 a_400_62400# 0.07fF
C10844 VN.n9803 a_400_62400# 2.51fF
C10845 VN.n9804 a_400_62400# 3.58fF
C10846 VN.t638 a_400_62400# 0.03fF
C10847 VN.n9805 a_400_62400# 0.32fF
C10848 VN.n9806 a_400_62400# 0.48fF
C10849 VN.n9807 a_400_62400# 0.81fF
C10850 VN.n9808 a_400_62400# 0.16fF
C10851 VN.t2009 a_400_62400# 0.03fF
C10852 VN.n9809 a_400_62400# 0.19fF
C10853 VN.n9811 a_400_62400# 7.29fF
C10854 VN.t141 a_400_62400# 0.03fF
C10855 VN.n9812 a_400_62400# 0.16fF
C10856 VN.n9813 a_400_62400# 0.19fF
C10857 VN.t2218 a_400_62400# 0.03fF
C10858 VN.n9815 a_400_62400# 0.32fF
C10859 VN.n9816 a_400_62400# 1.22fF
C10860 VN.n9817 a_400_62400# 0.07fF
C10861 VN.t125 a_400_62400# 64.17fF
C10862 VN.t1351 a_400_62400# 0.03fF
C10863 VN.n9818 a_400_62400# 1.60fF
C10864 VN.n9819 a_400_62400# 0.07fF
C10865 VN.t1936 a_400_62400# 0.03fF
C10866 VN.n9820 a_400_62400# 0.02fF
C10867 VN.n9821 a_400_62400# 0.34fF
C10868 VN.n9823 a_400_62400# 2.01fF
C10869 VN.n9824 a_400_62400# 1.75fF
C10870 VN.n9825 a_400_62400# 0.37fF
C10871 VN.n9826 a_400_62400# 0.33fF
C10872 VN.n9827 a_400_62400# 5.88fF
C10873 VN.n9828 a_400_62400# 0.02fF
C10874 VN.n9829 a_400_62400# 0.02fF
C10875 VN.n9830 a_400_62400# 0.03fF
C10876 VN.n9831 a_400_62400# 0.05fF
C10877 VN.n9832 a_400_62400# 0.23fF
C10878 VN.n9833 a_400_62400# 0.02fF
C10879 VN.n9834 a_400_62400# 0.03fF
C10880 VN.n9835 a_400_62400# 0.01fF
C10881 VN.n9836 a_400_62400# 0.01fF
C10882 VN.n9837 a_400_62400# 0.01fF
C10883 VN.n9838 a_400_62400# 0.02fF
C10884 VN.n9839 a_400_62400# 0.03fF
C10885 VN.n9840 a_400_62400# 0.06fF
C10886 VN.n9841 a_400_62400# 0.05fF
C10887 VN.n9842 a_400_62400# 0.15fF
C10888 VN.n9843 a_400_62400# 0.51fF
C10889 VN.n9844 a_400_62400# 0.27fF
C10890 VN.n9845 a_400_62400# 37.46fF
C10891 VN.n9846 a_400_62400# 37.46fF
C10892 VN.n9847 a_400_62400# 37.46fF
C10893 VN.n9848 a_400_62400# 37.46fF
C10894 VN.n9849 a_400_62400# 0.79fF
C10895 VN.n9850 a_400_62400# 0.23fF
C10896 VN.n9851 a_400_62400# 1.18fF
C10897 VN.t350 a_400_62400# 28.64fF
C10898 VN.n9852 a_400_62400# 0.79fF
C10899 VN.n9853 a_400_62400# 0.11fF
C10900 VN.n9854 a_400_62400# 4.98fF
C10901 VN.n9855 a_400_62400# 0.80fF
C10902 VN.n9856 a_400_62400# 0.29fF
C10903 VN.n9857 a_400_62400# 1.96fF
C10904 VN.n9859 a_400_62400# 25.18fF
C10905 VN.n9861 a_400_62400# 1.87fF
C10906 VN.n9862 a_400_62400# 5.36fF
C10907 VN.n9863 a_400_62400# 1.81fF
C10908 VN.t610 a_400_62400# 0.03fF
C10909 VN.n9864 a_400_62400# 0.85fF
C10910 VN.n9865 a_400_62400# 0.81fF
C10911 VN.n9866 a_400_62400# 2.53fF
C10912 VN.n9867 a_400_62400# 0.08fF
C10913 VN.n9868 a_400_62400# 0.04fF
C10914 VN.n9869 a_400_62400# 0.05fF
C10915 VN.n9870 a_400_62400# 1.33fF
C10916 VN.n9871 a_400_62400# 0.03fF
C10917 VN.n9872 a_400_62400# 0.01fF
C10918 VN.n9873 a_400_62400# 0.02fF
C10919 VN.n9874 a_400_62400# 0.11fF
C10920 VN.n9875 a_400_62400# 0.48fF
C10921 VN.n9876 a_400_62400# 2.48fF
C10922 VN.t426 a_400_62400# 0.03fF
C10923 VN.n9877 a_400_62400# 0.32fF
C10924 VN.n9878 a_400_62400# 0.48fF
C10925 VN.n9879 a_400_62400# 0.81fF
C10926 VN.n9880 a_400_62400# 0.16fF
C10927 VN.t1918 a_400_62400# 0.03fF
C10928 VN.n9881 a_400_62400# 0.19fF
C10929 VN.n9883 a_400_62400# 0.93fF
C10930 VN.n9884 a_400_62400# 0.30fF
C10931 VN.n9885 a_400_62400# 0.34fF
C10932 VN.n9886 a_400_62400# 0.12fF
C10933 VN.n9887 a_400_62400# 0.30fF
C10934 VN.n9888 a_400_62400# 0.93fF
C10935 VN.n9889 a_400_62400# 1.55fF
C10936 VN.n9890 a_400_62400# 0.29fF
C10937 VN.n9891 a_400_62400# 0.34fF
C10938 VN.n9892 a_400_62400# 0.12fF
C10939 VN.n9893 a_400_62400# 2.52fF
C10940 VN.t1534 a_400_62400# 0.03fF
C10941 VN.n9894 a_400_62400# 0.32fF
C10942 VN.n9895 a_400_62400# 1.22fF
C10943 VN.n9896 a_400_62400# 0.07fF
C10944 VN.t2588 a_400_62400# 0.03fF
C10945 VN.n9897 a_400_62400# 0.16fF
C10946 VN.n9898 a_400_62400# 0.19fF
C10947 VN.n9900 a_400_62400# 0.33fF
C10948 VN.n9901 a_400_62400# 0.12fF
C10949 VN.n9902 a_400_62400# 0.28fF
C10950 VN.n9903 a_400_62400# 1.23fF
C10951 VN.n9904 a_400_62400# 0.59fF
C10952 VN.n9905 a_400_62400# 2.51fF
C10953 VN.n9906 a_400_62400# 0.16fF
C10954 VN.t1042 a_400_62400# 0.03fF
C10955 VN.n9907 a_400_62400# 0.19fF
C10956 VN.t2201 a_400_62400# 0.03fF
C10957 VN.n9909 a_400_62400# 0.32fF
C10958 VN.n9910 a_400_62400# 0.48fF
C10959 VN.n9911 a_400_62400# 0.81fF
C10960 VN.n9912 a_400_62400# 0.03fF
C10961 VN.n9913 a_400_62400# 0.01fF
C10962 VN.n9914 a_400_62400# 0.02fF
C10963 VN.n9915 a_400_62400# 0.11fF
C10964 VN.n9916 a_400_62400# 0.08fF
C10965 VN.n9917 a_400_62400# 0.04fF
C10966 VN.n9918 a_400_62400# 0.05fF
C10967 VN.n9919 a_400_62400# 1.34fF
C10968 VN.n9920 a_400_62400# 0.48fF
C10969 VN.n9921 a_400_62400# 2.51fF
C10970 VN.n9922 a_400_62400# 2.67fF
C10971 VN.t784 a_400_62400# 0.03fF
C10972 VN.n9923 a_400_62400# 0.32fF
C10973 VN.n9924 a_400_62400# 1.22fF
C10974 VN.n9925 a_400_62400# 0.07fF
C10975 VN.t1718 a_400_62400# 0.03fF
C10976 VN.n9926 a_400_62400# 0.16fF
C10977 VN.n9927 a_400_62400# 0.19fF
C10978 VN.n9929 a_400_62400# 2.53fF
C10979 VN.n9930 a_400_62400# 0.08fF
C10980 VN.n9931 a_400_62400# 0.04fF
C10981 VN.n9932 a_400_62400# 0.05fF
C10982 VN.n9933 a_400_62400# 1.33fF
C10983 VN.n9934 a_400_62400# 0.03fF
C10984 VN.n9935 a_400_62400# 0.01fF
C10985 VN.n9936 a_400_62400# 0.02fF
C10986 VN.n9937 a_400_62400# 0.11fF
C10987 VN.n9938 a_400_62400# 0.48fF
C10988 VN.n9939 a_400_62400# 2.48fF
C10989 VN.t1334 a_400_62400# 0.03fF
C10990 VN.n9940 a_400_62400# 0.32fF
C10991 VN.n9941 a_400_62400# 0.48fF
C10992 VN.n9942 a_400_62400# 0.81fF
C10993 VN.n9943 a_400_62400# 0.16fF
C10994 VN.t172 a_400_62400# 0.03fF
C10995 VN.n9944 a_400_62400# 0.19fF
C10996 VN.n9946 a_400_62400# 0.93fF
C10997 VN.n9947 a_400_62400# 0.30fF
C10998 VN.n9948 a_400_62400# 0.34fF
C10999 VN.n9949 a_400_62400# 0.12fF
C11000 VN.n9950 a_400_62400# 0.30fF
C11001 VN.n9951 a_400_62400# 0.93fF
C11002 VN.n9952 a_400_62400# 1.55fF
C11003 VN.n9953 a_400_62400# 0.29fF
C11004 VN.n9954 a_400_62400# 0.34fF
C11005 VN.n9955 a_400_62400# 0.12fF
C11006 VN.n9956 a_400_62400# 2.52fF
C11007 VN.t2437 a_400_62400# 0.03fF
C11008 VN.n9957 a_400_62400# 0.32fF
C11009 VN.n9958 a_400_62400# 1.22fF
C11010 VN.n9959 a_400_62400# 0.07fF
C11011 VN.t845 a_400_62400# 0.03fF
C11012 VN.n9960 a_400_62400# 0.16fF
C11013 VN.n9961 a_400_62400# 0.19fF
C11014 VN.n9963 a_400_62400# 0.33fF
C11015 VN.n9964 a_400_62400# 0.12fF
C11016 VN.n9965 a_400_62400# 0.28fF
C11017 VN.n9966 a_400_62400# 1.72fF
C11018 VN.n9967 a_400_62400# 0.71fF
C11019 VN.n9968 a_400_62400# 2.51fF
C11020 VN.n9969 a_400_62400# 0.16fF
C11021 VN.t668 a_400_62400# 0.03fF
C11022 VN.n9970 a_400_62400# 0.19fF
C11023 VN.t1793 a_400_62400# 0.03fF
C11024 VN.n9972 a_400_62400# 0.32fF
C11025 VN.n9973 a_400_62400# 0.48fF
C11026 VN.n9974 a_400_62400# 0.81fF
C11027 VN.n9975 a_400_62400# 0.03fF
C11028 VN.n9976 a_400_62400# 0.01fF
C11029 VN.n9977 a_400_62400# 0.02fF
C11030 VN.n9978 a_400_62400# 0.11fF
C11031 VN.n9979 a_400_62400# 0.08fF
C11032 VN.n9980 a_400_62400# 0.04fF
C11033 VN.n9981 a_400_62400# 0.05fF
C11034 VN.n9982 a_400_62400# 1.34fF
C11035 VN.n9983 a_400_62400# 0.48fF
C11036 VN.n9984 a_400_62400# 2.51fF
C11037 VN.n9985 a_400_62400# 2.67fF
C11038 VN.t410 a_400_62400# 0.03fF
C11039 VN.n9986 a_400_62400# 0.32fF
C11040 VN.n9987 a_400_62400# 1.22fF
C11041 VN.n9988 a_400_62400# 0.07fF
C11042 VN.t2509 a_400_62400# 0.03fF
C11043 VN.n9989 a_400_62400# 0.16fF
C11044 VN.n9990 a_400_62400# 0.19fF
C11045 VN.n9992 a_400_62400# 2.53fF
C11046 VN.n9993 a_400_62400# 0.08fF
C11047 VN.n9994 a_400_62400# 0.04fF
C11048 VN.n9995 a_400_62400# 0.05fF
C11049 VN.n9996 a_400_62400# 1.33fF
C11050 VN.n9997 a_400_62400# 0.03fF
C11051 VN.n9998 a_400_62400# 0.01fF
C11052 VN.n9999 a_400_62400# 0.02fF
C11053 VN.n10000 a_400_62400# 0.11fF
C11054 VN.n10001 a_400_62400# 0.48fF
C11055 VN.n10002 a_400_62400# 2.48fF
C11056 VN.t918 a_400_62400# 0.03fF
C11057 VN.n10003 a_400_62400# 0.32fF
C11058 VN.n10004 a_400_62400# 0.48fF
C11059 VN.n10005 a_400_62400# 0.81fF
C11060 VN.n10006 a_400_62400# 0.16fF
C11061 VN.t2328 a_400_62400# 0.03fF
C11062 VN.n10007 a_400_62400# 0.19fF
C11063 VN.n10009 a_400_62400# 0.93fF
C11064 VN.n10010 a_400_62400# 0.30fF
C11065 VN.n10011 a_400_62400# 0.34fF
C11066 VN.n10012 a_400_62400# 0.12fF
C11067 VN.n10013 a_400_62400# 0.30fF
C11068 VN.n10014 a_400_62400# 0.93fF
C11069 VN.n10015 a_400_62400# 1.55fF
C11070 VN.n10016 a_400_62400# 0.29fF
C11071 VN.n10017 a_400_62400# 0.34fF
C11072 VN.n10018 a_400_62400# 0.12fF
C11073 VN.n10019 a_400_62400# 2.52fF
C11074 VN.t2059 a_400_62400# 0.03fF
C11075 VN.n10020 a_400_62400# 0.32fF
C11076 VN.n10021 a_400_62400# 1.22fF
C11077 VN.n10022 a_400_62400# 0.07fF
C11078 VN.t488 a_400_62400# 0.03fF
C11079 VN.n10023 a_400_62400# 0.16fF
C11080 VN.n10024 a_400_62400# 0.19fF
C11081 VN.n10026 a_400_62400# 0.33fF
C11082 VN.n10027 a_400_62400# 0.12fF
C11083 VN.n10028 a_400_62400# 0.28fF
C11084 VN.n10029 a_400_62400# 1.23fF
C11085 VN.n10030 a_400_62400# 0.59fF
C11086 VN.n10031 a_400_62400# 2.51fF
C11087 VN.n10032 a_400_62400# 0.16fF
C11088 VN.t1463 a_400_62400# 0.03fF
C11089 VN.n10033 a_400_62400# 0.19fF
C11090 VN.t2580 a_400_62400# 0.03fF
C11091 VN.n10035 a_400_62400# 0.32fF
C11092 VN.n10036 a_400_62400# 0.48fF
C11093 VN.n10037 a_400_62400# 0.81fF
C11094 VN.n10038 a_400_62400# 0.03fF
C11095 VN.n10039 a_400_62400# 0.01fF
C11096 VN.n10040 a_400_62400# 0.02fF
C11097 VN.n10041 a_400_62400# 0.11fF
C11098 VN.n10042 a_400_62400# 0.08fF
C11099 VN.n10043 a_400_62400# 0.04fF
C11100 VN.n10044 a_400_62400# 0.05fF
C11101 VN.n10045 a_400_62400# 1.34fF
C11102 VN.n10046 a_400_62400# 0.48fF
C11103 VN.n10047 a_400_62400# 2.51fF
C11104 VN.n10048 a_400_62400# 2.67fF
C11105 VN.t1188 a_400_62400# 0.03fF
C11106 VN.n10049 a_400_62400# 0.32fF
C11107 VN.n10050 a_400_62400# 1.22fF
C11108 VN.n10051 a_400_62400# 0.07fF
C11109 VN.t2142 a_400_62400# 0.03fF
C11110 VN.n10052 a_400_62400# 0.16fF
C11111 VN.n10053 a_400_62400# 0.19fF
C11112 VN.n10055 a_400_62400# 2.53fF
C11113 VN.n10056 a_400_62400# 0.08fF
C11114 VN.n10057 a_400_62400# 0.04fF
C11115 VN.n10058 a_400_62400# 0.05fF
C11116 VN.n10059 a_400_62400# 1.33fF
C11117 VN.n10060 a_400_62400# 0.03fF
C11118 VN.n10061 a_400_62400# 0.01fF
C11119 VN.n10062 a_400_62400# 0.02fF
C11120 VN.n10063 a_400_62400# 0.11fF
C11121 VN.n10064 a_400_62400# 0.48fF
C11122 VN.n10065 a_400_62400# 2.48fF
C11123 VN.t1711 a_400_62400# 0.03fF
C11124 VN.n10066 a_400_62400# 0.32fF
C11125 VN.n10067 a_400_62400# 0.48fF
C11126 VN.n10068 a_400_62400# 0.81fF
C11127 VN.n10069 a_400_62400# 0.16fF
C11128 VN.t591 a_400_62400# 0.03fF
C11129 VN.n10070 a_400_62400# 0.19fF
C11130 VN.n10072 a_400_62400# 0.93fF
C11131 VN.n10073 a_400_62400# 0.30fF
C11132 VN.n10074 a_400_62400# 0.34fF
C11133 VN.n10075 a_400_62400# 0.12fF
C11134 VN.n10076 a_400_62400# 0.30fF
C11135 VN.n10077 a_400_62400# 0.93fF
C11136 VN.n10078 a_400_62400# 1.55fF
C11137 VN.n10079 a_400_62400# 0.29fF
C11138 VN.n10080 a_400_62400# 0.34fF
C11139 VN.n10081 a_400_62400# 0.12fF
C11140 VN.n10082 a_400_62400# 2.52fF
C11141 VN.t319 a_400_62400# 0.03fF
C11142 VN.n10083 a_400_62400# 0.32fF
C11143 VN.n10084 a_400_62400# 1.22fF
C11144 VN.n10085 a_400_62400# 0.07fF
C11145 VN.t1392 a_400_62400# 0.03fF
C11146 VN.n10086 a_400_62400# 0.16fF
C11147 VN.n10087 a_400_62400# 0.19fF
C11148 VN.n10089 a_400_62400# 0.33fF
C11149 VN.n10090 a_400_62400# 0.12fF
C11150 VN.n10091 a_400_62400# 0.28fF
C11151 VN.n10092 a_400_62400# 1.23fF
C11152 VN.n10093 a_400_62400# 0.59fF
C11153 VN.n10094 a_400_62400# 2.51fF
C11154 VN.n10095 a_400_62400# 0.16fF
C11155 VN.t2244 a_400_62400# 0.03fF
C11156 VN.n10096 a_400_62400# 0.19fF
C11157 VN.t839 a_400_62400# 0.03fF
C11158 VN.n10098 a_400_62400# 0.32fF
C11159 VN.n10099 a_400_62400# 0.48fF
C11160 VN.n10100 a_400_62400# 0.81fF
C11161 VN.n10101 a_400_62400# 0.03fF
C11162 VN.n10102 a_400_62400# 0.01fF
C11163 VN.n10103 a_400_62400# 0.02fF
C11164 VN.n10104 a_400_62400# 0.11fF
C11165 VN.n10105 a_400_62400# 0.08fF
C11166 VN.n10106 a_400_62400# 0.04fF
C11167 VN.n10107 a_400_62400# 0.05fF
C11168 VN.n10108 a_400_62400# 1.34fF
C11169 VN.n10109 a_400_62400# 0.48fF
C11170 VN.n10110 a_400_62400# 2.51fF
C11171 VN.n10111 a_400_62400# 2.67fF
C11172 VN.t1968 a_400_62400# 0.03fF
C11173 VN.n10112 a_400_62400# 0.32fF
C11174 VN.n10113 a_400_62400# 1.22fF
C11175 VN.n10114 a_400_62400# 0.07fF
C11176 VN.t527 a_400_62400# 0.03fF
C11177 VN.n10115 a_400_62400# 0.16fF
C11178 VN.n10116 a_400_62400# 0.19fF
C11179 VN.n10118 a_400_62400# 2.53fF
C11180 VN.n10119 a_400_62400# 0.08fF
C11181 VN.n10120 a_400_62400# 0.04fF
C11182 VN.n10121 a_400_62400# 0.05fF
C11183 VN.n10122 a_400_62400# 1.33fF
C11184 VN.n10123 a_400_62400# 0.03fF
C11185 VN.n10124 a_400_62400# 0.01fF
C11186 VN.n10125 a_400_62400# 0.02fF
C11187 VN.n10126 a_400_62400# 0.11fF
C11188 VN.n10127 a_400_62400# 0.48fF
C11189 VN.n10128 a_400_62400# 2.48fF
C11190 VN.t2502 a_400_62400# 0.03fF
C11191 VN.n10129 a_400_62400# 0.32fF
C11192 VN.n10130 a_400_62400# 0.48fF
C11193 VN.n10131 a_400_62400# 0.81fF
C11194 VN.n10132 a_400_62400# 0.16fF
C11195 VN.t1382 a_400_62400# 0.03fF
C11196 VN.n10133 a_400_62400# 0.19fF
C11197 VN.n10135 a_400_62400# 0.93fF
C11198 VN.n10136 a_400_62400# 0.30fF
C11199 VN.n10137 a_400_62400# 0.34fF
C11200 VN.n10138 a_400_62400# 0.12fF
C11201 VN.n10139 a_400_62400# 0.30fF
C11202 VN.n10140 a_400_62400# 0.93fF
C11203 VN.n10141 a_400_62400# 1.55fF
C11204 VN.n10142 a_400_62400# 0.29fF
C11205 VN.n10143 a_400_62400# 0.34fF
C11206 VN.n10144 a_400_62400# 0.12fF
C11207 VN.n10145 a_400_62400# 2.52fF
C11208 VN.t1101 a_400_62400# 0.03fF
C11209 VN.n10146 a_400_62400# 0.32fF
C11210 VN.n10147 a_400_62400# 1.22fF
C11211 VN.n10148 a_400_62400# 0.07fF
C11212 VN.t2181 a_400_62400# 0.03fF
C11213 VN.n10149 a_400_62400# 0.16fF
C11214 VN.n10150 a_400_62400# 0.19fF
C11215 VN.n10152 a_400_62400# 0.33fF
C11216 VN.n10153 a_400_62400# 0.12fF
C11217 VN.n10154 a_400_62400# 0.28fF
C11218 VN.n10155 a_400_62400# 1.23fF
C11219 VN.n10156 a_400_62400# 0.59fF
C11220 VN.n10157 a_400_62400# 2.51fF
C11221 VN.n10158 a_400_62400# 0.16fF
C11222 VN.t516 a_400_62400# 0.03fF
C11223 VN.n10159 a_400_62400# 0.19fF
C11224 VN.t1640 a_400_62400# 0.03fF
C11225 VN.n10161 a_400_62400# 0.32fF
C11226 VN.n10162 a_400_62400# 0.48fF
C11227 VN.n10163 a_400_62400# 0.81fF
C11228 VN.n10164 a_400_62400# 0.03fF
C11229 VN.n10165 a_400_62400# 0.01fF
C11230 VN.n10166 a_400_62400# 0.02fF
C11231 VN.n10167 a_400_62400# 0.11fF
C11232 VN.n10168 a_400_62400# 0.08fF
C11233 VN.n10169 a_400_62400# 0.04fF
C11234 VN.n10170 a_400_62400# 0.05fF
C11235 VN.n10171 a_400_62400# 1.34fF
C11236 VN.n10172 a_400_62400# 0.48fF
C11237 VN.n10173 a_400_62400# 2.45fF
C11238 VN.n10174 a_400_62400# 2.67fF
C11239 VN.t234 a_400_62400# 0.03fF
C11240 VN.n10175 a_400_62400# 0.32fF
C11241 VN.n10176 a_400_62400# 1.22fF
C11242 VN.n10177 a_400_62400# 0.07fF
C11243 VN.t1313 a_400_62400# 0.03fF
C11244 VN.n10178 a_400_62400# 0.16fF
C11245 VN.n10179 a_400_62400# 0.19fF
C11246 VN.n10181 a_400_62400# 2.53fF
C11247 VN.n10182 a_400_62400# 0.85fF
C11248 VN.n10183 a_400_62400# 0.05fF
C11249 VN.n10184 a_400_62400# 0.09fF
C11250 VN.n10185 a_400_62400# 0.07fF
C11251 VN.n10186 a_400_62400# 1.16fF
C11252 VN.n10187 a_400_62400# 0.01fF
C11253 VN.n10188 a_400_62400# 0.01fF
C11254 VN.n10189 a_400_62400# 0.01fF
C11255 VN.n10190 a_400_62400# 0.09fF
C11256 VN.n10191 a_400_62400# 0.91fF
C11257 VN.n10192 a_400_62400# 0.18fF
C11258 VN.t768 a_400_62400# 0.03fF
C11259 VN.n10193 a_400_62400# 0.32fF
C11260 VN.n10194 a_400_62400# 0.48fF
C11261 VN.n10195 a_400_62400# 0.81fF
C11262 VN.n10196 a_400_62400# 0.16fF
C11263 VN.t2285 a_400_62400# 0.03fF
C11264 VN.n10197 a_400_62400# 0.19fF
C11265 VN.n10199 a_400_62400# 0.93fF
C11266 VN.n10200 a_400_62400# 0.30fF
C11267 VN.n10201 a_400_62400# 0.34fF
C11268 VN.n10202 a_400_62400# 0.12fF
C11269 VN.n10203 a_400_62400# 0.30fF
C11270 VN.n10204 a_400_62400# 0.93fF
C11271 VN.n10205 a_400_62400# 1.55fF
C11272 VN.n10206 a_400_62400# 0.29fF
C11273 VN.n10207 a_400_62400# 0.34fF
C11274 VN.n10208 a_400_62400# 0.12fF
C11275 VN.n10209 a_400_62400# 3.10fF
C11276 VN.t1881 a_400_62400# 0.03fF
C11277 VN.n10210 a_400_62400# 0.32fF
C11278 VN.n10211 a_400_62400# 1.22fF
C11279 VN.n10212 a_400_62400# 0.07fF
C11280 VN.t452 a_400_62400# 0.03fF
C11281 VN.n10213 a_400_62400# 0.16fF
C11282 VN.n10214 a_400_62400# 0.19fF
C11283 VN.n10216 a_400_62400# 2.51fF
C11284 VN.n10217 a_400_62400# 0.61fF
C11285 VN.n10218 a_400_62400# 0.30fF
C11286 VN.n10219 a_400_62400# 0.51fF
C11287 VN.n10220 a_400_62400# 0.21fF
C11288 VN.n10221 a_400_62400# 0.38fF
C11289 VN.n10222 a_400_62400# 0.29fF
C11290 VN.n10223 a_400_62400# 0.40fF
C11291 VN.n10224 a_400_62400# 0.28fF
C11292 VN.t2543 a_400_62400# 0.03fF
C11293 VN.n10225 a_400_62400# 0.32fF
C11294 VN.n10226 a_400_62400# 0.48fF
C11295 VN.n10227 a_400_62400# 0.81fF
C11296 VN.n10228 a_400_62400# 0.16fF
C11297 VN.t1416 a_400_62400# 0.03fF
C11298 VN.n10229 a_400_62400# 0.19fF
C11299 VN.n10231 a_400_62400# 0.06fF
C11300 VN.n10232 a_400_62400# 0.04fF
C11301 VN.n10233 a_400_62400# 0.04fF
C11302 VN.n10234 a_400_62400# 0.14fF
C11303 VN.n10235 a_400_62400# 0.48fF
C11304 VN.n10236 a_400_62400# 0.50fF
C11305 VN.n10237 a_400_62400# 0.14fF
C11306 VN.n10238 a_400_62400# 0.16fF
C11307 VN.n10239 a_400_62400# 0.09fF
C11308 VN.n10240 a_400_62400# 0.16fF
C11309 VN.n10241 a_400_62400# 0.24fF
C11310 VN.n10242 a_400_62400# 5.35fF
C11311 VN.t1147 a_400_62400# 0.03fF
C11312 VN.n10243 a_400_62400# 0.32fF
C11313 VN.n10244 a_400_62400# 1.22fF
C11314 VN.n10245 a_400_62400# 0.07fF
C11315 VN.t2098 a_400_62400# 0.03fF
C11316 VN.n10246 a_400_62400# 0.16fF
C11317 VN.n10247 a_400_62400# 0.19fF
C11318 VN.n10249 a_400_62400# 0.33fF
C11319 VN.n10250 a_400_62400# 0.12fF
C11320 VN.n10251 a_400_62400# 0.28fF
C11321 VN.n10252 a_400_62400# 1.72fF
C11322 VN.n10253 a_400_62400# 0.71fF
C11323 VN.n10254 a_400_62400# 2.51fF
C11324 VN.n10255 a_400_62400# 0.16fF
C11325 VN.t423 a_400_62400# 0.03fF
C11326 VN.n10256 a_400_62400# 0.19fF
C11327 VN.t1559 a_400_62400# 0.03fF
C11328 VN.n10258 a_400_62400# 0.32fF
C11329 VN.n10259 a_400_62400# 0.48fF
C11330 VN.n10260 a_400_62400# 0.81fF
C11331 VN.n10261 a_400_62400# 0.95fF
C11332 VN.n10262 a_400_62400# 2.11fF
C11333 VN.n10263 a_400_62400# 3.28fF
C11334 VN.t608 a_400_62400# 0.03fF
C11335 VN.n10264 a_400_62400# 0.32fF
C11336 VN.n10265 a_400_62400# 1.22fF
C11337 VN.n10266 a_400_62400# 0.07fF
C11338 VN.t1221 a_400_62400# 0.03fF
C11339 VN.n10267 a_400_62400# 0.16fF
C11340 VN.n10268 a_400_62400# 0.19fF
C11341 VN.n10270 a_400_62400# 2.53fF
C11342 VN.n10271 a_400_62400# 0.08fF
C11343 VN.n10272 a_400_62400# 0.04fF
C11344 VN.n10273 a_400_62400# 0.05fF
C11345 VN.n10274 a_400_62400# 1.33fF
C11346 VN.n10275 a_400_62400# 0.03fF
C11347 VN.n10276 a_400_62400# 0.01fF
C11348 VN.n10277 a_400_62400# 0.02fF
C11349 VN.n10278 a_400_62400# 0.11fF
C11350 VN.n10279 a_400_62400# 0.48fF
C11351 VN.n10280 a_400_62400# 2.48fF
C11352 VN.t688 a_400_62400# 0.03fF
C11353 VN.n10281 a_400_62400# 0.32fF
C11354 VN.n10282 a_400_62400# 0.48fF
C11355 VN.n10283 a_400_62400# 0.81fF
C11356 VN.n10284 a_400_62400# 0.16fF
C11357 VN.t2070 a_400_62400# 0.03fF
C11358 VN.n10285 a_400_62400# 0.19fF
C11359 VN.n10287 a_400_62400# 0.93fF
C11360 VN.n10288 a_400_62400# 0.30fF
C11361 VN.n10289 a_400_62400# 0.34fF
C11362 VN.n10290 a_400_62400# 0.12fF
C11363 VN.n10291 a_400_62400# 0.30fF
C11364 VN.n10292 a_400_62400# 0.93fF
C11365 VN.n10293 a_400_62400# 1.55fF
C11366 VN.n10294 a_400_62400# 0.29fF
C11367 VN.n10295 a_400_62400# 0.34fF
C11368 VN.n10296 a_400_62400# 0.12fF
C11369 VN.n10297 a_400_62400# 2.52fF
C11370 VN.t2262 a_400_62400# 0.03fF
C11371 VN.n10298 a_400_62400# 0.32fF
C11372 VN.n10299 a_400_62400# 1.22fF
C11373 VN.n10300 a_400_62400# 0.07fF
C11374 VN.t207 a_400_62400# 0.03fF
C11375 VN.n10301 a_400_62400# 0.16fF
C11376 VN.n10302 a_400_62400# 0.19fF
C11377 VN.n10304 a_400_62400# 27.83fF
C11378 VN.n10305 a_400_62400# 0.09fF
C11379 VN.n10306 a_400_62400# 0.27fF
C11380 VN.n10307 a_400_62400# 0.12fF
C11381 VN.n10308 a_400_62400# 0.28fF
C11382 VN.n10309 a_400_62400# 0.13fF
C11383 VN.n10310 a_400_62400# 0.40fF
C11384 VN.n10311 a_400_62400# 0.93fF
C11385 VN.n10312 a_400_62400# 0.60fF
C11386 VN.n10313 a_400_62400# 3.12fF
C11387 VN.n10314 a_400_62400# 0.16fF
C11388 VN.t121 a_400_62400# 0.03fF
C11389 VN.n10315 a_400_62400# 0.19fF
C11390 VN.t1293 a_400_62400# 0.03fF
C11391 VN.n10317 a_400_62400# 0.32fF
C11392 VN.n10318 a_400_62400# 0.48fF
C11393 VN.n10319 a_400_62400# 0.81fF
C11394 VN.n10320 a_400_62400# 2.54fF
C11395 VN.n10321 a_400_62400# 0.23fF
C11396 VN.n10322 a_400_62400# 1.02fF
C11397 VN.n10323 a_400_62400# 0.42fF
C11398 VN.n10324 a_400_62400# 0.34fF
C11399 VN.n10325 a_400_62400# 0.40fF
C11400 VN.n10326 a_400_62400# 0.63fF
C11401 VN.n10327 a_400_62400# 0.21fF
C11402 VN.n10328 a_400_62400# 2.58fF
C11403 VN.t925 a_400_62400# 0.03fF
C11404 VN.n10329 a_400_62400# 0.16fF
C11405 VN.n10330 a_400_62400# 0.19fF
C11406 VN.t2403 a_400_62400# 0.03fF
C11407 VN.n10332 a_400_62400# 0.32fF
C11408 VN.n10333 a_400_62400# 1.22fF
C11409 VN.n10334 a_400_62400# 0.07fF
C11410 VN.n10335 a_400_62400# 2.51fF
C11411 VN.n10336 a_400_62400# 0.16fF
C11412 VN.t2564 a_400_62400# 0.03fF
C11413 VN.n10337 a_400_62400# 0.19fF
C11414 VN.t673 a_400_62400# 0.03fF
C11415 VN.n10339 a_400_62400# 1.63fF
C11416 VN.n10340 a_400_62400# 0.81fF
C11417 VN.n10341 a_400_62400# 1.21fF
C11418 VN.n10342 a_400_62400# 1.54fF
C11419 VN.n10343 a_400_62400# 4.06fF
C11420 VN.t148 a_400_62400# 28.64fF
C11421 VN.n10344 a_400_62400# 28.43fF
C11422 VN.n10346 a_400_62400# 0.50fF
C11423 VN.n10347 a_400_62400# 0.31fF
C11424 VN.n10348 a_400_62400# 3.88fF
C11425 VN.n10349 a_400_62400# 3.29fF
C11426 VN.n10350 a_400_62400# 2.62fF
C11427 VN.n10351 a_400_62400# 5.27fF
C11428 VN.n10352 a_400_62400# 0.34fF
C11429 VN.n10353 a_400_62400# 0.02fF
C11430 VN.t2066 a_400_62400# 0.03fF
C11431 VN.n10354 a_400_62400# 0.34fF
C11432 VN.t2368 a_400_62400# 0.03fF
C11433 VN.n10355 a_400_62400# 1.28fF
C11434 VN.n10356 a_400_62400# 0.94fF
C11435 VN.n10357 a_400_62400# 1.04fF
C11436 VN.n10358 a_400_62400# 2.58fF
C11437 VN.n10359 a_400_62400# 2.51fF
C11438 VN.n10360 a_400_62400# 0.16fF
C11439 VN.t1196 a_400_62400# 0.03fF
C11440 VN.n10361 a_400_62400# 0.19fF
C11441 VN.t2332 a_400_62400# 0.03fF
C11442 VN.n10363 a_400_62400# 0.32fF
C11443 VN.n10364 a_400_62400# 0.48fF
C11444 VN.n10365 a_400_62400# 0.81fF
C11445 VN.n10366 a_400_62400# 2.03fF
C11446 VN.n10367 a_400_62400# 4.01fF
C11447 VN.t1496 a_400_62400# 0.03fF
C11448 VN.n10368 a_400_62400# 0.32fF
C11449 VN.n10369 a_400_62400# 1.22fF
C11450 VN.n10370 a_400_62400# 0.07fF
C11451 VN.t1272 a_400_62400# 0.03fF
C11452 VN.n10371 a_400_62400# 0.16fF
C11453 VN.n10372 a_400_62400# 0.19fF
C11454 VN.n10374 a_400_62400# 2.53fF
C11455 VN.n10375 a_400_62400# 2.51fF
C11456 VN.t1468 a_400_62400# 0.03fF
C11457 VN.n10376 a_400_62400# 0.32fF
C11458 VN.n10377 a_400_62400# 0.48fF
C11459 VN.n10378 a_400_62400# 0.81fF
C11460 VN.n10379 a_400_62400# 0.16fF
C11461 VN.t327 a_400_62400# 0.03fF
C11462 VN.n10380 a_400_62400# 0.19fF
C11463 VN.n10382 a_400_62400# 0.93fF
C11464 VN.n10383 a_400_62400# 1.55fF
C11465 VN.n10384 a_400_62400# 0.29fF
C11466 VN.n10385 a_400_62400# 2.52fF
C11467 VN.t630 a_400_62400# 0.03fF
C11468 VN.n10386 a_400_62400# 0.32fF
C11469 VN.n10387 a_400_62400# 1.22fF
C11470 VN.n10388 a_400_62400# 0.07fF
C11471 VN.t528 a_400_62400# 0.03fF
C11472 VN.n10389 a_400_62400# 0.16fF
C11473 VN.n10390 a_400_62400# 0.19fF
C11474 VN.n10392 a_400_62400# 1.04fF
C11475 VN.n10393 a_400_62400# 2.60fF
C11476 VN.n10394 a_400_62400# 2.51fF
C11477 VN.n10395 a_400_62400# 0.16fF
C11478 VN.t1972 a_400_62400# 0.03fF
C11479 VN.n10396 a_400_62400# 0.19fF
C11480 VN.t598 a_400_62400# 0.03fF
C11481 VN.n10398 a_400_62400# 0.32fF
C11482 VN.n10399 a_400_62400# 0.48fF
C11483 VN.n10400 a_400_62400# 0.81fF
C11484 VN.n10401 a_400_62400# 2.46fF
C11485 VN.n10402 a_400_62400# 4.01fF
C11486 VN.t2287 a_400_62400# 0.03fF
C11487 VN.n10403 a_400_62400# 0.32fF
C11488 VN.n10404 a_400_62400# 1.22fF
C11489 VN.n10405 a_400_62400# 0.07fF
C11490 VN.t2183 a_400_62400# 0.03fF
C11491 VN.n10406 a_400_62400# 0.16fF
C11492 VN.n10407 a_400_62400# 0.19fF
C11493 VN.n10409 a_400_62400# 2.53fF
C11494 VN.n10410 a_400_62400# 2.51fF
C11495 VN.t2253 a_400_62400# 0.03fF
C11496 VN.n10411 a_400_62400# 0.32fF
C11497 VN.n10412 a_400_62400# 0.48fF
C11498 VN.n10413 a_400_62400# 0.81fF
C11499 VN.n10414 a_400_62400# 0.16fF
C11500 VN.t1104 a_400_62400# 0.03fF
C11501 VN.n10415 a_400_62400# 0.19fF
C11502 VN.n10417 a_400_62400# 0.93fF
C11503 VN.n10418 a_400_62400# 1.55fF
C11504 VN.n10419 a_400_62400# 0.29fF
C11505 VN.n10420 a_400_62400# 2.52fF
C11506 VN.t1418 a_400_62400# 0.03fF
C11507 VN.n10421 a_400_62400# 0.32fF
C11508 VN.n10422 a_400_62400# 1.22fF
C11509 VN.n10423 a_400_62400# 0.07fF
C11510 VN.t1317 a_400_62400# 0.03fF
C11511 VN.n10424 a_400_62400# 0.16fF
C11512 VN.n10425 a_400_62400# 0.19fF
C11513 VN.n10427 a_400_62400# 1.05fF
C11514 VN.n10428 a_400_62400# 3.07fF
C11515 VN.n10429 a_400_62400# 2.51fF
C11516 VN.n10430 a_400_62400# 0.16fF
C11517 VN.t1588 a_400_62400# 0.03fF
C11518 VN.n10431 a_400_62400# 0.19fF
C11519 VN.t191 a_400_62400# 0.03fF
C11520 VN.n10433 a_400_62400# 0.32fF
C11521 VN.n10434 a_400_62400# 0.48fF
C11522 VN.n10435 a_400_62400# 0.81fF
C11523 VN.n10436 a_400_62400# 2.46fF
C11524 VN.n10437 a_400_62400# 2.91fF
C11525 VN.t1885 a_400_62400# 0.03fF
C11526 VN.n10438 a_400_62400# 0.32fF
C11527 VN.n10439 a_400_62400# 1.22fF
C11528 VN.n10440 a_400_62400# 0.07fF
C11529 VN.t1770 a_400_62400# 0.03fF
C11530 VN.n10441 a_400_62400# 0.16fF
C11531 VN.n10442 a_400_62400# 0.19fF
C11532 VN.n10444 a_400_62400# 2.53fF
C11533 VN.n10445 a_400_62400# 2.51fF
C11534 VN.t1849 a_400_62400# 0.03fF
C11535 VN.n10446 a_400_62400# 0.32fF
C11536 VN.n10447 a_400_62400# 0.48fF
C11537 VN.n10448 a_400_62400# 0.81fF
C11538 VN.n10449 a_400_62400# 0.16fF
C11539 VN.t723 a_400_62400# 0.03fF
C11540 VN.n10450 a_400_62400# 0.19fF
C11541 VN.n10452 a_400_62400# 0.93fF
C11542 VN.n10453 a_400_62400# 1.55fF
C11543 VN.n10454 a_400_62400# 0.29fF
C11544 VN.n10455 a_400_62400# 2.52fF
C11545 VN.t1013 a_400_62400# 0.03fF
C11546 VN.n10456 a_400_62400# 0.32fF
C11547 VN.n10457 a_400_62400# 1.22fF
C11548 VN.n10458 a_400_62400# 0.07fF
C11549 VN.t898 a_400_62400# 0.03fF
C11550 VN.n10459 a_400_62400# 0.16fF
C11551 VN.n10460 a_400_62400# 0.19fF
C11552 VN.n10462 a_400_62400# 1.04fF
C11553 VN.n10463 a_400_62400# 2.60fF
C11554 VN.n10464 a_400_62400# 2.51fF
C11555 VN.n10465 a_400_62400# 0.16fF
C11556 VN.t2495 a_400_62400# 0.03fF
C11557 VN.n10466 a_400_62400# 0.19fF
C11558 VN.t977 a_400_62400# 0.03fF
C11559 VN.n10468 a_400_62400# 0.32fF
C11560 VN.n10469 a_400_62400# 0.48fF
C11561 VN.n10470 a_400_62400# 0.81fF
C11562 VN.n10471 a_400_62400# 2.46fF
C11563 VN.n10472 a_400_62400# 4.01fF
C11564 VN.t139 a_400_62400# 0.03fF
C11565 VN.n10473 a_400_62400# 0.32fF
C11566 VN.n10474 a_400_62400# 1.22fF
C11567 VN.n10475 a_400_62400# 0.07fF
C11568 VN.t2561 a_400_62400# 0.03fF
C11569 VN.n10476 a_400_62400# 0.16fF
C11570 VN.n10477 a_400_62400# 0.19fF
C11571 VN.n10479 a_400_62400# 2.53fF
C11572 VN.n10480 a_400_62400# 2.51fF
C11573 VN.t244 a_400_62400# 0.03fF
C11574 VN.n10481 a_400_62400# 0.32fF
C11575 VN.n10482 a_400_62400# 0.48fF
C11576 VN.n10483 a_400_62400# 0.81fF
C11577 VN.n10484 a_400_62400# 0.16fF
C11578 VN.t1631 a_400_62400# 0.03fF
C11579 VN.n10485 a_400_62400# 0.19fF
C11580 VN.n10487 a_400_62400# 0.93fF
C11581 VN.n10488 a_400_62400# 1.55fF
C11582 VN.n10489 a_400_62400# 0.29fF
C11583 VN.n10490 a_400_62400# 2.52fF
C11584 VN.t1934 a_400_62400# 0.03fF
C11585 VN.n10491 a_400_62400# 0.32fF
C11586 VN.n10492 a_400_62400# 1.22fF
C11587 VN.n10493 a_400_62400# 0.07fF
C11588 VN.t1693 a_400_62400# 0.03fF
C11589 VN.n10494 a_400_62400# 0.16fF
C11590 VN.n10495 a_400_62400# 0.19fF
C11591 VN.n10497 a_400_62400# 1.04fF
C11592 VN.n10498 a_400_62400# 2.60fF
C11593 VN.n10499 a_400_62400# 2.51fF
C11594 VN.n10500 a_400_62400# 0.16fF
C11595 VN.t760 a_400_62400# 0.03fF
C11596 VN.n10501 a_400_62400# 0.19fF
C11597 VN.t1892 a_400_62400# 0.03fF
C11598 VN.n10503 a_400_62400# 0.32fF
C11599 VN.n10504 a_400_62400# 0.48fF
C11600 VN.n10505 a_400_62400# 0.81fF
C11601 VN.n10506 a_400_62400# 2.46fF
C11602 VN.n10507 a_400_62400# 4.01fF
C11603 VN.t1061 a_400_62400# 0.03fF
C11604 VN.n10508 a_400_62400# 0.32fF
C11605 VN.n10509 a_400_62400# 1.22fF
C11606 VN.n10510 a_400_62400# 0.07fF
C11607 VN.t823 a_400_62400# 0.03fF
C11608 VN.n10511 a_400_62400# 0.16fF
C11609 VN.n10512 a_400_62400# 0.19fF
C11610 VN.n10514 a_400_62400# 2.53fF
C11611 VN.n10515 a_400_62400# 2.51fF
C11612 VN.t1019 a_400_62400# 0.03fF
C11613 VN.n10516 a_400_62400# 0.32fF
C11614 VN.n10517 a_400_62400# 0.48fF
C11615 VN.n10518 a_400_62400# 0.81fF
C11616 VN.n10519 a_400_62400# 0.16fF
C11617 VN.t2416 a_400_62400# 0.03fF
C11618 VN.n10520 a_400_62400# 0.19fF
C11619 VN.n10522 a_400_62400# 0.93fF
C11620 VN.n10523 a_400_62400# 1.55fF
C11621 VN.n10524 a_400_62400# 0.29fF
C11622 VN.n10525 a_400_62400# 2.52fF
C11623 VN.t187 a_400_62400# 0.03fF
C11624 VN.n10526 a_400_62400# 0.32fF
C11625 VN.n10527 a_400_62400# 1.22fF
C11626 VN.n10528 a_400_62400# 0.07fF
C11627 VN.t2483 a_400_62400# 0.03fF
C11628 VN.n10529 a_400_62400# 0.16fF
C11629 VN.n10530 a_400_62400# 0.19fF
C11630 VN.n10532 a_400_62400# 1.04fF
C11631 VN.n10533 a_400_62400# 2.60fF
C11632 VN.n10534 a_400_62400# 2.51fF
C11633 VN.n10535 a_400_62400# 0.16fF
C11634 VN.t1554 a_400_62400# 0.03fF
C11635 VN.n10536 a_400_62400# 0.19fF
C11636 VN.t149 a_400_62400# 0.03fF
C11637 VN.n10538 a_400_62400# 0.32fF
C11638 VN.n10539 a_400_62400# 0.48fF
C11639 VN.n10540 a_400_62400# 0.81fF
C11640 VN.n10541 a_400_62400# 0.04fF
C11641 VN.n10542 a_400_62400# 0.08fF
C11642 VN.n10543 a_400_62400# 1.20fF
C11643 VN.n10544 a_400_62400# 1.48fF
C11644 VN.n10545 a_400_62400# 3.99fF
C11645 VN.t1845 a_400_62400# 0.03fF
C11646 VN.n10546 a_400_62400# 0.32fF
C11647 VN.n10547 a_400_62400# 1.22fF
C11648 VN.n10548 a_400_62400# 0.07fF
C11649 VN.t1619 a_400_62400# 0.03fF
C11650 VN.n10549 a_400_62400# 0.16fF
C11651 VN.n10550 a_400_62400# 0.19fF
C11652 VN.n10552 a_400_62400# 0.93fF
C11653 VN.n10553 a_400_62400# 1.55fF
C11654 VN.n10554 a_400_62400# 0.29fF
C11655 VN.n10555 a_400_62400# 2.53fF
C11656 VN.n10556 a_400_62400# 0.16fF
C11657 VN.t680 a_400_62400# 0.03fF
C11658 VN.n10557 a_400_62400# 0.19fF
C11659 VN.t1812 a_400_62400# 0.03fF
C11660 VN.n10559 a_400_62400# 0.32fF
C11661 VN.n10560 a_400_62400# 0.48fF
C11662 VN.n10561 a_400_62400# 0.81fF
C11663 VN.n10562 a_400_62400# 1.47fF
C11664 VN.n10563 a_400_62400# 0.91fF
C11665 VN.n10564 a_400_62400# 0.73fF
C11666 VN.n10565 a_400_62400# 0.42fF
C11667 VN.n10566 a_400_62400# 2.45fF
C11668 VN.t973 a_400_62400# 0.03fF
C11669 VN.n10567 a_400_62400# 0.32fF
C11670 VN.n10568 a_400_62400# 1.22fF
C11671 VN.n10569 a_400_62400# 0.07fF
C11672 VN.t859 a_400_62400# 0.03fF
C11673 VN.n10570 a_400_62400# 0.16fF
C11674 VN.n10571 a_400_62400# 0.19fF
C11675 VN.n10573 a_400_62400# 2.51fF
C11676 VN.n10574 a_400_62400# 0.56fF
C11677 VN.n10575 a_400_62400# 0.64fF
C11678 VN.n10576 a_400_62400# 0.12fF
C11679 VN.n10577 a_400_62400# 0.44fF
C11680 VN.n10578 a_400_62400# 0.40fF
C11681 VN.n10579 a_400_62400# 1.03fF
C11682 VN.n10580 a_400_62400# 0.79fF
C11683 VN.t937 a_400_62400# 0.03fF
C11684 VN.n10581 a_400_62400# 0.32fF
C11685 VN.n10582 a_400_62400# 0.48fF
C11686 VN.n10583 a_400_62400# 0.81fF
C11687 VN.n10584 a_400_62400# 0.16fF
C11688 VN.t2340 a_400_62400# 0.03fF
C11689 VN.n10585 a_400_62400# 0.19fF
C11690 VN.n10587 a_400_62400# 3.50fF
C11691 VN.n10588 a_400_62400# 2.89fF
C11692 VN.t79 a_400_62400# 0.03fF
C11693 VN.n10589 a_400_62400# 0.32fF
C11694 VN.n10590 a_400_62400# 1.22fF
C11695 VN.n10591 a_400_62400# 0.07fF
C11696 VN.t2521 a_400_62400# 0.03fF
C11697 VN.n10592 a_400_62400# 0.16fF
C11698 VN.n10593 a_400_62400# 0.19fF
C11699 VN.n10595 a_400_62400# 2.51fF
C11700 VN.n10596 a_400_62400# 0.56fF
C11701 VN.n10597 a_400_62400# 0.64fF
C11702 VN.n10598 a_400_62400# 0.47fF
C11703 VN.n10599 a_400_62400# 0.40fF
C11704 VN.n10600 a_400_62400# 1.70fF
C11705 VN.t428 a_400_62400# 0.03fF
C11706 VN.n10601 a_400_62400# 0.32fF
C11707 VN.n10602 a_400_62400# 0.48fF
C11708 VN.n10603 a_400_62400# 0.81fF
C11709 VN.n10604 a_400_62400# 0.16fF
C11710 VN.t1776 a_400_62400# 0.03fF
C11711 VN.n10605 a_400_62400# 0.19fF
C11712 VN.n10607 a_400_62400# 1.05fF
C11713 VN.n10608 a_400_62400# 3.07fF
C11714 VN.n10609 a_400_62400# 2.71fF
C11715 VN.t2220 a_400_62400# 0.03fF
C11716 VN.n10610 a_400_62400# 0.32fF
C11717 VN.n10611 a_400_62400# 1.22fF
C11718 VN.n10612 a_400_62400# 0.07fF
C11719 VN.t1976 a_400_62400# 0.03fF
C11720 VN.n10613 a_400_62400# 0.16fF
C11721 VN.n10614 a_400_62400# 0.19fF
C11722 VN.n10616 a_400_62400# 2.53fF
C11723 VN.n10617 a_400_62400# 3.57fF
C11724 VN.t2074 a_400_62400# 0.03fF
C11725 VN.n10618 a_400_62400# 0.32fF
C11726 VN.n10619 a_400_62400# 0.48fF
C11727 VN.n10620 a_400_62400# 0.81fF
C11728 VN.n10621 a_400_62400# 0.16fF
C11729 VN.t903 a_400_62400# 0.03fF
C11730 VN.n10622 a_400_62400# 0.19fF
C11731 VN.n10624 a_400_62400# 0.93fF
C11732 VN.n10625 a_400_62400# 1.55fF
C11733 VN.n10626 a_400_62400# 0.29fF
C11734 VN.n10627 a_400_62400# 2.52fF
C11735 VN.t1352 a_400_62400# 0.03fF
C11736 VN.n10628 a_400_62400# 0.32fF
C11737 VN.n10629 a_400_62400# 1.22fF
C11738 VN.n10630 a_400_62400# 0.07fF
C11739 VN.t1109 a_400_62400# 0.03fF
C11740 VN.n10631 a_400_62400# 0.16fF
C11741 VN.n10632 a_400_62400# 0.19fF
C11742 VN.n10634 a_400_62400# 27.83fF
C11743 VN.n10635 a_400_62400# 3.65fF
C11744 VN.n10636 a_400_62400# 2.12fF
C11745 VN.n10637 a_400_62400# 0.16fF
C11746 VN.t1822 a_400_62400# 0.03fF
C11747 VN.n10638 a_400_62400# 0.19fF
C11748 VN.t336 a_400_62400# 0.03fF
C11749 VN.n10640 a_400_62400# 0.32fF
C11750 VN.n10641 a_400_62400# 0.48fF
C11751 VN.n10642 a_400_62400# 0.81fF
C11752 VN.n10643 a_400_62400# 3.17fF
C11753 VN.n10644 a_400_62400# 3.08fF
C11754 VN.t1890 a_400_62400# 0.03fF
C11755 VN.n10645 a_400_62400# 0.16fF
C11756 VN.n10646 a_400_62400# 0.19fF
C11757 VN.t2139 a_400_62400# 0.03fF
C11758 VN.n10648 a_400_62400# 0.32fF
C11759 VN.n10649 a_400_62400# 1.22fF
C11760 VN.n10650 a_400_62400# 0.07fF
C11761 VN.t241 a_400_62400# 64.69fF
C11762 VN.t242 a_400_62400# 0.03fF
C11763 VN.n10651 a_400_62400# 0.16fF
C11764 VN.n10652 a_400_62400# 0.19fF
C11765 VN.t484 a_400_62400# 0.03fF
C11766 VN.n10654 a_400_62400# 0.32fF
C11767 VN.n10655 a_400_62400# 1.22fF
C11768 VN.n10656 a_400_62400# 0.07fF
C11769 VN.t1202 a_400_62400# 0.03fF
C11770 VN.n10657 a_400_62400# 0.32fF
C11771 VN.n10658 a_400_62400# 0.48fF
C11772 VN.n10659 a_400_62400# 0.81fF
C11773 VN.n10660 a_400_62400# 2.07fF
C11774 VN.n10661 a_400_62400# 0.21fF
C11775 VN.n10662 a_400_62400# 6.66fF
C11776 VN.n10663 a_400_62400# 2.51fF
C11777 VN.n10664 a_400_62400# 0.16fF
C11778 VN.t1198 a_400_62400# 0.03fF
C11779 VN.n10665 a_400_62400# 0.19fF
C11780 VN.t2346 a_400_62400# 0.03fF
C11781 VN.n10667 a_400_62400# 0.32fF
C11782 VN.n10668 a_400_62400# 0.48fF
C11783 VN.n10669 a_400_62400# 0.81fF
C11784 VN.n10670 a_400_62400# 1.24fF
C11785 VN.n10671 a_400_62400# 0.43fF
C11786 VN.n10672 a_400_62400# 0.43fF
C11787 VN.n10673 a_400_62400# 1.24fF
C11788 VN.n10674 a_400_62400# 1.46fF
C11789 VN.n10675 a_400_62400# 0.21fF
C11790 VN.n10676 a_400_62400# 6.27fF
C11791 VN.t1860 a_400_62400# 0.03fF
C11792 VN.n10677 a_400_62400# 0.16fF
C11793 VN.n10678 a_400_62400# 0.19fF
C11794 VN.t1397 a_400_62400# 0.03fF
C11795 VN.n10680 a_400_62400# 0.32fF
C11796 VN.n10681 a_400_62400# 1.22fF
C11797 VN.n10682 a_400_62400# 0.07fF
C11798 VN.n10683 a_400_62400# 2.51fF
C11799 VN.n10684 a_400_62400# 3.58fF
C11800 VN.t1478 a_400_62400# 0.03fF
C11801 VN.n10685 a_400_62400# 0.32fF
C11802 VN.n10686 a_400_62400# 0.48fF
C11803 VN.n10687 a_400_62400# 0.81fF
C11804 VN.n10688 a_400_62400# 0.16fF
C11805 VN.t330 a_400_62400# 0.03fF
C11806 VN.n10689 a_400_62400# 0.19fF
C11807 VN.n10691 a_400_62400# 7.31fF
C11808 VN.t991 a_400_62400# 0.03fF
C11809 VN.n10692 a_400_62400# 0.16fF
C11810 VN.n10693 a_400_62400# 0.19fF
C11811 VN.t535 a_400_62400# 0.03fF
C11812 VN.n10695 a_400_62400# 0.32fF
C11813 VN.n10696 a_400_62400# 1.22fF
C11814 VN.n10697 a_400_62400# 0.07fF
C11815 VN.t120 a_400_62400# 64.17fF
C11816 VN.t2190 a_400_62400# 0.03fF
C11817 VN.n10698 a_400_62400# 1.60fF
C11818 VN.n10699 a_400_62400# 0.07fF
C11819 VN.t255 a_400_62400# 0.03fF
C11820 VN.n10700 a_400_62400# 0.02fF
C11821 VN.n10701 a_400_62400# 0.34fF
C11822 VN.n10703 a_400_62400# 2.01fF
C11823 VN.n10704 a_400_62400# 1.75fF
C11824 VN.n10705 a_400_62400# 0.37fF
C11825 VN.n10706 a_400_62400# 0.33fF
C11826 VN.n10707 a_400_62400# 5.88fF
C11827 VN.n10708 a_400_62400# 0.33fF
C11828 VN.n10709 a_400_62400# 0.79fF
C11829 VN.n10710 a_400_62400# 0.23fF
C11830 VN.n10711 a_400_62400# 1.18fF
C11831 VN.t78 a_400_62400# 28.64fF
C11832 VN.n10712 a_400_62400# 0.79fF
C11833 VN.n10713 a_400_62400# 0.11fF
C11834 VN.n10714 a_400_62400# 4.98fF
C11835 VN.n10715 a_400_62400# 0.80fF
C11836 VN.n10716 a_400_62400# 0.29fF
C11837 VN.n10717 a_400_62400# 1.96fF
C11838 VN.n10719 a_400_62400# 25.18fF
C11839 VN.n10721 a_400_62400# 1.87fF
C11840 VN.n10722 a_400_62400# 5.36fF
C11841 VN.n10723 a_400_62400# 2.01fF
C11842 VN.n10724 a_400_62400# 1.75fF
C11843 VN.n10725 a_400_62400# 0.37fF
C11844 VN.n10726 a_400_62400# 2.51fF
C11845 VN.n10727 a_400_62400# 0.33fF
C11846 VN.n10728 a_400_62400# 0.12fF
C11847 VN.n10729 a_400_62400# 0.28fF
C11848 VN.n10730 a_400_62400# 1.06fF
C11849 VN.n10731 a_400_62400# 0.59fF
C11850 VN.n10732 a_400_62400# 0.16fF
C11851 VN.t2487 a_400_62400# 0.03fF
C11852 VN.n10733 a_400_62400# 0.19fF
C11853 VN.t696 a_400_62400# 0.03fF
C11854 VN.n10735 a_400_62400# 0.32fF
C11855 VN.n10736 a_400_62400# 0.48fF
C11856 VN.n10737 a_400_62400# 0.81fF
C11857 VN.n10738 a_400_62400# 0.03fF
C11858 VN.n10739 a_400_62400# 0.01fF
C11859 VN.n10740 a_400_62400# 0.02fF
C11860 VN.n10741 a_400_62400# 0.11fF
C11861 VN.n10742 a_400_62400# 0.08fF
C11862 VN.n10743 a_400_62400# 0.04fF
C11863 VN.n10744 a_400_62400# 0.05fF
C11864 VN.n10745 a_400_62400# 1.34fF
C11865 VN.n10746 a_400_62400# 0.48fF
C11866 VN.n10747 a_400_62400# 2.48fF
C11867 VN.n10748 a_400_62400# 2.66fF
C11868 VN.t1806 a_400_62400# 0.03fF
C11869 VN.n10749 a_400_62400# 0.32fF
C11870 VN.n10750 a_400_62400# 1.22fF
C11871 VN.n10751 a_400_62400# 0.07fF
C11872 VN.t645 a_400_62400# 0.03fF
C11873 VN.n10752 a_400_62400# 0.16fF
C11874 VN.n10753 a_400_62400# 0.19fF
C11875 VN.n10755 a_400_62400# 2.53fF
C11876 VN.n10756 a_400_62400# 0.08fF
C11877 VN.n10757 a_400_62400# 0.04fF
C11878 VN.n10758 a_400_62400# 0.05fF
C11879 VN.n10759 a_400_62400# 1.33fF
C11880 VN.n10760 a_400_62400# 0.03fF
C11881 VN.n10761 a_400_62400# 0.01fF
C11882 VN.n10762 a_400_62400# 0.02fF
C11883 VN.n10763 a_400_62400# 0.11fF
C11884 VN.n10764 a_400_62400# 0.48fF
C11885 VN.n10765 a_400_62400# 2.48fF
C11886 VN.t2472 a_400_62400# 0.03fF
C11887 VN.n10766 a_400_62400# 0.32fF
C11888 VN.n10767 a_400_62400# 0.48fF
C11889 VN.n10768 a_400_62400# 0.81fF
C11890 VN.n10769 a_400_62400# 0.16fF
C11891 VN.t1623 a_400_62400# 0.03fF
C11892 VN.n10770 a_400_62400# 0.19fF
C11893 VN.n10772 a_400_62400# 0.29fF
C11894 VN.n10773 a_400_62400# 1.27fF
C11895 VN.n10774 a_400_62400# 0.79fF
C11896 VN.n10775 a_400_62400# 0.34fF
C11897 VN.n10776 a_400_62400# 0.12fF
C11898 VN.n10777 a_400_62400# 2.52fF
C11899 VN.t1066 a_400_62400# 0.03fF
C11900 VN.n10778 a_400_62400# 0.32fF
C11901 VN.n10779 a_400_62400# 1.22fF
C11902 VN.n10780 a_400_62400# 0.07fF
C11903 VN.t2303 a_400_62400# 0.03fF
C11904 VN.n10781 a_400_62400# 0.16fF
C11905 VN.n10782 a_400_62400# 0.19fF
C11906 VN.n10784 a_400_62400# 2.51fF
C11907 VN.n10785 a_400_62400# 0.33fF
C11908 VN.n10786 a_400_62400# 0.12fF
C11909 VN.n10787 a_400_62400# 0.28fF
C11910 VN.n10788 a_400_62400# 1.06fF
C11911 VN.n10789 a_400_62400# 0.59fF
C11912 VN.n10790 a_400_62400# 0.16fF
C11913 VN.t751 a_400_62400# 0.03fF
C11914 VN.n10791 a_400_62400# 0.19fF
C11915 VN.t1610 a_400_62400# 0.03fF
C11916 VN.n10793 a_400_62400# 0.32fF
C11917 VN.n10794 a_400_62400# 0.48fF
C11918 VN.n10795 a_400_62400# 0.81fF
C11919 VN.n10796 a_400_62400# 0.03fF
C11920 VN.n10797 a_400_62400# 0.01fF
C11921 VN.n10798 a_400_62400# 0.02fF
C11922 VN.n10799 a_400_62400# 0.11fF
C11923 VN.n10800 a_400_62400# 0.08fF
C11924 VN.n10801 a_400_62400# 0.04fF
C11925 VN.n10802 a_400_62400# 0.05fF
C11926 VN.n10803 a_400_62400# 1.34fF
C11927 VN.n10804 a_400_62400# 0.48fF
C11928 VN.n10805 a_400_62400# 2.48fF
C11929 VN.n10806 a_400_62400# 2.66fF
C11930 VN.t192 a_400_62400# 0.03fF
C11931 VN.n10807 a_400_62400# 0.32fF
C11932 VN.n10808 a_400_62400# 1.22fF
C11933 VN.n10809 a_400_62400# 0.07fF
C11934 VN.t1430 a_400_62400# 0.03fF
C11935 VN.n10810 a_400_62400# 0.16fF
C11936 VN.n10811 a_400_62400# 0.19fF
C11937 VN.n10813 a_400_62400# 2.53fF
C11938 VN.n10814 a_400_62400# 0.08fF
C11939 VN.n10815 a_400_62400# 0.04fF
C11940 VN.n10816 a_400_62400# 0.05fF
C11941 VN.n10817 a_400_62400# 1.33fF
C11942 VN.n10818 a_400_62400# 0.03fF
C11943 VN.n10819 a_400_62400# 0.01fF
C11944 VN.n10820 a_400_62400# 0.02fF
C11945 VN.n10821 a_400_62400# 0.11fF
C11946 VN.n10822 a_400_62400# 0.48fF
C11947 VN.n10823 a_400_62400# 2.48fF
C11948 VN.t2101 a_400_62400# 0.03fF
C11949 VN.n10824 a_400_62400# 0.32fF
C11950 VN.n10825 a_400_62400# 0.48fF
C11951 VN.n10826 a_400_62400# 0.81fF
C11952 VN.n10827 a_400_62400# 0.16fF
C11953 VN.t1238 a_400_62400# 0.03fF
C11954 VN.n10828 a_400_62400# 0.19fF
C11955 VN.n10830 a_400_62400# 0.29fF
C11956 VN.n10831 a_400_62400# 1.27fF
C11957 VN.n10832 a_400_62400# 0.79fF
C11958 VN.n10833 a_400_62400# 0.34fF
C11959 VN.n10834 a_400_62400# 0.12fF
C11960 VN.n10835 a_400_62400# 2.52fF
C11961 VN.t682 a_400_62400# 0.03fF
C11962 VN.n10836 a_400_62400# 0.32fF
C11963 VN.n10837 a_400_62400# 1.22fF
C11964 VN.n10838 a_400_62400# 0.07fF
C11965 VN.t564 a_400_62400# 0.03fF
C11966 VN.n10839 a_400_62400# 0.16fF
C11967 VN.n10840 a_400_62400# 0.19fF
C11968 VN.n10842 a_400_62400# 0.33fF
C11969 VN.n10843 a_400_62400# 0.12fF
C11970 VN.n10844 a_400_62400# 0.28fF
C11971 VN.n10845 a_400_62400# 1.72fF
C11972 VN.n10846 a_400_62400# 0.71fF
C11973 VN.n10847 a_400_62400# 2.51fF
C11974 VN.n10848 a_400_62400# 0.16fF
C11975 VN.t373 a_400_62400# 0.03fF
C11976 VN.n10849 a_400_62400# 0.19fF
C11977 VN.t1224 a_400_62400# 0.03fF
C11978 VN.n10851 a_400_62400# 0.32fF
C11979 VN.n10852 a_400_62400# 0.48fF
C11980 VN.n10853 a_400_62400# 0.81fF
C11981 VN.n10854 a_400_62400# 0.03fF
C11982 VN.n10855 a_400_62400# 0.01fF
C11983 VN.n10856 a_400_62400# 0.02fF
C11984 VN.n10857 a_400_62400# 0.11fF
C11985 VN.n10858 a_400_62400# 0.08fF
C11986 VN.n10859 a_400_62400# 0.04fF
C11987 VN.n10860 a_400_62400# 0.05fF
C11988 VN.n10861 a_400_62400# 1.34fF
C11989 VN.n10862 a_400_62400# 0.48fF
C11990 VN.n10863 a_400_62400# 2.51fF
C11991 VN.n10864 a_400_62400# 2.67fF
C11992 VN.t2342 a_400_62400# 0.03fF
C11993 VN.n10865 a_400_62400# 0.32fF
C11994 VN.n10866 a_400_62400# 1.22fF
C11995 VN.n10867 a_400_62400# 0.07fF
C11996 VN.t1026 a_400_62400# 0.03fF
C11997 VN.n10868 a_400_62400# 0.16fF
C11998 VN.n10869 a_400_62400# 0.19fF
C11999 VN.n10871 a_400_62400# 2.53fF
C12000 VN.n10872 a_400_62400# 0.08fF
C12001 VN.n10873 a_400_62400# 0.04fF
C12002 VN.n10874 a_400_62400# 0.05fF
C12003 VN.n10875 a_400_62400# 1.33fF
C12004 VN.n10876 a_400_62400# 0.03fF
C12005 VN.n10877 a_400_62400# 0.01fF
C12006 VN.n10878 a_400_62400# 0.02fF
C12007 VN.n10879 a_400_62400# 0.11fF
C12008 VN.n10880 a_400_62400# 0.48fF
C12009 VN.n10881 a_400_62400# 2.48fF
C12010 VN.t359 a_400_62400# 0.03fF
C12011 VN.n10882 a_400_62400# 0.32fF
C12012 VN.n10883 a_400_62400# 0.48fF
C12013 VN.n10884 a_400_62400# 0.81fF
C12014 VN.n10885 a_400_62400# 0.16fF
C12015 VN.t2026 a_400_62400# 0.03fF
C12016 VN.n10886 a_400_62400# 0.19fF
C12017 VN.n10888 a_400_62400# 0.29fF
C12018 VN.n10889 a_400_62400# 1.27fF
C12019 VN.n10890 a_400_62400# 0.79fF
C12020 VN.n10891 a_400_62400# 0.34fF
C12021 VN.n10892 a_400_62400# 0.12fF
C12022 VN.n10893 a_400_62400# 2.52fF
C12023 VN.t1474 a_400_62400# 0.03fF
C12024 VN.n10894 a_400_62400# 0.32fF
C12025 VN.n10895 a_400_62400# 1.22fF
C12026 VN.n10896 a_400_62400# 0.07fF
C12027 VN.t153 a_400_62400# 0.03fF
C12028 VN.n10897 a_400_62400# 0.16fF
C12029 VN.n10898 a_400_62400# 0.19fF
C12030 VN.n10900 a_400_62400# 2.51fF
C12031 VN.n10901 a_400_62400# 0.33fF
C12032 VN.n10902 a_400_62400# 0.12fF
C12033 VN.n10903 a_400_62400# 0.28fF
C12034 VN.n10904 a_400_62400# 1.06fF
C12035 VN.n10905 a_400_62400# 0.59fF
C12036 VN.n10906 a_400_62400# 0.16fF
C12037 VN.t1151 a_400_62400# 0.03fF
C12038 VN.n10907 a_400_62400# 0.19fF
C12039 VN.t2008 a_400_62400# 0.03fF
C12040 VN.n10909 a_400_62400# 0.32fF
C12041 VN.n10910 a_400_62400# 0.48fF
C12042 VN.n10911 a_400_62400# 0.81fF
C12043 VN.n10912 a_400_62400# 0.03fF
C12044 VN.n10913 a_400_62400# 0.01fF
C12045 VN.n10914 a_400_62400# 0.02fF
C12046 VN.n10915 a_400_62400# 0.11fF
C12047 VN.n10916 a_400_62400# 0.08fF
C12048 VN.n10917 a_400_62400# 0.04fF
C12049 VN.n10918 a_400_62400# 0.05fF
C12050 VN.n10919 a_400_62400# 1.34fF
C12051 VN.n10920 a_400_62400# 0.48fF
C12052 VN.n10921 a_400_62400# 2.48fF
C12053 VN.n10922 a_400_62400# 2.66fF
C12054 VN.t607 a_400_62400# 0.03fF
C12055 VN.n10923 a_400_62400# 0.32fF
C12056 VN.n10924 a_400_62400# 1.22fF
C12057 VN.n10925 a_400_62400# 0.07fF
C12058 VN.t1952 a_400_62400# 0.03fF
C12059 VN.n10926 a_400_62400# 0.16fF
C12060 VN.n10927 a_400_62400# 0.19fF
C12061 VN.n10929 a_400_62400# 2.53fF
C12062 VN.n10930 a_400_62400# 0.08fF
C12063 VN.n10931 a_400_62400# 0.04fF
C12064 VN.n10932 a_400_62400# 0.05fF
C12065 VN.n10933 a_400_62400# 1.33fF
C12066 VN.n10934 a_400_62400# 0.03fF
C12067 VN.n10935 a_400_62400# 0.01fF
C12068 VN.n10936 a_400_62400# 0.02fF
C12069 VN.n10937 a_400_62400# 0.11fF
C12070 VN.n10938 a_400_62400# 0.48fF
C12071 VN.n10939 a_400_62400# 2.48fF
C12072 VN.t1135 a_400_62400# 0.03fF
C12073 VN.n10940 a_400_62400# 0.32fF
C12074 VN.n10941 a_400_62400# 0.48fF
C12075 VN.n10942 a_400_62400# 0.81fF
C12076 VN.n10943 a_400_62400# 0.16fF
C12077 VN.t284 a_400_62400# 0.03fF
C12078 VN.n10944 a_400_62400# 0.19fF
C12079 VN.n10946 a_400_62400# 0.29fF
C12080 VN.n10947 a_400_62400# 1.27fF
C12081 VN.n10948 a_400_62400# 0.79fF
C12082 VN.n10949 a_400_62400# 0.34fF
C12083 VN.n10950 a_400_62400# 0.12fF
C12084 VN.n10951 a_400_62400# 2.52fF
C12085 VN.t2260 a_400_62400# 0.03fF
C12086 VN.n10952 a_400_62400# 0.32fF
C12087 VN.n10953 a_400_62400# 1.22fF
C12088 VN.n10954 a_400_62400# 0.07fF
C12089 VN.t1083 a_400_62400# 0.03fF
C12090 VN.n10955 a_400_62400# 0.16fF
C12091 VN.n10956 a_400_62400# 0.19fF
C12092 VN.n10958 a_400_62400# 2.51fF
C12093 VN.n10959 a_400_62400# 0.33fF
C12094 VN.n10960 a_400_62400# 0.12fF
C12095 VN.n10961 a_400_62400# 0.28fF
C12096 VN.n10962 a_400_62400# 1.06fF
C12097 VN.n10963 a_400_62400# 0.59fF
C12098 VN.n10964 a_400_62400# 0.16fF
C12099 VN.t1935 a_400_62400# 0.03fF
C12100 VN.n10965 a_400_62400# 0.19fF
C12101 VN.t272 a_400_62400# 0.03fF
C12102 VN.n10967 a_400_62400# 0.32fF
C12103 VN.n10968 a_400_62400# 0.48fF
C12104 VN.n10969 a_400_62400# 0.81fF
C12105 VN.n10970 a_400_62400# 0.03fF
C12106 VN.n10971 a_400_62400# 0.01fF
C12107 VN.n10972 a_400_62400# 0.02fF
C12108 VN.n10973 a_400_62400# 0.11fF
C12109 VN.n10974 a_400_62400# 0.08fF
C12110 VN.n10975 a_400_62400# 0.04fF
C12111 VN.n10976 a_400_62400# 0.05fF
C12112 VN.n10977 a_400_62400# 1.34fF
C12113 VN.n10978 a_400_62400# 0.48fF
C12114 VN.n10979 a_400_62400# 2.48fF
C12115 VN.n10980 a_400_62400# 2.66fF
C12116 VN.t1395 a_400_62400# 0.03fF
C12117 VN.n10981 a_400_62400# 0.32fF
C12118 VN.n10982 a_400_62400# 1.22fF
C12119 VN.n10983 a_400_62400# 0.07fF
C12120 VN.t209 a_400_62400# 0.03fF
C12121 VN.n10984 a_400_62400# 0.16fF
C12122 VN.n10985 a_400_62400# 0.19fF
C12123 VN.n10987 a_400_62400# 2.53fF
C12124 VN.n10988 a_400_62400# 0.08fF
C12125 VN.n10989 a_400_62400# 0.04fF
C12126 VN.n10990 a_400_62400# 0.05fF
C12127 VN.n10991 a_400_62400# 1.33fF
C12128 VN.n10992 a_400_62400# 0.03fF
C12129 VN.n10993 a_400_62400# 0.01fF
C12130 VN.n10994 a_400_62400# 0.02fF
C12131 VN.n10995 a_400_62400# 0.11fF
C12132 VN.n10996 a_400_62400# 0.48fF
C12133 VN.n10997 a_400_62400# 2.48fF
C12134 VN.t1922 a_400_62400# 0.03fF
C12135 VN.n10998 a_400_62400# 0.32fF
C12136 VN.n10999 a_400_62400# 0.48fF
C12137 VN.n11000 a_400_62400# 0.81fF
C12138 VN.n11001 a_400_62400# 0.16fF
C12139 VN.t1062 a_400_62400# 0.03fF
C12140 VN.n11002 a_400_62400# 0.19fF
C12141 VN.n11004 a_400_62400# 0.29fF
C12142 VN.n11005 a_400_62400# 1.27fF
C12143 VN.n11006 a_400_62400# 0.79fF
C12144 VN.n11007 a_400_62400# 0.34fF
C12145 VN.n11008 a_400_62400# 0.12fF
C12146 VN.n11009 a_400_62400# 2.52fF
C12147 VN.t533 a_400_62400# 0.03fF
C12148 VN.n11010 a_400_62400# 0.32fF
C12149 VN.n11011 a_400_62400# 1.22fF
C12150 VN.n11012 a_400_62400# 0.07fF
C12151 VN.t1862 a_400_62400# 0.03fF
C12152 VN.n11013 a_400_62400# 0.16fF
C12153 VN.n11014 a_400_62400# 0.19fF
C12154 VN.n11016 a_400_62400# 2.51fF
C12155 VN.n11017 a_400_62400# 0.33fF
C12156 VN.n11018 a_400_62400# 0.12fF
C12157 VN.n11019 a_400_62400# 0.28fF
C12158 VN.n11020 a_400_62400# 1.06fF
C12159 VN.n11021 a_400_62400# 0.59fF
C12160 VN.n11022 a_400_62400# 0.16fF
C12161 VN.t334 a_400_62400# 0.03fF
C12162 VN.n11023 a_400_62400# 0.19fF
C12163 VN.t1047 a_400_62400# 0.03fF
C12164 VN.n11025 a_400_62400# 0.32fF
C12165 VN.n11026 a_400_62400# 0.48fF
C12166 VN.n11027 a_400_62400# 0.81fF
C12167 VN.n11028 a_400_62400# 0.03fF
C12168 VN.n11029 a_400_62400# 0.01fF
C12169 VN.n11030 a_400_62400# 0.02fF
C12170 VN.n11031 a_400_62400# 0.11fF
C12171 VN.n11032 a_400_62400# 0.05fF
C12172 VN.n11033 a_400_62400# 1.36fF
C12173 VN.n11034 a_400_62400# 0.48fF
C12174 VN.n11035 a_400_62400# 2.48fF
C12175 VN.n11036 a_400_62400# 2.66fF
C12176 VN.t2187 a_400_62400# 0.03fF
C12177 VN.n11037 a_400_62400# 0.32fF
C12178 VN.n11038 a_400_62400# 1.22fF
C12179 VN.n11039 a_400_62400# 0.07fF
C12180 VN.t992 a_400_62400# 0.03fF
C12181 VN.n11040 a_400_62400# 0.16fF
C12182 VN.n11041 a_400_62400# 0.19fF
C12183 VN.n11043 a_400_62400# 0.34fF
C12184 VN.n11044 a_400_62400# 0.12fF
C12185 VN.n11045 a_400_62400# 0.30fF
C12186 VN.n11046 a_400_62400# 1.27fF
C12187 VN.n11047 a_400_62400# 0.79fF
C12188 VN.n11048 a_400_62400# 2.53fF
C12189 VN.n11049 a_400_62400# 0.16fF
C12190 VN.t1979 a_400_62400# 0.03fF
C12191 VN.n11050 a_400_62400# 0.19fF
C12192 VN.t315 a_400_62400# 0.03fF
C12193 VN.n11052 a_400_62400# 0.32fF
C12194 VN.n11053 a_400_62400# 0.48fF
C12195 VN.n11054 a_400_62400# 0.81fF
C12196 VN.n11055 a_400_62400# 0.24fF
C12197 VN.n11056 a_400_62400# 0.29fF
C12198 VN.n11057 a_400_62400# 0.63fF
C12199 VN.n11058 a_400_62400# 0.44fF
C12200 VN.n11059 a_400_62400# 0.01fF
C12201 VN.n11060 a_400_62400# 0.01fF
C12202 VN.n11061 a_400_62400# 0.01fF
C12203 VN.n11062 a_400_62400# 0.09fF
C12204 VN.n11063 a_400_62400# 0.05fF
C12205 VN.n11064 a_400_62400# 0.09fF
C12206 VN.n11065 a_400_62400# 0.07fF
C12207 VN.n11066 a_400_62400# 0.55fF
C12208 VN.n11067 a_400_62400# 0.77fF
C12209 VN.n11068 a_400_62400# 0.25fF
C12210 VN.n11069 a_400_62400# 2.64fF
C12211 VN.t1436 a_400_62400# 0.03fF
C12212 VN.n11070 a_400_62400# 0.32fF
C12213 VN.n11071 a_400_62400# 1.22fF
C12214 VN.n11072 a_400_62400# 0.07fF
C12215 VN.t107 a_400_62400# 0.03fF
C12216 VN.n11073 a_400_62400# 0.16fF
C12217 VN.n11074 a_400_62400# 0.19fF
C12218 VN.n11076 a_400_62400# 0.06fF
C12219 VN.n11077 a_400_62400# 0.04fF
C12220 VN.n11078 a_400_62400# 0.04fF
C12221 VN.n11079 a_400_62400# 0.14fF
C12222 VN.n11080 a_400_62400# 0.48fF
C12223 VN.n11081 a_400_62400# 0.50fF
C12224 VN.n11082 a_400_62400# 0.14fF
C12225 VN.n11083 a_400_62400# 0.16fF
C12226 VN.n11084 a_400_62400# 0.09fF
C12227 VN.n11085 a_400_62400# 0.16fF
C12228 VN.n11086 a_400_62400# 0.24fF
C12229 VN.n11087 a_400_62400# 2.51fF
C12230 VN.n11088 a_400_62400# 0.16fF
C12231 VN.t59 a_400_62400# 0.03fF
C12232 VN.n11089 a_400_62400# 0.19fF
C12233 VN.n11091 a_400_62400# 2.62fF
C12234 VN.n11092 a_400_62400# 0.16fF
C12235 VN.t135 a_400_62400# 0.03fF
C12236 VN.n11093 a_400_62400# 0.19fF
C12237 VN.t1178 a_400_62400# 0.03fF
C12238 VN.n11095 a_400_62400# 0.32fF
C12239 VN.n11096 a_400_62400# 0.48fF
C12240 VN.n11097 a_400_62400# 0.81fF
C12241 VN.n11098 a_400_62400# 2.09fF
C12242 VN.n11099 a_400_62400# 0.37fF
C12243 VN.n11100 a_400_62400# 2.82fF
C12244 VN.t2127 a_400_62400# 0.03fF
C12245 VN.n11101 a_400_62400# 0.32fF
C12246 VN.n11102 a_400_62400# 1.22fF
C12247 VN.n11103 a_400_62400# 0.07fF
C12248 VN.t214 a_400_62400# 0.03fF
C12249 VN.n11104 a_400_62400# 0.16fF
C12250 VN.n11105 a_400_62400# 0.19fF
C12251 VN.n11107 a_400_62400# 27.83fF
C12252 VN.n11108 a_400_62400# 2.53fF
C12253 VN.n11109 a_400_62400# 3.68fF
C12254 VN.t2046 a_400_62400# 0.03fF
C12255 VN.n11110 a_400_62400# 0.32fF
C12256 VN.n11111 a_400_62400# 0.48fF
C12257 VN.n11112 a_400_62400# 0.81fF
C12258 VN.n11113 a_400_62400# 0.16fF
C12259 VN.t877 a_400_62400# 0.03fF
C12260 VN.n11114 a_400_62400# 0.19fF
C12261 VN.n11116 a_400_62400# 1.55fF
C12262 VN.n11117 a_400_62400# 0.29fF
C12263 VN.n11118 a_400_62400# 2.52fF
C12264 VN.t1087 a_400_62400# 0.03fF
C12265 VN.n11119 a_400_62400# 0.16fF
C12266 VN.n11120 a_400_62400# 0.19fF
C12267 VN.t473 a_400_62400# 0.03fF
C12268 VN.n11122 a_400_62400# 0.32fF
C12269 VN.n11123 a_400_62400# 1.22fF
C12270 VN.n11124 a_400_62400# 0.07fF
C12271 VN.n11125 a_400_62400# 1.05fF
C12272 VN.n11126 a_400_62400# 3.07fF
C12273 VN.n11127 a_400_62400# 2.51fF
C12274 VN.n11128 a_400_62400# 0.16fF
C12275 VN.t1751 a_400_62400# 0.03fF
C12276 VN.n11129 a_400_62400# 0.19fF
C12277 VN.t396 a_400_62400# 0.03fF
C12278 VN.n11131 a_400_62400# 0.32fF
C12279 VN.n11132 a_400_62400# 0.48fF
C12280 VN.n11133 a_400_62400# 0.81fF
C12281 VN.n11134 a_400_62400# 1.03fF
C12282 VN.n11135 a_400_62400# 0.65fF
C12283 VN.n11136 a_400_62400# 0.12fF
C12284 VN.n11137 a_400_62400# 0.44fF
C12285 VN.n11138 a_400_62400# 2.71fF
C12286 VN.t1955 a_400_62400# 0.03fF
C12287 VN.n11139 a_400_62400# 0.16fF
C12288 VN.n11140 a_400_62400# 0.19fF
C12289 VN.t1337 a_400_62400# 0.03fF
C12290 VN.n11142 a_400_62400# 0.32fF
C12291 VN.n11143 a_400_62400# 1.22fF
C12292 VN.n11144 a_400_62400# 0.07fF
C12293 VN.n11145 a_400_62400# 3.55fF
C12294 VN.n11146 a_400_62400# 2.53fF
C12295 VN.n11147 a_400_62400# 0.16fF
C12296 VN.t36 a_400_62400# 0.03fF
C12297 VN.n11148 a_400_62400# 0.19fF
C12298 VN.t1244 a_400_62400# 0.03fF
C12299 VN.n11150 a_400_62400# 0.32fF
C12300 VN.n11151 a_400_62400# 0.48fF
C12301 VN.n11152 a_400_62400# 0.81fF
C12302 VN.n11153 a_400_62400# 3.00fF
C12303 VN.n11154 a_400_62400# 3.61fF
C12304 VN.t297 a_400_62400# 0.03fF
C12305 VN.n11155 a_400_62400# 0.16fF
C12306 VN.n11156 a_400_62400# 0.19fF
C12307 VN.t690 a_400_62400# 0.03fF
C12308 VN.n11158 a_400_62400# 0.32fF
C12309 VN.n11159 a_400_62400# 1.22fF
C12310 VN.n11160 a_400_62400# 0.07fF
C12311 VN.n11161 a_400_62400# 1.03fF
C12312 VN.n11162 a_400_62400# 1.66fF
C12313 VN.n11163 a_400_62400# 1.71fF
C12314 VN.n11164 a_400_62400# 2.51fF
C12315 VN.n11165 a_400_62400# 0.16fF
C12316 VN.t953 a_400_62400# 0.03fF
C12317 VN.n11166 a_400_62400# 0.19fF
C12318 VN.t2120 a_400_62400# 0.03fF
C12319 VN.n11168 a_400_62400# 0.32fF
C12320 VN.n11169 a_400_62400# 0.48fF
C12321 VN.n11170 a_400_62400# 0.81fF
C12322 VN.n11171 a_400_62400# 3.68fF
C12323 VN.n11172 a_400_62400# 2.90fF
C12324 VN.t1166 a_400_62400# 0.03fF
C12325 VN.n11173 a_400_62400# 0.16fF
C12326 VN.n11174 a_400_62400# 0.19fF
C12327 VN.t1560 a_400_62400# 0.03fF
C12328 VN.n11176 a_400_62400# 0.32fF
C12329 VN.n11177 a_400_62400# 1.22fF
C12330 VN.n11178 a_400_62400# 0.07fF
C12331 VN.n11179 a_400_62400# 3.68fF
C12332 VN.t469 a_400_62400# 0.03fF
C12333 VN.n11180 a_400_62400# 0.32fF
C12334 VN.n11181 a_400_62400# 0.48fF
C12335 VN.n11182 a_400_62400# 0.81fF
C12336 VN.n11183 a_400_62400# 0.16fF
C12337 VN.t1830 a_400_62400# 0.03fF
C12338 VN.n11184 a_400_62400# 0.19fF
C12339 VN.n11186 a_400_62400# 2.42fF
C12340 VN.n11187 a_400_62400# 2.53fF
C12341 VN.n11188 a_400_62400# 2.75fF
C12342 VN.t1894 a_400_62400# 0.03fF
C12343 VN.n11189 a_400_62400# 0.16fF
C12344 VN.n11190 a_400_62400# 0.19fF
C12345 VN.t2422 a_400_62400# 0.03fF
C12346 VN.n11192 a_400_62400# 0.32fF
C12347 VN.n11193 a_400_62400# 1.22fF
C12348 VN.n11194 a_400_62400# 0.07fF
C12349 VN.n11195 a_400_62400# 1.03fF
C12350 VN.n11196 a_400_62400# 1.66fF
C12351 VN.n11197 a_400_62400# 1.71fF
C12352 VN.n11198 a_400_62400# 2.51fF
C12353 VN.n11199 a_400_62400# 0.16fF
C12354 VN.t169 a_400_62400# 0.03fF
C12355 VN.n11200 a_400_62400# 0.19fF
C12356 VN.t1331 a_400_62400# 0.03fF
C12357 VN.n11202 a_400_62400# 0.32fF
C12358 VN.n11203 a_400_62400# 0.48fF
C12359 VN.n11204 a_400_62400# 0.81fF
C12360 VN.n11205 a_400_62400# 3.68fF
C12361 VN.n11206 a_400_62400# 2.90fF
C12362 VN.t247 a_400_62400# 0.03fF
C12363 VN.n11207 a_400_62400# 0.16fF
C12364 VN.n11208 a_400_62400# 0.19fF
C12365 VN.t771 a_400_62400# 0.03fF
C12366 VN.n11210 a_400_62400# 0.32fF
C12367 VN.n11211 a_400_62400# 1.22fF
C12368 VN.n11212 a_400_62400# 0.07fF
C12369 VN.n11213 a_400_62400# 3.68fF
C12370 VN.t2200 a_400_62400# 0.03fF
C12371 VN.n11214 a_400_62400# 0.32fF
C12372 VN.n11215 a_400_62400# 0.48fF
C12373 VN.n11216 a_400_62400# 0.81fF
C12374 VN.n11217 a_400_62400# 0.16fF
C12375 VN.t1041 a_400_62400# 0.03fF
C12376 VN.n11218 a_400_62400# 0.19fF
C12377 VN.n11220 a_400_62400# 2.42fF
C12378 VN.n11221 a_400_62400# 2.53fF
C12379 VN.n11222 a_400_62400# 2.75fF
C12380 VN.t1111 a_400_62400# 0.03fF
C12381 VN.n11223 a_400_62400# 0.16fF
C12382 VN.n11224 a_400_62400# 0.19fF
C12383 VN.t1642 a_400_62400# 0.03fF
C12384 VN.n11226 a_400_62400# 0.32fF
C12385 VN.n11227 a_400_62400# 1.22fF
C12386 VN.n11228 a_400_62400# 0.07fF
C12387 VN.n11229 a_400_62400# 1.03fF
C12388 VN.n11230 a_400_62400# 1.66fF
C12389 VN.n11231 a_400_62400# 1.71fF
C12390 VN.n11232 a_400_62400# 2.51fF
C12391 VN.n11233 a_400_62400# 0.16fF
C12392 VN.t1916 a_400_62400# 0.03fF
C12393 VN.n11234 a_400_62400# 0.19fF
C12394 VN.t544 a_400_62400# 0.03fF
C12395 VN.n11236 a_400_62400# 0.32fF
C12396 VN.n11237 a_400_62400# 0.48fF
C12397 VN.n11238 a_400_62400# 0.81fF
C12398 VN.n11239 a_400_62400# 3.68fF
C12399 VN.n11240 a_400_62400# 2.90fF
C12400 VN.t1985 a_400_62400# 0.03fF
C12401 VN.n11241 a_400_62400# 0.16fF
C12402 VN.n11242 a_400_62400# 0.19fF
C12403 VN.t2505 a_400_62400# 0.03fF
C12404 VN.n11244 a_400_62400# 0.32fF
C12405 VN.n11245 a_400_62400# 1.22fF
C12406 VN.n11246 a_400_62400# 0.07fF
C12407 VN.n11247 a_400_62400# 3.68fF
C12408 VN.t1289 a_400_62400# 0.03fF
C12409 VN.n11248 a_400_62400# 0.32fF
C12410 VN.n11249 a_400_62400# 0.48fF
C12411 VN.n11250 a_400_62400# 0.81fF
C12412 VN.n11251 a_400_62400# 0.16fF
C12413 VN.t265 a_400_62400# 0.03fF
C12414 VN.n11252 a_400_62400# 0.19fF
C12415 VN.n11254 a_400_62400# 2.42fF
C12416 VN.n11255 a_400_62400# 2.53fF
C12417 VN.n11256 a_400_62400# 2.75fF
C12418 VN.t341 a_400_62400# 0.03fF
C12419 VN.n11257 a_400_62400# 0.16fF
C12420 VN.n11258 a_400_62400# 0.19fF
C12421 VN.t729 a_400_62400# 0.03fF
C12422 VN.n11260 a_400_62400# 0.32fF
C12423 VN.n11261 a_400_62400# 1.22fF
C12424 VN.n11262 a_400_62400# 0.07fF
C12425 VN.n11263 a_400_62400# 1.03fF
C12426 VN.n11264 a_400_62400# 3.07fF
C12427 VN.n11265 a_400_62400# 2.51fF
C12428 VN.n11266 a_400_62400# 0.16fF
C12429 VN.t996 a_400_62400# 0.03fF
C12430 VN.n11267 a_400_62400# 0.19fF
C12431 VN.t2158 a_400_62400# 0.03fF
C12432 VN.n11269 a_400_62400# 0.32fF
C12433 VN.n11270 a_400_62400# 0.48fF
C12434 VN.n11271 a_400_62400# 0.81fF
C12435 VN.n11272 a_400_62400# 3.30fF
C12436 VN.n11273 a_400_62400# 2.91fF
C12437 VN.t1205 a_400_62400# 0.03fF
C12438 VN.n11274 a_400_62400# 0.16fF
C12439 VN.n11275 a_400_62400# 0.19fF
C12440 VN.t1594 a_400_62400# 0.03fF
C12441 VN.n11277 a_400_62400# 0.32fF
C12442 VN.n11278 a_400_62400# 1.22fF
C12443 VN.n11279 a_400_62400# 0.07fF
C12444 VN.n11280 a_400_62400# 2.53fF
C12445 VN.n11281 a_400_62400# 3.68fF
C12446 VN.t503 a_400_62400# 0.03fF
C12447 VN.n11282 a_400_62400# 0.32fF
C12448 VN.n11283 a_400_62400# 0.48fF
C12449 VN.n11284 a_400_62400# 0.81fF
C12450 VN.n11285 a_400_62400# 0.16fF
C12451 VN.t1866 a_400_62400# 0.03fF
C12452 VN.n11286 a_400_62400# 0.19fF
C12453 VN.n11288 a_400_62400# 2.97fF
C12454 VN.n11289 a_400_62400# 2.75fF
C12455 VN.t2077 a_400_62400# 0.03fF
C12456 VN.n11290 a_400_62400# 0.16fF
C12457 VN.n11291 a_400_62400# 0.19fF
C12458 VN.t2459 a_400_62400# 0.03fF
C12459 VN.n11293 a_400_62400# 0.32fF
C12460 VN.n11294 a_400_62400# 1.22fF
C12461 VN.n11295 a_400_62400# 0.07fF
C12462 VN.n11296 a_400_62400# 1.03fF
C12463 VN.n11297 a_400_62400# 1.66fF
C12464 VN.n11298 a_400_62400# 1.71fF
C12465 VN.n11299 a_400_62400# 2.51fF
C12466 VN.n11300 a_400_62400# 0.16fF
C12467 VN.t1399 a_400_62400# 0.03fF
C12468 VN.n11301 a_400_62400# 0.19fF
C12469 VN.t2523 a_400_62400# 0.03fF
C12470 VN.n11303 a_400_62400# 0.32fF
C12471 VN.n11304 a_400_62400# 0.48fF
C12472 VN.n11305 a_400_62400# 0.81fF
C12473 VN.n11306 a_400_62400# 3.68fF
C12474 VN.n11307 a_400_62400# 2.90fF
C12475 VN.t1589 a_400_62400# 0.03fF
C12476 VN.n11308 a_400_62400# 0.16fF
C12477 VN.n11309 a_400_62400# 0.19fF
C12478 VN.t1980 a_400_62400# 0.03fF
C12479 VN.n11311 a_400_62400# 0.32fF
C12480 VN.n11312 a_400_62400# 1.22fF
C12481 VN.n11313 a_400_62400# 0.07fF
C12482 VN.n11314 a_400_62400# 3.68fF
C12483 VN.t861 a_400_62400# 0.03fF
C12484 VN.n11315 a_400_62400# 0.32fF
C12485 VN.n11316 a_400_62400# 0.48fF
C12486 VN.n11317 a_400_62400# 0.81fF
C12487 VN.n11318 a_400_62400# 0.16fF
C12488 VN.t2264 a_400_62400# 0.03fF
C12489 VN.n11319 a_400_62400# 0.19fF
C12490 VN.n11321 a_400_62400# 2.42fF
C12491 VN.n11322 a_400_62400# 2.53fF
C12492 VN.n11323 a_400_62400# 2.75fF
C12493 VN.t2452 a_400_62400# 0.03fF
C12494 VN.n11324 a_400_62400# 0.16fF
C12495 VN.n11325 a_400_62400# 0.19fF
C12496 VN.t337 a_400_62400# 0.03fF
C12497 VN.n11327 a_400_62400# 0.32fF
C12498 VN.n11328 a_400_62400# 1.22fF
C12499 VN.n11329 a_400_62400# 0.07fF
C12500 VN.n11330 a_400_62400# 1.03fF
C12501 VN.n11331 a_400_62400# 1.66fF
C12502 VN.n11332 a_400_62400# 1.71fF
C12503 VN.n11333 a_400_62400# 2.51fF
C12504 VN.n11334 a_400_62400# 0.16fF
C12505 VN.t613 a_400_62400# 0.03fF
C12506 VN.n11335 a_400_62400# 0.19fF
C12507 VN.t1735 a_400_62400# 0.03fF
C12508 VN.n11337 a_400_62400# 0.32fF
C12509 VN.n11338 a_400_62400# 0.48fF
C12510 VN.n11339 a_400_62400# 0.81fF
C12511 VN.n11340 a_400_62400# 3.68fF
C12512 VN.n11341 a_400_62400# 2.90fF
C12513 VN.t797 a_400_62400# 0.03fF
C12514 VN.n11342 a_400_62400# 0.16fF
C12515 VN.n11343 a_400_62400# 0.19fF
C12516 VN.t1203 a_400_62400# 0.03fF
C12517 VN.n11345 a_400_62400# 0.32fF
C12518 VN.n11346 a_400_62400# 1.22fF
C12519 VN.n11347 a_400_62400# 0.07fF
C12520 VN.n11348 a_400_62400# 3.68fF
C12521 VN.t21 a_400_62400# 0.03fF
C12522 VN.n11349 a_400_62400# 0.32fF
C12523 VN.n11350 a_400_62400# 0.48fF
C12524 VN.n11351 a_400_62400# 0.81fF
C12525 VN.n11352 a_400_62400# 0.16fF
C12526 VN.t1481 a_400_62400# 0.03fF
C12527 VN.n11353 a_400_62400# 0.19fF
C12528 VN.n11355 a_400_62400# 2.40fF
C12529 VN.n11356 a_400_62400# 2.53fF
C12530 VN.n11357 a_400_62400# 2.75fF
C12531 VN.t1546 a_400_62400# 0.03fF
C12532 VN.n11358 a_400_62400# 0.16fF
C12533 VN.n11359 a_400_62400# 0.19fF
C12534 VN.t2075 a_400_62400# 0.03fF
C12535 VN.n11361 a_400_62400# 0.32fF
C12536 VN.n11362 a_400_62400# 1.22fF
C12537 VN.n11363 a_400_62400# 0.07fF
C12538 VN.t430 a_400_62400# 0.03fF
C12539 VN.n11364 a_400_62400# 1.28fF
C12540 VN.n11365 a_400_62400# 0.94fF
C12541 VN.t945 a_400_62400# 0.03fF
C12542 VN.n11366 a_400_62400# 1.63fF
C12543 VN.n11367 a_400_62400# 0.81fF
C12544 VN.n11368 a_400_62400# 1.21fF
C12545 VN.n11369 a_400_62400# 1.54fF
C12546 VN.n11370 a_400_62400# 4.06fF
C12547 VN.t20 a_400_62400# 28.64fF
C12548 VN.n11371 a_400_62400# 28.43fF
C12549 VN.n11373 a_400_62400# 0.50fF
C12550 VN.n11374 a_400_62400# 0.31fF
C12551 VN.n11375 a_400_62400# 3.87fF
C12552 VN.n11376 a_400_62400# 3.29fF
C12553 VN.n11377 a_400_62400# 1.06fF
C12554 VN.n11378 a_400_62400# 3.07fF
C12555 VN.n11379 a_400_62400# 5.74fF
C12556 VN.n11380 a_400_62400# 0.34fF
C12557 VN.n11381 a_400_62400# 0.02fF
C12558 VN.t2348 a_400_62400# 0.03fF
C12559 VN.n11382 a_400_62400# 0.34fF
C12560 VN.t35 a_400_62400# 64.69fF
C12561 VN.t306 a_400_62400# 0.03fF
C12562 VN.n11383 a_400_62400# 0.16fF
C12563 VN.n11384 a_400_62400# 0.19fF
C12564 VN.t2205 a_400_62400# 0.03fF
C12565 VN.n11386 a_400_62400# 0.32fF
C12566 VN.n11387 a_400_62400# 1.22fF
C12567 VN.n11388 a_400_62400# 0.07fF
C12568 VN.t1264 a_400_62400# 0.03fF
C12569 VN.n11389 a_400_62400# 0.32fF
C12570 VN.n11390 a_400_62400# 0.48fF
C12571 VN.n11391 a_400_62400# 0.81fF
C12572 VN.n11392 a_400_62400# 1.21fF
C12573 VN.n11393 a_400_62400# 1.03fF
C12574 VN.n11394 a_400_62400# 1.30fF
C12575 VN.n11395 a_400_62400# 0.12fF
C12576 VN.n11396 a_400_62400# 0.44fF
C12577 VN.n11397 a_400_62400# 2.89fF
C12578 VN.n11398 a_400_62400# 3.50fF
C12579 VN.n11399 a_400_62400# 2.51fF
C12580 VN.n11400 a_400_62400# 0.16fF
C12581 VN.t406 a_400_62400# 0.03fF
C12582 VN.n11401 a_400_62400# 0.19fF
C12583 VN.t2404 a_400_62400# 0.03fF
C12584 VN.n11403 a_400_62400# 0.32fF
C12585 VN.n11404 a_400_62400# 0.48fF
C12586 VN.n11405 a_400_62400# 0.81fF
C12587 VN.n11406 a_400_62400# 0.28fF
C12588 VN.n11407 a_400_62400# 0.21fF
C12589 VN.n11408 a_400_62400# 0.38fF
C12590 VN.n11409 a_400_62400# 0.29fF
C12591 VN.n11410 a_400_62400# 1.05fF
C12592 VN.n11411 a_400_62400# 0.42fF
C12593 VN.n11412 a_400_62400# 0.30fF
C12594 VN.n11413 a_400_62400# 0.51fF
C12595 VN.n11414 a_400_62400# 4.83fF
C12596 VN.t1456 a_400_62400# 0.03fF
C12597 VN.n11415 a_400_62400# 0.32fF
C12598 VN.n11416 a_400_62400# 1.22fF
C12599 VN.n11417 a_400_62400# 0.07fF
C12600 VN.t1777 a_400_62400# 0.03fF
C12601 VN.n11418 a_400_62400# 0.16fF
C12602 VN.n11419 a_400_62400# 0.19fF
C12603 VN.n11421 a_400_62400# 0.33fF
C12604 VN.n11422 a_400_62400# 0.12fF
C12605 VN.n11423 a_400_62400# 0.28fF
C12606 VN.n11424 a_400_62400# 1.72fF
C12607 VN.n11425 a_400_62400# 0.71fF
C12608 VN.n11426 a_400_62400# 2.51fF
C12609 VN.n11427 a_400_62400# 0.16fF
C12610 VN.t2056 a_400_62400# 0.03fF
C12611 VN.n11428 a_400_62400# 0.19fF
C12612 VN.t1536 a_400_62400# 0.03fF
C12613 VN.n11430 a_400_62400# 0.32fF
C12614 VN.n11431 a_400_62400# 0.48fF
C12615 VN.n11432 a_400_62400# 0.81fF
C12616 VN.n11433 a_400_62400# 0.28fF
C12617 VN.n11434 a_400_62400# 0.21fF
C12618 VN.n11435 a_400_62400# 0.38fF
C12619 VN.n11436 a_400_62400# 0.29fF
C12620 VN.n11437 a_400_62400# 0.40fF
C12621 VN.n11438 a_400_62400# 0.48fF
C12622 VN.n11439 a_400_62400# 0.30fF
C12623 VN.n11440 a_400_62400# 0.51fF
C12624 VN.n11441 a_400_62400# 3.24fF
C12625 VN.t586 a_400_62400# 0.03fF
C12626 VN.n11442 a_400_62400# 0.32fF
C12627 VN.n11443 a_400_62400# 1.22fF
C12628 VN.n11444 a_400_62400# 0.07fF
C12629 VN.t188 a_400_62400# 0.03fF
C12630 VN.n11445 a_400_62400# 0.16fF
C12631 VN.n11446 a_400_62400# 0.19fF
C12632 VN.n11448 a_400_62400# 2.53fF
C12633 VN.n11449 a_400_62400# 3.57fF
C12634 VN.t664 a_400_62400# 0.03fF
C12635 VN.n11450 a_400_62400# 0.32fF
C12636 VN.n11451 a_400_62400# 0.48fF
C12637 VN.n11452 a_400_62400# 0.81fF
C12638 VN.n11453 a_400_62400# 0.16fF
C12639 VN.t1186 a_400_62400# 0.03fF
C12640 VN.n11454 a_400_62400# 0.19fF
C12641 VN.n11456 a_400_62400# 0.30fF
C12642 VN.n11457 a_400_62400# 0.34fF
C12643 VN.n11458 a_400_62400# 0.12fF
C12644 VN.n11459 a_400_62400# 0.30fF
C12645 VN.n11460 a_400_62400# 0.93fF
C12646 VN.n11461 a_400_62400# 1.55fF
C12647 VN.n11462 a_400_62400# 0.29fF
C12648 VN.n11463 a_400_62400# 0.34fF
C12649 VN.n11464 a_400_62400# 0.12fF
C12650 VN.n11465 a_400_62400# 2.52fF
C12651 VN.t2242 a_400_62400# 0.03fF
C12652 VN.n11466 a_400_62400# 0.32fF
C12653 VN.n11467 a_400_62400# 1.22fF
C12654 VN.n11468 a_400_62400# 0.07fF
C12655 VN.t1846 a_400_62400# 0.03fF
C12656 VN.n11469 a_400_62400# 0.16fF
C12657 VN.n11470 a_400_62400# 0.19fF
C12658 VN.n11472 a_400_62400# 27.83fF
C12659 VN.n11473 a_400_62400# 2.30fF
C12660 VN.n11474 a_400_62400# 4.08fF
C12661 VN.t1566 a_400_62400# 0.03fF
C12662 VN.n11475 a_400_62400# 0.32fF
C12663 VN.n11476 a_400_62400# 0.48fF
C12664 VN.n11477 a_400_62400# 0.81fF
C12665 VN.n11478 a_400_62400# 0.16fF
C12666 VN.t713 a_400_62400# 0.03fF
C12667 VN.n11479 a_400_62400# 0.19fF
C12668 VN.n11481 a_400_62400# 0.37fF
C12669 VN.n11482 a_400_62400# 0.99fF
C12670 VN.n11483 a_400_62400# 0.80fF
C12671 VN.n11484 a_400_62400# 0.28fF
C12672 VN.n11485 a_400_62400# 0.27fF
C12673 VN.n11486 a_400_62400# 0.09fF
C12674 VN.n11487 a_400_62400# 0.12fF
C12675 VN.n11488 a_400_62400# 0.13fF
C12676 VN.n11489 a_400_62400# 2.66fF
C12677 VN.t1513 a_400_62400# 0.03fF
C12678 VN.n11490 a_400_62400# 0.16fF
C12679 VN.n11491 a_400_62400# 0.19fF
C12680 VN.t143 a_400_62400# 0.03fF
C12681 VN.n11493 a_400_62400# 0.32fF
C12682 VN.n11494 a_400_62400# 1.22fF
C12683 VN.n11495 a_400_62400# 0.07fF
C12684 VN.n11496 a_400_62400# 3.65fF
C12685 VN.n11497 a_400_62400# 2.51fF
C12686 VN.n11498 a_400_62400# 0.16fF
C12687 VN.t317 a_400_62400# 0.03fF
C12688 VN.n11499 a_400_62400# 0.19fF
C12689 VN.t2326 a_400_62400# 0.03fF
C12690 VN.n11501 a_400_62400# 0.32fF
C12691 VN.n11502 a_400_62400# 0.48fF
C12692 VN.n11503 a_400_62400# 0.81fF
C12693 VN.n11504 a_400_62400# 0.94fF
C12694 VN.n11505 a_400_62400# 1.71fF
C12695 VN.n11506 a_400_62400# 7.99fF
C12696 VN.t976 a_400_62400# 0.03fF
C12697 VN.n11507 a_400_62400# 0.16fF
C12698 VN.n11508 a_400_62400# 0.19fF
C12699 VN.t1379 a_400_62400# 0.03fF
C12700 VN.n11510 a_400_62400# 0.32fF
C12701 VN.n11511 a_400_62400# 1.22fF
C12702 VN.n11512 a_400_62400# 0.07fF
C12703 VN.t106 a_400_62400# 64.17fF
C12704 VN.t243 a_400_62400# 0.03fF
C12705 VN.n11513 a_400_62400# 0.02fF
C12706 VN.n11514 a_400_62400# 0.34fF
C12707 VN.t514 a_400_62400# 0.03fF
C12708 VN.n11516 a_400_62400# 1.60fF
C12709 VN.n11517 a_400_62400# 0.07fF
C12710 VN.t1460 a_400_62400# 0.03fF
C12711 VN.n11518 a_400_62400# 0.85fF
C12712 VN.n11519 a_400_62400# 0.81fF
C12713 VN.n11520 a_400_62400# 2.01fF
C12714 VN.n11521 a_400_62400# 0.47fF
C12715 VN.n11522 a_400_62400# 1.74fF
C12716 VN.n11523 a_400_62400# 0.21fF
C12717 VN.n11524 a_400_62400# 2.23fF
C12718 VN.n11525 a_400_62400# 3.54fF
C12719 VN.n11526 a_400_62400# 1.52fF
C12720 VN.n11527 a_400_62400# 145.00fF
C12721 VN.n11528 a_400_62400# 145.00fF
C12722 VN.n11529 a_400_62400# 0.28fF
C12723 VN.n11530 a_400_62400# 1.89fF
C12724 VN.t110 a_400_62400# 28.64fF
C12725 VN.n11531 a_400_62400# 1.18fF
C12726 VN.n11532 a_400_62400# 0.11fF
C12727 VN.n11533 a_400_62400# 1.18fF
C12728 VN.n11534 a_400_62400# 4.98fF
C12729 VN.n11535 a_400_62400# 0.80fF
C12730 VN.n11536 a_400_62400# 0.29fF
C12731 VN.n11537 a_400_62400# 1.96fF
C12732 VN.n11539 a_400_62400# 25.18fF
C12733 VN.n11541 a_400_62400# 1.87fF
C12734 VN.n11542 a_400_62400# 5.69fF
C12735 VN.n11543 a_400_62400# 2.41fF
C12736 VN.t1440 a_400_62400# 0.03fF
C12737 VN.n11544 a_400_62400# 0.85fF
C12738 VN.n11545 a_400_62400# 0.81fF
C12739 VN.n11546 a_400_62400# 0.32fF
C12740 VN.t464 a_400_62400# 0.03fF
C12741 VN.n11547 a_400_62400# 0.48fF
C12742 VN.n11548 a_400_62400# 0.48fF
C12743 VN.n11549 a_400_62400# 0.90fF
C12744 VN.n11550 a_400_62400# 0.28fF
C12745 VN.n11551 a_400_62400# 0.27fF
C12746 VN.n11552 a_400_62400# 0.09fF
C12747 VN.n11553 a_400_62400# 0.12fF
C12748 VN.n11554 a_400_62400# 0.13fF
C12749 VN.n11555 a_400_62400# 0.58fF
C12750 VN.n11556 a_400_62400# 0.34fF
C12751 VN.n11557 a_400_62400# 1.25fF
C12752 VN.n11558 a_400_62400# 0.28fF
C12753 VN.n11559 a_400_62400# 0.60fF
C12754 VN.n11560 a_400_62400# 3.51fF
C12755 VN.n11561 a_400_62400# 2.62fF
C12756 VN.n11562 a_400_62400# 0.28fF
C12757 VN.n11563 a_400_62400# 1.64fF
C12758 VN.n11564 a_400_62400# 0.59fF
C12759 VN.n11565 a_400_62400# 0.33fF
C12760 VN.n11566 a_400_62400# 0.12fF
C12761 VN.n11567 a_400_62400# 0.75fF
C12762 VN.n11568 a_400_62400# 0.32fF
C12763 VN.t2148 a_400_62400# 0.03fF
C12764 VN.n11569 a_400_62400# 0.48fF
C12765 VN.n11570 a_400_62400# 0.84fF
C12766 VN.n11571 a_400_62400# 0.53fF
C12767 VN.n11572 a_400_62400# 0.53fF
C12768 VN.n11573 a_400_62400# 0.16fF
C12769 VN.t987 a_400_62400# 0.03fF
C12770 VN.n11574 a_400_62400# 0.19fF
C12771 VN.t1788 a_400_62400# 0.03fF
C12772 VN.n11576 a_400_62400# 0.16fF
C12773 VN.n11577 a_400_62400# 0.19fF
C12774 VN.n11579 a_400_62400# 0.87fF
C12775 VN.n11580 a_400_62400# 0.51fF
C12776 VN.n11581 a_400_62400# 0.59fF
C12777 VN.n11582 a_400_62400# 2.16fF
C12778 VN.n11583 a_400_62400# 0.67fF
C12779 VN.n11584 a_400_62400# 0.62fF
C12780 VN.n11585 a_400_62400# 0.60fF
C12781 VN.n11586 a_400_62400# 2.47fF
C12782 VN.n11587 a_400_62400# 0.16fF
C12783 VN.t252 a_400_62400# 0.03fF
C12784 VN.n11588 a_400_62400# 0.19fF
C12785 VN.t1278 a_400_62400# 0.03fF
C12786 VN.n11590 a_400_62400# 0.32fF
C12787 VN.n11591 a_400_62400# 0.48fF
C12788 VN.n11592 a_400_62400# 0.81fF
C12789 VN.n11593 a_400_62400# 3.34fF
C12790 VN.n11594 a_400_62400# 2.71fF
C12791 VN.t2114 a_400_62400# 0.03fF
C12792 VN.n11595 a_400_62400# 0.32fF
C12793 VN.n11596 a_400_62400# 1.22fF
C12794 VN.n11597 a_400_62400# 0.07fF
C12795 VN.t913 a_400_62400# 0.03fF
C12796 VN.n11598 a_400_62400# 0.16fF
C12797 VN.n11599 a_400_62400# 0.19fF
C12798 VN.n11601 a_400_62400# 0.24fF
C12799 VN.n11602 a_400_62400# 0.13fF
C12800 VN.n11603 a_400_62400# 1.27fF
C12801 VN.n11604 a_400_62400# 0.62fF
C12802 VN.n11605 a_400_62400# 0.28fF
C12803 VN.n11606 a_400_62400# 0.48fF
C12804 VN.n11607 a_400_62400# 0.71fF
C12805 VN.n11608 a_400_62400# 3.52fF
C12806 VN.n11609 a_400_62400# 2.00fF
C12807 VN.n11610 a_400_62400# 0.16fF
C12808 VN.t1902 a_400_62400# 0.03fF
C12809 VN.n11611 a_400_62400# 0.19fF
C12810 VN.t536 a_400_62400# 0.03fF
C12811 VN.n11613 a_400_62400# 0.32fF
C12812 VN.n11614 a_400_62400# 0.48fF
C12813 VN.n11615 a_400_62400# 0.81fF
C12814 VN.n11616 a_400_62400# 3.32fF
C12815 VN.n11617 a_400_62400# 2.63fF
C12816 VN.t1370 a_400_62400# 0.03fF
C12817 VN.n11618 a_400_62400# 0.32fF
C12818 VN.n11619 a_400_62400# 1.22fF
C12819 VN.n11620 a_400_62400# 0.07fF
C12820 VN.t2575 a_400_62400# 0.03fF
C12821 VN.n11621 a_400_62400# 0.16fF
C12822 VN.n11622 a_400_62400# 0.19fF
C12823 VN.n11624 a_400_62400# 0.87fF
C12824 VN.n11625 a_400_62400# 0.51fF
C12825 VN.n11626 a_400_62400# 0.59fF
C12826 VN.n11627 a_400_62400# 2.16fF
C12827 VN.n11628 a_400_62400# 0.67fF
C12828 VN.n11629 a_400_62400# 0.62fF
C12829 VN.n11630 a_400_62400# 0.60fF
C12830 VN.n11631 a_400_62400# 2.47fF
C12831 VN.n11632 a_400_62400# 0.16fF
C12832 VN.t1027 a_400_62400# 0.03fF
C12833 VN.n11633 a_400_62400# 0.19fF
C12834 VN.t2191 a_400_62400# 0.03fF
C12835 VN.n11635 a_400_62400# 0.32fF
C12836 VN.n11636 a_400_62400# 0.48fF
C12837 VN.n11637 a_400_62400# 0.81fF
C12838 VN.n11638 a_400_62400# 3.34fF
C12839 VN.n11639 a_400_62400# 2.71fF
C12840 VN.t504 a_400_62400# 0.03fF
C12841 VN.n11640 a_400_62400# 0.32fF
C12842 VN.n11641 a_400_62400# 1.22fF
C12843 VN.n11642 a_400_62400# 0.07fF
C12844 VN.t1703 a_400_62400# 0.03fF
C12845 VN.n11643 a_400_62400# 0.16fF
C12846 VN.n11644 a_400_62400# 0.19fF
C12847 VN.n11646 a_400_62400# 0.24fF
C12848 VN.n11647 a_400_62400# 0.13fF
C12849 VN.n11648 a_400_62400# 1.27fF
C12850 VN.n11649 a_400_62400# 0.62fF
C12851 VN.n11650 a_400_62400# 0.28fF
C12852 VN.n11651 a_400_62400# 0.48fF
C12853 VN.n11652 a_400_62400# 0.71fF
C12854 VN.n11653 a_400_62400# 41.70fF
C12855 VN.n11654 a_400_62400# 41.70fF
C12856 VN.n11655 a_400_62400# 7.09fF
C12857 VN.n11656 a_400_62400# 1.28fF
C12858 VN.n11657 a_400_62400# 0.46fF
C12859 VN.n11658 a_400_62400# 0.45fF
C12860 VN.n11659 a_400_62400# 7.20fF
C12861 VN.n11660 a_400_62400# 2.75fF
C12862 VN.n11661 a_400_62400# 0.46fF
C12863 VN.n11662 a_400_62400# 0.40fF
C12864 VN.n11663 a_400_62400# 1.28fF
C12865 VN.t1823 a_400_62400# 0.03fF
C12866 VN.n11664 a_400_62400# 1.20fF
C12867 VN.n11665 a_400_62400# 0.02fF
C12868 VN.t387 a_400_62400# 0.03fF
C12869 VN.n11666 a_400_62400# 0.49fF
C12870 VN.t1754 a_400_62400# 0.03fF
C12871 VN.n11667 a_400_62400# 1.19fF
C12872 VN.n11668 a_400_62400# 2.17fF
C12873 VN.n11669 a_400_62400# 4.37fF
C12874 VN.n11670 a_400_62400# 135.89fF
C12875 VN.n11671 a_400_62400# 135.89fF
C12876 VN.n11672 a_400_62400# 7.74fF
C12877 VN.n11673 a_400_62400# 2.62fF
C12878 VN.t1053 a_400_62400# 0.03fF
C12879 VN.n11674 a_400_62400# 1.20fF
C12880 VN.n11675 a_400_62400# 0.02fF
C12881 VN.t2020 a_400_62400# 0.03fF
C12882 VN.n11676 a_400_62400# 0.49fF
C12883 VN.t983 a_400_62400# 0.03fF
C12884 VN.n11677 a_400_62400# 1.19fF
C12885 VN.n11678 a_400_62400# 41.70fF
C12886 VN.n11679 a_400_62400# 41.70fF
C12887 VN.n11680 a_400_62400# 7.48fF
C12888 VN.n11681 a_400_62400# 2.02fF
C12889 VN.n11682 a_400_62400# 2.16fF
C12890 VN.t1928 a_400_62400# 0.03fF
C12891 VN.n11683 a_400_62400# 1.20fF
C12892 VN.n11684 a_400_62400# 0.02fF
C12893 VN.t367 a_400_62400# 0.03fF
C12894 VN.n11685 a_400_62400# 0.49fF
C12895 VN.t1727 a_400_62400# 0.03fF
C12896 VN.n11686 a_400_62400# 1.19fF
C12897 VN.n11687 a_400_62400# 1.52fF
C12898 VN.n11688 a_400_62400# 0.00fF
C12899 VN.n11689 a_400_62400# 0.53fF
C12900 VN.n11690 a_400_62400# 41.70fF
C12901 VN.n11691 a_400_62400# 41.70fF
C12902 VN.n11692 a_400_62400# 7.59fF
C12903 VN.n11693 a_400_62400# 2.38fF
C12904 VN.n11694 a_400_62400# 0.50fF
C12905 VN.n11695 a_400_62400# 1.11fF
C12906 VN.t278 a_400_62400# 0.03fF
C12907 VN.n11696 a_400_62400# 1.20fF
C12908 VN.n11697 a_400_62400# 0.02fF
C12909 VN.t1232 a_400_62400# 0.03fF
C12910 VN.n11698 a_400_62400# 0.49fF
C12911 VN.t9 a_400_62400# 0.03fF
C12912 VN.n11699 a_400_62400# 1.19fF
C12913 VN.n11700 a_400_62400# 1.41fF
C12914 VN.n11701 a_400_62400# 0.56fF
C12915 VN.n11702 a_400_62400# 0.36fF
C12916 VN.n11703 a_400_62400# 4.37fF
C12917 VN.n11704 a_400_62400# 0.41fF
C12918 VN.n11705 a_400_62400# 41.70fF
C12919 VN.n11706 a_400_62400# 41.70fF
C12920 VN.n11707 a_400_62400# 7.02fF
C12921 VN.n11708 a_400_62400# 1.34fF
C12922 VN.t1142 a_400_62400# 0.03fF
C12923 VN.n11709 a_400_62400# 1.20fF
C12924 VN.n11710 a_400_62400# 0.02fF
C12925 VN.t2109 a_400_62400# 0.03fF
C12926 VN.n11711 a_400_62400# 0.49fF
C12927 VN.t933 a_400_62400# 0.03fF
C12928 VN.n11712 a_400_62400# 1.19fF
C12929 VN.n11713 a_400_62400# 41.70fF
C12930 VN.n11714 a_400_62400# 41.70fF
C12931 VN.n11715 a_400_62400# 7.32fF
C12932 VN.n11716 a_400_62400# 2.62fF
C12933 VN.n11717 a_400_62400# 4.37fF
C12934 VN.n11718 a_400_62400# 0.41fF
C12935 VN.n11719 a_400_62400# 1.34fF
C12936 VN.t1461 a_400_62400# 0.03fF
C12937 VN.n11720 a_400_62400# 1.20fF
C12938 VN.n11721 a_400_62400# 0.02fF
C12939 VN.t2398 a_400_62400# 0.03fF
C12940 VN.n11722 a_400_62400# 0.49fF
C12941 VN.t1266 a_400_62400# 0.03fF
C12942 VN.n11723 a_400_62400# 1.19fF
C12943 VN.n11724 a_400_62400# 41.70fF
C12944 VN.n11725 a_400_62400# 41.70fF
C12945 VN.n11726 a_400_62400# 7.32fF
C12946 VN.n11727 a_400_62400# 2.62fF
C12947 VN.n11728 a_400_62400# 4.37fF
C12948 VN.n11729 a_400_62400# 0.41fF
C12949 VN.n11730 a_400_62400# 1.34fF
C12950 VN.t547 a_400_62400# 0.03fF
C12951 VN.n11731 a_400_62400# 1.20fF
C12952 VN.n11732 a_400_62400# 0.02fF
C12953 VN.t1607 a_400_62400# 0.03fF
C12954 VN.n11733 a_400_62400# 0.49fF
C12955 VN.t486 a_400_62400# 0.03fF
C12956 VN.n11734 a_400_62400# 1.19fF
C12957 VN.n11735 a_400_62400# 41.70fF
C12958 VN.n11736 a_400_62400# 41.70fF
C12959 VN.n11737 a_400_62400# 7.41fF
C12960 VN.n11738 a_400_62400# 2.62fF
C12961 VN.n11739 a_400_62400# 4.37fF
C12962 VN.n11740 a_400_62400# 0.41fF
C12963 VN.n11741 a_400_62400# 1.34fF
C12964 VN.t2277 a_400_62400# 0.03fF
C12965 VN.n11742 a_400_62400# 1.20fF
C12966 VN.n11743 a_400_62400# 0.02fF
C12967 VN.t813 a_400_62400# 0.03fF
C12968 VN.n11744 a_400_62400# 0.49fF
C12969 VN.t2219 a_400_62400# 0.03fF
C12970 VN.n11745 a_400_62400# 1.19fF
C12971 VN.n11746 a_400_62400# 41.70fF
C12972 VN.n11747 a_400_62400# 41.70fF
C12973 VN.n11748 a_400_62400# 7.32fF
C12974 VN.n11749 a_400_62400# 2.62fF
C12975 VN.n11750 a_400_62400# 4.37fF
C12976 VN.n11751 a_400_62400# 0.41fF
C12977 VN.n11752 a_400_62400# 1.34fF
C12978 VN.t1490 a_400_62400# 0.03fF
C12979 VN.n11753 a_400_62400# 1.20fF
C12980 VN.n11754 a_400_62400# 0.02fF
C12981 VN.t2426 a_400_62400# 0.03fF
C12982 VN.n11755 a_400_62400# 0.49fF
C12983 VN.t1307 a_400_62400# 0.03fF
C12984 VN.n11756 a_400_62400# 1.19fF
C12985 VN.n11757 a_400_62400# 41.70fF
C12986 VN.n11758 a_400_62400# 41.70fF
C12987 VN.n11759 a_400_62400# 7.32fF
C12988 VN.n11760 a_400_62400# 2.62fF
C12989 VN.n11761 a_400_62400# 4.37fF
C12990 VN.n11762 a_400_62400# 0.41fF
C12991 VN.n11763 a_400_62400# 1.34fF
C12992 VN.t1867 a_400_62400# 0.03fF
C12993 VN.n11764 a_400_62400# 1.20fF
C12994 VN.n11765 a_400_62400# 0.02fF
C12995 VN.t300 a_400_62400# 0.03fF
C12996 VN.n11766 a_400_62400# 0.49fF
C12997 VN.t1674 a_400_62400# 0.03fF
C12998 VN.n11767 a_400_62400# 1.19fF
C12999 VN.n11768 a_400_62400# 7.36fF
C13000 VN.n11769 a_400_62400# 2.62fF
C13001 VN.n11770 a_400_62400# 4.37fF
C13002 VN.n11771 a_400_62400# 0.41fF
C13003 VN.n11772 a_400_62400# 1.34fF
C13004 VN.t1088 a_400_62400# 0.03fF
C13005 VN.n11773 a_400_62400# 1.20fF
C13006 VN.n11774 a_400_62400# 0.02fF
C13007 VN.t2041 a_400_62400# 0.03fF
C13008 VN.n11775 a_400_62400# 0.49fF
C13009 VN.t880 a_400_62400# 0.03fF
C13010 VN.n11776 a_400_62400# 1.19fF
C13011 VN.t60 a_400_62400# 0.03fF
C13012 VN.n11777 a_400_62400# 0.59fF
C13013 VN.n11778 a_400_62400# 72.42fF
C13014 VN.n11779 a_400_62400# 2.97fF
C13015 VN.n11780 a_400_62400# 1.20fF
C13016 VN.n11781 a_400_62400# 0.70fF
C13017 VN.n11782 a_400_62400# 4.93fF
C13018 VN.n11783 a_400_62400# 41.70fF
C13019 VN.n11784 a_400_62400# 65.40fF
C13020 VN.n11785 a_400_62400# 41.70fF
C13021 VN.n11786 a_400_62400# 65.40fF
C13022 VN.n11787 a_400_62400# 17.08fF
C13023 VN.n11788 a_400_62400# 2.54fF
C13024 VN.n11789 a_400_62400# 12.03fF
C13025 VN.t1256 a_400_62400# 0.03fF
C13026 VN.n11790 a_400_62400# 1.75fF
C13027 VN.n11791 a_400_62400# 0.42fF
C13028 VN.n11792 a_400_62400# 1.28fF
C13029 VN.n11793 a_400_62400# 0.46fF
C13030 VN.n11794 a_400_62400# 0.45fF
C13031 VN.n11795 a_400_62400# 41.70fF
C13032 VN.n11796 a_400_62400# 41.70fF
C13033 VN.n11797 a_400_62400# 7.28fF
C13034 VN.n11798 a_400_62400# 2.91fF
C13035 VN.t216 a_400_62400# 0.03fF
C13036 VN.n11799 a_400_62400# 1.20fF
C13037 VN.n11800 a_400_62400# 0.02fF
C13038 VN.t1169 a_400_62400# 0.03fF
C13039 VN.n11801 a_400_62400# 0.49fF
C13040 VN.t2539 a_400_62400# 0.03fF
C13041 VN.n11802 a_400_62400# 1.19fF
C13042 VN.n11803 a_400_62400# 1.28fF
C13043 VN.n11804 a_400_62400# 0.46fF
C13044 VN.n11805 a_400_62400# 0.45fF
C13045 VN.n11806 a_400_62400# 41.70fF
C13046 VN.n11807 a_400_62400# 41.70fF
C13047 VN.n11808 a_400_62400# 7.28fF
C13048 VN.n11809 a_400_62400# 2.91fF
C13049 VN.t2358 a_400_62400# 0.03fF
C13050 VN.n11810 a_400_62400# 1.20fF
C13051 VN.n11811 a_400_62400# 0.02fF
C13052 VN.t776 a_400_62400# 0.03fF
C13053 VN.n11812 a_400_62400# 0.49fF
C13054 VN.t2174 a_400_62400# 0.03fF
C13055 VN.n11813 a_400_62400# 1.19fF
C13056 VN.n11814 a_400_62400# 1.28fF
C13057 VN.n11815 a_400_62400# 0.46fF
C13058 VN.n11816 a_400_62400# 0.45fF
C13059 VN.n11817 a_400_62400# 41.70fF
C13060 VN.n11818 a_400_62400# 41.70fF
C13061 VN.n11819 a_400_62400# 7.28fF
C13062 VN.n11820 a_400_62400# 2.91fF
C13063 VN.t1407 a_400_62400# 0.03fF
C13064 VN.n11821 a_400_62400# 1.20fF
C13065 VN.n11822 a_400_62400# 0.02fF
C13066 VN.t2470 a_400_62400# 0.03fF
C13067 VN.n11823 a_400_62400# 0.49fF
C13068 VN.t1354 a_400_62400# 0.03fF
C13069 VN.n11824 a_400_62400# 1.19fF
C13070 VN.n11825 a_400_62400# 1.28fF
C13071 VN.n11826 a_400_62400# 0.46fF
C13072 VN.n11827 a_400_62400# 0.45fF
C13073 VN.n11828 a_400_62400# 41.70fF
C13074 VN.n11829 a_400_62400# 41.70fF
C13075 VN.n11830 a_400_62400# 7.28fF
C13076 VN.n11831 a_400_62400# 2.91fF
C13077 VN.t2202 a_400_62400# 0.03fF
C13078 VN.n11832 a_400_62400# 1.20fF
C13079 VN.n11833 a_400_62400# 0.02fF
C13080 VN.t741 a_400_62400# 0.03fF
C13081 VN.n11834 a_400_62400# 0.49fF
C13082 VN.t2140 a_400_62400# 0.03fF
C13083 VN.n11835 a_400_62400# 1.19fF
C13084 VN.n11836 a_400_62400# 1.28fF
C13085 VN.n11837 a_400_62400# 0.46fF
C13086 VN.n11838 a_400_62400# 0.45fF
C13087 VN.n11839 a_400_62400# 41.70fF
C13088 VN.n11840 a_400_62400# 41.70fF
C13089 VN.n11841 a_400_62400# 5.49fF
C13090 VN.n11842 a_400_62400# 5.49fF
C13091 VN.n11843 a_400_62400# 5.44fF
C13092 VN.n11844 a_400_62400# 5.49fF
C13093 VN.n11845 a_400_62400# 5.49fF
C13094 VN.n11846 a_400_62400# 5.56fF
C13095 VN.n11847 a_400_62400# 5.73fF
C13096 VN.n11848 a_400_62400# 5.74fF
C13097 VN.n11849 a_400_62400# 6.30fF
C13098 VN.n11850 a_400_62400# 2.95fF
C13099 VN.n11851 a_400_62400# 5.53fF
C13100 VN.n11852 a_400_62400# 169.21fF
C13101 VN.n11853 a_400_62400# 5.56fF
C13102 VN.n11854 a_400_62400# 7.21fF
C13103 VN.n11855 a_400_62400# 2.91fF
C13104 VN.t590 a_400_62400# 0.03fF
C13105 VN.n11856 a_400_62400# 1.20fF
C13106 VN.n11857 a_400_62400# 0.02fF
C13107 VN.t1529 a_400_62400# 0.03fF
C13108 VN.n11858 a_400_62400# 0.49fF
C13109 VN.t397 a_400_62400# 0.03fF
C13110 VN.n11859 a_400_62400# 1.19fF
C13111 VN.n11860 a_400_62400# 0.02fF
C13112 VN.t1563 a_400_62400# 0.03fF
C13113 VN.n11861 a_400_62400# 0.49fF
C13114 VN.t625 a_400_62400# 0.03fF
C13115 VN.n11862 a_400_62400# 1.20fF
C13116 VN.t560 a_400_62400# 0.03fF
C13117 VN.n11863 a_400_62400# 1.19fF
C13118 VN.n11864 a_400_62400# 0.46fF
C13119 VN.n11865 a_400_62400# 0.40fF
C13120 VN.n11866 a_400_62400# 1.28fF
C13121 VN.t8 a_400_62400# 171.82fF
C13122 VN.n11867 a_400_62400# 3.52fF
C13123 VN.n11868 a_400_62400# 2.00fF
C13124 VN.n11869 a_400_62400# 0.16fF
C13125 VN.t1523 a_400_62400# 0.03fF
C13126 VN.n11870 a_400_62400# 0.19fF
C13127 VN.t111 a_400_62400# 0.03fF
C13128 VN.n11872 a_400_62400# 0.32fF
C13129 VN.n11873 a_400_62400# 0.48fF
C13130 VN.n11874 a_400_62400# 0.81fF
C13131 VN.n11875 a_400_62400# 3.32fF
C13132 VN.n11876 a_400_62400# 2.63fF
C13133 VN.t956 a_400_62400# 0.03fF
C13134 VN.n11877 a_400_62400# 0.32fF
C13135 VN.n11878 a_400_62400# 1.22fF
C13136 VN.n11879 a_400_62400# 0.07fF
C13137 VN.t832 a_400_62400# 0.03fF
C13138 VN.n11880 a_400_62400# 0.16fF
C13139 VN.n11881 a_400_62400# 0.19fF
C13140 VN.n11883 a_400_62400# 0.87fF
C13141 VN.n11884 a_400_62400# 0.51fF
C13142 VN.n11885 a_400_62400# 0.59fF
C13143 VN.n11886 a_400_62400# 1.79fF
C13144 VN.n11887 a_400_62400# 0.62fF
C13145 VN.n11888 a_400_62400# 0.60fF
C13146 VN.n11889 a_400_62400# 2.47fF
C13147 VN.n11890 a_400_62400# 0.16fF
C13148 VN.t653 a_400_62400# 0.03fF
C13149 VN.n11891 a_400_62400# 0.19fF
C13150 VN.t1779 a_400_62400# 0.03fF
C13151 VN.n11893 a_400_62400# 0.32fF
C13152 VN.n11894 a_400_62400# 0.48fF
C13153 VN.n11895 a_400_62400# 0.81fF
C13154 VN.n11896 a_400_62400# 3.34fF
C13155 VN.n11897 a_400_62400# 2.71fF
C13156 VN.t44 a_400_62400# 0.03fF
C13157 VN.n11898 a_400_62400# 0.32fF
C13158 VN.n11899 a_400_62400# 1.22fF
C13159 VN.n11900 a_400_62400# 0.07fF
C13160 VN.t1340 a_400_62400# 0.03fF
C13161 VN.n11901 a_400_62400# 0.16fF
C13162 VN.n11902 a_400_62400# 0.19fF
C13163 VN.n11904 a_400_62400# 0.24fF
C13164 VN.n11905 a_400_62400# 0.13fF
C13165 VN.n11906 a_400_62400# 1.27fF
C13166 VN.n11907 a_400_62400# 0.62fF
C13167 VN.n11908 a_400_62400# 0.28fF
C13168 VN.n11909 a_400_62400# 0.48fF
C13169 VN.n11910 a_400_62400# 0.71fF
C13170 VN.n11911 a_400_62400# 3.51fF
C13171 VN.n11912 a_400_62400# 2.01fF
C13172 VN.n11913 a_400_62400# 0.16fF
C13173 VN.t2312 a_400_62400# 0.03fF
C13174 VN.n11914 a_400_62400# 0.19fF
C13175 VN.t904 a_400_62400# 0.03fF
C13176 VN.n11916 a_400_62400# 0.32fF
C13177 VN.n11917 a_400_62400# 0.48fF
C13178 VN.n11918 a_400_62400# 0.81fF
C13179 VN.n11919 a_400_62400# 1.27fF
C13180 VN.n11920 a_400_62400# 0.58fF
C13181 VN.n11921 a_400_62400# 0.73fF
C13182 VN.n11922 a_400_62400# 0.44fF
C13183 VN.n11923 a_400_62400# 1.56fF
C13184 VN.n11924 a_400_62400# 2.58fF
C13185 VN.t1744 a_400_62400# 0.03fF
C13186 VN.n11925 a_400_62400# 0.32fF
C13187 VN.n11926 a_400_62400# 1.22fF
C13188 VN.n11927 a_400_62400# 0.07fF
C13189 VN.t475 a_400_62400# 0.03fF
C13190 VN.n11928 a_400_62400# 0.16fF
C13191 VN.n11929 a_400_62400# 0.19fF
C13192 VN.n11931 a_400_62400# 0.87fF
C13193 VN.n11932 a_400_62400# 0.51fF
C13194 VN.n11933 a_400_62400# 0.59fF
C13195 VN.n11934 a_400_62400# 2.16fF
C13196 VN.n11935 a_400_62400# 0.67fF
C13197 VN.n11936 a_400_62400# 0.62fF
C13198 VN.n11937 a_400_62400# 0.60fF
C13199 VN.n11938 a_400_62400# 2.47fF
C13200 VN.n11939 a_400_62400# 0.16fF
C13201 VN.t1442 a_400_62400# 0.03fF
C13202 VN.n11940 a_400_62400# 0.19fF
C13203 VN.t2566 a_400_62400# 0.03fF
C13204 VN.n11942 a_400_62400# 0.32fF
C13205 VN.n11943 a_400_62400# 0.48fF
C13206 VN.n11944 a_400_62400# 0.81fF
C13207 VN.n11945 a_400_62400# 3.34fF
C13208 VN.n11946 a_400_62400# 2.71fF
C13209 VN.t873 a_400_62400# 0.03fF
C13210 VN.n11947 a_400_62400# 0.32fF
C13211 VN.n11948 a_400_62400# 1.22fF
C13212 VN.n11949 a_400_62400# 0.07fF
C13213 VN.t2247 a_400_62400# 0.03fF
C13214 VN.n11950 a_400_62400# 0.16fF
C13215 VN.n11951 a_400_62400# 0.19fF
C13216 VN.n11953 a_400_62400# 0.24fF
C13217 VN.n11954 a_400_62400# 0.13fF
C13218 VN.n11955 a_400_62400# 1.27fF
C13219 VN.n11956 a_400_62400# 0.62fF
C13220 VN.n11957 a_400_62400# 0.28fF
C13221 VN.n11958 a_400_62400# 0.48fF
C13222 VN.n11959 a_400_62400# 0.71fF
C13223 VN.n11960 a_400_62400# 3.52fF
C13224 VN.n11961 a_400_62400# 2.00fF
C13225 VN.n11962 a_400_62400# 0.16fF
C13226 VN.t574 a_400_62400# 0.03fF
C13227 VN.n11963 a_400_62400# 0.19fF
C13228 VN.t1696 a_400_62400# 0.03fF
C13229 VN.n11965 a_400_62400# 0.32fF
C13230 VN.n11966 a_400_62400# 0.48fF
C13231 VN.n11967 a_400_62400# 0.81fF
C13232 VN.n11968 a_400_62400# 3.32fF
C13233 VN.n11969 a_400_62400# 2.63fF
C13234 VN.t2532 a_400_62400# 0.03fF
C13235 VN.n11970 a_400_62400# 0.32fF
C13236 VN.n11971 a_400_62400# 1.22fF
C13237 VN.n11972 a_400_62400# 0.07fF
C13238 VN.t1385 a_400_62400# 0.03fF
C13239 VN.n11973 a_400_62400# 0.16fF
C13240 VN.n11974 a_400_62400# 0.19fF
C13241 VN.n11976 a_400_62400# 0.87fF
C13242 VN.n11977 a_400_62400# 0.51fF
C13243 VN.n11978 a_400_62400# 0.59fF
C13244 VN.n11979 a_400_62400# 2.16fF
C13245 VN.n11980 a_400_62400# 0.67fF
C13246 VN.n11981 a_400_62400# 0.62fF
C13247 VN.n11982 a_400_62400# 0.60fF
C13248 VN.n11983 a_400_62400# 2.47fF
C13249 VN.n11984 a_400_62400# 0.16fF
C13250 VN.t2232 a_400_62400# 0.03fF
C13251 VN.n11985 a_400_62400# 0.19fF
C13252 VN.t826 a_400_62400# 0.03fF
C13253 VN.n11987 a_400_62400# 0.32fF
C13254 VN.n11988 a_400_62400# 0.48fF
C13255 VN.n11989 a_400_62400# 0.81fF
C13256 VN.n11990 a_400_62400# 3.34fF
C13257 VN.n11991 a_400_62400# 2.71fF
C13258 VN.t1668 a_400_62400# 0.03fF
C13259 VN.n11992 a_400_62400# 0.32fF
C13260 VN.n11993 a_400_62400# 1.22fF
C13261 VN.n11994 a_400_62400# 0.07fF
C13262 VN.t519 a_400_62400# 0.03fF
C13263 VN.n11995 a_400_62400# 0.16fF
C13264 VN.n11996 a_400_62400# 0.19fF
C13265 VN.n11998 a_400_62400# 0.24fF
C13266 VN.n11999 a_400_62400# 0.13fF
C13267 VN.n12000 a_400_62400# 1.27fF
C13268 VN.n12001 a_400_62400# 0.62fF
C13269 VN.n12002 a_400_62400# 0.28fF
C13270 VN.n12003 a_400_62400# 0.48fF
C13271 VN.n12004 a_400_62400# 0.71fF
C13272 VN.n12005 a_400_62400# 3.52fF
C13273 VN.n12006 a_400_62400# 2.00fF
C13274 VN.n12007 a_400_62400# 0.16fF
C13275 VN.t1367 a_400_62400# 0.03fF
C13276 VN.n12008 a_400_62400# 0.19fF
C13277 VN.t2490 a_400_62400# 0.03fF
C13278 VN.n12010 a_400_62400# 0.32fF
C13279 VN.n12011 a_400_62400# 0.48fF
C13280 VN.n12012 a_400_62400# 0.81fF
C13281 VN.n12013 a_400_62400# 3.32fF
C13282 VN.n12014 a_400_62400# 2.63fF
C13283 VN.t803 a_400_62400# 0.03fF
C13284 VN.n12015 a_400_62400# 0.32fF
C13285 VN.n12016 a_400_62400# 1.22fF
C13286 VN.n12017 a_400_62400# 0.07fF
C13287 VN.t2170 a_400_62400# 0.03fF
C13288 VN.n12018 a_400_62400# 0.16fF
C13289 VN.n12019 a_400_62400# 0.19fF
C13290 VN.n12021 a_400_62400# 0.87fF
C13291 VN.n12022 a_400_62400# 0.51fF
C13292 VN.n12023 a_400_62400# 0.59fF
C13293 VN.n12024 a_400_62400# 2.16fF
C13294 VN.n12025 a_400_62400# 0.67fF
C13295 VN.n12026 a_400_62400# 0.62fF
C13296 VN.n12027 a_400_62400# 0.60fF
C13297 VN.n12028 a_400_62400# 2.47fF
C13298 VN.n12029 a_400_62400# 0.16fF
C13299 VN.t621 a_400_62400# 0.03fF
C13300 VN.n12030 a_400_62400# 0.19fF
C13301 VN.t1625 a_400_62400# 0.03fF
C13302 VN.n12032 a_400_62400# 0.32fF
C13303 VN.n12033 a_400_62400# 0.48fF
C13304 VN.n12034 a_400_62400# 0.81fF
C13305 VN.n12035 a_400_62400# 3.34fF
C13306 VN.n12036 a_400_62400# 2.71fF
C13307 VN.t2456 a_400_62400# 0.03fF
C13308 VN.n12037 a_400_62400# 0.32fF
C13309 VN.n12038 a_400_62400# 1.22fF
C13310 VN.n12039 a_400_62400# 0.07fF
C13311 VN.t1303 a_400_62400# 0.03fF
C13312 VN.n12040 a_400_62400# 0.16fF
C13313 VN.n12041 a_400_62400# 0.19fF
C13314 VN.n12043 a_400_62400# 0.24fF
C13315 VN.n12044 a_400_62400# 0.13fF
C13316 VN.n12045 a_400_62400# 1.27fF
C13317 VN.n12046 a_400_62400# 0.62fF
C13318 VN.n12047 a_400_62400# 0.28fF
C13319 VN.n12048 a_400_62400# 0.48fF
C13320 VN.n12049 a_400_62400# 0.71fF
C13321 VN.n12050 a_400_62400# 3.52fF
C13322 VN.n12051 a_400_62400# 2.00fF
C13323 VN.n12052 a_400_62400# 0.16fF
C13324 VN.t2272 a_400_62400# 0.03fF
C13325 VN.n12053 a_400_62400# 0.19fF
C13326 VN.t867 a_400_62400# 0.03fF
C13327 VN.n12055 a_400_62400# 0.32fF
C13328 VN.n12056 a_400_62400# 0.48fF
C13329 VN.n12057 a_400_62400# 0.81fF
C13330 VN.n12058 a_400_62400# 3.32fF
C13331 VN.n12059 a_400_62400# 2.63fF
C13332 VN.t1710 a_400_62400# 0.03fF
C13333 VN.n12060 a_400_62400# 0.32fF
C13334 VN.n12061 a_400_62400# 1.22fF
C13335 VN.n12062 a_400_62400# 0.07fF
C13336 VN.t439 a_400_62400# 0.03fF
C13337 VN.n12063 a_400_62400# 0.16fF
C13338 VN.n12064 a_400_62400# 0.19fF
C13339 VN.n12066 a_400_62400# 1.53fF
C13340 VN.n12067 a_400_62400# 3.17fF
C13341 VN.n12068 a_400_62400# 2.47fF
C13342 VN.n12069 a_400_62400# 0.16fF
C13343 VN.t1245 a_400_62400# 0.03fF
C13344 VN.n12070 a_400_62400# 0.19fF
C13345 VN.t2387 a_400_62400# 0.03fF
C13346 VN.n12072 a_400_62400# 0.32fF
C13347 VN.n12073 a_400_62400# 0.48fF
C13348 VN.n12074 a_400_62400# 0.81fF
C13349 VN.n12075 a_400_62400# 0.47fF
C13350 VN.n12076 a_400_62400# 0.54fF
C13351 VN.n12077 a_400_62400# 0.89fF
C13352 VN.n12078 a_400_62400# 0.73fF
C13353 VN.n12079 a_400_62400# 0.44fF
C13354 VN.n12080 a_400_62400# 1.44fF
C13355 VN.n12081 a_400_62400# 2.85fF
C13356 VN.t2297 a_400_62400# 0.03fF
C13357 VN.n12082 a_400_62400# 0.32fF
C13358 VN.n12083 a_400_62400# 1.22fF
C13359 VN.n12084 a_400_62400# 0.07fF
C13360 VN.t2084 a_400_62400# 0.03fF
C13361 VN.n12085 a_400_62400# 0.16fF
C13362 VN.n12086 a_400_62400# 0.19fF
C13363 VN.n12088 a_400_62400# 0.04fF
C13364 VN.n12089 a_400_62400# 0.04fF
C13365 VN.n12090 a_400_62400# 0.14fF
C13366 VN.n12091 a_400_62400# 0.48fF
C13367 VN.n12092 a_400_62400# 0.50fF
C13368 VN.n12093 a_400_62400# 0.14fF
C13369 VN.n12094 a_400_62400# 0.16fF
C13370 VN.n12095 a_400_62400# 0.04fF
C13371 VN.n12096 a_400_62400# 0.09fF
C13372 VN.n12097 a_400_62400# 1.88fF
C13373 VN.n12098 a_400_62400# 0.06fF
C13374 VN.n12099 a_400_62400# 0.65fF
C13375 VN.n12100 a_400_62400# 0.51fF
C13376 VN.n12101 a_400_62400# 3.52fF
C13377 VN.n12102 a_400_62400# 2.00fF
C13378 VN.n12103 a_400_62400# 0.16fF
C13379 VN.t378 a_400_62400# 0.03fF
C13380 VN.n12104 a_400_62400# 0.19fF
C13381 VN.t1518 a_400_62400# 0.03fF
C13382 VN.n12106 a_400_62400# 0.32fF
C13383 VN.n12107 a_400_62400# 0.48fF
C13384 VN.n12108 a_400_62400# 0.81fF
C13385 VN.n12109 a_400_62400# 0.47fF
C13386 VN.n12110 a_400_62400# 0.72fF
C13387 VN.n12111 a_400_62400# 0.51fF
C13388 VN.n12112 a_400_62400# 0.24fF
C13389 VN.n12113 a_400_62400# 0.34fF
C13390 VN.n12114 a_400_62400# 0.12fF
C13391 VN.n12115 a_400_62400# 2.63fF
C13392 VN.t1426 a_400_62400# 0.03fF
C13393 VN.n12116 a_400_62400# 0.32fF
C13394 VN.n12117 a_400_62400# 1.22fF
C13395 VN.n12118 a_400_62400# 0.07fF
C13396 VN.t1031 a_400_62400# 0.03fF
C13397 VN.n12119 a_400_62400# 0.16fF
C13398 VN.n12120 a_400_62400# 0.19fF
C13399 VN.n12122 a_400_62400# 3.52fF
C13400 VN.n12123 a_400_62400# 2.01fF
C13401 VN.n12124 a_400_62400# 0.33fF
C13402 VN.n12125 a_400_62400# 0.12fF
C13403 VN.n12126 a_400_62400# 0.28fF
C13404 VN.n12127 a_400_62400# 2.32fF
C13405 VN.n12128 a_400_62400# 0.59fF
C13406 VN.n12129 a_400_62400# 0.16fF
C13407 VN.t2032 a_400_62400# 0.03fF
C13408 VN.n12130 a_400_62400# 0.19fF
C13409 VN.t651 a_400_62400# 0.03fF
C13410 VN.n12132 a_400_62400# 0.32fF
C13411 VN.n12133 a_400_62400# 0.48fF
C13412 VN.n12134 a_400_62400# 0.81fF
C13413 VN.n12135 a_400_62400# 1.11fF
C13414 VN.n12136 a_400_62400# 0.42fF
C13415 VN.n12137 a_400_62400# 0.39fF
C13416 VN.n12138 a_400_62400# 0.34fF
C13417 VN.n12139 a_400_62400# 0.29fF
C13418 VN.n12140 a_400_62400# 0.81fF
C13419 VN.n12141 a_400_62400# 0.37fF
C13420 VN.n12142 a_400_62400# 0.19fF
C13421 VN.n12143 a_400_62400# 2.33fF
C13422 VN.n12144 a_400_62400# 2.59fF
C13423 VN.t561 a_400_62400# 0.03fF
C13424 VN.n12145 a_400_62400# 0.32fF
C13425 VN.n12146 a_400_62400# 1.22fF
C13426 VN.n12147 a_400_62400# 0.07fF
C13427 VN.t161 a_400_62400# 0.03fF
C13428 VN.n12148 a_400_62400# 0.16fF
C13429 VN.n12149 a_400_62400# 0.19fF
C13430 VN.n12151 a_400_62400# 2.47fF
C13431 VN.n12152 a_400_62400# 3.34fF
C13432 VN.t2310 a_400_62400# 0.03fF
C13433 VN.n12153 a_400_62400# 0.32fF
C13434 VN.n12154 a_400_62400# 0.48fF
C13435 VN.n12155 a_400_62400# 0.81fF
C13436 VN.n12156 a_400_62400# 0.16fF
C13437 VN.t1158 a_400_62400# 0.03fF
C13438 VN.n12157 a_400_62400# 0.19fF
C13439 VN.n12159 a_400_62400# 0.91fF
C13440 VN.n12160 a_400_62400# 0.37fF
C13441 VN.n12161 a_400_62400# 2.33fF
C13442 VN.n12162 a_400_62400# 0.28fF
C13443 VN.n12163 a_400_62400# 0.25fF
C13444 VN.n12164 a_400_62400# 0.13fF
C13445 VN.n12165 a_400_62400# 2.49fF
C13446 VN.t2221 a_400_62400# 0.03fF
C13447 VN.n12166 a_400_62400# 0.32fF
C13448 VN.n12167 a_400_62400# 1.22fF
C13449 VN.n12168 a_400_62400# 0.07fF
C13450 VN.t1825 a_400_62400# 0.03fF
C13451 VN.n12169 a_400_62400# 0.16fF
C13452 VN.n12170 a_400_62400# 0.19fF
C13453 VN.t43 a_400_62400# 32.18fF
C13454 VN.n12172 a_400_62400# 27.83fF
C13455 VN.t160 a_400_62400# 64.17fF
C13456 VN.t1355 a_400_62400# 0.03fF
C13457 VN.n12173 a_400_62400# 1.60fF
C13458 VN.n12174 a_400_62400# 0.07fF
C13459 VN.t1091 a_400_62400# 0.03fF
C13460 VN.n12175 a_400_62400# 0.02fF
C13461 VN.n12176 a_400_62400# 0.34fF
C13462 VN.n12178 a_400_62400# 1.62fF
C13463 VN.n12179 a_400_62400# 0.49fF
C13464 VN.n12180 a_400_62400# 1.58fF
C13465 VN.n12181 a_400_62400# 0.51fF
C13466 VN.n12182 a_400_62400# 5.67fF
C13467 VN.n12183 a_400_62400# 70.60fF
C13468 VN.n12184 a_400_62400# 42.32fF
C13469 VN.n12185 a_400_62400# 42.32fF
C13470 VN.n12186 a_400_62400# 42.32fF
C13471 VN.n12187 a_400_62400# 42.32fF
C13472 VN.n12188 a_400_62400# 42.32fF
C13473 VN.n12189 a_400_62400# 42.32fF
C13474 VN.n12190 a_400_62400# 42.32fF
C13475 VN.n12191 a_400_62400# 42.32fF
C13476 VN.n12192 a_400_62400# 42.32fF
C13477 VN.n12193 a_400_62400# 42.32fF
C13478 VN.n12194 a_400_62400# 42.32fF
C13479 VN.n12195 a_400_62400# 42.32fF
C13480 VN.n12196 a_400_62400# 42.32fF
C13481 VN.n12197 a_400_62400# 42.32fF
C13482 VN.n12198 a_400_62400# 42.32fF
C13483 VN.n12199 a_400_62400# 134.35fF
C13484 VN.n12200 a_400_62400# 145.11fF
C13485 VN.n12201 a_400_62400# 37.96fF
C13486 VN.n12202 a_400_62400# 37.88fF
C13487 VN.n12203 a_400_62400# 37.88fF
C13488 VN.n12204 a_400_62400# 37.88fF
C13489 VN.n12205 a_400_62400# 37.88fF
C13490 VN.n12206 a_400_62400# 37.88fF
C13491 VN.n12207 a_400_62400# 37.88fF
C13492 VN.n12208 a_400_62400# 37.88fF
C13493 VN.n12209 a_400_62400# 37.88fF
C13494 VN.n12210 a_400_62400# 37.88fF
C13495 VN.n12211 a_400_62400# 37.88fF
C13496 VN.n12212 a_400_62400# 37.88fF
C13497 VN.n12213 a_400_62400# 37.88fF
C13498 VN.n12214 a_400_62400# 37.88fF
C13499 VN.n12215 a_400_62400# 37.88fF
C13500 VN.n12216 a_400_62400# 3.75fF
C13501 VN.t1439 a_400_62400# 0.03fF
C13502 VN.n12217 a_400_62400# 0.32fF
C13503 VN.n12218 a_400_62400# 1.22fF
C13504 VN.n12219 a_400_62400# 0.07fF
C13505 VN.n12220 a_400_62400# 0.33fF
C13506 VN.n12221 a_400_62400# 0.12fF
C13507 VN.n12222 a_400_62400# 0.27fF
C13508 VN.n12223 a_400_62400# 1.04fF
C13509 VN.n12224 a_400_62400# 2.59fF
C13510 VN.n12225 a_400_62400# 2.51fF
C13511 VN.n12226 a_400_62400# 0.16fF
C13512 VN.t1246 a_400_62400# 0.03fF
C13513 VN.n12227 a_400_62400# 0.19fF
C13514 VN.t2390 a_400_62400# 0.03fF
C13515 VN.n12229 a_400_62400# 0.32fF
C13516 VN.n12230 a_400_62400# 0.48fF
C13517 VN.n12231 a_400_62400# 0.81fF
C13518 VN.n12232 a_400_62400# 3.56fF
C13519 VN.n12233 a_400_62400# 4.01fF
C13520 VN.t1907 a_400_62400# 0.03fF
C13521 VN.n12234 a_400_62400# 0.16fF
C13522 VN.n12235 a_400_62400# 0.19fF
C13523 VN.n12237 a_400_62400# 27.83fF
C13524 VN.n12238 a_400_62400# 2.36fF
C13525 VN.n12239 a_400_62400# 4.08fF
C13526 VN.t1084 a_400_62400# 0.03fF
C13527 VN.n12240 a_400_62400# 0.32fF
C13528 VN.n12241 a_400_62400# 0.48fF
C13529 VN.n12242 a_400_62400# 0.81fF
C13530 VN.n12243 a_400_62400# 0.16fF
C13531 VN.t2466 a_400_62400# 0.03fF
C13532 VN.n12244 a_400_62400# 0.19fF
C13533 VN.n12246 a_400_62400# 0.24fF
C13534 VN.n12247 a_400_62400# 0.27fF
C13535 VN.n12248 a_400_62400# 0.34fF
C13536 VN.n12249 a_400_62400# 0.12fF
C13537 VN.n12250 a_400_62400# 0.30fF
C13538 VN.n12251 a_400_62400# 0.88fF
C13539 VN.n12252 a_400_62400# 1.21fF
C13540 VN.n12253 a_400_62400# 0.30fF
C13541 VN.n12254 a_400_62400# 0.13fF
C13542 VN.n12255 a_400_62400# 0.28fF
C13543 VN.n12256 a_400_62400# 0.09fF
C13544 VN.n12257 a_400_62400# 0.08fF
C13545 VN.n12258 a_400_62400# 0.09fF
C13546 VN.n12259 a_400_62400# 2.66fF
C13547 VN.t747 a_400_62400# 0.03fF
C13548 VN.n12260 a_400_62400# 0.16fF
C13549 VN.n12261 a_400_62400# 0.19fF
C13550 VN.t2217 a_400_62400# 0.03fF
C13551 VN.n12263 a_400_62400# 0.32fF
C13552 VN.n12264 a_400_62400# 1.22fF
C13553 VN.n12265 a_400_62400# 0.07fF
C13554 VN.n12266 a_400_62400# 2.60fF
C13555 VN.n12267 a_400_62400# 0.16fF
C13556 VN.t716 a_400_62400# 0.03fF
C13557 VN.n12268 a_400_62400# 0.19fF
C13558 VN.t781 a_400_62400# 0.03fF
C13559 VN.n12270 a_400_62400# 0.16fF
C13560 VN.n12271 a_400_62400# 0.19fF
C13561 VN.t1004 a_400_62400# 0.03fF
C13562 VN.n12273 a_400_62400# 0.32fF
C13563 VN.n12274 a_400_62400# 1.22fF
C13564 VN.n12275 a_400_62400# 0.07fF
C13565 VN.t1567 a_400_62400# 0.03fF
C13566 VN.n12276 a_400_62400# 0.32fF
C13567 VN.n12277 a_400_62400# 0.48fF
C13568 VN.n12278 a_400_62400# 0.81fF
C13569 VN.n12279 a_400_62400# 0.40fF
C13570 VN.n12280 a_400_62400# 1.46fF
C13571 VN.n12281 a_400_62400# 0.21fF
C13572 VN.n12282 a_400_62400# 2.81fF
C13573 VN.n12283 a_400_62400# 2.39fF
C13574 VN.n12284 a_400_62400# 2.51fF
C13575 VN.n12285 a_400_62400# 0.16fF
C13576 VN.t102 a_400_62400# 0.03fF
C13577 VN.n12286 a_400_62400# 0.19fF
C13578 VN.t328 a_400_62400# 0.03fF
C13579 VN.n12288 a_400_62400# 0.16fF
C13580 VN.n12289 a_400_62400# 0.19fF
C13581 VN.t454 a_400_62400# 0.03fF
C13582 VN.n12291 a_400_62400# 0.32fF
C13583 VN.n12292 a_400_62400# 1.22fF
C13584 VN.n12293 a_400_62400# 0.07fF
C13585 VN.t1282 a_400_62400# 0.03fF
C13586 VN.n12294 a_400_62400# 0.32fF
C13587 VN.n12295 a_400_62400# 0.48fF
C13588 VN.n12296 a_400_62400# 0.81fF
C13589 VN.n12297 a_400_62400# 1.46fF
C13590 VN.n12298 a_400_62400# 0.21fF
C13591 VN.n12299 a_400_62400# 2.81fF
C13592 VN.n12300 a_400_62400# 3.93fF
C13593 VN.n12301 a_400_62400# 2.51fF
C13594 VN.n12302 a_400_62400# 0.16fF
C13595 VN.t1720 a_400_62400# 0.03fF
C13596 VN.n12303 a_400_62400# 0.19fF
C13597 VN.t211 a_400_62400# 0.03fF
C13598 VN.n12305 a_400_62400# 0.32fF
C13599 VN.n12306 a_400_62400# 0.48fF
C13600 VN.n12307 a_400_62400# 0.81fF
C13601 VN.n12308 a_400_62400# 1.24fF
C13602 VN.n12309 a_400_62400# 0.43fF
C13603 VN.n12310 a_400_62400# 0.43fF
C13604 VN.n12311 a_400_62400# 1.24fF
C13605 VN.n12312 a_400_62400# 1.46fF
C13606 VN.n12313 a_400_62400# 0.21fF
C13607 VN.n12314 a_400_62400# 6.64fF
C13608 VN.t2406 a_400_62400# 0.03fF
C13609 VN.n12315 a_400_62400# 0.16fF
C13610 VN.n12316 a_400_62400# 0.19fF
C13611 VN.t1350 a_400_62400# 0.03fF
C13612 VN.n12318 a_400_62400# 0.32fF
C13613 VN.n12319 a_400_62400# 1.22fF
C13614 VN.n12320 a_400_62400# 0.07fF
C13615 VN.n12321 a_400_62400# 2.51fF
C13616 VN.n12322 a_400_62400# 3.57fF
C13617 VN.t1996 a_400_62400# 0.03fF
C13618 VN.n12323 a_400_62400# 0.32fF
C13619 VN.n12324 a_400_62400# 0.48fF
C13620 VN.n12325 a_400_62400# 0.81fF
C13621 VN.n12326 a_400_62400# 0.16fF
C13622 VN.t847 a_400_62400# 0.03fF
C13623 VN.n12327 a_400_62400# 0.19fF
C13624 VN.n12329 a_400_62400# 2.51fF
C13625 VN.n12330 a_400_62400# 3.57fF
C13626 VN.t414 a_400_62400# 0.03fF
C13627 VN.n12331 a_400_62400# 0.32fF
C13628 VN.n12332 a_400_62400# 0.48fF
C13629 VN.n12333 a_400_62400# 0.81fF
C13630 VN.t2102 a_400_62400# 0.03fF
C13631 VN.n12334 a_400_62400# 0.32fF
C13632 VN.n12335 a_400_62400# 1.22fF
C13633 VN.n12336 a_400_62400# 0.07fF
C13634 VN.t1974 a_400_62400# 0.03fF
C13635 VN.n12337 a_400_62400# 0.16fF
C13636 VN.n12338 a_400_62400# 0.19fF
C13637 VN.n12340 a_400_62400# 0.16fF
C13638 VN.t1773 a_400_62400# 0.03fF
C13639 VN.n12341 a_400_62400# 0.19fF
C13640 VN.n12343 a_400_62400# 3.08fF
C13641 VN.n12344 a_400_62400# 3.93fF
C13642 VN.n12345 a_400_62400# 2.60fF
C13643 VN.n12346 a_400_62400# 3.40fF
C13644 VN.t697 a_400_62400# 0.03fF
C13645 VN.n12347 a_400_62400# 0.32fF
C13646 VN.n12348 a_400_62400# 0.48fF
C13647 VN.n12349 a_400_62400# 0.81fF
C13648 VN.t2428 a_400_62400# 0.03fF
C13649 VN.n12350 a_400_62400# 1.63fF
C13650 VN.n12351 a_400_62400# 2.62fF
C13651 VN.n12352 a_400_62400# 0.08fF
C13652 VN.n12353 a_400_62400# 0.13fF
C13653 VN.n12354 a_400_62400# 0.81fF
C13654 VN.n12355 a_400_62400# 1.54fF
C13655 VN.n12356 a_400_62400# 4.06fF
C13656 VN.n12357 a_400_62400# 1.13fF
C13657 VN.n12358 a_400_62400# 0.02fF
C13658 VN.n12359 a_400_62400# 1.30fF
C13659 VN.t178 a_400_62400# 28.64fF
C13660 VN.n12360 a_400_62400# 27.84fF
C13661 VN.n12362 a_400_62400# 0.50fF
C13662 VN.n12363 a_400_62400# 1.93fF
C13663 VN.n12364 a_400_62400# 3.88fF
C13664 VN.n12365 a_400_62400# 3.24fF
C13665 VN.n12366 a_400_62400# 5.16fF
C13666 VN.n12367 a_400_62400# 0.34fF
C13667 VN.n12368 a_400_62400# 0.02fF
C13668 VN.t1581 a_400_62400# 0.03fF
C13669 VN.n12369 a_400_62400# 0.34fF
C13670 VN.t1874 a_400_62400# 0.03fF
C13671 VN.n12370 a_400_62400# 1.28fF
C13672 VN.n12371 a_400_62400# 0.94fF
C13673 VN.n12372 a_400_62400# 0.34fF
C13674 VN.n12373 a_400_62400# 0.16fF
C13675 VN.n12374 a_400_62400# 0.07fF
C13676 VN.n12375 a_400_62400# 0.23fF
C13677 VN.n12376 a_400_62400# 1.68fF
C13678 VN.n12377 a_400_62400# 3.71fF
C13679 VN.n12378 a_400_62400# 0.16fF
C13680 VN.t83 a_400_62400# 0.03fF
C13681 VN.n12379 a_400_62400# 0.19fF
C13682 VN.t2138 a_400_62400# 0.03fF
C13683 VN.n12381 a_400_62400# 0.32fF
C13684 VN.n12382 a_400_62400# 0.48fF
C13685 VN.n12383 a_400_62400# 0.81fF
C13686 VN.n12384 a_400_62400# 3.54fF
C13687 VN.n12385 a_400_62400# 2.75fF
C13688 VN.t550 a_400_62400# 0.03fF
C13689 VN.n12386 a_400_62400# 0.32fF
C13690 VN.n12387 a_400_62400# 1.22fF
C13691 VN.n12388 a_400_62400# 0.07fF
C13692 VN.t316 a_400_62400# 0.03fF
C13693 VN.n12389 a_400_62400# 0.16fF
C13694 VN.n12390 a_400_62400# 0.19fF
C13695 VN.n12392 a_400_62400# 3.45fF
C13696 VN.n12393 a_400_62400# 2.50fF
C13697 VN.n12394 a_400_62400# 0.07fF
C13698 VN.n12395 a_400_62400# 0.18fF
C13699 VN.n12396 a_400_62400# 1.67fF
C13700 VN.n12397 a_400_62400# 0.34fF
C13701 VN.n12398 a_400_62400# 0.16fF
C13702 VN.n12399 a_400_62400# 0.32fF
C13703 VN.t1265 a_400_62400# 0.03fF
C13704 VN.n12400 a_400_62400# 0.48fF
C13705 VN.n12401 a_400_62400# 0.81fF
C13706 VN.n12402 a_400_62400# 0.32fF
C13707 VN.t2207 a_400_62400# 0.03fF
C13708 VN.n12403 a_400_62400# 1.18fF
C13709 VN.n12404 a_400_62400# 0.11fF
C13710 VN.n12405 a_400_62400# 2.64fF
C13711 VN.n12406 a_400_62400# 0.16fF
C13712 VN.t1891 a_400_62400# 0.03fF
C13713 VN.n12407 a_400_62400# 0.19fF
C13714 VN.t1965 a_400_62400# 0.03fF
C13715 VN.n12409 a_400_62400# 0.16fF
C13716 VN.n12410 a_400_62400# 0.19fF
C13717 VN.n12412 a_400_62400# 27.83fF
C13718 VN.n12413 a_400_62400# 2.60fF
C13719 VN.n12414 a_400_62400# 3.40fF
C13720 VN.t2356 a_400_62400# 0.03fF
C13721 VN.n12415 a_400_62400# 0.32fF
C13722 VN.n12416 a_400_62400# 0.48fF
C13723 VN.n12417 a_400_62400# 0.81fF
C13724 VN.n12418 a_400_62400# 0.16fF
C13725 VN.t1502 a_400_62400# 0.03fF
C13726 VN.n12419 a_400_62400# 0.19fF
C13727 VN.n12421 a_400_62400# 3.23fF
C13728 VN.n12422 a_400_62400# 3.08fF
C13729 VN.t1684 a_400_62400# 0.03fF
C13730 VN.n12423 a_400_62400# 0.16fF
C13731 VN.n12424 a_400_62400# 0.19fF
C13732 VN.t1795 a_400_62400# 0.03fF
C13733 VN.n12426 a_400_62400# 0.32fF
C13734 VN.n12427 a_400_62400# 1.22fF
C13735 VN.n12428 a_400_62400# 0.07fF
C13736 VN.n12429 a_400_62400# 2.60fF
C13737 VN.n12430 a_400_62400# 3.40fF
C13738 VN.t1488 a_400_62400# 0.03fF
C13739 VN.n12431 a_400_62400# 0.32fF
C13740 VN.n12432 a_400_62400# 0.48fF
C13741 VN.n12433 a_400_62400# 0.81fF
C13742 VN.n12434 a_400_62400# 0.16fF
C13743 VN.t635 a_400_62400# 0.03fF
C13744 VN.n12435 a_400_62400# 0.19fF
C13745 VN.n12437 a_400_62400# 3.23fF
C13746 VN.n12438 a_400_62400# 3.08fF
C13747 VN.t818 a_400_62400# 0.03fF
C13748 VN.n12439 a_400_62400# 0.16fF
C13749 VN.n12440 a_400_62400# 0.19fF
C13750 VN.t920 a_400_62400# 0.03fF
C13751 VN.n12442 a_400_62400# 0.32fF
C13752 VN.n12443 a_400_62400# 1.22fF
C13753 VN.n12444 a_400_62400# 0.07fF
C13754 VN.n12445 a_400_62400# 2.60fF
C13755 VN.n12446 a_400_62400# 3.40fF
C13756 VN.t1960 a_400_62400# 0.03fF
C13757 VN.n12447 a_400_62400# 0.32fF
C13758 VN.n12448 a_400_62400# 0.48fF
C13759 VN.n12449 a_400_62400# 0.81fF
C13760 VN.n12450 a_400_62400# 0.16fF
C13761 VN.t1106 a_400_62400# 0.03fF
C13762 VN.n12451 a_400_62400# 0.19fF
C13763 VN.n12453 a_400_62400# 3.23fF
C13764 VN.n12454 a_400_62400# 3.08fF
C13765 VN.t1320 a_400_62400# 0.03fF
C13766 VN.n12455 a_400_62400# 0.16fF
C13767 VN.n12456 a_400_62400# 0.19fF
C13768 VN.t1419 a_400_62400# 0.03fF
C13769 VN.n12458 a_400_62400# 0.32fF
C13770 VN.n12459 a_400_62400# 1.22fF
C13771 VN.n12460 a_400_62400# 0.07fF
C13772 VN.n12461 a_400_62400# 2.60fF
C13773 VN.n12462 a_400_62400# 3.40fF
C13774 VN.t1092 a_400_62400# 0.03fF
C13775 VN.n12463 a_400_62400# 0.32fF
C13776 VN.n12464 a_400_62400# 0.48fF
C13777 VN.n12465 a_400_62400# 0.81fF
C13778 VN.n12466 a_400_62400# 0.16fF
C13779 VN.t239 a_400_62400# 0.03fF
C13780 VN.n12467 a_400_62400# 0.19fF
C13781 VN.n12469 a_400_62400# 3.23fF
C13782 VN.n12470 a_400_62400# 3.08fF
C13783 VN.t457 a_400_62400# 0.03fF
C13784 VN.n12471 a_400_62400# 0.16fF
C13785 VN.n12472 a_400_62400# 0.19fF
C13786 VN.t555 a_400_62400# 0.03fF
C13787 VN.n12474 a_400_62400# 0.32fF
C13788 VN.n12475 a_400_62400# 1.22fF
C13789 VN.n12476 a_400_62400# 0.07fF
C13790 VN.n12477 a_400_62400# 2.60fF
C13791 VN.n12478 a_400_62400# 3.40fF
C13792 VN.t222 a_400_62400# 0.03fF
C13793 VN.n12479 a_400_62400# 0.32fF
C13794 VN.n12480 a_400_62400# 0.48fF
C13795 VN.n12481 a_400_62400# 0.81fF
C13796 VN.n12482 a_400_62400# 0.16fF
C13797 VN.t2028 a_400_62400# 0.03fF
C13798 VN.n12483 a_400_62400# 0.19fF
C13799 VN.n12485 a_400_62400# 3.23fF
C13800 VN.n12486 a_400_62400# 3.08fF
C13801 VN.t2105 a_400_62400# 0.03fF
C13802 VN.n12487 a_400_62400# 0.16fF
C13803 VN.n12488 a_400_62400# 0.19fF
C13804 VN.t2213 a_400_62400# 0.03fF
C13805 VN.n12490 a_400_62400# 0.32fF
C13806 VN.n12491 a_400_62400# 1.22fF
C13807 VN.n12492 a_400_62400# 0.07fF
C13808 VN.n12493 a_400_62400# 2.60fF
C13809 VN.n12494 a_400_62400# 3.40fF
C13810 VN.t2010 a_400_62400# 0.03fF
C13811 VN.n12495 a_400_62400# 0.32fF
C13812 VN.n12496 a_400_62400# 0.48fF
C13813 VN.n12497 a_400_62400# 0.81fF
C13814 VN.n12498 a_400_62400# 0.16fF
C13815 VN.t1153 a_400_62400# 0.03fF
C13816 VN.n12499 a_400_62400# 0.19fF
C13817 VN.n12501 a_400_62400# 3.23fF
C13818 VN.n12502 a_400_62400# 3.08fF
C13819 VN.t1228 a_400_62400# 0.03fF
C13820 VN.n12503 a_400_62400# 0.16fF
C13821 VN.n12504 a_400_62400# 0.19fF
C13822 VN.t1466 a_400_62400# 0.03fF
C13823 VN.n12506 a_400_62400# 0.32fF
C13824 VN.n12507 a_400_62400# 1.22fF
C13825 VN.n12508 a_400_62400# 0.07fF
C13826 VN.n12509 a_400_62400# 2.60fF
C13827 VN.n12510 a_400_62400# 3.40fF
C13828 VN.t1137 a_400_62400# 0.03fF
C13829 VN.n12511 a_400_62400# 0.32fF
C13830 VN.n12512 a_400_62400# 0.48fF
C13831 VN.n12513 a_400_62400# 0.81fF
C13832 VN.n12514 a_400_62400# 0.16fF
C13833 VN.t286 a_400_62400# 0.03fF
C13834 VN.n12515 a_400_62400# 0.19fF
C13835 VN.n12517 a_400_62400# 3.23fF
C13836 VN.n12518 a_400_62400# 3.08fF
C13837 VN.t362 a_400_62400# 0.03fF
C13838 VN.n12519 a_400_62400# 0.16fF
C13839 VN.n12520 a_400_62400# 0.19fF
C13840 VN.t595 a_400_62400# 0.03fF
C13841 VN.n12522 a_400_62400# 0.32fF
C13842 VN.n12523 a_400_62400# 1.22fF
C13843 VN.n12524 a_400_62400# 0.07fF
C13844 VN.n12525 a_400_62400# 2.60fF
C13845 VN.n12526 a_400_62400# 3.40fF
C13846 VN.t274 a_400_62400# 0.03fF
C13847 VN.n12527 a_400_62400# 0.32fF
C13848 VN.n12528 a_400_62400# 0.48fF
C13849 VN.n12529 a_400_62400# 0.81fF
C13850 VN.n12530 a_400_62400# 0.16fF
C13851 VN.t1938 a_400_62400# 0.03fF
C13852 VN.n12531 a_400_62400# 0.19fF
C13853 VN.n12533 a_400_62400# 3.23fF
C13854 VN.n12534 a_400_62400# 3.08fF
C13855 VN.t2012 a_400_62400# 0.03fF
C13856 VN.n12535 a_400_62400# 0.16fF
C13857 VN.n12536 a_400_62400# 0.19fF
C13858 VN.t2250 a_400_62400# 0.03fF
C13859 VN.n12538 a_400_62400# 0.32fF
C13860 VN.n12539 a_400_62400# 1.22fF
C13861 VN.n12540 a_400_62400# 0.07fF
C13862 VN.n12541 a_400_62400# 2.60fF
C13863 VN.n12542 a_400_62400# 3.40fF
C13864 VN.t1924 a_400_62400# 0.03fF
C13865 VN.n12543 a_400_62400# 0.32fF
C13866 VN.n12544 a_400_62400# 0.48fF
C13867 VN.n12545 a_400_62400# 0.81fF
C13868 VN.n12546 a_400_62400# 0.16fF
C13869 VN.t1065 a_400_62400# 0.03fF
C13870 VN.n12547 a_400_62400# 0.19fF
C13871 VN.n12549 a_400_62400# 3.23fF
C13872 VN.n12550 a_400_62400# 3.08fF
C13873 VN.t1139 a_400_62400# 0.03fF
C13874 VN.n12551 a_400_62400# 0.16fF
C13875 VN.n12552 a_400_62400# 0.19fF
C13876 VN.t1389 a_400_62400# 0.03fF
C13877 VN.n12554 a_400_62400# 0.32fF
C13878 VN.n12555 a_400_62400# 1.22fF
C13879 VN.n12556 a_400_62400# 0.07fF
C13880 VN.n12557 a_400_62400# 2.60fF
C13881 VN.n12558 a_400_62400# 3.40fF
C13882 VN.t1049 a_400_62400# 0.03fF
C13883 VN.n12559 a_400_62400# 0.32fF
C13884 VN.n12560 a_400_62400# 0.48fF
C13885 VN.n12561 a_400_62400# 0.81fF
C13886 VN.n12562 a_400_62400# 0.16fF
C13887 VN.t190 a_400_62400# 0.03fF
C13888 VN.n12563 a_400_62400# 0.19fF
C13889 VN.n12565 a_400_62400# 3.23fF
C13890 VN.n12566 a_400_62400# 3.08fF
C13891 VN.t409 a_400_62400# 0.03fF
C13892 VN.n12567 a_400_62400# 0.16fF
C13893 VN.n12568 a_400_62400# 0.19fF
C13894 VN.t523 a_400_62400# 0.03fF
C13895 VN.n12570 a_400_62400# 0.32fF
C13896 VN.n12571 a_400_62400# 1.22fF
C13897 VN.n12572 a_400_62400# 0.07fF
C13898 VN.n12573 a_400_62400# 2.60fF
C13899 VN.n12574 a_400_62400# 3.40fF
C13900 VN.t179 a_400_62400# 0.03fF
C13901 VN.n12575 a_400_62400# 0.32fF
C13902 VN.n12576 a_400_62400# 0.48fF
C13903 VN.n12577 a_400_62400# 0.81fF
C13904 VN.n12578 a_400_62400# 0.16fF
C13905 VN.t1848 a_400_62400# 0.03fF
C13906 VN.n12579 a_400_62400# 0.19fF
C13907 VN.n12581 a_400_62400# 3.23fF
C13908 VN.n12582 a_400_62400# 3.08fF
C13909 VN.t2058 a_400_62400# 0.03fF
C13910 VN.n12583 a_400_62400# 0.16fF
C13911 VN.n12584 a_400_62400# 0.19fF
C13912 VN.t2177 a_400_62400# 0.03fF
C13913 VN.n12586 a_400_62400# 0.32fF
C13914 VN.n12587 a_400_62400# 1.22fF
C13915 VN.n12588 a_400_62400# 0.07fF
C13916 VN.n12589 a_400_62400# 2.60fF
C13917 VN.n12590 a_400_62400# 3.40fF
C13918 VN.t1353 a_400_62400# 0.03fF
C13919 VN.n12591 a_400_62400# 0.32fF
C13920 VN.n12592 a_400_62400# 0.48fF
C13921 VN.n12593 a_400_62400# 0.81fF
C13922 VN.n12594 a_400_62400# 0.16fF
C13923 VN.t1847 a_400_62400# 0.03fF
C13924 VN.n12595 a_400_62400# 0.19fF
C13925 VN.n12597 a_400_62400# 3.23fF
C13926 VN.n12598 a_400_62400# 3.08fF
C13927 VN.t2055 a_400_62400# 0.03fF
C13928 VN.n12599 a_400_62400# 0.16fF
C13929 VN.n12600 a_400_62400# 0.19fF
C13930 VN.t2280 a_400_62400# 0.03fF
C13931 VN.n12602 a_400_62400# 0.32fF
C13932 VN.n12603 a_400_62400# 1.22fF
C13933 VN.n12604 a_400_62400# 0.07fF
C13934 VN.n12605 a_400_62400# 3.22fF
C13935 VN.n12606 a_400_62400# 2.65fF
C13936 VN.n12607 a_400_62400# 0.16fF
C13937 VN.t975 a_400_62400# 0.03fF
C13938 VN.n12608 a_400_62400# 0.19fF
C13939 VN.t485 a_400_62400# 0.03fF
C13940 VN.n12610 a_400_62400# 0.32fF
C13941 VN.n12611 a_400_62400# 0.48fF
C13942 VN.n12612 a_400_62400# 0.81fF
C13943 VN.n12613 a_400_62400# 3.42fF
C13944 VN.n12614 a_400_62400# 3.09fF
C13945 VN.t1187 a_400_62400# 0.03fF
C13946 VN.n12615 a_400_62400# 0.16fF
C13947 VN.n12616 a_400_62400# 0.19fF
C13948 VN.t1410 a_400_62400# 0.03fF
C13949 VN.n12618 a_400_62400# 0.32fF
C13950 VN.n12619 a_400_62400# 1.22fF
C13951 VN.n12620 a_400_62400# 0.07fF
C13952 VN.t82 a_400_62400# 64.69fF
C13953 VN.t130 a_400_62400# 0.03fF
C13954 VN.n12621 a_400_62400# 0.32fF
C13955 VN.n12622 a_400_62400# 1.22fF
C13956 VN.n12623 a_400_62400# 0.07fF
C13957 VN.t2552 a_400_62400# 0.03fF
C13958 VN.n12624 a_400_62400# 0.16fF
C13959 VN.n12625 a_400_62400# 0.19fF
C13960 VN.n12627 a_400_62400# 0.16fF
C13961 VN.t2371 a_400_62400# 0.03fF
C13962 VN.n12628 a_400_62400# 0.19fF
C13963 VN.n12630 a_400_62400# 3.08fF
C13964 VN.n12631 a_400_62400# 2.37fF
C13965 VN.n12632 a_400_62400# 6.91fF
C13966 VN.t1539 a_400_62400# 0.03fF
C13967 VN.n12633 a_400_62400# 0.16fF
C13968 VN.n12634 a_400_62400# 0.19fF
C13969 VN.t601 a_400_62400# 0.03fF
C13970 VN.n12636 a_400_62400# 0.32fF
C13971 VN.n12637 a_400_62400# 1.22fF
C13972 VN.n12638 a_400_62400# 0.07fF
C13973 VN.n12639 a_400_62400# 2.51fF
C13974 VN.n12640 a_400_62400# 3.57fF
C13975 VN.t1124 a_400_62400# 0.03fF
C13976 VN.n12641 a_400_62400# 0.32fF
C13977 VN.n12642 a_400_62400# 0.48fF
C13978 VN.n12643 a_400_62400# 0.81fF
C13979 VN.n12644 a_400_62400# 0.16fF
C13980 VN.t2512 a_400_62400# 0.03fF
C13981 VN.n12645 a_400_62400# 0.19fF
C13982 VN.n12647 a_400_62400# 2.51fF
C13983 VN.n12648 a_400_62400# 3.57fF
C13984 VN.t2062 a_400_62400# 0.03fF
C13985 VN.n12649 a_400_62400# 0.32fF
C13986 VN.n12650 a_400_62400# 0.48fF
C13987 VN.n12651 a_400_62400# 0.81fF
C13988 VN.t1225 a_400_62400# 0.03fF
C13989 VN.n12652 a_400_62400# 0.32fF
C13990 VN.n12653 a_400_62400# 1.22fF
C13991 VN.n12654 a_400_62400# 0.07fF
C13992 VN.t1107 a_400_62400# 0.03fF
C13993 VN.n12655 a_400_62400# 0.16fF
C13994 VN.n12656 a_400_62400# 0.19fF
C13995 VN.n12658 a_400_62400# 0.16fF
C13996 VN.t900 a_400_62400# 0.03fF
C13997 VN.n12659 a_400_62400# 0.19fF
C13998 VN.n12661 a_400_62400# 3.08fF
C13999 VN.n12662 a_400_62400# 3.75fF
C14000 VN.n12663 a_400_62400# 6.92fF
C14001 VN.t669 a_400_62400# 0.03fF
C14002 VN.n12664 a_400_62400# 0.16fF
C14003 VN.n12665 a_400_62400# 0.19fF
C14004 VN.t2255 a_400_62400# 0.03fF
C14005 VN.n12667 a_400_62400# 0.32fF
C14006 VN.n12668 a_400_62400# 1.22fF
C14007 VN.n12669 a_400_62400# 0.07fF
C14008 VN.n12670 a_400_62400# 2.51fF
C14009 VN.n12671 a_400_62400# 3.57fF
C14010 VN.t1611 a_400_62400# 0.03fF
C14011 VN.n12672 a_400_62400# 0.32fF
C14012 VN.n12673 a_400_62400# 0.48fF
C14013 VN.n12674 a_400_62400# 0.81fF
C14014 VN.n12675 a_400_62400# 0.16fF
C14015 VN.t489 a_400_62400# 0.03fF
C14016 VN.n12676 a_400_62400# 0.19fF
C14017 VN.n12678 a_400_62400# 2.51fF
C14018 VN.n12679 a_400_62400# 3.57fF
C14019 VN.t2525 a_400_62400# 0.03fF
C14020 VN.n12680 a_400_62400# 0.32fF
C14021 VN.n12681 a_400_62400# 0.48fF
C14022 VN.n12682 a_400_62400# 0.81fF
C14023 VN.t493 a_400_62400# 0.03fF
C14024 VN.n12683 a_400_62400# 1.63fF
C14025 VN.n12684 a_400_62400# 0.08fF
C14026 VN.n12685 a_400_62400# 0.13fF
C14027 VN.n12686 a_400_62400# 0.81fF
C14028 VN.n12687 a_400_62400# 1.21fF
C14029 VN.n12688 a_400_62400# 1.54fF
C14030 VN.n12689 a_400_62400# 4.06fF
C14031 VN.t88 a_400_62400# 28.64fF
C14032 VN.n12690 a_400_62400# 28.43fF
C14033 VN.n12692 a_400_62400# 0.50fF
C14034 VN.n12693 a_400_62400# 0.31fF
C14035 VN.n12694 a_400_62400# 3.88fF
C14036 VN.n12695 a_400_62400# 3.24fF
C14037 VN.n12696 a_400_62400# 3.31fF
C14038 VN.n12697 a_400_62400# 5.74fF
C14039 VN.n12698 a_400_62400# 0.34fF
C14040 VN.n12699 a_400_62400# 0.02fF
C14041 VN.t1856 a_400_62400# 0.03fF
C14042 VN.n12700 a_400_62400# 0.34fF
C14043 VN.t2182 a_400_62400# 0.03fF
C14044 VN.n12701 a_400_62400# 1.28fF
C14045 VN.n12702 a_400_62400# 0.94fF
C14046 VN.n12703 a_400_62400# 2.53fF
C14047 VN.n12704 a_400_62400# 2.51fF
C14048 VN.t2150 a_400_62400# 0.03fF
C14049 VN.n12705 a_400_62400# 0.32fF
C14050 VN.n12706 a_400_62400# 0.48fF
C14051 VN.n12707 a_400_62400# 0.81fF
C14052 VN.n12708 a_400_62400# 0.16fF
C14053 VN.t989 a_400_62400# 0.03fF
C14054 VN.n12709 a_400_62400# 0.19fF
C14055 VN.n12711 a_400_62400# 1.55fF
C14056 VN.n12712 a_400_62400# 0.29fF
C14057 VN.n12713 a_400_62400# 2.52fF
C14058 VN.t1316 a_400_62400# 0.03fF
C14059 VN.n12714 a_400_62400# 0.32fF
C14060 VN.n12715 a_400_62400# 1.22fF
C14061 VN.n12716 a_400_62400# 0.07fF
C14062 VN.t1059 a_400_62400# 0.03fF
C14063 VN.n12717 a_400_62400# 0.16fF
C14064 VN.n12718 a_400_62400# 0.19fF
C14065 VN.n12720 a_400_62400# 2.13fF
C14066 VN.n12721 a_400_62400# 0.96fF
C14067 VN.n12722 a_400_62400# 0.76fF
C14068 VN.n12723 a_400_62400# 0.16fF
C14069 VN.t218 a_400_62400# 0.03fF
C14070 VN.n12724 a_400_62400# 0.19fF
C14071 VN.t1250 a_400_62400# 0.03fF
C14072 VN.n12726 a_400_62400# 0.32fF
C14073 VN.n12727 a_400_62400# 0.48fF
C14074 VN.n12728 a_400_62400# 0.81fF
C14075 VN.n12729 a_400_62400# 0.02fF
C14076 VN.n12730 a_400_62400# 0.09fF
C14077 VN.n12731 a_400_62400# 0.01fF
C14078 VN.n12732 a_400_62400# 0.02fF
C14079 VN.n12733 a_400_62400# 0.02fF
C14080 VN.n12734 a_400_62400# 0.32fF
C14081 VN.n12735 a_400_62400# 1.56fF
C14082 VN.n12736 a_400_62400# 1.81fF
C14083 VN.n12737 a_400_62400# 2.66fF
C14084 VN.t526 a_400_62400# 0.03fF
C14085 VN.n12738 a_400_62400# 0.32fF
C14086 VN.n12739 a_400_62400# 1.22fF
C14087 VN.n12740 a_400_62400# 0.07fF
C14088 VN.t289 a_400_62400# 0.03fF
C14089 VN.n12741 a_400_62400# 0.16fF
C14090 VN.n12742 a_400_62400# 0.19fF
C14091 VN.n12744 a_400_62400# 27.83fF
C14092 VN.n12745 a_400_62400# 0.13fF
C14093 VN.n12746 a_400_62400# 0.16fF
C14094 VN.n12747 a_400_62400# 0.24fF
C14095 VN.n12748 a_400_62400# 2.51fF
C14096 VN.n12749 a_400_62400# 0.16fF
C14097 VN.t949 a_400_62400# 0.03fF
C14098 VN.n12750 a_400_62400# 0.19fF
C14099 VN.t2126 a_400_62400# 0.03fF
C14100 VN.n12752 a_400_62400# 0.32fF
C14101 VN.n12753 a_400_62400# 0.48fF
C14102 VN.n12754 a_400_62400# 0.81fF
C14103 VN.n12755 a_400_62400# 3.56fF
C14104 VN.n12756 a_400_62400# 4.39fF
C14105 VN.t1157 a_400_62400# 0.03fF
C14106 VN.n12757 a_400_62400# 0.16fF
C14107 VN.n12758 a_400_62400# 0.19fF
C14108 VN.t1391 a_400_62400# 0.03fF
C14109 VN.n12760 a_400_62400# 0.32fF
C14110 VN.n12761 a_400_62400# 1.22fF
C14111 VN.n12762 a_400_62400# 0.07fF
C14112 VN.t101 a_400_62400# 64.69fF
C14113 VN.t1691 a_400_62400# 0.03fF
C14114 VN.n12763 a_400_62400# 0.32fF
C14115 VN.n12764 a_400_62400# 1.22fF
C14116 VN.n12765 a_400_62400# 0.07fF
C14117 VN.t1592 a_400_62400# 0.03fF
C14118 VN.n12766 a_400_62400# 0.16fF
C14119 VN.n12767 a_400_62400# 0.19fF
C14120 VN.n12769 a_400_62400# 0.16fF
C14121 VN.t1402 a_400_62400# 0.03fF
C14122 VN.n12770 a_400_62400# 0.19fF
C14123 VN.n12772 a_400_62400# 3.08fF
C14124 VN.n12773 a_400_62400# 3.75fF
C14125 VN.n12774 a_400_62400# 6.92fF
C14126 VN.t2329 a_400_62400# 0.03fF
C14127 VN.n12775 a_400_62400# 0.16fF
C14128 VN.n12776 a_400_62400# 0.19fF
C14129 VN.t195 a_400_62400# 0.03fF
C14130 VN.n12778 a_400_62400# 0.32fF
C14131 VN.n12779 a_400_62400# 1.22fF
C14132 VN.n12780 a_400_62400# 0.07fF
C14133 VN.n12781 a_400_62400# 2.51fF
C14134 VN.n12782 a_400_62400# 3.57fF
C14135 VN.t744 a_400_62400# 0.03fF
C14136 VN.n12783 a_400_62400# 0.32fF
C14137 VN.n12784 a_400_62400# 0.48fF
C14138 VN.n12785 a_400_62400# 0.81fF
C14139 VN.t1851 a_400_62400# 0.03fF
C14140 VN.n12786 a_400_62400# 0.32fF
C14141 VN.n12787 a_400_62400# 1.22fF
C14142 VN.n12788 a_400_62400# 0.07fF
C14143 VN.n12789 a_400_62400# 0.16fF
C14144 VN.t2143 a_400_62400# 0.03fF
C14145 VN.n12790 a_400_62400# 0.19fF
C14146 VN.n12792 a_400_62400# 2.51fF
C14147 VN.n12793 a_400_62400# 3.57fF
C14148 VN.t1662 a_400_62400# 0.03fF
C14149 VN.n12794 a_400_62400# 0.32fF
C14150 VN.n12795 a_400_62400# 0.48fF
C14151 VN.n12796 a_400_62400# 0.81fF
C14152 VN.t822 a_400_62400# 0.03fF
C14153 VN.n12797 a_400_62400# 0.32fF
C14154 VN.n12798 a_400_62400# 1.22fF
C14155 VN.n12799 a_400_62400# 0.07fF
C14156 VN.t726 a_400_62400# 0.03fF
C14157 VN.n12800 a_400_62400# 0.16fF
C14158 VN.n12801 a_400_62400# 0.19fF
C14159 VN.n12803 a_400_62400# 0.16fF
C14160 VN.t541 a_400_62400# 0.03fF
C14161 VN.n12804 a_400_62400# 0.19fF
C14162 VN.n12806 a_400_62400# 3.08fF
C14163 VN.n12807 a_400_62400# 3.75fF
C14164 VN.n12808 a_400_62400# 6.92fF
C14165 VN.t281 a_400_62400# 0.03fF
C14166 VN.n12809 a_400_62400# 0.16fF
C14167 VN.n12810 a_400_62400# 0.19fF
C14168 VN.n12812 a_400_62400# 2.51fF
C14169 VN.n12813 a_400_62400# 3.57fF
C14170 VN.t2401 a_400_62400# 0.03fF
C14171 VN.n12814 a_400_62400# 0.32fF
C14172 VN.n12815 a_400_62400# 0.48fF
C14173 VN.n12816 a_400_62400# 0.81fF
C14174 VN.t980 a_400_62400# 0.03fF
C14175 VN.n12817 a_400_62400# 0.32fF
C14176 VN.n12818 a_400_62400# 1.22fF
C14177 VN.n12819 a_400_62400# 0.07fF
C14178 VN.n12820 a_400_62400# 0.16fF
C14179 VN.t1271 a_400_62400# 0.03fF
C14180 VN.n12821 a_400_62400# 0.19fF
C14181 VN.n12823 a_400_62400# 2.51fF
C14182 VN.n12824 a_400_62400# 3.57fF
C14183 VN.t794 a_400_62400# 0.03fF
C14184 VN.n12825 a_400_62400# 0.32fF
C14185 VN.n12826 a_400_62400# 0.48fF
C14186 VN.n12827 a_400_62400# 0.81fF
C14187 VN.t2482 a_400_62400# 0.03fF
C14188 VN.n12828 a_400_62400# 0.32fF
C14189 VN.n12829 a_400_62400# 1.22fF
C14190 VN.n12830 a_400_62400# 0.07fF
C14191 VN.t2379 a_400_62400# 0.03fF
C14192 VN.n12831 a_400_62400# 0.16fF
C14193 VN.n12832 a_400_62400# 0.19fF
C14194 VN.n12834 a_400_62400# 0.16fF
C14195 VN.t2314 a_400_62400# 0.03fF
C14196 VN.n12835 a_400_62400# 0.19fF
C14197 VN.n12837 a_400_62400# 3.08fF
C14198 VN.n12838 a_400_62400# 3.75fF
C14199 VN.n12839 a_400_62400# 6.92fF
C14200 VN.t1932 a_400_62400# 0.03fF
C14201 VN.n12840 a_400_62400# 0.16fF
C14202 VN.n12841 a_400_62400# 0.19fF
C14203 VN.n12843 a_400_62400# 2.51fF
C14204 VN.n12844 a_400_62400# 3.57fF
C14205 VN.t1532 a_400_62400# 0.03fF
C14206 VN.n12845 a_400_62400# 0.32fF
C14207 VN.n12846 a_400_62400# 0.48fF
C14208 VN.n12847 a_400_62400# 0.81fF
C14209 VN.n12848 a_400_62400# 0.16fF
C14210 VN.t402 a_400_62400# 0.03fF
C14211 VN.n12849 a_400_62400# 0.19fF
C14212 VN.n12851 a_400_62400# 2.51fF
C14213 VN.n12852 a_400_62400# 3.57fF
C14214 VN.t2568 a_400_62400# 0.03fF
C14215 VN.n12853 a_400_62400# 0.32fF
C14216 VN.n12854 a_400_62400# 0.48fF
C14217 VN.n12855 a_400_62400# 0.81fF
C14218 VN.t1733 a_400_62400# 0.03fF
C14219 VN.n12856 a_400_62400# 0.32fF
C14220 VN.n12857 a_400_62400# 1.22fF
C14221 VN.n12858 a_400_62400# 0.07fF
C14222 VN.t1511 a_400_62400# 0.03fF
C14223 VN.n12859 a_400_62400# 0.16fF
C14224 VN.n12860 a_400_62400# 0.19fF
C14225 VN.n12862 a_400_62400# 0.16fF
C14226 VN.t1444 a_400_62400# 0.03fF
C14227 VN.n12863 a_400_62400# 0.19fF
C14228 VN.n12865 a_400_62400# 3.08fF
C14229 VN.n12866 a_400_62400# 3.75fF
C14230 VN.n12867 a_400_62400# 6.92fF
C14231 VN.t1194 a_400_62400# 0.03fF
C14232 VN.n12868 a_400_62400# 0.16fF
C14233 VN.n12869 a_400_62400# 0.19fF
C14234 VN.t89 a_400_62400# 0.03fF
C14235 VN.n12871 a_400_62400# 0.32fF
C14236 VN.n12872 a_400_62400# 1.22fF
C14237 VN.n12873 a_400_62400# 0.07fF
C14238 VN.n12874 a_400_62400# 2.51fF
C14239 VN.n12875 a_400_62400# 3.57fF
C14240 VN.t661 a_400_62400# 0.03fF
C14241 VN.n12876 a_400_62400# 0.32fF
C14242 VN.n12877 a_400_62400# 0.48fF
C14243 VN.n12878 a_400_62400# 0.81fF
C14244 VN.n12879 a_400_62400# 0.16fF
C14245 VN.t2050 a_400_62400# 0.03fF
C14246 VN.n12880 a_400_62400# 0.19fF
C14247 VN.n12882 a_400_62400# 2.51fF
C14248 VN.n12883 a_400_62400# 3.57fF
C14249 VN.t1697 a_400_62400# 0.03fF
C14250 VN.n12884 a_400_62400# 0.32fF
C14251 VN.n12885 a_400_62400# 0.48fF
C14252 VN.n12886 a_400_62400# 0.81fF
C14253 VN.t858 a_400_62400# 0.03fF
C14254 VN.n12887 a_400_62400# 0.32fF
C14255 VN.n12888 a_400_62400# 1.22fF
C14256 VN.n12889 a_400_62400# 0.07fF
C14257 VN.t642 a_400_62400# 0.03fF
C14258 VN.n12890 a_400_62400# 0.16fF
C14259 VN.n12891 a_400_62400# 0.19fF
C14260 VN.n12893 a_400_62400# 0.16fF
C14261 VN.t575 a_400_62400# 0.03fF
C14262 VN.n12894 a_400_62400# 0.19fF
C14263 VN.n12896 a_400_62400# 3.08fF
C14264 VN.n12897 a_400_62400# 3.75fF
C14265 VN.n12898 a_400_62400# 6.92fF
C14266 VN.t325 a_400_62400# 0.03fF
C14267 VN.n12899 a_400_62400# 0.16fF
C14268 VN.n12900 a_400_62400# 0.19fF
C14269 VN.t1767 a_400_62400# 0.03fF
C14270 VN.n12902 a_400_62400# 0.32fF
C14271 VN.n12903 a_400_62400# 1.22fF
C14272 VN.n12904 a_400_62400# 0.07fF
C14273 VN.n12905 a_400_62400# 2.51fF
C14274 VN.n12906 a_400_62400# 3.57fF
C14275 VN.t2321 a_400_62400# 0.03fF
C14276 VN.n12907 a_400_62400# 0.32fF
C14277 VN.n12908 a_400_62400# 0.48fF
C14278 VN.n12909 a_400_62400# 0.81fF
C14279 VN.n12910 a_400_62400# 0.16fF
C14280 VN.t1181 a_400_62400# 0.03fF
C14281 VN.n12911 a_400_62400# 0.19fF
C14282 VN.n12913 a_400_62400# 2.51fF
C14283 VN.n12914 a_400_62400# 3.57fF
C14284 VN.t827 a_400_62400# 0.03fF
C14285 VN.n12915 a_400_62400# 0.32fF
C14286 VN.n12916 a_400_62400# 0.48fF
C14287 VN.n12917 a_400_62400# 0.81fF
C14288 VN.t2520 a_400_62400# 0.03fF
C14289 VN.n12918 a_400_62400# 0.32fF
C14290 VN.n12919 a_400_62400# 1.22fF
C14291 VN.n12920 a_400_62400# 0.07fF
C14292 VN.t2301 a_400_62400# 0.03fF
C14293 VN.n12921 a_400_62400# 0.16fF
C14294 VN.n12922 a_400_62400# 0.19fF
C14295 VN.n12924 a_400_62400# 0.16fF
C14296 VN.t2233 a_400_62400# 0.03fF
C14297 VN.n12925 a_400_62400# 0.19fF
C14298 VN.n12927 a_400_62400# 3.08fF
C14299 VN.n12928 a_400_62400# 3.75fF
C14300 VN.n12929 a_400_62400# 6.92fF
C14301 VN.t1971 a_400_62400# 0.03fF
C14302 VN.n12930 a_400_62400# 0.16fF
C14303 VN.n12931 a_400_62400# 0.19fF
C14304 VN.t896 a_400_62400# 0.03fF
C14305 VN.n12933 a_400_62400# 0.32fF
C14306 VN.n12934 a_400_62400# 1.22fF
C14307 VN.n12935 a_400_62400# 0.07fF
C14308 VN.n12936 a_400_62400# 2.51fF
C14309 VN.n12937 a_400_62400# 3.57fF
C14310 VN.t1453 a_400_62400# 0.03fF
C14311 VN.n12938 a_400_62400# 0.32fF
C14312 VN.n12939 a_400_62400# 0.48fF
C14313 VN.n12940 a_400_62400# 0.81fF
C14314 VN.n12941 a_400_62400# 0.16fF
C14315 VN.t311 a_400_62400# 0.03fF
C14316 VN.n12942 a_400_62400# 0.19fF
C14317 VN.n12944 a_400_62400# 2.51fF
C14318 VN.n12945 a_400_62400# 3.57fF
C14319 VN.t2492 a_400_62400# 0.03fF
C14320 VN.n12946 a_400_62400# 0.32fF
C14321 VN.n12947 a_400_62400# 0.48fF
C14322 VN.n12948 a_400_62400# 0.81fF
C14323 VN.t1660 a_400_62400# 0.03fF
C14324 VN.n12949 a_400_62400# 0.32fF
C14325 VN.n12950 a_400_62400# 1.22fF
C14326 VN.n12951 a_400_62400# 0.07fF
C14327 VN.t1428 a_400_62400# 0.03fF
C14328 VN.n12952 a_400_62400# 0.16fF
C14329 VN.n12953 a_400_62400# 0.19fF
C14330 VN.n12955 a_400_62400# 0.16fF
C14331 VN.t1369 a_400_62400# 0.03fF
C14332 VN.n12956 a_400_62400# 0.19fF
C14333 VN.n12958 a_400_62400# 3.08fF
C14334 VN.n12959 a_400_62400# 3.75fF
C14335 VN.n12960 a_400_62400# 6.92fF
C14336 VN.t1103 a_400_62400# 0.03fF
C14337 VN.n12961 a_400_62400# 0.16fF
C14338 VN.n12962 a_400_62400# 0.19fF
C14339 VN.t2558 a_400_62400# 0.03fF
C14340 VN.n12964 a_400_62400# 0.32fF
C14341 VN.n12965 a_400_62400# 1.22fF
C14342 VN.n12966 a_400_62400# 0.07fF
C14343 VN.n12967 a_400_62400# 2.51fF
C14344 VN.n12968 a_400_62400# 3.57fF
C14345 VN.t584 a_400_62400# 0.03fF
C14346 VN.n12969 a_400_62400# 0.32fF
C14347 VN.n12970 a_400_62400# 0.48fF
C14348 VN.n12971 a_400_62400# 0.81fF
C14349 VN.n12972 a_400_62400# 0.16fF
C14350 VN.t2100 a_400_62400# 0.03fF
C14351 VN.n12973 a_400_62400# 0.19fF
C14352 VN.n12975 a_400_62400# 2.51fF
C14353 VN.n12976 a_400_62400# 3.57fF
C14354 VN.t1627 a_400_62400# 0.03fF
C14355 VN.n12977 a_400_62400# 0.32fF
C14356 VN.n12978 a_400_62400# 0.48fF
C14357 VN.n12979 a_400_62400# 0.81fF
C14358 VN.t792 a_400_62400# 0.03fF
C14359 VN.n12980 a_400_62400# 0.32fF
C14360 VN.n12981 a_400_62400# 1.22fF
C14361 VN.n12982 a_400_62400# 0.07fF
C14362 VN.t681 a_400_62400# 0.03fF
C14363 VN.n12983 a_400_62400# 0.16fF
C14364 VN.n12984 a_400_62400# 0.19fF
C14365 VN.n12986 a_400_62400# 0.16fF
C14366 VN.t502 a_400_62400# 0.03fF
C14367 VN.n12987 a_400_62400# 0.19fF
C14368 VN.n12989 a_400_62400# 3.08fF
C14369 VN.n12990 a_400_62400# 3.75fF
C14370 VN.n12991 a_400_62400# 6.92fF
C14371 VN.t237 a_400_62400# 0.03fF
C14372 VN.n12992 a_400_62400# 0.16fF
C14373 VN.n12993 a_400_62400# 0.19fF
C14374 VN.t1688 a_400_62400# 0.03fF
C14375 VN.n12995 a_400_62400# 0.32fF
C14376 VN.n12996 a_400_62400# 1.22fF
C14377 VN.n12997 a_400_62400# 0.07fF
C14378 VN.n12998 a_400_62400# 2.51fF
C14379 VN.n12999 a_400_62400# 3.57fF
C14380 VN.t2363 a_400_62400# 0.03fF
C14381 VN.n13000 a_400_62400# 0.32fF
C14382 VN.n13001 a_400_62400# 0.48fF
C14383 VN.n13002 a_400_62400# 0.81fF
C14384 VN.n13003 a_400_62400# 0.16fF
C14385 VN.t1223 a_400_62400# 0.03fF
C14386 VN.n13004 a_400_62400# 0.19fF
C14387 VN.n13006 a_400_62400# 2.51fF
C14388 VN.n13007 a_400_62400# 3.57fF
C14389 VN.t755 a_400_62400# 0.03fF
C14390 VN.n13008 a_400_62400# 0.32fF
C14391 VN.n13009 a_400_62400# 0.48fF
C14392 VN.n13010 a_400_62400# 0.81fF
C14393 VN.t2446 a_400_62400# 0.03fF
C14394 VN.n13011 a_400_62400# 0.32fF
C14395 VN.n13012 a_400_62400# 1.22fF
C14396 VN.n13013 a_400_62400# 0.07fF
C14397 VN.t2341 a_400_62400# 0.03fF
C14398 VN.n13014 a_400_62400# 0.16fF
C14399 VN.n13015 a_400_62400# 0.19fF
C14400 VN.n13017 a_400_62400# 0.16fF
C14401 VN.t2157 a_400_62400# 0.03fF
C14402 VN.n13018 a_400_62400# 0.19fF
C14403 VN.n13020 a_400_62400# 3.08fF
C14404 VN.n13021 a_400_62400# 3.75fF
C14405 VN.n13022 a_400_62400# 6.92fF
C14406 VN.t1884 a_400_62400# 0.03fF
C14407 VN.n13023 a_400_62400# 0.16fF
C14408 VN.n13024 a_400_62400# 0.19fF
C14409 VN.t939 a_400_62400# 0.03fF
C14410 VN.n13026 a_400_62400# 0.32fF
C14411 VN.n13027 a_400_62400# 1.22fF
C14412 VN.n13028 a_400_62400# 0.07fF
C14413 VN.n13029 a_400_62400# 2.51fF
C14414 VN.n13030 a_400_62400# 3.57fF
C14415 VN.t2467 a_400_62400# 0.03fF
C14416 VN.n13031 a_400_62400# 0.32fF
C14417 VN.n13032 a_400_62400# 0.48fF
C14418 VN.n13033 a_400_62400# 0.81fF
C14419 VN.n13034 a_400_62400# 0.16fF
C14420 VN.t1333 a_400_62400# 0.03fF
C14421 VN.n13035 a_400_62400# 0.19fF
C14422 VN.n13037 a_400_62400# 2.51fF
C14423 VN.n13038 a_400_62400# 3.57fF
C14424 VN.t1338 a_400_62400# 0.03fF
C14425 VN.n13039 a_400_62400# 0.32fF
C14426 VN.n13040 a_400_62400# 0.48fF
C14427 VN.n13041 a_400_62400# 0.81fF
C14428 VN.t602 a_400_62400# 0.03fF
C14429 VN.n13042 a_400_62400# 0.32fF
C14430 VN.n13043 a_400_62400# 1.22fF
C14431 VN.n13044 a_400_62400# 0.07fF
C14432 VN.t379 a_400_62400# 0.03fF
C14433 VN.n13045 a_400_62400# 0.16fF
C14434 VN.n13046 a_400_62400# 0.19fF
C14435 VN.n13048 a_400_62400# 0.16fF
C14436 VN.t162 a_400_62400# 0.03fF
C14437 VN.n13049 a_400_62400# 0.19fF
C14438 VN.n13051 a_400_62400# 3.08fF
C14439 VN.n13052 a_400_62400# 3.75fF
C14440 VN.n13053 a_400_62400# 6.92fF
C14441 VN.t1012 a_400_62400# 0.03fF
C14442 VN.n13054 a_400_62400# 0.16fF
C14443 VN.n13055 a_400_62400# 0.19fF
C14444 VN.t1519 a_400_62400# 0.03fF
C14445 VN.n13057 a_400_62400# 0.32fF
C14446 VN.n13058 a_400_62400# 1.22fF
C14447 VN.n13059 a_400_62400# 0.07fF
C14448 VN.n13060 a_400_62400# 2.51fF
C14449 VN.n13061 a_400_62400# 3.57fF
C14450 VN.t1599 a_400_62400# 0.03fF
C14451 VN.n13062 a_400_62400# 0.32fF
C14452 VN.n13063 a_400_62400# 0.48fF
C14453 VN.n13064 a_400_62400# 0.81fF
C14454 VN.n13065 a_400_62400# 0.16fF
C14455 VN.t471 a_400_62400# 0.03fF
C14456 VN.n13066 a_400_62400# 0.19fF
C14457 VN.n13068 a_400_62400# 2.51fF
C14458 VN.n13069 a_400_62400# 3.57fF
C14459 VN.t474 a_400_62400# 0.03fF
C14460 VN.n13070 a_400_62400# 0.32fF
C14461 VN.n13071 a_400_62400# 0.48fF
C14462 VN.n13072 a_400_62400# 0.81fF
C14463 VN.t2256 a_400_62400# 0.03fF
C14464 VN.n13073 a_400_62400# 0.32fF
C14465 VN.n13074 a_400_62400# 1.22fF
C14466 VN.n13075 a_400_62400# 0.07fF
C14467 VN.t2033 a_400_62400# 0.03fF
C14468 VN.n13076 a_400_62400# 0.16fF
C14469 VN.n13077 a_400_62400# 0.19fF
C14470 VN.n13079 a_400_62400# 0.16fF
C14471 VN.t1824 a_400_62400# 0.03fF
C14472 VN.n13080 a_400_62400# 0.19fF
C14473 VN.n13082 a_400_62400# 3.08fF
C14474 VN.n13083 a_400_62400# 3.75fF
C14475 VN.n13084 a_400_62400# 6.92fF
C14476 VN.t1119 a_400_62400# 0.03fF
C14477 VN.n13085 a_400_62400# 0.16fF
C14478 VN.n13086 a_400_62400# 0.19fF
C14479 VN.t650 a_400_62400# 0.03fF
C14480 VN.n13088 a_400_62400# 0.32fF
C14481 VN.n13089 a_400_62400# 1.22fF
C14482 VN.n13090 a_400_62400# 0.07fF
C14483 VN.n13091 a_400_62400# 0.16fF
C14484 VN.n13092 a_400_62400# 0.14fF
C14485 VN.n13093 a_400_62400# 0.48fF
C14486 VN.n13094 a_400_62400# 0.62fF
C14487 VN.n13095 a_400_62400# 1.52fF
C14488 VN.n13096 a_400_62400# 2.51fF
C14489 VN.n13097 a_400_62400# 0.16fF
C14490 VN.t2121 a_400_62400# 0.03fF
C14491 VN.n13098 a_400_62400# 0.19fF
C14492 VN.t735 a_400_62400# 0.03fF
C14493 VN.n13100 a_400_62400# 0.32fF
C14494 VN.n13101 a_400_62400# 0.48fF
C14495 VN.n13102 a_400_62400# 0.81fF
C14496 VN.n13103 a_400_62400# 3.57fF
C14497 VN.n13104 a_400_62400# 5.26fF
C14498 VN.t256 a_400_62400# 0.03fF
C14499 VN.n13105 a_400_62400# 0.16fF
C14500 VN.n13106 a_400_62400# 0.19fF
C14501 VN.t2309 a_400_62400# 0.03fF
C14502 VN.n13108 a_400_62400# 0.32fF
C14503 VN.n13109 a_400_62400# 1.22fF
C14504 VN.n13110 a_400_62400# 0.07fF
C14505 VN.t236 a_400_62400# 64.17fF
C14506 VN.t1177 a_400_62400# 0.03fF
C14507 VN.n13111 a_400_62400# 0.02fF
C14508 VN.n13112 a_400_62400# 0.34fF
C14509 VN.t571 a_400_62400# 0.03fF
C14510 VN.n13114 a_400_62400# 1.60fF
C14511 VN.n13115 a_400_62400# 0.07fF
C14512 VN.t1521 a_400_62400# 0.03fF
C14513 VN.n13116 a_400_62400# 0.85fF
C14514 VN.n13117 a_400_62400# 0.81fF
C14515 VN.n13118 a_400_62400# 37.46fF
C14516 VN.n13119 a_400_62400# 54.05fF
C14517 VN.n13120 a_400_62400# 37.46fF
C14518 VN.n13121 a_400_62400# 54.05fF
C14519 VN.n13122 a_400_62400# 0.79fF
C14520 VN.n13123 a_400_62400# 0.23fF
C14521 VN.n13124 a_400_62400# 1.18fF
C14522 VN.t129 a_400_62400# 28.64fF
C14523 VN.n13125 a_400_62400# 0.79fF
C14524 VN.n13126 a_400_62400# 0.11fF
C14525 VN.n13127 a_400_62400# 4.98fF
C14526 VN.n13128 a_400_62400# 0.80fF
C14527 VN.n13129 a_400_62400# 0.29fF
C14528 VN.n13130 a_400_62400# 1.96fF
C14529 VN.n13132 a_400_62400# 25.18fF
C14530 VN.n13134 a_400_62400# 1.88fF
C14531 VN.n13135 a_400_62400# 6.03fF
C14532 VN.n13136 a_400_62400# 3.12fF
C14533 VN.n13137 a_400_62400# 7.48fF
C14534 VN.n13138 a_400_62400# 35.55fF
.ends

