magic
tech sky130A
timestamp 1677073009
<< checkpaint >>
rect -6555 -6605 18705 18655
<< dnwell >>
rect -3475 -3525 15625 15575
<< nwell >>
rect -5925 13225 18075 18025
rect -5925 -1175 -1125 13225
rect 13275 -1175 18075 13225
rect -5925 -5975 18075 -1175
<< pwell >>
rect -1125 12100 0 13225
rect 12100 12100 13275 13225
rect -1125 -1175 0 0
rect 12100 -1175 13275 0
<< mvnmos >>
rect 12100 12131 12150 12569
rect -469 -50 -31 0
rect 12181 -50 12619 0
rect 12100 -519 12150 -81
<< mvndiff >>
rect 12179 12569 12621 12571
rect -29 12563 0 12569
rect -29 12164 -23 12563
rect -64 12137 -23 12164
rect -6 12137 0 12563
rect -64 12131 0 12137
rect 12097 12131 12100 12569
rect 12150 12563 12621 12569
rect 12150 12137 12156 12563
rect 12173 12515 12621 12563
rect 12173 12185 12235 12515
rect 12565 12185 12621 12515
rect 12173 12137 12621 12185
rect 12150 12131 12621 12137
rect -64 12129 -31 12131
rect -469 12123 -31 12129
rect -469 12106 -463 12123
rect -37 12106 -31 12123
rect -469 12100 -31 12106
rect 12179 12129 12621 12131
rect 12181 12123 12619 12129
rect 12181 12106 12187 12123
rect 12613 12106 12619 12123
rect 12181 12100 12619 12106
rect -469 0 -31 3
rect 12181 0 12619 3
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 12181 -56 12619 -50
rect 12181 -73 12187 -56
rect 12613 -73 12619 -56
rect 12181 -79 12619 -73
rect 12181 -81 12214 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 12097 -519 12100 -81
rect 12150 -87 12214 -81
rect 12150 -513 12156 -87
rect 12173 -114 12214 -87
rect 12173 -513 12179 -114
rect 12150 -519 12179 -513
rect -471 -521 -29 -519
<< mvndiffc >>
rect -23 12137 -6 12563
rect 12156 12137 12173 12563
rect -463 12106 -37 12123
rect 12187 12106 12613 12123
rect -463 -73 -37 -56
rect 12187 -73 12613 -56
rect -23 -513 -6 -87
rect 12156 -513 12173 -87
<< mvpsubdiff >>
rect -1025 13113 0 13125
rect -1025 12117 -1013 13113
rect -19 12837 0 13113
rect -737 12825 0 12837
rect 12100 13113 13175 13125
rect 12100 12825 12887 12837
rect -737 12117 -725 12825
rect -1025 12100 -725 12117
rect 12235 12503 12565 12515
rect 12235 12197 12247 12503
rect 12553 12197 12565 12503
rect 12235 12185 12565 12197
rect 12875 12117 12887 12825
rect 13163 12117 13175 13113
rect 12875 12100 13175 12117
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 12875 -775 12887 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 12100 -787 12887 -775
rect 13163 -1063 13175 0
rect 12100 -1075 13175 -1063
<< mvnsubdiff >>
rect -5525 17613 17675 17625
rect -5525 -5563 -5513 17613
rect -1537 13625 13687 13637
rect -1537 -1575 -1525 13625
rect 13675 -1575 13687 13625
rect -1537 -1587 13687 -1575
rect 17663 -5563 17675 17613
rect -5525 -5575 17675 -5563
<< mvpsubdiffcont >>
rect -1013 12837 -19 13113
rect -1013 12117 -737 12837
rect 12100 12837 13163 13113
rect 12247 12197 12553 12503
rect 12887 12117 13163 12837
rect -1013 -787 -737 0
rect -403 -453 -97 -147
rect -1013 -1063 -17 -787
rect 12887 -787 13163 0
rect 12100 -1063 13163 -787
<< mvnsubdiffcont >>
rect -5513 13637 17663 17613
rect -5513 -1587 -1537 13637
rect 13687 -1587 17663 13637
rect -5513 -5563 17663 -1587
<< poly >>
rect -550 12642 0 12650
rect -550 12608 -542 12642
rect -508 12608 0 12642
rect -550 12600 0 12608
rect 12100 12642 12700 12650
rect 12100 12608 12108 12642
rect 12142 12608 12658 12642
rect 12692 12608 12700 12642
rect 12100 12600 12700 12608
rect -550 12100 -500 12600
rect 12100 12569 12150 12600
rect 12100 12100 12150 12131
rect 12650 12100 12700 12600
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -50 0 0
rect 12100 -8 12181 0
rect 12100 -42 12108 -8
rect 12142 -42 12181 -8
rect 12100 -50 12181 -42
rect 12619 -8 12700 0
rect 12619 -42 12658 -8
rect 12692 -42 12700 -8
rect 12619 -50 12700 -42
rect -550 -550 -500 -50
rect 12100 -81 12150 -50
rect 12100 -550 12150 -519
rect 12650 -550 12700 -50
rect -550 -558 0 -550
rect -550 -592 -542 -558
rect -508 -592 0 -558
rect -550 -600 0 -592
rect 12100 -558 12700 -550
rect 12100 -592 12108 -558
rect 12142 -592 12658 -558
rect 12692 -592 12700 -558
rect 12100 -600 12700 -592
<< polycont >>
rect -542 12608 -508 12642
rect 12108 12608 12142 12642
rect 12658 12608 12692 12642
rect -542 -42 -508 -8
rect 12108 -42 12142 -8
rect 12658 -42 12692 -8
rect -542 -592 -508 -558
rect 12108 -592 12142 -558
rect 12658 -592 12692 -558
<< locali >>
rect -5525 17613 17675 17625
rect -5525 -5563 -5513 17613
rect -1537 13625 13687 13637
rect -1537 -1575 -1525 13625
rect -1025 13113 0 13125
rect -1025 12117 -1013 13113
rect -19 12837 0 13113
rect -737 12825 0 12837
rect 12100 13113 13175 13125
rect 12100 12825 12887 12837
rect -737 12117 -725 12825
rect -550 12642 -500 12650
rect -550 12608 -542 12642
rect -508 12608 -500 12642
rect -550 12600 -500 12608
rect 12100 12642 12150 12650
rect 12100 12608 12108 12642
rect 12142 12608 12150 12642
rect 12100 12600 12150 12608
rect 12650 12642 12700 12650
rect 12650 12608 12658 12642
rect 12692 12608 12700 12642
rect 12650 12600 12700 12608
rect 12173 12571 12627 12577
rect -23 12563 -6 12571
rect -64 12137 -23 12164
rect -64 12129 -6 12137
rect 12156 12563 12627 12571
rect 12173 12515 12627 12563
rect 12173 12185 12235 12515
rect 12565 12185 12627 12515
rect 12173 12137 12627 12185
rect 12156 12129 12627 12137
rect -64 12123 -29 12129
rect 12173 12123 12627 12129
rect -1025 12100 -725 12117
rect -471 12106 -463 12123
rect -37 12106 -29 12123
rect 12179 12106 12187 12123
rect 12613 12106 12621 12123
rect 12875 12117 12887 12825
rect 13163 12117 13175 13113
rect 12875 12100 13175 12117
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 12100 -8 12150 0
rect 12100 -42 12108 -8
rect 12142 -42 12150 -8
rect 12100 -50 12150 -42
rect 12650 -8 12700 0
rect 12650 -42 12658 -8
rect 12692 -42 12700 -8
rect 12650 -50 12700 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 12179 -73 12187 -56
rect 12613 -73 12621 -56
rect -477 -79 -23 -73
rect 12179 -79 12214 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 12156 -87 12214 -79
rect 12173 -114 12214 -87
rect 12156 -521 12173 -513
rect -477 -527 -23 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 12100 -558 12150 -550
rect 12100 -592 12108 -558
rect 12142 -592 12150 -558
rect 12100 -600 12150 -592
rect 12650 -558 12700 -550
rect 12650 -592 12658 -558
rect 12692 -592 12700 -558
rect 12650 -600 12700 -592
rect 12875 -775 12887 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 12100 -787 12887 -775
rect 13163 -1063 13175 0
rect 12100 -1075 13175 -1063
rect 13675 -1575 13687 13625
rect -1537 -1587 13687 -1575
rect 17663 -5563 17675 17613
rect -5525 -5575 17675 -5563
<< viali >>
rect -5513 13637 17663 17613
rect -5513 -1587 -1537 13637
rect -1013 12837 -19 13113
rect -1013 12119 -737 12837
rect 12100 12837 13163 13113
rect -542 12608 -508 12642
rect 12108 12608 12142 12642
rect 12658 12608 12692 12642
rect -23 12137 -6 12563
rect 12156 12137 12173 12563
rect 12235 12503 12565 12515
rect 12235 12197 12247 12503
rect 12247 12197 12553 12503
rect 12553 12197 12565 12503
rect 12235 12185 12565 12197
rect -463 12106 -37 12123
rect 12187 12106 12613 12123
rect 12887 12119 13163 12837
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 12108 -42 12142 -8
rect 12658 -42 12692 -8
rect -463 -73 -37 -56
rect 12187 -73 12613 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 12156 -513 12173 -87
rect -542 -592 -508 -558
rect 12108 -592 12142 -558
rect 12658 -592 12692 -558
rect -1013 -1063 -19 -787
rect 12887 -787 13163 0
rect 12100 -1063 13163 -787
rect 13687 -1587 17663 13637
rect -5513 -5563 17663 -1587
<< metal1 >>
rect -5525 17613 17675 17625
rect -5525 -5563 -5513 17613
rect -1537 13625 13687 13637
rect -1537 -1575 -1525 13625
rect -1025 13113 0 13125
rect -1025 12119 -1013 13113
rect -19 12837 0 13113
rect -737 12825 0 12837
rect 12100 13113 13175 13125
rect 12100 12825 12887 12837
rect -737 12119 -725 12825
rect -550 12642 -500 12650
rect -550 12608 -542 12642
rect -508 12608 -500 12642
rect -550 12600 -500 12608
rect 12100 12642 12150 12650
rect 12100 12608 12108 12642
rect 12142 12608 12150 12642
rect 12100 12600 12150 12608
rect 12650 12642 12700 12650
rect 12650 12608 12658 12642
rect 12692 12608 12700 12642
rect 12650 12600 12700 12608
rect -474 12569 -26 12574
rect 12176 12569 12624 12574
rect -474 12563 -3 12569
rect -474 12515 -23 12563
rect -474 12185 -415 12515
rect -85 12185 -23 12515
rect -474 12137 -23 12185
rect -6 12137 -3 12563
rect -474 12131 -3 12137
rect 12153 12563 12624 12569
rect 12153 12137 12156 12563
rect 12173 12515 12624 12563
rect 12173 12185 12235 12515
rect 12565 12185 12624 12515
rect 12173 12137 12624 12185
rect 12153 12131 12624 12137
rect -474 12126 -26 12131
rect 12176 12126 12624 12131
rect -1025 12100 -725 12119
rect -469 12123 -31 12126
rect -469 12106 -463 12123
rect -37 12106 -31 12123
rect -469 12103 -31 12106
rect 12181 12123 12619 12126
rect 12181 12106 12187 12123
rect 12613 12106 12619 12123
rect 12181 12103 12619 12106
rect 12875 12119 12887 12825
rect 13163 12119 13175 13113
rect 12875 12100 13175 12119
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 12100 -8 12150 0
rect 12100 -42 12108 -8
rect 12142 -42 12150 -8
rect 12100 -50 12150 -42
rect 12650 -8 12700 0
rect 12650 -42 12658 -8
rect 12692 -42 12700 -8
rect 12650 -50 12700 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 12181 -56 12619 -53
rect 12181 -73 12187 -56
rect 12613 -73 12619 -56
rect 12181 -76 12619 -73
rect -474 -81 -26 -76
rect 12176 -81 12624 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 12153 -87 12624 -81
rect 12153 -513 12156 -87
rect 12173 -135 12624 -87
rect 12173 -465 12235 -135
rect 12565 -465 12624 -135
rect 12173 -513 12624 -465
rect 12153 -519 12624 -513
rect -474 -524 -26 -519
rect 12176 -524 12624 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 12100 -558 12150 -550
rect 12100 -592 12108 -558
rect 12142 -592 12150 -558
rect 12100 -600 12150 -592
rect 12650 -558 12700 -550
rect 12650 -592 12658 -558
rect 12692 -592 12700 -558
rect 12650 -600 12700 -592
rect 12875 -775 12887 0
rect -737 -787 0 -775
rect -19 -1063 0 -787
rect -1025 -1075 0 -1063
rect 12100 -787 12887 -775
rect 13163 -1063 13175 0
rect 12100 -1075 13175 -1063
rect 13675 -1575 13687 13625
rect -1537 -1587 13687 -1575
rect 17663 -5563 17675 17613
rect -5525 -5575 17675 -5563
<< via1 >>
rect -5513 13637 17663 17613
rect -5513 1117 -1537 13625
rect 12188 12925 12288 13025
rect -542 12608 -508 12642
rect 12108 12608 12142 12642
rect 12658 12608 12692 12642
rect -415 12185 -85 12515
rect 12235 12185 12565 12515
rect 12975 12138 13075 12238
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 12108 -42 12142 -8
rect 12658 -42 12692 -8
rect -415 -465 -85 -135
rect 12235 -465 12565 -135
rect -542 -592 -508 -558
rect 12108 -592 12142 -558
rect 12658 -592 12692 -558
rect -138 -975 -38 -875
rect 13687 -1587 17663 13637
rect -495 -5563 17663 -1587
<< metal2 >>
rect -5525 17613 17675 17625
rect -5525 13637 -5513 17613
rect -5525 13625 13687 13637
rect -5525 1117 -5513 13625
rect -1537 1117 -1525 13625
rect 12178 13025 12298 13035
rect 12178 12925 12188 13025
rect 12288 12925 12298 13025
rect 12178 12915 12298 12925
rect -725 12642 0 12825
rect -725 12608 -542 12642
rect -508 12608 0 12642
rect -725 12600 0 12608
rect 12100 12642 12875 12825
rect 12100 12608 12108 12642
rect 12142 12608 12658 12642
rect 12692 12608 12875 12642
rect 12100 12600 12875 12608
rect -725 12100 -500 12600
rect -425 12515 -75 12525
rect -425 12185 -415 12515
rect -85 12185 -75 12515
rect -425 12175 -75 12185
rect 12100 12100 12150 12600
rect 12225 12515 12575 12525
rect 12225 12185 12235 12515
rect 12565 12185 12575 12515
rect 12225 12175 12575 12185
rect 12650 12100 12875 12600
rect 12965 12238 13085 12248
rect 12965 12138 12975 12238
rect 13075 12138 13085 12238
rect 12965 12128 13085 12138
rect -725 -8 0 0
rect -725 -42 -542 -8
rect -508 -42 0 -8
rect -725 -50 0 -42
rect 12100 -8 12875 0
rect 12100 -42 12108 -8
rect 12142 -42 12658 -8
rect 12692 -42 12875 -8
rect 12100 -50 12875 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 12100 -550 12150 -50
rect 12225 -135 12575 -125
rect 12225 -465 12235 -135
rect 12565 -465 12575 -135
rect 12225 -475 12575 -465
rect 12650 -550 12875 -50
rect -725 -558 0 -550
rect -725 -592 -542 -558
rect -508 -592 0 -558
rect -725 -775 0 -592
rect 12100 -558 12875 -550
rect 12100 -592 12108 -558
rect 12142 -592 12658 -558
rect 12692 -592 12875 -558
rect 12100 -775 12875 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
rect 13675 -1575 13687 13625
rect -507 -1587 13687 -1575
rect -507 -5563 -495 -1587
rect 17663 -5563 17675 17613
rect -507 -5575 17675 -5563
<< via2 >>
rect 12188 12925 12288 13025
rect -310 12290 -190 12410
rect 12340 12290 12460 12410
rect 12975 12138 13075 12238
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 12340 -360 12460 -240
rect -138 -975 -38 -875
<< metal3 >>
rect -2525 13625 12675 14625
rect -2525 12738 -1525 13625
rect -638 12738 -186 13625
rect -2525 12414 -186 12738
rect -88 12512 0 13125
tri -186 12414 -88 12512 sw
tri -88 12424 0 12512 ne
rect 12100 13025 12464 13125
rect 12100 12925 12188 13025
rect 12288 12925 12464 13025
rect 12100 12424 12464 12925
rect -2525 12410 -88 12414
rect -2525 12290 -310 12410
rect -190 12326 -88 12410
tri -88 12326 0 12414 sw
rect -190 12290 0 12326
rect -2525 12286 0 12290
rect -2525 -575 -1525 12286
tri -412 12188 -314 12286 ne
rect -314 12188 0 12286
rect -1025 12100 -412 12188
tri -412 12100 -324 12188 sw
tri -314 12100 -226 12188 ne
rect -226 12100 0 12188
tri 12100 12326 12198 12424 ne
rect 12198 12414 12464 12424
tri 12464 12414 12562 12512 sw
rect 13675 12414 14675 12625
rect 12198 12410 14675 12414
rect 12198 12326 12340 12410
tri 12100 12238 12188 12326 sw
tri 12198 12238 12286 12326 ne
rect 12286 12290 12340 12326
rect 12460 12290 14675 12410
rect 12286 12238 14675 12290
rect 12100 12158 12188 12238
tri 12188 12158 12268 12238 sw
tri 12286 12158 12366 12238 ne
rect 12366 12158 12975 12238
rect 12100 12100 12268 12158
tri 12268 12100 12326 12158 sw
tri 12366 12100 12424 12158 ne
rect 12424 12138 12975 12158
rect 13075 12138 14675 12238
rect 12424 12100 14675 12138
rect 13675 0 14675 12100
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 12100 -40 12326 0
tri 12326 -40 12366 0 sw
tri 12424 -40 12464 0 ne
rect 12464 -40 14675 0
rect 12100 -138 12366 -40
tri 12366 -138 12464 -40 sw
tri 12464 -138 12562 -40 ne
rect 12562 -138 14675 -40
rect 12100 -226 12464 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 12100 -324 12198 -226 ne
rect 12198 -236 12464 -226
tri 12464 -236 12562 -138 sw
rect 12198 -240 13175 -236
rect 12198 -324 12340 -240
tri 12100 -364 12140 -324 sw
tri 12198 -364 12238 -324 ne
rect 12238 -360 12340 -324
rect 12460 -360 13175 -240
rect 12238 -364 13175 -360
rect 12100 -462 12140 -364
tri 12140 -462 12238 -364 sw
tri 12238 -462 12336 -364 ne
rect 12100 -1575 12238 -462
rect 12336 -688 13175 -364
rect 12336 -1075 12788 -688
rect 13675 -1575 14675 -138
rect -525 -2575 14675 -1575
<< via3 >>
rect 12188 12925 12288 13025
rect -310 12290 -190 12410
rect 12340 12290 12460 12410
rect 12975 12138 13075 12238
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect -138 -975 -38 -875
rect 12340 -360 12460 -240
<< metal4 >>
rect -2525 13625 12675 14625
rect -2525 12738 -1525 13625
rect -638 12738 -186 13625
rect -2525 12414 -186 12738
rect -88 12512 0 13125
tri -186 12414 -88 12512 sw
tri -88 12424 0 12512 ne
rect 12100 13025 12464 13125
rect 12100 12925 12188 13025
rect 12288 12925 12464 13025
rect 12100 12424 12464 12925
rect -2525 12410 -88 12414
rect -2525 12290 -310 12410
rect -190 12326 -88 12410
tri -88 12326 0 12414 sw
rect -190 12290 0 12326
rect -2525 12286 0 12290
rect -2525 -575 -1525 12286
tri -412 12188 -314 12286 ne
rect -314 12188 0 12286
rect -1025 12100 -412 12188
tri -412 12100 -324 12188 sw
tri -314 12100 -226 12188 ne
rect -226 12100 0 12188
tri 12100 12326 12198 12424 ne
rect 12198 12414 12464 12424
tri 12464 12414 12562 12512 sw
rect 13675 12414 14675 12625
rect 12198 12410 14675 12414
rect 12198 12326 12340 12410
tri 12100 12238 12188 12326 sw
tri 12198 12238 12286 12326 ne
rect 12286 12290 12340 12326
rect 12460 12290 14675 12410
rect 12286 12238 14675 12290
rect 12100 12158 12188 12238
tri 12188 12158 12268 12238 sw
tri 12286 12158 12366 12238 ne
rect 12366 12158 12975 12238
rect 12100 12100 12268 12158
tri 12268 12100 12326 12158 sw
tri 12366 12100 12424 12158 ne
rect 12424 12138 12975 12158
rect 13075 12138 14675 12238
rect 12424 12100 14675 12138
rect 13675 0 14675 12100
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 12100 -40 12326 0
tri 12326 -40 12366 0 sw
tri 12424 -40 12464 0 ne
rect 12464 -40 14675 0
rect 12100 -138 12366 -40
tri 12366 -138 12464 -40 sw
tri 12464 -138 12562 -40 ne
rect 12562 -138 14675 -40
rect 12100 -226 12464 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 12100 -324 12198 -226 ne
rect 12198 -236 12464 -226
tri 12464 -236 12562 -138 sw
rect 12198 -240 13175 -236
rect 12198 -324 12340 -240
tri 12100 -364 12140 -324 sw
tri 12198 -364 12238 -324 ne
rect 12238 -360 12340 -324
rect 12460 -360 13175 -240
rect 12238 -364 13175 -360
rect 12100 -462 12140 -364
tri 12140 -462 12238 -364 sw
tri 12238 -462 12336 -364 ne
rect 12100 -1575 12238 -462
rect 12336 -688 13175 -364
rect 12336 -1075 12788 -688
rect 13675 -1575 14675 -138
rect -525 -2575 14675 -1575
<< via4 >>
rect -310 12290 -190 12410
rect 12340 12290 12460 12410
rect -310 -360 -190 -240
rect 12340 -360 12460 -240
<< metal5 >>
rect -2525 13625 12675 14625
rect -2525 12703 -1525 13625
rect -603 12703 -292 13625
rect -2525 12410 -292 12703
tri -292 12410 -154 12548 sw
rect -53 12547 0 13125
tri -53 12494 0 12547 ne
rect 12100 12494 12358 13125
rect -2525 12392 -310 12410
rect -2525 -575 -1525 12392
tri -448 12290 -346 12392 ne
rect -346 12290 -310 12392
rect -190 12290 -154 12410
rect -1025 12100 -447 12153
tri -447 12100 -394 12153 sw
tri -346 12100 -156 12290 ne
rect -156 12256 -154 12290
tri -154 12256 0 12410 sw
rect -156 12100 0 12256
tri 12100 12256 12338 12494 ne
rect 12338 12410 12358 12494
tri 12358 12410 12496 12548 sw
rect 12338 12290 12340 12410
rect 12460 12308 12496 12410
tri 12496 12308 12598 12410 sw
rect 13675 12308 14675 12625
rect 12460 12290 14675 12308
rect 12338 12256 14675 12290
tri 12100 12100 12256 12256 sw
tri 12338 12100 12494 12256 ne
rect 12494 12100 14675 12256
rect 13675 0 14675 12100
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 0 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -156 0 -103 ne
rect 12100 -103 12256 0
tri 12256 -103 12359 0 sw
tri 12494 -103 12597 0 ne
rect 12597 -103 14675 0
rect 12100 -156 12359 -103
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
rect -208 -1575 0 -394
tri 12100 -394 12338 -156 ne
rect 12338 -240 12359 -156
tri 12359 -240 12496 -103 sw
rect 12338 -360 12340 -240
rect 12460 -342 12496 -240
tri 12496 -342 12598 -240 sw
rect 12460 -360 13175 -342
rect 12338 -394 13175 -360
tri 12100 -497 12203 -394 sw
rect 12100 -1575 12203 -497
tri 12338 -498 12442 -394 ne
rect 12442 -653 13175 -394
rect 12442 -1075 12753 -653
rect 13675 -1575 14675 -103
rect -525 -2575 14675 -1575
use nmos_drain_frame_lt  nmos_drain_frame_lt_0 mag_files
timestamp 1675431365
transform 1 0 -550 0 1 0
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_1
timestamp 1675431365
transform 0 -1 1100 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_2
timestamp 1675431365
transform 1 0 -550 0 1 1100
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_3
timestamp 1675431365
transform 0 -1 2200 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_4
timestamp 1675431365
transform 1 0 -550 0 1 2200
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_5
timestamp 1675431365
transform 0 -1 3300 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_6
timestamp 1675431365
transform 1 0 -550 0 1 3300
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_7
timestamp 1675431365
transform 0 -1 4400 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_8
timestamp 1675431365
transform 1 0 -550 0 1 4400
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_9
timestamp 1675431365
transform 0 -1 5500 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_10
timestamp 1675431365
transform 1 0 -550 0 1 5500
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_11
timestamp 1675431365
transform 0 -1 6600 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_12
timestamp 1675431365
transform 1 0 -550 0 1 6600
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_13
timestamp 1675431365
transform 0 -1 7700 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_14
timestamp 1675431365
transform 1 0 -550 0 1 7700
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_15
timestamp 1675431365
transform 0 -1 8800 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_16
timestamp 1675431365
transform 1 0 -550 0 1 8800
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_17
timestamp 1675431365
transform 0 -1 9900 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_18
timestamp 1675431365
transform 1 0 -550 0 1 9900
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_19
timestamp 1675431365
transform 0 -1 11000 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_20
timestamp 1675431365
transform 1 0 -550 0 1 11000
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_21
timestamp 1675431365
transform 0 -1 12100 -1 0 12650
box -975 -113 663 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_0 mag_files
timestamp 1675431051
transform 0 -1 550 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_1
timestamp 1675431051
transform 1 0 12100 0 1 550
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_2
timestamp 1675431051
transform 0 -1 1650 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_3
timestamp 1675431051
transform 1 0 12100 0 1 1650
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_4
timestamp 1675431051
transform 0 -1 2750 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_5
timestamp 1675431051
transform 1 0 12100 0 1 2750
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_6
timestamp 1675431051
transform 0 -1 3850 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_7
timestamp 1675431051
transform 1 0 12100 0 1 3850
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_8
timestamp 1675431051
transform 0 -1 4950 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_9
timestamp 1675431051
transform 1 0 12100 0 1 4950
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_10
timestamp 1675431051
transform 0 -1 6050 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_11
timestamp 1675431051
transform 1 0 12100 0 1 6050
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_12
timestamp 1675431051
transform 0 -1 7150 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_13
timestamp 1675431051
transform 1 0 12100 0 1 7150
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_14
timestamp 1675431051
transform 0 -1 8250 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_15
timestamp 1675431051
transform 1 0 12100 0 1 8250
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_16
timestamp 1675431051
transform 0 -1 9350 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_17
timestamp 1675431051
transform 1 0 12100 0 1 9350
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_18
timestamp 1675431051
transform 0 -1 10450 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_19
timestamp 1675431051
transform 1 0 12100 0 1 10450
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_20
timestamp 1675431051
transform 0 -1 11550 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_21
timestamp 1675431051
transform 1 0 12100 0 1 11550
box -113 -113 1575 663
use nmos_drain_in  nmos_drain_in_0 mag_files
timestamp 1675431861
transform 1 0 0 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_1
timestamp 1675431861
transform 1 0 0 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_2
timestamp 1675431861
transform 1 0 0 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_3
timestamp 1675431861
transform 1 0 0 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_4
timestamp 1675431861
transform 1 0 0 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_5
timestamp 1675431861
transform 1 0 0 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_6
timestamp 1675431861
transform 1 0 0 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_7
timestamp 1675431861
transform 1 0 0 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_8
timestamp 1675431861
transform 1 0 0 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_9
timestamp 1675431861
transform 1 0 0 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_10
timestamp 1675431861
transform 1 0 0 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_11
timestamp 1675431861
transform 1 0 550 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_12
timestamp 1675431861
transform 1 0 550 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_13
timestamp 1675431861
transform 1 0 550 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_14
timestamp 1675431861
transform 1 0 550 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_15
timestamp 1675431861
transform 1 0 550 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_16
timestamp 1675431861
transform 1 0 550 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_17
timestamp 1675431861
transform 1 0 550 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_18
timestamp 1675431861
transform 1 0 550 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_19
timestamp 1675431861
transform 1 0 550 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_20
timestamp 1675431861
transform 1 0 550 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_21
timestamp 1675431861
transform 1 0 550 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_22
timestamp 1675431861
transform 1 0 1100 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_23
timestamp 1675431861
transform 1 0 1100 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_24
timestamp 1675431861
transform 1 0 1100 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_25
timestamp 1675431861
transform 1 0 1100 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_26
timestamp 1675431861
transform 1 0 1100 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_27
timestamp 1675431861
transform 1 0 1100 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_28
timestamp 1675431861
transform 1 0 1100 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_29
timestamp 1675431861
transform 1 0 1100 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_30
timestamp 1675431861
transform 1 0 1100 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_31
timestamp 1675431861
transform 1 0 1100 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_32
timestamp 1675431861
transform 1 0 1100 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_33
timestamp 1675431861
transform 1 0 1650 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_34
timestamp 1675431861
transform 1 0 1650 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_35
timestamp 1675431861
transform 1 0 1650 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_36
timestamp 1675431861
transform 1 0 1650 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_37
timestamp 1675431861
transform 1 0 1650 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_38
timestamp 1675431861
transform 1 0 1650 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_39
timestamp 1675431861
transform 1 0 1650 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_40
timestamp 1675431861
transform 1 0 1650 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_41
timestamp 1675431861
transform 1 0 1650 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_42
timestamp 1675431861
transform 1 0 1650 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_43
timestamp 1675431861
transform 1 0 1650 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_44
timestamp 1675431861
transform 1 0 2200 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_45
timestamp 1675431861
transform 1 0 2200 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_46
timestamp 1675431861
transform 1 0 2200 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_47
timestamp 1675431861
transform 1 0 2200 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_48
timestamp 1675431861
transform 1 0 2200 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_49
timestamp 1675431861
transform 1 0 2200 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_50
timestamp 1675431861
transform 1 0 2200 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_51
timestamp 1675431861
transform 1 0 2200 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_52
timestamp 1675431861
transform 1 0 2200 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_53
timestamp 1675431861
transform 1 0 2200 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_54
timestamp 1675431861
transform 1 0 2200 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_55
timestamp 1675431861
transform 1 0 2750 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_56
timestamp 1675431861
transform 1 0 2750 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_57
timestamp 1675431861
transform 1 0 2750 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_58
timestamp 1675431861
transform 1 0 2750 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_59
timestamp 1675431861
transform 1 0 2750 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_60
timestamp 1675431861
transform 1 0 2750 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_61
timestamp 1675431861
transform 1 0 2750 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_62
timestamp 1675431861
transform 1 0 2750 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_63
timestamp 1675431861
transform 1 0 2750 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_64
timestamp 1675431861
transform 1 0 2750 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_65
timestamp 1675431861
transform 1 0 2750 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_66
timestamp 1675431861
transform 1 0 3300 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_67
timestamp 1675431861
transform 1 0 3300 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_68
timestamp 1675431861
transform 1 0 3300 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_69
timestamp 1675431861
transform 1 0 3300 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_70
timestamp 1675431861
transform 1 0 3300 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_71
timestamp 1675431861
transform 1 0 3300 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_72
timestamp 1675431861
transform 1 0 3300 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_73
timestamp 1675431861
transform 1 0 3300 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_74
timestamp 1675431861
transform 1 0 3300 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_75
timestamp 1675431861
transform 1 0 3300 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_76
timestamp 1675431861
transform 1 0 3300 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_77
timestamp 1675431861
transform 1 0 3850 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_78
timestamp 1675431861
transform 1 0 3850 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_79
timestamp 1675431861
transform 1 0 3850 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_80
timestamp 1675431861
transform 1 0 3850 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_81
timestamp 1675431861
transform 1 0 3850 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_82
timestamp 1675431861
transform 1 0 3850 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_83
timestamp 1675431861
transform 1 0 3850 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_84
timestamp 1675431861
transform 1 0 3850 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_85
timestamp 1675431861
transform 1 0 3850 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_86
timestamp 1675431861
transform 1 0 3850 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_87
timestamp 1675431861
transform 1 0 3850 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_88
timestamp 1675431861
transform 1 0 4400 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_89
timestamp 1675431861
transform 1 0 4400 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_90
timestamp 1675431861
transform 1 0 4400 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_91
timestamp 1675431861
transform 1 0 4400 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_92
timestamp 1675431861
transform 1 0 4400 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_93
timestamp 1675431861
transform 1 0 4400 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_94
timestamp 1675431861
transform 1 0 4400 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_95
timestamp 1675431861
transform 1 0 4400 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_96
timestamp 1675431861
transform 1 0 4400 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_97
timestamp 1675431861
transform 1 0 4400 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_98
timestamp 1675431861
transform 1 0 4400 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_99
timestamp 1675431861
transform 1 0 4950 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_100
timestamp 1675431861
transform 1 0 4950 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_101
timestamp 1675431861
transform 1 0 4950 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_102
timestamp 1675431861
transform 1 0 4950 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_103
timestamp 1675431861
transform 1 0 4950 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_104
timestamp 1675431861
transform 1 0 4950 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_105
timestamp 1675431861
transform 1 0 4950 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_106
timestamp 1675431861
transform 1 0 4950 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_107
timestamp 1675431861
transform 1 0 4950 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_108
timestamp 1675431861
transform 1 0 4950 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_109
timestamp 1675431861
transform 1 0 4950 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_110
timestamp 1675431861
transform 1 0 5500 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_111
timestamp 1675431861
transform 1 0 5500 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_112
timestamp 1675431861
transform 1 0 5500 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_113
timestamp 1675431861
transform 1 0 5500 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_114
timestamp 1675431861
transform 1 0 5500 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_115
timestamp 1675431861
transform 1 0 5500 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_116
timestamp 1675431861
transform 1 0 5500 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_117
timestamp 1675431861
transform 1 0 5500 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_118
timestamp 1675431861
transform 1 0 5500 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_119
timestamp 1675431861
transform 1 0 5500 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_120
timestamp 1675431861
transform 1 0 5500 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_121
timestamp 1675431861
transform 1 0 6050 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_122
timestamp 1675431861
transform 1 0 6050 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_123
timestamp 1675431861
transform 1 0 6050 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_124
timestamp 1675431861
transform 1 0 6050 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_125
timestamp 1675431861
transform 1 0 6050 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_126
timestamp 1675431861
transform 1 0 6050 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_127
timestamp 1675431861
transform 1 0 6050 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_128
timestamp 1675431861
transform 1 0 6050 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_129
timestamp 1675431861
transform 1 0 6050 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_130
timestamp 1675431861
transform 1 0 6050 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_131
timestamp 1675431861
transform 1 0 6050 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_132
timestamp 1675431861
transform 1 0 6600 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_133
timestamp 1675431861
transform 1 0 6600 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_134
timestamp 1675431861
transform 1 0 6600 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_135
timestamp 1675431861
transform 1 0 6600 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_136
timestamp 1675431861
transform 1 0 6600 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_137
timestamp 1675431861
transform 1 0 6600 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_138
timestamp 1675431861
transform 1 0 6600 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_139
timestamp 1675431861
transform 1 0 6600 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_140
timestamp 1675431861
transform 1 0 6600 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_141
timestamp 1675431861
transform 1 0 6600 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_142
timestamp 1675431861
transform 1 0 6600 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_143
timestamp 1675431861
transform 1 0 7150 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_144
timestamp 1675431861
transform 1 0 7150 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_145
timestamp 1675431861
transform 1 0 7150 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_146
timestamp 1675431861
transform 1 0 7150 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_147
timestamp 1675431861
transform 1 0 7150 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_148
timestamp 1675431861
transform 1 0 7150 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_149
timestamp 1675431861
transform 1 0 7150 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_150
timestamp 1675431861
transform 1 0 7150 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_151
timestamp 1675431861
transform 1 0 7150 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_152
timestamp 1675431861
transform 1 0 7150 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_153
timestamp 1675431861
transform 1 0 7150 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_154
timestamp 1675431861
transform 1 0 7700 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_155
timestamp 1675431861
transform 1 0 7700 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_156
timestamp 1675431861
transform 1 0 7700 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_157
timestamp 1675431861
transform 1 0 7700 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_158
timestamp 1675431861
transform 1 0 7700 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_159
timestamp 1675431861
transform 1 0 7700 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_160
timestamp 1675431861
transform 1 0 7700 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_161
timestamp 1675431861
transform 1 0 7700 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_162
timestamp 1675431861
transform 1 0 7700 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_163
timestamp 1675431861
transform 1 0 7700 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_164
timestamp 1675431861
transform 1 0 7700 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_165
timestamp 1675431861
transform 1 0 8250 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_166
timestamp 1675431861
transform 1 0 8250 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_167
timestamp 1675431861
transform 1 0 8250 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_168
timestamp 1675431861
transform 1 0 8250 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_169
timestamp 1675431861
transform 1 0 8250 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_170
timestamp 1675431861
transform 1 0 8250 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_171
timestamp 1675431861
transform 1 0 8250 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_172
timestamp 1675431861
transform 1 0 8250 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_173
timestamp 1675431861
transform 1 0 8250 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_174
timestamp 1675431861
transform 1 0 8250 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_175
timestamp 1675431861
transform 1 0 8250 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_176
timestamp 1675431861
transform 1 0 8800 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_177
timestamp 1675431861
transform 1 0 8800 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_178
timestamp 1675431861
transform 1 0 8800 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_179
timestamp 1675431861
transform 1 0 8800 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_180
timestamp 1675431861
transform 1 0 8800 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_181
timestamp 1675431861
transform 1 0 8800 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_182
timestamp 1675431861
transform 1 0 8800 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_183
timestamp 1675431861
transform 1 0 8800 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_184
timestamp 1675431861
transform 1 0 8800 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_185
timestamp 1675431861
transform 1 0 8800 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_186
timestamp 1675431861
transform 1 0 8800 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_187
timestamp 1675431861
transform 1 0 9350 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_188
timestamp 1675431861
transform 1 0 9350 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_189
timestamp 1675431861
transform 1 0 9350 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_190
timestamp 1675431861
transform 1 0 9350 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_191
timestamp 1675431861
transform 1 0 9350 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_192
timestamp 1675431861
transform 1 0 9350 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_193
timestamp 1675431861
transform 1 0 9350 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_194
timestamp 1675431861
transform 1 0 9350 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_195
timestamp 1675431861
transform 1 0 9350 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_196
timestamp 1675431861
transform 1 0 9350 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_197
timestamp 1675431861
transform 1 0 9350 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_198
timestamp 1675431861
transform 1 0 9900 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_199
timestamp 1675431861
transform 1 0 9900 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_200
timestamp 1675431861
transform 1 0 9900 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_201
timestamp 1675431861
transform 1 0 9900 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_202
timestamp 1675431861
transform 1 0 9900 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_203
timestamp 1675431861
transform 1 0 9900 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_204
timestamp 1675431861
transform 1 0 9900 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_205
timestamp 1675431861
transform 1 0 9900 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_206
timestamp 1675431861
transform 1 0 9900 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_207
timestamp 1675431861
transform 1 0 9900 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_208
timestamp 1675431861
transform 1 0 9900 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_209
timestamp 1675431861
transform 1 0 10450 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_210
timestamp 1675431861
transform 1 0 10450 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_211
timestamp 1675431861
transform 1 0 10450 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_212
timestamp 1675431861
transform 1 0 10450 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_213
timestamp 1675431861
transform 1 0 10450 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_214
timestamp 1675431861
transform 1 0 10450 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_215
timestamp 1675431861
transform 1 0 10450 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_216
timestamp 1675431861
transform 1 0 10450 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_217
timestamp 1675431861
transform 1 0 10450 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_218
timestamp 1675431861
transform 1 0 10450 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_219
timestamp 1675431861
transform 1 0 10450 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_220
timestamp 1675431861
transform 1 0 11000 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_221
timestamp 1675431861
transform 1 0 11000 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_222
timestamp 1675431861
transform 1 0 11000 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_223
timestamp 1675431861
transform 1 0 11000 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_224
timestamp 1675431861
transform 1 0 11000 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_225
timestamp 1675431861
transform 1 0 11000 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_226
timestamp 1675431861
transform 1 0 11000 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_227
timestamp 1675431861
transform 1 0 11000 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_228
timestamp 1675431861
transform 1 0 11000 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_229
timestamp 1675431861
transform 1 0 11000 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_230
timestamp 1675431861
transform 1 0 11000 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_231
timestamp 1675431861
transform 1 0 11550 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_232
timestamp 1675431861
transform 1 0 11550 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_233
timestamp 1675431861
transform 1 0 11550 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_234
timestamp 1675431861
transform 1 0 11550 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_235
timestamp 1675431861
transform 1 0 11550 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_236
timestamp 1675431861
transform 1 0 11550 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_237
timestamp 1675431861
transform 1 0 11550 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_238
timestamp 1675431861
transform 1 0 11550 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_239
timestamp 1675431861
transform 1 0 11550 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_240
timestamp 1675431861
transform 1 0 11550 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_241
timestamp 1675431861
transform 1 0 11550 0 1 11000
box -113 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_0 mag_files
timestamp 1675431308
transform 0 -1 550 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_1
timestamp 1675431308
transform 1 0 -550 0 1 550
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_2
timestamp 1675431308
transform 0 -1 1650 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_3
timestamp 1675431308
transform 1 0 -550 0 1 1650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_4
timestamp 1675431308
transform 0 -1 2750 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_5
timestamp 1675431308
transform 1 0 -550 0 1 2750
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_6
timestamp 1675431308
transform 0 -1 3850 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_7
timestamp 1675431308
transform 1 0 -550 0 1 3850
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_8
timestamp 1675431308
transform 0 -1 4950 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_9
timestamp 1675431308
transform 1 0 -550 0 1 4950
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_10
timestamp 1675431308
transform 0 -1 6050 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_11
timestamp 1675431308
transform 1 0 -550 0 1 6050
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_12
timestamp 1675431308
transform 0 -1 7150 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_13
timestamp 1675431308
transform 1 0 -550 0 1 7150
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_14
timestamp 1675431308
transform 0 -1 8250 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_15
timestamp 1675431308
transform 1 0 -550 0 1 8250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_16
timestamp 1675431308
transform 0 -1 9350 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_17
timestamp 1675431308
transform 1 0 -550 0 1 9350
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_18
timestamp 1675431308
transform 0 -1 10450 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_19
timestamp 1675431308
transform 1 0 -550 0 1 10450
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_20
timestamp 1675431308
transform 0 -1 11550 -1 0 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_21
timestamp 1675431308
transform 1 0 -550 0 1 11550
box -975 -113 663 663
use nmos_source_frame_rb  nmos_source_frame_rb_0 mag_files
timestamp 1675430904
transform 1 0 12100 0 1 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_1
timestamp 1675430904
transform 0 -1 1100 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_2
timestamp 1675430904
transform 1 0 12100 0 1 1100
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_3
timestamp 1675430904
transform 0 -1 2200 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_4
timestamp 1675430904
transform 1 0 12100 0 1 2200
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_5
timestamp 1675430904
transform 0 -1 3300 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_6
timestamp 1675430904
transform 1 0 12100 0 1 3300
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_7
timestamp 1675430904
transform 0 -1 4400 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_8
timestamp 1675430904
transform 1 0 12100 0 1 4400
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_9
timestamp 1675430904
transform 0 -1 5500 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_10
timestamp 1675430904
transform 1 0 12100 0 1 5500
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_11
timestamp 1675430904
transform 0 -1 6600 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_12
timestamp 1675430904
transform 1 0 12100 0 1 6600
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_13
timestamp 1675430904
transform 0 -1 7700 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_14
timestamp 1675430904
transform 1 0 12100 0 1 7700
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_15
timestamp 1675430904
transform 0 -1 8800 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_16
timestamp 1675430904
transform 1 0 12100 0 1 8800
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_17
timestamp 1675430904
transform 0 -1 9900 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_18
timestamp 1675430904
transform 1 0 12100 0 1 9900
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_19
timestamp 1675430904
transform 0 -1 11000 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_20
timestamp 1675430904
transform 1 0 12100 0 1 11000
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_21
timestamp 1675430904
transform 0 -1 12100 -1 0 0
box -113 -113 1575 663
use nmos_source_in  nmos_source_in_0 mag_files
timestamp 1675431769
transform 1 0 0 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_1
timestamp 1675431769
transform 1 0 0 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_2
timestamp 1675431769
transform 1 0 0 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_3
timestamp 1675431769
transform 1 0 0 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_4
timestamp 1675431769
transform 1 0 0 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_5
timestamp 1675431769
transform 1 0 0 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_6
timestamp 1675431769
transform 1 0 0 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_7
timestamp 1675431769
transform 1 0 0 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_8
timestamp 1675431769
transform 1 0 0 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_9
timestamp 1675431769
transform 1 0 0 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_10
timestamp 1675431769
transform 1 0 0 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_11
timestamp 1675431769
transform 1 0 550 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_12
timestamp 1675431769
transform 1 0 550 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_13
timestamp 1675431769
transform 1 0 550 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_14
timestamp 1675431769
transform 1 0 550 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_15
timestamp 1675431769
transform 1 0 550 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_16
timestamp 1675431769
transform 1 0 550 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_17
timestamp 1675431769
transform 1 0 550 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_18
timestamp 1675431769
transform 1 0 550 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_19
timestamp 1675431769
transform 1 0 550 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_20
timestamp 1675431769
transform 1 0 550 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_21
timestamp 1675431769
transform 1 0 550 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_22
timestamp 1675431769
transform 1 0 1100 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_23
timestamp 1675431769
transform 1 0 1100 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_24
timestamp 1675431769
transform 1 0 1100 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_25
timestamp 1675431769
transform 1 0 1100 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_26
timestamp 1675431769
transform 1 0 1100 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_27
timestamp 1675431769
transform 1 0 1100 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_28
timestamp 1675431769
transform 1 0 1100 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_29
timestamp 1675431769
transform 1 0 1100 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_30
timestamp 1675431769
transform 1 0 1100 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_31
timestamp 1675431769
transform 1 0 1100 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_32
timestamp 1675431769
transform 1 0 1100 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_33
timestamp 1675431769
transform 1 0 1650 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_34
timestamp 1675431769
transform 1 0 1650 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_35
timestamp 1675431769
transform 1 0 1650 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_36
timestamp 1675431769
transform 1 0 1650 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_37
timestamp 1675431769
transform 1 0 1650 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_38
timestamp 1675431769
transform 1 0 1650 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_39
timestamp 1675431769
transform 1 0 1650 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_40
timestamp 1675431769
transform 1 0 1650 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_41
timestamp 1675431769
transform 1 0 1650 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_42
timestamp 1675431769
transform 1 0 1650 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_43
timestamp 1675431769
transform 1 0 1650 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_44
timestamp 1675431769
transform 1 0 2200 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_45
timestamp 1675431769
transform 1 0 2200 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_46
timestamp 1675431769
transform 1 0 2200 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_47
timestamp 1675431769
transform 1 0 2200 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_48
timestamp 1675431769
transform 1 0 2200 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_49
timestamp 1675431769
transform 1 0 2200 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_50
timestamp 1675431769
transform 1 0 2200 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_51
timestamp 1675431769
transform 1 0 2200 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_52
timestamp 1675431769
transform 1 0 2200 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_53
timestamp 1675431769
transform 1 0 2200 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_54
timestamp 1675431769
transform 1 0 2200 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_55
timestamp 1675431769
transform 1 0 2750 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_56
timestamp 1675431769
transform 1 0 2750 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_57
timestamp 1675431769
transform 1 0 2750 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_58
timestamp 1675431769
transform 1 0 2750 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_59
timestamp 1675431769
transform 1 0 2750 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_60
timestamp 1675431769
transform 1 0 2750 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_61
timestamp 1675431769
transform 1 0 2750 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_62
timestamp 1675431769
transform 1 0 2750 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_63
timestamp 1675431769
transform 1 0 2750 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_64
timestamp 1675431769
transform 1 0 2750 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_65
timestamp 1675431769
transform 1 0 2750 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_66
timestamp 1675431769
transform 1 0 3300 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_67
timestamp 1675431769
transform 1 0 3300 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_68
timestamp 1675431769
transform 1 0 3300 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_69
timestamp 1675431769
transform 1 0 3300 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_70
timestamp 1675431769
transform 1 0 3300 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_71
timestamp 1675431769
transform 1 0 3300 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_72
timestamp 1675431769
transform 1 0 3300 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_73
timestamp 1675431769
transform 1 0 3300 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_74
timestamp 1675431769
transform 1 0 3300 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_75
timestamp 1675431769
transform 1 0 3300 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_76
timestamp 1675431769
transform 1 0 3300 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_77
timestamp 1675431769
transform 1 0 3850 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_78
timestamp 1675431769
transform 1 0 3850 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_79
timestamp 1675431769
transform 1 0 3850 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_80
timestamp 1675431769
transform 1 0 3850 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_81
timestamp 1675431769
transform 1 0 3850 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_82
timestamp 1675431769
transform 1 0 3850 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_83
timestamp 1675431769
transform 1 0 3850 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_84
timestamp 1675431769
transform 1 0 3850 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_85
timestamp 1675431769
transform 1 0 3850 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_86
timestamp 1675431769
transform 1 0 3850 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_87
timestamp 1675431769
transform 1 0 3850 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_88
timestamp 1675431769
transform 1 0 4400 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_89
timestamp 1675431769
transform 1 0 4400 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_90
timestamp 1675431769
transform 1 0 4400 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_91
timestamp 1675431769
transform 1 0 4400 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_92
timestamp 1675431769
transform 1 0 4400 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_93
timestamp 1675431769
transform 1 0 4400 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_94
timestamp 1675431769
transform 1 0 4400 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_95
timestamp 1675431769
transform 1 0 4400 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_96
timestamp 1675431769
transform 1 0 4400 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_97
timestamp 1675431769
transform 1 0 4400 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_98
timestamp 1675431769
transform 1 0 4400 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_99
timestamp 1675431769
transform 1 0 4950 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_100
timestamp 1675431769
transform 1 0 4950 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_101
timestamp 1675431769
transform 1 0 4950 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_102
timestamp 1675431769
transform 1 0 4950 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_103
timestamp 1675431769
transform 1 0 4950 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_104
timestamp 1675431769
transform 1 0 4950 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_105
timestamp 1675431769
transform 1 0 4950 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_106
timestamp 1675431769
transform 1 0 4950 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_107
timestamp 1675431769
transform 1 0 4950 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_108
timestamp 1675431769
transform 1 0 4950 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_109
timestamp 1675431769
transform 1 0 4950 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_110
timestamp 1675431769
transform 1 0 5500 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_111
timestamp 1675431769
transform 1 0 5500 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_112
timestamp 1675431769
transform 1 0 5500 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_113
timestamp 1675431769
transform 1 0 5500 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_114
timestamp 1675431769
transform 1 0 5500 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_115
timestamp 1675431769
transform 1 0 5500 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_116
timestamp 1675431769
transform 1 0 5500 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_117
timestamp 1675431769
transform 1 0 5500 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_118
timestamp 1675431769
transform 1 0 5500 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_119
timestamp 1675431769
transform 1 0 5500 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_120
timestamp 1675431769
transform 1 0 5500 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_121
timestamp 1675431769
transform 1 0 6050 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_122
timestamp 1675431769
transform 1 0 6050 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_123
timestamp 1675431769
transform 1 0 6050 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_124
timestamp 1675431769
transform 1 0 6050 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_125
timestamp 1675431769
transform 1 0 6050 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_126
timestamp 1675431769
transform 1 0 6050 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_127
timestamp 1675431769
transform 1 0 6050 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_128
timestamp 1675431769
transform 1 0 6050 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_129
timestamp 1675431769
transform 1 0 6050 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_130
timestamp 1675431769
transform 1 0 6050 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_131
timestamp 1675431769
transform 1 0 6050 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_132
timestamp 1675431769
transform 1 0 6600 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_133
timestamp 1675431769
transform 1 0 6600 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_134
timestamp 1675431769
transform 1 0 6600 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_135
timestamp 1675431769
transform 1 0 6600 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_136
timestamp 1675431769
transform 1 0 6600 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_137
timestamp 1675431769
transform 1 0 6600 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_138
timestamp 1675431769
transform 1 0 6600 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_139
timestamp 1675431769
transform 1 0 6600 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_140
timestamp 1675431769
transform 1 0 6600 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_141
timestamp 1675431769
transform 1 0 6600 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_142
timestamp 1675431769
transform 1 0 6600 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_143
timestamp 1675431769
transform 1 0 7150 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_144
timestamp 1675431769
transform 1 0 7150 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_145
timestamp 1675431769
transform 1 0 7150 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_146
timestamp 1675431769
transform 1 0 7150 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_147
timestamp 1675431769
transform 1 0 7150 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_148
timestamp 1675431769
transform 1 0 7150 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_149
timestamp 1675431769
transform 1 0 7150 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_150
timestamp 1675431769
transform 1 0 7150 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_151
timestamp 1675431769
transform 1 0 7150 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_152
timestamp 1675431769
transform 1 0 7150 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_153
timestamp 1675431769
transform 1 0 7150 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_154
timestamp 1675431769
transform 1 0 7700 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_155
timestamp 1675431769
transform 1 0 7700 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_156
timestamp 1675431769
transform 1 0 7700 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_157
timestamp 1675431769
transform 1 0 7700 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_158
timestamp 1675431769
transform 1 0 7700 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_159
timestamp 1675431769
transform 1 0 7700 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_160
timestamp 1675431769
transform 1 0 7700 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_161
timestamp 1675431769
transform 1 0 7700 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_162
timestamp 1675431769
transform 1 0 7700 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_163
timestamp 1675431769
transform 1 0 7700 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_164
timestamp 1675431769
transform 1 0 7700 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_165
timestamp 1675431769
transform 1 0 8250 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_166
timestamp 1675431769
transform 1 0 8250 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_167
timestamp 1675431769
transform 1 0 8250 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_168
timestamp 1675431769
transform 1 0 8250 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_169
timestamp 1675431769
transform 1 0 8250 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_170
timestamp 1675431769
transform 1 0 8250 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_171
timestamp 1675431769
transform 1 0 8250 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_172
timestamp 1675431769
transform 1 0 8250 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_173
timestamp 1675431769
transform 1 0 8250 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_174
timestamp 1675431769
transform 1 0 8250 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_175
timestamp 1675431769
transform 1 0 8250 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_176
timestamp 1675431769
transform 1 0 8800 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_177
timestamp 1675431769
transform 1 0 8800 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_178
timestamp 1675431769
transform 1 0 8800 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_179
timestamp 1675431769
transform 1 0 8800 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_180
timestamp 1675431769
transform 1 0 8800 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_181
timestamp 1675431769
transform 1 0 8800 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_182
timestamp 1675431769
transform 1 0 8800 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_183
timestamp 1675431769
transform 1 0 8800 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_184
timestamp 1675431769
transform 1 0 8800 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_185
timestamp 1675431769
transform 1 0 8800 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_186
timestamp 1675431769
transform 1 0 8800 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_187
timestamp 1675431769
transform 1 0 9350 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_188
timestamp 1675431769
transform 1 0 9350 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_189
timestamp 1675431769
transform 1 0 9350 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_190
timestamp 1675431769
transform 1 0 9350 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_191
timestamp 1675431769
transform 1 0 9350 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_192
timestamp 1675431769
transform 1 0 9350 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_193
timestamp 1675431769
transform 1 0 9350 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_194
timestamp 1675431769
transform 1 0 9350 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_195
timestamp 1675431769
transform 1 0 9350 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_196
timestamp 1675431769
transform 1 0 9350 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_197
timestamp 1675431769
transform 1 0 9350 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_198
timestamp 1675431769
transform 1 0 9900 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_199
timestamp 1675431769
transform 1 0 9900 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_200
timestamp 1675431769
transform 1 0 9900 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_201
timestamp 1675431769
transform 1 0 9900 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_202
timestamp 1675431769
transform 1 0 9900 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_203
timestamp 1675431769
transform 1 0 9900 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_204
timestamp 1675431769
transform 1 0 9900 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_205
timestamp 1675431769
transform 1 0 9900 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_206
timestamp 1675431769
transform 1 0 9900 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_207
timestamp 1675431769
transform 1 0 9900 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_208
timestamp 1675431769
transform 1 0 9900 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_209
timestamp 1675431769
transform 1 0 10450 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_210
timestamp 1675431769
transform 1 0 10450 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_211
timestamp 1675431769
transform 1 0 10450 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_212
timestamp 1675431769
transform 1 0 10450 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_213
timestamp 1675431769
transform 1 0 10450 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_214
timestamp 1675431769
transform 1 0 10450 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_215
timestamp 1675431769
transform 1 0 10450 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_216
timestamp 1675431769
transform 1 0 10450 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_217
timestamp 1675431769
transform 1 0 10450 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_218
timestamp 1675431769
transform 1 0 10450 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_219
timestamp 1675431769
transform 1 0 10450 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_220
timestamp 1675431769
transform 1 0 11000 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_221
timestamp 1675431769
transform 1 0 11000 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_222
timestamp 1675431769
transform 1 0 11000 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_223
timestamp 1675431769
transform 1 0 11000 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_224
timestamp 1675431769
transform 1 0 11000 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_225
timestamp 1675431769
transform 1 0 11000 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_226
timestamp 1675431769
transform 1 0 11000 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_227
timestamp 1675431769
transform 1 0 11000 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_228
timestamp 1675431769
transform 1 0 11000 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_229
timestamp 1675431769
transform 1 0 11000 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_230
timestamp 1675431769
transform 1 0 11000 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_231
timestamp 1675431769
transform 1 0 11550 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_232
timestamp 1675431769
transform 1 0 11550 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_233
timestamp 1675431769
transform 1 0 11550 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_234
timestamp 1675431769
transform 1 0 11550 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_235
timestamp 1675431769
transform 1 0 11550 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_236
timestamp 1675431769
transform 1 0 11550 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_237
timestamp 1675431769
transform 1 0 11550 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_238
timestamp 1675431769
transform 1 0 11550 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_239
timestamp 1675431769
transform 1 0 11550 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_240
timestamp 1675431769
transform 1 0 11550 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_241
timestamp 1675431769
transform 1 0 11550 0 1 11550
box -113 -113 663 663
<< properties >>
string MASKHINTS_HVI -140 24200 0 24340 -140 -140 0 0 24200 -140 24340 0 24200 24200 24340 24340
string MASKHINTS_HVNTM -1007 -1107 -21 -1079 -1007 -1079 -979 -121 24321 25179 25307 25207 25279 24221 25307 25179 -170 24230 -30 24370
<< end >>
