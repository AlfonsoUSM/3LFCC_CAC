* NGSPICE file created from mag_files/POSTLAYOUT/pmos_flat_24x24.ext - technology: sky130A

.subckt mag_files/POSTLAYOUT/pmos_flat_24x24 G D PW S
X0 D.t1103 G.t0 S.t1150 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1 S.t1149 G.t1 D.t1102 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 S.t1143 G.t2 D.t1101 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 S.t1148 G.t3 D.t1100 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 S.t1147 G.t4 D.t1099 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 S.t1146 G.t5 D.t1098 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 D.t1097 G.t6 S.t1145 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 D.t1096 G.t7 S.t1144 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 D.t1095 G.t8 S.t1142 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 D.t1094 G.t9 S.t1141 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 S.t1090 G.t10 D.t1093 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 D.t1092 G.t11 S.t1139 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 D.t1091 G.t12 S.t1138 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 S.t1140 G.t13 D.t1090 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 D.t1089 G.t14 S.t1137 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D.t1088 G.t15 S.t1088 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 S.t1087 G.t16 D.t1087 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 D.t1086 G.t17 S.t1091 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 D.t1085 G.t18 S.t1136 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 S.t1135 G.t19 D.t1084 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 S.t1134 G.t20 D.t1083 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 S.t1133 G.t21 D.t1082 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 S.t1132 G.t22 D.t1081 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D.t1080 G.t23 S.t1131 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 S.t1130 G.t24 D.t1079 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 S.t1129 G.t25 D.t1078 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D.t1077 G.t26 S.t1128 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 D.t1076 G.t27 S.t1127 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D.t1075 G.t28 S.t1126 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 D.t1074 G.t29 S.t1125 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 S.t1089 G.t30 D.t1073 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 S.t1124 G.t31 D.t1072 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 S.t1123 G.t32 D.t1071 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 D.t1070 G.t33 S.t1122 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 D.t1069 G.t34 S.t1094 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 S.t1121 G.t35 D.t1068 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 D.t1067 G.t36 S.t1120 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t1119 G.t37 D.t1066 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 D.t1065 G.t38 S.t1118 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 S.t1117 G.t39 D.t1064 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D.t1063 G.t40 S.t1115 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 D.t1062 G.t41 S.t1116 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 D.t1061 G.t42 S.t1114 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 S.t1111 G.t43 D.t1060 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 D.t1059 G.t44 S.t1113 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 D.t1058 G.t45 S.t1112 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 D.t1057 G.t46 S.t1110 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 D.t1056 G.t47 S.t1109 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 S.t1108 G.t48 D.t1055 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 S.t1107 G.t49 D.t1054 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 D.t1053 G.t50 S.t1106 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D.t1052 G.t51 S.t1105 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 S.t1104 G.t52 D.t1051 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 S.t1103 G.t53 D.t1050 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 S.t1102 G.t54 D.t1049 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 D.t1048 G.t55 S.t1101 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 D.t1047 G.t56 S.t1083 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 D.t1046 G.t57 S.t1100 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 D.t1045 G.t58 S.t1086 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D.t1044 G.t59 S.t1099 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 D.t1043 G.t60 S.t1095 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 D.t1042 G.t61 S.t1098 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 D.t1041 G.t62 S.t1097 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 D.t1040 G.t63 S.t1096 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 D.t1039 G.t64 S.t1093 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 D.t1038 G.t65 S.t1092 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 D.t1037 G.t66 S.t1085 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 D.t1036 G.t67 S.t1084 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 D.t1035 G.t68 S.t1082 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 D.t1034 G.t69 S.t1081 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 D.t1033 G.t70 S.t1074 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D.t1032 G.t71 S.t1076 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 D.t1031 G.t72 S.t1075 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 S.t1080 G.t73 D.t1030 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 D.t1029 G.t74 S.t1079 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 D.t1028 G.t75 S.t1078 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 D.t1027 G.t76 S.t1077 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 D.t1026 G.t77 S.t1073 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 D.t1025 G.t78 S.t1072 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 S.t1071 G.t79 D.t1024 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 S.t1070 G.t80 D.t1023 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 D.t1022 G.t81 S.t1069 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 D.t1021 G.t82 S.t1068 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 D.t1020 G.t83 S.t1067 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 D.t1019 G.t84 S.t1066 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 D.t1018 G.t85 S.t1065 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 S.t1020 G.t86 D.t1017 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 D.t1016 G.t87 S.t1064 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 S.t1063 G.t88 D.t1015 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 D.t1014 G.t89 S.t1062 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D.t1013 G.t90 S.t1061 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 D.t1012 G.t91 S.t1060 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 S.t1059 G.t92 D.t1011 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 D.t1010 G.t93 S.t1058 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 D.t1009 G.t94 S.t1057 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 D.t1008 G.t95 S.t1056 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D.t1007 G.t96 S.t1055 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 D.t1006 G.t97 S.t1054 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 S.t1053 G.t98 D.t1005 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 S.t1015 G.t99 D.t1004 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 D.t1003 G.t100 S.t1014 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 S.t1052 G.t101 D.t1002 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 S.t1051 G.t102 D.t1001 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 S.t1021 G.t103 D.t1000 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 S.t1050 G.t104 D.t999 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 D.t998 G.t105 S.t1049 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 S.t1048 G.t106 D.t997 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 S.t1047 G.t107 D.t996 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 D.t995 G.t108 S.t1046 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 D.t994 G.t109 S.t1045 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D.t993 G.t110 S.t1044 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 S.t1043 G.t111 D.t992 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t1042 G.t112 D.t991 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 D.t990 G.t113 S.t1041 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 S.t1040 G.t114 D.t989 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 D.t988 G.t115 S.t1039 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 S.t1038 G.t116 D.t987 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 S.t1037 G.t117 D.t986 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 D.t985 G.t118 S.t1036 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 S.t1035 G.t119 D.t984 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 D.t983 G.t120 S.t1034 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 S.t1033 G.t121 D.t982 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 S.t1032 G.t122 D.t981 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 S.t1030 G.t123 D.t980 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 S.t1029 G.t124 D.t979 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 S.t1031 G.t125 D.t978 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 D.t977 G.t126 S.t1028 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 S.t1017 G.t127 D.t976 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 S.t1016 G.t128 D.t975 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 S.t1018 G.t129 D.t974 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 S.t1027 G.t130 D.t973 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 S.t1026 G.t131 D.t972 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 D.t971 G.t132 S.t1025 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t1024 G.t133 D.t970 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 D.t969 G.t134 S.t1023 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t1022 G.t135 D.t968 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 S.t1019 G.t136 D.t967 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 S.t1013 G.t137 D.t966 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 D.t965 G.t138 S.t1012 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 S.t1011 G.t139 D.t964 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 S.t1005 G.t140 D.t963 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 S.t1010 G.t141 D.t962 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 D.t961 G.t142 S.t1008 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 D.t960 G.t143 S.t1009 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 S.t1007 G.t144 D.t959 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 S.t1006 G.t145 D.t958 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 S.t1004 G.t146 D.t957 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 D.t956 G.t147 S.t1003 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 S.t999 G.t148 D.t955 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 D.t954 G.t149 S.t1001 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 D.t953 G.t150 S.t1000 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 S.t1002 G.t151 D.t952 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 D.t951 G.t152 S.t998 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 S.t997 G.t153 D.t950 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 S.t996 G.t154 D.t949 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 S.t982 G.t155 D.t948 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 S.t995 G.t156 D.t947 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 D.t946 G.t157 S.t994 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 S.t993 G.t158 D.t945 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 S.t992 G.t159 D.t944 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 S.t991 G.t160 D.t943 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 S.t990 G.t161 D.t942 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 S.t989 G.t162 D.t941 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 D.t940 G.t163 S.t988 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 S.t987 G.t164 D.t939 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 D.t938 G.t165 S.t986 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 S.t985 G.t166 D.t937 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 D.t936 G.t167 S.t984 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 S.t945 G.t168 D.t935 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 D.t934 G.t169 S.t983 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 D.t933 G.t170 S.t981 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 S.t980 G.t171 D.t932 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 S.t946 G.t172 D.t931 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 D.t930 G.t173 S.t979 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 D.t929 G.t174 S.t978 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 D.t928 G.t175 S.t977 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 D.t927 G.t176 S.t976 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 S.t975 G.t177 D.t926 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 S.t964 G.t178 D.t925 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 S.t966 G.t179 D.t924 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 D.t923 G.t180 S.t965 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 D.t922 G.t181 S.t967 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 S.t974 G.t182 D.t921 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 D.t920 G.t183 S.t973 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 S.t972 G.t184 D.t919 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 D.t918 G.t185 S.t971 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 S.t970 G.t186 D.t917 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 D.t916 G.t187 S.t969 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 S.t968 G.t188 D.t915 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 S.t963 G.t189 D.t914 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 S.t962 G.t190 D.t913 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 S.t961 G.t191 D.t912 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 S.t960 G.t192 D.t911 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 D.t910 G.t193 S.t959 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 S.t947 G.t194 D.t909 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 D.t908 G.t195 S.t958 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 S.t956 G.t196 D.t907 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 D.t906 G.t197 S.t957 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 D.t905 G.t198 S.t955 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 S.t954 G.t199 D.t904 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 S.t953 G.t200 D.t903 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 S.t952 G.t201 D.t902 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 S.t951 G.t202 D.t901 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 S.t950 G.t203 D.t900 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 S.t949 G.t204 D.t899 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 S.t948 G.t205 D.t898 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 S.t944 G.t206 D.t897 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 D.t896 G.t207 S.t943 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 S.t942 G.t208 D.t895 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 D.t894 G.t209 S.t938 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 S.t937 G.t210 D.t893 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 D.t892 G.t211 S.t941 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 S.t940 G.t212 D.t891 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 D.t890 G.t213 S.t939 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 S.t936 G.t214 D.t889 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 D.t888 G.t215 S.t935 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 S.t934 G.t216 D.t887 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 S.t933 G.t217 D.t886 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 S.t878 G.t218 D.t885 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 S.t932 G.t219 D.t884 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 S.t914 G.t220 D.t883 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 D.t882 G.t221 S.t931 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 S.t930 G.t222 D.t881 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 S.t929 G.t223 D.t880 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 D.t879 G.t224 S.t915 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 S.t928 G.t225 D.t878 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 S.t927 G.t226 D.t877 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 S.t926 G.t227 D.t876 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 D.t875 G.t228 S.t925 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 S.t924 G.t229 D.t874 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 D.t873 G.t230 S.t923 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 D.t872 G.t231 S.t922 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 D.t871 G.t232 S.t921 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 D.t870 G.t233 S.t920 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 D.t869 G.t234 S.t919 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 D.t868 G.t235 S.t877 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 D.t867 G.t236 S.t876 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 D.t866 G.t237 S.t918 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 S.t917 G.t238 D.t865 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 S.t916 G.t239 D.t864 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 S.t913 G.t240 D.t863 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 D.t862 G.t241 S.t881 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 D.t861 G.t242 S.t912 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 D.t860 G.t243 S.t911 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 S.t910 G.t244 D.t859 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 S.t909 G.t245 D.t858 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 D.t857 G.t246 S.t908 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 D.t856 G.t247 S.t907 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 D.t855 G.t248 S.t897 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 D.t854 G.t249 S.t906 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 D.t853 G.t250 S.t898 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 D.t852 G.t251 S.t905 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 S.t904 G.t252 D.t851 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 D.t850 G.t253 S.t903 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 D.t849 G.t254 S.t902 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 D.t848 G.t255 S.t901 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 S.t900 G.t256 D.t847 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 D.t846 G.t257 S.t899 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 D.t845 G.t258 S.t896 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 D.t844 G.t259 S.t895 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 D.t843 G.t260 S.t893 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 D.t842 G.t261 S.t894 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 D.t841 G.t262 S.t892 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 S.t890 G.t263 D.t840 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 D.t839 G.t264 S.t889 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 D.t838 G.t265 S.t891 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 S.t888 G.t266 D.t837 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 S.t880 G.t267 D.t836 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 S.t887 G.t268 D.t835 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 D.t834 G.t269 S.t886 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 S.t885 G.t270 D.t833 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 S.t884 G.t271 D.t832 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 D.t831 G.t272 S.t883 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 S.t882 G.t273 D.t830 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 D.t829 G.t274 S.t879 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 S.t875 G.t275 D.t828 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 D.t827 G.t276 S.t874 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 D.t826 G.t277 S.t873 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 D.t825 G.t278 S.t872 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 S.t871 G.t279 D.t824 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 D.t823 G.t280 S.t867 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 D.t822 G.t281 S.t870 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 D.t821 G.t282 S.t869 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D.t820 G.t283 S.t868 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 S.t866 G.t284 D.t819 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 D.t818 G.t285 S.t865 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 D.t817 G.t286 S.t864 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 S.t863 G.t287 D.t816 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 D.t815 G.t288 S.t862 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 D.t814 G.t289 S.t807 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 S.t861 G.t290 D.t813 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 D.t812 G.t291 S.t860 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 D.t811 G.t292 S.t859 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 D.t810 G.t293 S.t808 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 D.t809 G.t294 S.t858 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 D.t808 G.t295 S.t857 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 S.t856 G.t296 D.t807 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 S.t855 G.t297 D.t806 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 D.t805 G.t298 S.t854 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 S.t853 G.t299 D.t804 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 S.t852 G.t300 D.t803 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 S.t851 G.t301 D.t802 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 D.t801 G.t302 S.t850 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 D.t800 G.t303 S.t811 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 D.t799 G.t304 S.t847 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 D.t798 G.t305 S.t848 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 S.t849 G.t306 D.t797 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 D.t796 G.t307 S.t818 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 S.t846 G.t308 D.t795 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 D.t794 G.t309 S.t812 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 S.t819 G.t310 D.t793 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 S.t845 G.t311 D.t792 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 D.t791 G.t312 S.t844 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 S.t843 G.t313 D.t790 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 S.t842 G.t314 D.t789 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 S.t841 G.t315 D.t788 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 S.t830 G.t316 D.t787 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 S.t840 G.t317 D.t786 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 S.t839 G.t318 D.t785 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 D.t784 G.t319 S.t831 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 S.t838 G.t320 D.t783 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 D.t782 G.t321 S.t837 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 D.t781 G.t322 S.t836 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 D.t780 G.t323 S.t835 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 S.t834 G.t324 D.t779 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 D.t778 G.t325 S.t833 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 D.t777 G.t326 S.t832 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 D.t776 G.t327 S.t829 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 S.t828 G.t328 D.t775 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 D.t774 G.t329 S.t809 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 S.t827 G.t330 D.t773 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 S.t826 G.t331 D.t772 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 S.t810 G.t332 D.t771 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 S.t825 G.t333 D.t770 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 S.t824 G.t334 D.t769 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 D.t768 G.t335 S.t823 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 S.t817 G.t336 D.t767 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 D.t766 G.t337 S.t822 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 S.t821 G.t338 D.t765 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 D.t764 G.t339 S.t820 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 S.t816 G.t340 D.t763 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 D.t762 G.t341 S.t815 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 S.t814 G.t342 D.t761 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 S.t813 G.t343 D.t760 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 S.t806 G.t344 D.t759 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 S.t805 G.t345 D.t758 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 S.t804 G.t346 D.t757 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 S.t798 G.t347 D.t756 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 S.t803 G.t348 D.t755 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t799 G.t349 D.t754 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 S.t802 G.t350 D.t753 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 S.t801 G.t351 D.t752 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 S.t800 G.t352 D.t751 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 S.t797 G.t353 D.t750 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 D.t749 G.t354 S.t796 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 S.t795 G.t355 D.t748 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 S.t794 G.t356 D.t747 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 D.t746 G.t357 S.t740 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 D.t745 G.t358 S.t751 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 S.t793 G.t359 D.t744 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 S.t739 G.t360 D.t743 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 D.t742 G.t361 S.t743 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 S.t792 G.t362 D.t741 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 D.t740 G.t363 S.t791 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 S.t790 G.t364 D.t739 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 S.t789 G.t365 D.t738 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 S.t788 G.t366 D.t737 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 S.t787 G.t367 D.t736 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 S.t786 G.t368 D.t735 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 S.t785 G.t369 D.t734 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 S.t784 G.t370 D.t733 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 S.t783 G.t371 D.t732 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 D.t731 G.t372 S.t741 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 D.t730 G.t373 S.t782 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 S.t742 G.t374 D.t729 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 D.t728 G.t375 S.t746 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 S.t781 G.t376 D.t727 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 S.t744 G.t377 D.t726 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 S.t745 G.t378 D.t725 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 S.t766 G.t379 D.t724 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 D.t723 G.t380 S.t780 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 S.t779 G.t381 D.t722 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 D.t721 G.t382 S.t778 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 S.t777 G.t383 D.t720 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 S.t776 G.t384 D.t719 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 D.t718 G.t385 S.t774 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 S.t775 G.t386 D.t717 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 D.t716 G.t387 S.t773 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 S.t764 G.t388 D.t715 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 S.t772 G.t389 D.t714 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 S.t771 G.t390 D.t713 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 S.t770 G.t391 D.t712 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 D.t711 G.t392 S.t769 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 D.t710 G.t393 S.t768 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 D.t709 G.t394 S.t767 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 D.t708 G.t395 S.t765 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 D.t707 G.t396 S.t763 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 D.t706 G.t397 S.t762 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 D.t705 G.t398 S.t760 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 S.t761 G.t399 D.t704 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 D.t703 G.t400 S.t759 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 D.t702 G.t401 S.t758 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 D.t701 G.t402 S.t757 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 S.t756 G.t403 D.t700 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 D.t699 G.t404 S.t755 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 D.t698 G.t405 S.t738 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 S.t754 G.t406 D.t697 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 D.t696 G.t407 S.t753 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 S.t752 G.t408 D.t695 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 S.t750 G.t409 D.t694 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 S.t749 G.t410 D.t693 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 D.t692 G.t411 S.t748 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 S.t747 G.t412 D.t691 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 D.t690 G.t413 S.t737 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 D.t689 G.t414 S.t736 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 D.t688 G.t415 S.t729 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 S.t735 G.t416 D.t687 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 D.t686 G.t417 S.t734 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 S.t733 G.t418 D.t685 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 D.t684 G.t419 S.t732 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 D.t683 G.t420 S.t731 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 D.t682 G.t421 S.t730 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 S.t728 G.t422 D.t681 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 D.t680 G.t423 S.t727 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 D.t679 G.t424 S.t726 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 S.t706 G.t425 D.t678 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 D.t677 G.t426 S.t725 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 D.t676 G.t427 S.t708 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 D.t675 G.t428 S.t724 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 D.t674 G.t429 S.t670 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 S.t723 G.t430 D.t673 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 S.t709 G.t431 D.t672 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 D.t671 G.t432 S.t722 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 D.t670 G.t433 S.t721 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 D.t669 G.t434 S.t720 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 D.t668 G.t435 S.t719 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 D.t667 G.t436 S.t718 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 S.t717 G.t437 D.t666 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 D.t665 G.t438 S.t716 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 D.t664 G.t439 S.t715 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 S.t714 G.t440 D.t663 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 S.t669 G.t441 D.t662 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 D.t661 G.t442 S.t713 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 D.t660 G.t443 S.t707 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 D.t659 G.t444 S.t710 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 D.t658 G.t445 S.t711 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 D.t657 G.t446 S.t712 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 D.t656 G.t447 S.t705 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 D.t655 G.t448 S.t671 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 D.t654 G.t449 S.t704 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 S.t703 G.t450 D.t653 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 D.t652 G.t451 S.t702 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 D.t651 G.t452 S.t701 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 D.t650 G.t453 S.t700 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 D.t649 G.t454 S.t689 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 S.t690 G.t455 D.t648 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 D.t647 G.t456 S.t691 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 D.t646 G.t457 S.t692 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 S.t699 G.t458 D.t645 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 D.t644 G.t459 S.t698 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 D.t643 G.t460 S.t697 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 D.t642 G.t461 S.t696 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 S.t695 G.t462 D.t641 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t694 G.t463 D.t640 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 S.t693 G.t464 D.t639 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 D.t638 G.t465 S.t688 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 S.t687 G.t466 D.t637 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 D.t636 G.t467 S.t686 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 S.t673 G.t468 D.t635 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 S.t685 G.t469 D.t634 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 D.t633 G.t470 S.t676 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 D.t632 G.t471 S.t684 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 D.t631 G.t472 S.t674 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 S.t675 G.t473 D.t630 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 D.t629 G.t474 S.t677 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 S.t683 G.t475 D.t628 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 S.t682 G.t476 D.t627 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 S.t681 G.t477 D.t626 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 D.t625 G.t478 S.t680 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 D.t624 G.t479 S.t679 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 D.t623 G.t480 S.t678 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 S.t672 G.t481 D.t622 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 D.t621 G.t482 S.t668 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 S.t667 G.t483 D.t620 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 S.t666 G.t484 D.t619 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 D.t618 G.t485 S.t664 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 D.t617 G.t486 S.t665 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 D.t616 G.t487 S.t663 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 S.t662 G.t488 D.t615 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 S.t661 G.t489 D.t614 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 D.t613 G.t490 S.t660 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 S.t659 G.t491 D.t612 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 S.t658 G.t492 D.t611 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 S.t609 G.t493 D.t610 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t613 G.t494 D.t609 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 D.t608 G.t495 S.t614 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 S.t618 G.t496 D.t607 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 D.t606 G.t497 S.t646 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 S.t647 G.t498 D.t605 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 S.t617 G.t499 D.t604 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 S.t657 G.t500 D.t603 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 D.t602 G.t501 S.t656 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 S.t655 G.t502 D.t601 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 S.t654 G.t503 D.t600 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 D.t599 G.t504 S.t653 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 S.t652 G.t505 D.t598 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 S.t651 G.t506 D.t597 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 S.t650 G.t507 D.t596 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 D.t595 G.t508 S.t649 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 S.t648 G.t509 D.t594 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t602 G.t510 D.t593 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 S.t645 G.t511 D.t592 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 S.t603 G.t512 D.t591 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 S.t604 G.t513 D.t590 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 D.t589 G.t514 S.t644 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 D.t588 G.t515 S.t601 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 S.t600 G.t516 D.t587 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 S.t619 G.t517 D.t586 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 S.t643 G.t518 D.t585 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 D.t584 G.t519 S.t642 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 S.t641 G.t520 D.t583 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 S.t640 G.t521 D.t582 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 S.t639 G.t522 D.t581 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 S.t628 G.t523 D.t580 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 D.t579 G.t524 S.t629 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 S.t638 G.t525 D.t578 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 D.t577 G.t526 S.t630 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 D.t576 G.t527 S.t637 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 D.t575 G.t528 S.t636 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 S.t635 G.t529 D.t574 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 S.t634 G.t530 D.t573 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D.t572 G.t531 S.t633 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 S.t632 G.t532 D.t571 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 D.t570 G.t533 S.t631 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 D.t569 G.t534 S.t627 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 S.t626 G.t535 D.t568 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 S.t605 G.t536 D.t567 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 S.t606 G.t537 D.t566 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 D.t565 G.t538 S.t607 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 S.t608 G.t539 D.t564 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 D.t563 G.t540 S.t610 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 D.t562 G.t541 S.t611 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 D.t561 G.t542 S.t612 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 S.t615 G.t543 D.t560 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 D.t559 G.t544 S.t625 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t624 G.t545 D.t558 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 S.t623 G.t546 D.t557 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 D.t556 G.t547 S.t622 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 D.t555 G.t548 S.t621 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 D.t554 G.t549 S.t620 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 S.t616 G.t550 D.t553 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 S.t599 G.t551 D.t552 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 S.t598 G.t552 D.t551 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 D.t550 G.t553 S.t597 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 D.t549 G.t554 S.t592 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 S.t593 G.t555 D.t548 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 S.t594 G.t556 D.t547 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 S.t596 G.t557 D.t546 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 S.t595 G.t558 D.t545 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 S.t591 G.t559 D.t544 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 S.t590 G.t560 D.t543 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 S.t589 G.t561 D.t542 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 S.t588 G.t562 D.t541 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 D.t540 G.t563 S.t532 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 D.t539 G.t564 S.t587 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 S.t585 G.t565 D.t538 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 S.t533 G.t566 D.t537 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 D.t536 G.t567 S.t586 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 D.t535 G.t568 S.t584 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 S.t539 G.t569 D.t534 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 D.t533 G.t570 S.t583 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 S.t582 G.t571 D.t532 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 D.t531 G.t572 S.t581 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 D.t530 G.t573 S.t580 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 D.t529 G.t574 S.t579 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 S.t578 G.t575 D.t528 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 S.t577 G.t576 D.t527 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 D.t526 G.t577 S.t576 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 S.t575 G.t578 D.t525 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 S.t574 G.t579 D.t524 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 D.t523 G.t580 S.t540 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 S.t538 G.t581 D.t522 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 D.t521 G.t582 S.t552 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 S.t573 G.t583 D.t520 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 S.t548 G.t584 D.t519 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 S.t549 G.t585 D.t518 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 D.t517 G.t586 S.t553 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 S.t572 G.t587 D.t516 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 D.t515 G.t588 S.t571 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 S.t570 G.t589 D.t514 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 D.t513 G.t590 S.t569 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 S.t568 G.t591 D.t512 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 S.t557 G.t592 D.t511 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 D.t510 G.t593 S.t567 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 D.t509 G.t594 S.t558 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 S.t559 G.t595 D.t508 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 D.t507 G.t596 S.t566 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 S.t565 G.t597 D.t506 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 D.t505 G.t598 S.t564 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 D.t504 G.t599 S.t563 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 D.t503 G.t600 S.t562 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D.t502 G.t601 S.t561 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 D.t501 G.t602 S.t560 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 S.t556 G.t603 D.t500 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 D.t499 G.t604 S.t555 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 S.t531 G.t605 D.t498 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 D.t497 G.t606 S.t543 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 D.t496 G.t607 S.t541 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 D.t495 G.t608 S.t550 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 D.t494 G.t609 S.t554 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 D.t493 G.t610 S.t534 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 D.t492 G.t611 S.t535 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 D.t491 G.t612 S.t551 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 S.t547 G.t613 D.t490 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 D.t489 G.t614 S.t546 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 D.t488 G.t615 S.t545 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 D.t487 G.t616 S.t544 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 S.t542 G.t617 D.t486 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 D.t485 G.t618 S.t537 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 S.t536 G.t619 D.t484 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 D.t483 G.t620 S.t530 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 D.t482 G.t621 S.t529 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 S.t528 G.t622 D.t481 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 S.t523 G.t623 D.t480 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 D.t479 G.t624 S.t522 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 D.t478 G.t625 S.t524 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 S.t527 G.t626 D.t477 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 D.t476 G.t627 S.t526 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 D.t475 G.t628 S.t525 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 D.t474 G.t629 S.t521 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 S.t520 G.t630 D.t473 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 D.t472 G.t631 S.t519 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 S.t518 G.t632 D.t471 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 S.t517 G.t633 D.t470 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 D.t469 G.t634 S.t465 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 D.t468 G.t635 S.t516 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 D.t467 G.t636 S.t515 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 D.t466 G.t637 S.t514 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 D.t465 G.t638 S.t466 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 D.t464 G.t639 S.t513 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 D.t463 G.t640 S.t512 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 D.t462 G.t641 S.t511 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 D.t461 G.t642 S.t510 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 S.t509 G.t643 D.t460 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 S.t508 G.t644 D.t459 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 D.t458 G.t645 S.t507 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 S.t506 G.t646 D.t457 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 D.t456 G.t647 S.t505 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 D.t455 G.t648 S.t504 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 S.t503 G.t649 D.t454 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 S.t502 G.t650 D.t453 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 D.t452 G.t651 S.t462 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 S.t467 G.t652 D.t451 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 D.t450 G.t653 S.t470 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 D.t449 G.t654 S.t501 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 D.t448 G.t655 S.t498 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 D.t447 G.t656 S.t500 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 D.t446 G.t657 S.t499 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 D.t445 G.t658 S.t497 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 D.t444 G.t659 S.t496 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 S.t495 G.t660 D.t443 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 S.t494 G.t661 D.t442 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 D.t441 G.t662 S.t487 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 S.t493 G.t663 D.t440 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 D.t439 G.t664 S.t488 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 D.t438 G.t665 S.t492 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 S.t491 G.t666 D.t437 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 D.t436 G.t667 S.t490 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 D.t435 G.t668 S.t489 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 S.t486 G.t669 D.t434 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 S.t485 G.t670 D.t433 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 S.t484 G.t671 D.t432 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 D.t431 G.t672 S.t483 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 S.t482 G.t673 D.t430 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 D.t429 G.t674 S.t481 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 D.t428 G.t675 S.t469 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 D.t427 G.t676 S.t468 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 S.t471 G.t677 D.t426 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 D.t425 G.t678 S.t472 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 S.t480 G.t679 D.t424 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 S.t478 G.t680 D.t423 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 S.t479 G.t681 D.t422 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 S.t477 G.t682 D.t421 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 S.t476 G.t683 D.t420 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 S.t475 G.t684 D.t419 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 D.t418 G.t685 S.t474 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 D.t417 G.t686 S.t473 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 S.t464 G.t687 D.t416 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 S.t463 G.t688 D.t415 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 D.t414 G.t689 S.t461 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 S.t460 G.t690 D.t413 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 D.t412 G.t691 S.t459 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 D.t411 G.t692 S.t453 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 S.t458 G.t693 D.t410 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 S.t457 G.t694 D.t409 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 S.t456 G.t695 D.t408 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 S.t455 G.t696 D.t407 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 S.t454 G.t697 D.t406 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 D.t405 G.t698 S.t452 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 D.t404 G.t699 S.t451 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 S.t448 G.t700 D.t403 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 D.t402 G.t701 S.t450 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 S.t394 G.t702 D.t401 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 D.t400 G.t703 S.t449 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 S.t446 G.t704 D.t399 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 S.t447 G.t705 D.t398 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 D.t397 G.t706 S.t445 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 S.t395 G.t707 D.t396 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 S.t444 G.t708 D.t395 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 S.t443 G.t709 D.t394 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 D.t393 G.t710 S.t442 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 D.t392 G.t711 S.t441 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 S.t440 G.t712 D.t391 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 S.t439 G.t713 D.t390 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 S.t438 G.t714 D.t389 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 D.t388 G.t715 S.t437 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 S.t436 G.t716 D.t387 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 S.t435 G.t717 D.t386 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 S.t397 G.t718 D.t385 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 S.t393 G.t719 D.t384 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 D.t383 G.t720 S.t413 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 S.t412 G.t721 D.t382 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 S.t414 G.t722 D.t381 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 S.t398 G.t723 D.t380 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 D.t379 G.t724 S.t434 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 S.t433 G.t725 D.t378 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 S.t432 G.t726 D.t377 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 S.t431 G.t727 D.t376 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 S.t430 G.t728 D.t375 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 S.t429 G.t729 D.t374 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 S.t428 G.t730 D.t373 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 S.t427 G.t731 D.t372 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 D.t371 G.t732 S.t419 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 S.t420 G.t733 D.t370 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 S.t426 G.t734 D.t369 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 S.t425 G.t735 D.t368 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 D.t367 G.t736 S.t424 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 S.t423 G.t737 D.t366 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 D.t365 G.t738 S.t422 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 D.t364 G.t739 S.t421 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 S.t418 G.t740 D.t363 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 S.t417 G.t741 D.t362 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 S.t416 G.t742 D.t361 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 S.t415 G.t743 D.t360 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 D.t359 G.t744 S.t401 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 D.t358 G.t745 S.t402 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 D.t357 G.t746 S.t411 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 D.t356 G.t747 S.t396 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 S.t400 G.t748 D.t355 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 S.t399 G.t749 D.t354 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 S.t410 G.t750 D.t353 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 D.t352 G.t751 S.t409 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 S.t408 G.t752 D.t351 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 D.t350 G.t753 S.t407 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 S.t406 G.t754 D.t349 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 S.t405 G.t755 D.t348 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 S.t404 G.t756 D.t347 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 D.t346 G.t757 S.t403 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 D.t345 G.t758 S.t392 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 S.t391 G.t759 D.t344 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 D.t343 G.t760 S.t384 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 D.t342 G.t761 S.t385 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 S.t387 G.t762 D.t341 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 S.t390 G.t763 D.t340 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 D.t339 G.t764 S.t389 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 D.t338 G.t765 S.t388 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 D.t337 G.t766 S.t386 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 S.t383 G.t767 D.t336 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 D.t335 G.t768 S.t382 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 S.t324 G.t769 D.t334 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 S.t381 G.t770 D.t333 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 S.t380 G.t771 D.t332 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 D.t331 G.t772 S.t325 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 D.t330 G.t773 S.t326 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 D.t329 G.t774 S.t327 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 D.t328 G.t775 S.t328 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 D.t327 G.t776 S.t329 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 D.t326 G.t777 S.t379 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 D.t325 G.t778 S.t378 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 D.t324 G.t779 S.t377 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 S.t376 G.t780 D.t323 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 S.t375 G.t781 D.t322 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 S.t374 G.t782 D.t321 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 D.t320 G.t783 S.t373 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 D.t319 G.t784 S.t372 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 D.t318 G.t785 S.t371 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 D.t317 G.t786 S.t370 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 S.t369 G.t787 D.t316 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 D.t315 G.t788 S.t368 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 D.t314 G.t789 S.t331 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 D.t313 G.t790 S.t339 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 S.t340 G.t791 D.t312 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 D.t311 G.t792 S.t367 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 D.t310 G.t793 S.t341 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 D.t309 G.t794 S.t366 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 D.t308 G.t795 S.t365 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 D.t307 G.t796 S.t364 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 D.t306 G.t797 S.t363 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 D.t305 G.t798 S.t362 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 D.t304 G.t799 S.t351 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 S.t352 G.t800 D.t303 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 S.t353 G.t801 D.t302 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 D.t301 G.t802 S.t355 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 D.t300 G.t803 S.t361 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 D.t299 G.t804 S.t360 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 D.t298 G.t805 S.t359 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 D.t297 G.t806 S.t358 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 S.t357 G.t807 D.t296 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 D.t295 G.t808 S.t356 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 D.t294 G.t809 S.t354 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 D.t293 G.t810 S.t350 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 D.t292 G.t811 S.t349 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 D.t291 G.t812 S.t348 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 D.t290 G.t813 S.t330 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 S.t347 G.t814 D.t289 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 D.t288 G.t815 S.t346 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 D.t287 G.t816 S.t345 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 D.t286 G.t817 S.t332 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 D.t285 G.t818 S.t333 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 D.t284 G.t819 S.t334 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 D.t283 G.t820 S.t344 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 D.t282 G.t821 S.t343 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 S.t342 G.t822 D.t281 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 S.t338 G.t823 D.t280 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 D.t279 G.t824 S.t337 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 D.t278 G.t825 S.t336 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 D.t277 G.t826 S.t335 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 S.t323 G.t827 D.t276 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 S.t322 G.t828 D.t275 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 D.t274 G.t829 S.t316 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 S.t317 G.t830 D.t273 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 S.t315 G.t831 D.t272 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 D.t271 G.t832 S.t318 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 D.t270 G.t833 S.t321 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 S.t320 G.t834 D.t269 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 S.t319 G.t835 D.t268 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 D.t267 G.t836 S.t314 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 D.t266 G.t837 S.t313 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 S.t263 G.t838 D.t265 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 S.t311 G.t839 D.t264 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 D.t263 G.t840 S.t262 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 D.t262 G.t841 S.t312 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 D.t261 G.t842 S.t310 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 S.t265 G.t843 D.t260 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 S.t267 G.t844 D.t259 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 D.t258 G.t845 S.t268 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 S.t309 G.t846 D.t257 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 S.t308 G.t847 D.t256 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 S.t307 G.t848 D.t255 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 D.t254 G.t849 S.t306 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 D.t253 G.t850 S.t305 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 D.t252 G.t851 S.t304 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 D.t251 G.t852 S.t303 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 S.t302 G.t853 D.t250 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 S.t301 G.t854 D.t249 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 D.t248 G.t855 S.t300 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 S.t266 G.t856 D.t247 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 S.t259 G.t857 D.t246 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 S.t299 G.t858 D.t245 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 S.t269 G.t859 D.t244 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 D.t243 G.t860 S.t270 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 S.t298 G.t861 D.t242 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 S.t271 G.t862 D.t241 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 D.t240 G.t863 S.t297 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 D.t239 G.t864 S.t296 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 S.t295 G.t865 D.t238 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 S.t294 G.t866 D.t237 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 S.t293 G.t867 D.t236 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 S.t292 G.t868 D.t235 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 S.t291 G.t869 D.t234 S.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 S.t289 G.t870 D.t233 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 D.t232 G.t871 S.t281 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 S.t288 G.t872 D.t231 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 S.t287 G.t873 D.t230 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 S.t286 G.t874 D.t229 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 S.t285 G.t875 D.t228 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 S.t284 G.t876 D.t227 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 D.t226 G.t877 S.t283 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 S.t282 G.t878 D.t225 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 D.t224 G.t879 S.t280 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 S.t279 G.t880 D.t223 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 S.t278 G.t881 D.t222 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 D.t221 G.t882 S.t277 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 S.t276 G.t883 D.t220 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 S.t257 G.t884 D.t219 S.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 D.t218 G.t885 S.t255 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 S.t264 G.t886 D.t217 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 S.t258 G.t887 D.t216 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 S.t272 G.t888 D.t215 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 S.t275 G.t889 D.t214 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 S.t274 G.t890 D.t213 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 S.t273 G.t891 D.t212 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 S.t261 G.t892 D.t211 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 S.t260 G.t893 D.t210 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 D.t209 G.t894 S.t254 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 D.t208 G.t895 S.t253 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 S.t252 G.t896 D.t207 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 S.t251 G.t897 D.t206 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 D.t205 G.t898 S.t250 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 S.t244 G.t899 D.t204 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 S.t245 G.t900 D.t203 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 D.t202 G.t901 S.t246 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 S.t249 G.t902 D.t201 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 D.t200 G.t903 S.t248 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 D.t199 G.t904 S.t247 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 S.t243 G.t905 D.t198 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 S.t242 G.t906 D.t197 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 S.t239 G.t907 D.t196 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 S.t241 G.t908 D.t195 S.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 D.t194 G.t909 S.t238 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 D.t193 G.t910 S.t221 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 D.t192 G.t911 S.t237 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 D.t191 G.t912 S.t222 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 D.t190 G.t913 S.t236 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 D.t189 G.t914 S.t232 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 S.t235 G.t915 D.t188 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 S.t234 G.t916 D.t187 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 S.t233 G.t917 D.t186 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 S.t231 G.t918 D.t185 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 D.t184 G.t919 S.t230 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 S.t229 G.t920 D.t183 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 D.t182 G.t921 S.t228 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 S.t227 G.t922 D.t181 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 S.t226 G.t923 D.t180 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 S.t223 G.t924 D.t179 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 S.t225 G.t925 D.t178 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 S.t224 G.t926 D.t177 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 D.t176 G.t927 S.t220 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 S.t219 G.t928 D.t175 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 D.t174 G.t929 S.t218 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 S.t217 G.t930 D.t173 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 D.t172 G.t931 S.t181 S.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 S.t216 G.t932 D.t171 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 S.t215 G.t933 D.t170 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 D.t169 G.t934 S.t214 S.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 S.t212 G.t935 D.t168 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 S.t211 G.t936 D.t167 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 D.t166 G.t937 S.t210 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 S.t209 G.t938 D.t165 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 D.t164 G.t939 S.t208 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 S.t199 G.t940 D.t163 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 D.t162 G.t941 S.t207 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 S.t206 G.t942 D.t161 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 S.t205 G.t943 D.t160 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 D.t159 G.t944 S.t204 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 D.t158 G.t945 S.t203 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 D.t157 G.t946 S.t202 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 S.t201 G.t947 D.t156 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 S.t198 G.t948 D.t155 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 S.t197 G.t949 D.t154 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 S.t196 G.t950 D.t153 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 D.t152 G.t951 S.t192 S.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 S.t193 G.t952 D.t151 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 S.t194 G.t953 D.t150 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 D.t149 G.t954 S.t179 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 D.t148 G.t955 S.t195 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 S.t190 G.t956 D.t147 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 S.t182 G.t957 D.t146 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 D.t145 G.t958 S.t189 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 D.t144 G.t959 S.t188 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 S.t187 G.t960 D.t143 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 D.t142 G.t961 S.t186 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 S.t185 G.t962 D.t141 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 S.t184 G.t963 D.t140 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 D.t139 G.t964 S.t183 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 S.t178 G.t965 D.t138 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 S.t177 G.t966 D.t137 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 D.t136 G.t967 S.t176 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 S.t175 G.t968 D.t135 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 D.t134 G.t969 S.t170 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 S.t171 G.t970 D.t133 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 S.t174 G.t971 D.t132 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 D.t131 G.t972 S.t173 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 D.t130 G.t973 S.t172 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 S.t169 G.t974 D.t129 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 D.t128 G.t975 S.t168 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 D.t127 G.t976 S.t150 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 S.t152 G.t977 D.t126 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 D.t125 G.t978 S.t153 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 D.t124 G.t979 S.t154 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 D.t123 G.t980 S.t167 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 D.t122 G.t981 S.t155 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 D.t121 G.t982 S.t156 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 D.t120 G.t983 S.t157 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 S.t166 G.t984 D.t119 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 D.t118 G.t985 S.t165 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 D.t117 G.t986 S.t164 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 D.t116 G.t987 S.t163 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 D.t115 G.t988 S.t162 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 S.t161 G.t989 D.t114 S.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 D.t113 G.t990 S.t160 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 D.t112 G.t991 S.t159 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 D.t111 G.t992 S.t158 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 D.t110 G.t993 S.t149 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 D.t109 G.t994 S.t146 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 S.t148 G.t995 D.t108 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 S.t147 G.t996 D.t107 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 D.t106 G.t997 S.t108 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 D.t105 G.t998 S.t145 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 S.t144 G.t999 D.t104 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 S.t109 G.t1000 D.t103 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 D.t102 G.t1001 S.t143 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 D.t101 G.t1002 S.t142 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 S.t141 G.t1003 D.t100 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 D.t99 G.t1004 S.t140 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 D.t98 G.t1005 S.t139 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 S.t133 G.t1006 D.t97 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 S.t134 G.t1007 D.t96 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 D.t95 G.t1008 S.t128 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 S.t135 G.t1009 D.t94 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 D.t93 G.t1010 S.t138 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 D.t92 G.t1011 S.t137 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 D.t91 G.t1012 S.t136 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 D.t90 G.t1013 S.t132 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 D.t89 G.t1014 S.t131 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 S.t130 G.t1015 D.t88 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 D.t87 G.t1016 S.t129 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 S.t127 G.t1017 D.t86 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 D.t85 G.t1018 S.t126 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 D.t84 G.t1019 S.t125 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 S.t111 G.t1020 D.t83 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 S.t124 G.t1021 D.t82 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 D.t81 G.t1022 S.t123 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 D.t80 G.t1023 S.t110 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 D.t79 G.t1024 S.t122 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 D.t78 G.t1025 S.t121 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 D.t77 G.t1026 S.t115 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 D.t76 G.t1027 S.t120 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 D.t75 G.t1028 S.t119 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 S.t118 G.t1029 D.t74 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 D.t73 G.t1030 S.t117 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 S.t116 G.t1031 D.t72 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 D.t71 G.t1032 S.t114 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 D.t70 G.t1033 S.t113 S.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 S.t107 G.t1034 D.t69 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 S.t106 G.t1035 D.t68 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 D.t67 G.t1036 S.t104 S.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 D.t66 G.t1037 S.t105 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 S.t102 G.t1038 D.t65 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 S.t97 G.t1039 D.t64 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 S.t101 G.t1040 D.t63 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 D.t62 G.t1041 S.t100 S.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 S.t98 G.t1042 D.t61 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 D.t60 G.t1043 S.t96 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 D.t59 G.t1044 S.t94 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 S.t93 G.t1045 D.t58 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 D.t57 G.t1046 S.t11 S.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 D.t56 G.t1047 S.t91 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 S.t92 G.t1048 D.t55 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 S.t7 G.t1049 D.t54 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 S.t9 G.t1050 D.t53 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 D.t52 G.t1051 S.t90 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 S.t71 G.t1052 D.t51 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 S.t89 G.t1053 D.t50 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 S.t88 G.t1054 D.t49 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 S.t87 G.t1055 D.t48 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 D.t47 G.t1056 S.t86 S.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 D.t46 G.t1057 S.t84 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 S.t83 G.t1058 D.t45 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 D.t44 G.t1059 S.t82 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 S.t80 G.t1060 D.t43 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 D.t42 G.t1061 S.t79 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 D.t41 G.t1062 S.t78 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 S.t76 G.t1063 D.t40 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 S.t74 G.t1064 D.t39 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 S.t3 G.t1065 D.t38 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 S.t73 G.t1066 D.t37 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 S.t72 G.t1067 D.t36 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 S.t70 G.t1068 D.t35 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 S.t13 G.t1069 D.t34 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 S.t69 G.t1070 D.t33 S.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 S.t67 G.t1071 D.t32 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 S.t66 G.t1072 D.t31 S.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 S.t64 G.t1073 D.t30 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 S.t63 G.t1074 D.t29 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 D.t28 G.t1075 S.t61 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 S.t48 G.t1076 D.t27 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 D.t26 G.t1077 S.t59 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 S.t51 G.t1078 D.t25 S.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 S.t57 G.t1079 D.t24 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 S.t55 G.t1080 D.t23 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 S.t54 G.t1081 D.t22 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 S.t53 G.t1082 D.t21 S.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 D.t20 G.t1083 S.t49 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 S.t46 G.t1084 D.t19 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 S.t44 G.t1085 D.t18 S.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 S.t43 G.t1086 D.t17 S.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 D.t16 G.t1087 S.t41 S.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 S.t39 G.t1088 D.t15 S.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 D.t14 G.t1089 S.t37 S.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 D.t13 G.t1090 S.t35 S.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 D.t12 G.t1091 S.t29 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 S.t33 G.t1092 D.t11 S.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 D.t10 G.t1093 S.t31 S.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 S.t28 G.t1094 D.t9 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 S.t5 G.t1095 D.t8 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 S.t26 G.t1096 D.t7 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 S.t25 G.t1097 D.t6 S.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 S.t23 G.t1098 D.t5 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 D.t4 G.t1099 S.t21 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 D.t3 G.t1100 S.t19 S.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 S.t17 G.t1101 D.t2 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 S.t15 G.t1102 D.t1 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 S.t1 G.t1103 D.t0 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 G.n563 G.t935 132.223
R1 G.n888 G.t467 132.223
R2 G.n892 G.t137 132.223
R3 G.n566 G.t611 132.223
R4 G.n570 G.t552 132.223
R5 G.n899 G.t163 132.223
R6 G.n909 G.t908 132.223
R7 G.n577 G.t207 132.223
R8 G.n584 G.t178 132.223
R9 G.n922 G.t895 132.223
R10 G.n938 G.t536 132.223
R11 G.n594 G.t929 132.223
R12 G.n604 G.t906 132.223
R13 G.n957 G.t524 132.223
R14 G.n979 G.t161 132.223
R15 G.n617 G.t548 132.223
R16 G.n632 G.t535 132.223
R17 G.n1004 G.t147 132.223
R18 G.n1029 G.t891 132.223
R19 G.n648 G.t174 132.223
R20 G.n667 G.t160 132.223
R21 G.n1057 G.t879 132.223
R22 G.n1088 G.t543 132.223
R23 G.n686 G.t951 132.223
R24 G.n708 G.t889 132.223
R25 G.n1122 G.t501 132.223
R26 G.n1159 G.t171 132.223
R27 G.n730 G.t564 132.223
R28 G.n754 G.t517 132.223
R29 G.n1197 G.t118 132.223
R30 G.n1230 G.t899 132.223
R31 G.n775 G.t187 132.223
R32 G.n793 G.t141 132.223
R33 G.n1260 G.t841 132.223
R34 G.n1284 G.t529 132.223
R35 G.n808 G.t912 132.223
R36 G.n820 G.t870 132.223
R37 G.n1305 G.t460 132.223
R38 G.n1332 G.t703 132.223
R39 G.n1320 G.t801 132.223
R40 G.n829 G.t519 132.223
R41 G.n836 G.t431 132.223
R42 G.n1341 G.t380 132.223
R43 G.n1338 G.t418 132.223
R44 G.n840 G.t143 132.223
R45 G.n841 G.t114 132.223
R46 G.n557 G.t969 132.208
R47 G.n548 G.t476 132.208
R48 G.n534 G.t504 132.208
R49 G.n514 G.t239 132.208
R50 G.n490 G.t1100 132.208
R51 G.n460 G.t874 132.208
R52 G.n425 G.t582 132.208
R53 G.n384 G.t342 132.208
R54 G.n341 G.t120 132.208
R55 G.n298 G.t918 132.208
R56 G.n255 G.t691 132.208
R57 G.n215 G.t458 132.208
R58 G.n178 G.t176 132.208
R59 G.n144 G.t1035 132.208
R60 G.n113 G.t1062 132.208
R61 G.n88 G.t532 132.208
R62 G.n66 G.t544 132.208
R63 G.n47 G.t24 132.208
R64 G.n31 G.t61 132.208
R65 G.n18 G.t603 132.208
R66 G.n8 G.t281 132.208
R67 G.n1 G.t154 132.208
R68 G.n890 G.t909 132.208
R69 G.n5 G.t1055 132.208
R70 G.n15 G.t298 132.208
R71 G.n28 G.t858 132.208
R72 G.n44 G.t819 132.208
R73 G.n63 G.t216 132.208
R74 G.n85 G.t185 132.208
R75 G.n110 G.t730 132.208
R76 G.n141 G.t706 132.208
R77 G.n175 G.t947 132.208
R78 G.n212 G.t132 132.208
R79 G.n252 G.t365 132.208
R80 G.n295 G.t594 132.208
R81 G.n338 G.t884 132.208
R82 G.n381 G.t9 132.208
R83 G.n422 G.t273 132.208
R84 G.n457 G.t528 132.208
R85 G.n487 G.t780 132.208
R86 G.n511 G.t1028 132.208
R87 G.n531 G.t156 132.208
R88 G.n545 G.t142 132.208
R89 G.n554 G.t650 132.208
R90 G.n568 G.t973 132.208
R91 G.n542 G.t920 132.208
R92 G.n528 G.t235 132.208
R93 G.n508 G.t43 132.208
R94 G.n484 G.t850 132.208
R95 G.n454 G.t416 132.208
R96 G.n419 G.t109 132.208
R97 G.n378 G.t782 132.208
R98 G.n335 G.t486 132.208
R99 G.n292 G.t48 132.208
R100 G.n249 G.t855 132.208
R101 G.n209 G.t422 132.208
R102 G.n172 G.t113 132.208
R103 G.n138 G.t787 132.208
R104 G.n107 G.t105 132.208
R105 G.n82 G.t53 132.208
R106 G.n60 G.t482 132.208
R107 G.n41 G.t425 132.208
R108 G.n25 G.t851 132.208
R109 G.n12 G.t791 132.208
R110 G.n895 G.t514 132.208
R111 G.n897 G.t102 132.208
R112 G.n907 G.t860 132.208
R113 G.n905 G.t151 132.208
R114 G.n903 G.t447 132.208
R115 G.n22 G.t498 132.208
R116 G.n38 G.t77 132.208
R117 G.n57 G.t129 132.208
R118 G.n79 G.t816 132.208
R119 G.n104 G.t866 132.208
R120 G.n135 G.t445 132.208
R121 G.n169 G.t872 132.208
R122 G.n206 G.t75 132.208
R123 G.n246 G.t505 132.208
R124 G.n289 G.t812 132.208
R125 G.n332 G.t133 132.208
R126 G.n375 G.t444 132.208
R127 G.n416 G.t869 132.208
R128 G.n451 G.t72 132.208
R129 G.n481 G.t503 132.208
R130 G.n505 G.t809 132.208
R131 G.n525 G.t995 132.208
R132 G.n573 G.t570 132.208
R133 G.n575 G.t622 132.208
R134 G.n582 G.t586 132.208
R135 G.n580 G.t546 132.208
R136 G.n522 G.t958 132.208
R137 G.n502 G.t763 132.208
R138 G.n478 G.t471 132.208
R139 G.n448 G.t30 132.208
R140 G.n413 G.t837 132.208
R141 G.n372 G.t403 132.208
R142 G.n329 G.t100 132.208
R143 G.n286 G.t767 132.208
R144 G.n243 G.t474 132.208
R145 G.n203 G.t35 132.208
R146 G.n166 G.t840 132.208
R147 G.n132 G.t406 132.208
R148 G.n101 G.t833 132.208
R149 G.n76 G.t771 132.208
R150 G.n54 G.t97 132.208
R151 G.n35 G.t37 132.208
R152 G.n914 G.t472 132.208
R153 G.n916 G.t408 132.208
R154 G.n918 G.t138 132.208
R155 G.n920 G.t823 132.208
R156 G.n936 G.t480 132.208
R157 G.n934 G.t881 132.208
R158 G.n932 G.t62 132.208
R159 G.n930 G.t116 132.208
R160 G.n928 G.t799 132.208
R161 G.n51 G.t859 132.208
R162 G.n73 G.t433 132.208
R163 G.n98 G.t489 132.208
R164 G.n129 G.t60 132.208
R165 G.n163 G.t492 132.208
R166 G.n200 G.t796 132.208
R167 G.n240 G.t122 132.208
R168 G.n283 G.t429 132.208
R169 G.n326 G.t861 132.208
R170 G.n369 G.t57 132.208
R171 G.n410 G.t491 132.208
R172 G.n445 G.t793 132.208
R173 G.n475 G.t121 132.208
R174 G.n499 G.t427 132.208
R175 G.n588 G.t605 132.208
R176 G.n590 G.t197 132.208
R177 G.n592 G.t244 132.208
R178 G.n602 G.t209 132.208
R179 G.n600 G.t172 132.208
R180 G.n598 G.t572 132.208
R181 G.n496 G.t384 132.208
R182 G.n472 G.t82 132.208
R183 G.n442 G.t748 132.208
R184 G.n407 G.t454 132.208
R185 G.n366 G.t13 132.208
R186 G.n323 G.t824 132.208
R187 G.n280 G.t386 132.208
R188 G.n237 G.t84 132.208
R189 G.n197 G.t752 132.208
R190 G.n160 G.t459 132.208
R191 G.n126 G.t16 132.208
R192 G.n95 G.t446 132.208
R193 G.n70 G.t391 132.208
R194 G.n945 G.t817 132.208
R195 G.n947 G.t754 132.208
R196 G.n949 G.t78 132.208
R197 G.n951 G.t19 132.208
R198 G.n953 G.t863 132.208
R199 G.n955 G.t441 132.208
R200 G.n977 G.t93 132.208
R201 G.n975 G.t511 132.208
R202 G.n973 G.t783 132.208
R203 G.n971 G.t844 132.208
R204 G.n969 G.t417 132.208
R205 G.n967 G.t477 132.208
R206 G.n965 G.t44 132.208
R207 G.n92 G.t103 132.208
R208 G.n123 G.t777 132.208
R209 G.n157 G.t106 132.208
R210 G.n194 G.t413 132.208
R211 G.n234 G.t847 132.208
R212 G.n277 G.t41 132.208
R213 G.n320 G.t481 132.208
R214 G.n363 G.t775 132.208
R215 G.n404 G.t104 132.208
R216 G.n439 G.t411 132.208
R217 G.n469 G.t846 132.208
R218 G.n609 G.t40 132.208
R219 G.n611 G.t227 132.208
R220 G.n613 G.t913 132.208
R221 G.n615 G.t963 132.208
R222 G.n630 G.t927 132.208
R223 G.n628 G.t900 132.208
R224 G.n626 G.t193 132.208
R225 G.n624 G.t1102 132.208
R226 G.n466 G.t803 132.208
R227 G.n436 G.t374 132.208
R228 G.n401 G.t67 132.208
R229 G.n360 G.t737 132.208
R230 G.n317 G.t439 132.208
R231 G.n274 G.t3 132.208
R232 G.n231 G.t805 132.208
R233 G.n191 G.t376 132.208
R234 G.n154 G.t69 132.208
R235 G.n120 G.t740 132.208
R236 G.n988 G.t58 132.208
R237 G.n990 G.t5 132.208
R238 G.n992 G.t432 132.208
R239 G.n994 G.t378 132.208
R240 G.n996 G.t798 132.208
R241 G.n998 G.t741 132.208
R242 G.n1000 G.t485 132.208
R243 G.n1002 G.t52 132.208
R244 G.n1027 G.t815 132.208
R245 G.n1025 G.t131 132.208
R246 G.n1023 G.t398 132.208
R247 G.n1021 G.t462 132.208
R248 G.n1019 G.t26 132.208
R249 G.n1017 G.t88 132.208
R250 G.n1015 G.t758 132.208
R251 G.n1013 G.t827 132.208
R252 G.n117 G.t395 132.208
R253 G.n151 G.t831 132.208
R254 G.n188 G.t23 132.208
R255 G.n228 G.t466 132.208
R256 G.n271 G.t757 132.208
R257 G.n314 G.t92 132.208
R258 G.n357 G.t394 132.208
R259 G.n398 G.t830 132.208
R260 G.n433 G.t17 132.208
R261 G.n638 G.t463 132.208
R262 G.n640 G.t753 132.208
R263 G.n642 G.t952 132.208
R264 G.n644 G.t540 132.208
R265 G.n646 G.t579 132.208
R266 G.n665 G.t549 132.208
R267 G.n663 G.t530 132.208
R268 G.n661 G.t914 132.208
R269 G.n659 G.t722 132.208
R270 G.n657 G.t421 132.208
R271 G.n655 G.t1092 132.208
R272 G.n395 G.t786 132.208
R273 G.n354 G.t362 132.208
R274 G.n311 G.t51 132.208
R275 G.n268 G.t727 132.208
R276 G.n225 G.t424 132.208
R277 G.n185 G.t1094 132.208
R278 G.n148 G.t789 132.208
R279 G.n1039 G.t364 132.208
R280 G.n1041 G.t776 132.208
R281 G.n1043 G.t728 132.208
R282 G.n1045 G.t42 132.208
R283 G.n1047 G.t1095 132.208
R284 G.n1049 G.t415 132.208
R285 G.n1051 G.t367 132.208
R286 G.n1053 G.t95 132.208
R287 G.n1055 G.t769 132.208
R288 G.n1086 G.t497 132.208
R289 G.n1084 G.t892 132.208
R290 G.n1082 G.t91 132.208
R291 G.n1080 G.t136 132.208
R292 G.n1078 G.t829 132.208
R293 G.n1076 G.t873 132.208
R294 G.n1074 G.t461 132.208
R295 G.n1072 G.t506 132.208
R296 G.n1070 G.t87 132.208
R297 G.n1068 G.t510 132.208
R298 G.n182 G.t826 132.208
R299 G.n222 G.t140 132.208
R300 G.n265 G.t457 132.208
R301 G.n308 G.t878 132.208
R302 G.n351 G.t83 132.208
R303 G.n392 G.t509 132.208
R304 G.n674 G.t821 132.208
R305 G.n676 G.t139 132.208
R306 G.n678 G.t451 132.208
R307 G.n680 G.t633 132.208
R308 G.n682 G.t215 132.208
R309 G.n684 G.t271 132.208
R310 G.n706 G.t175 132.208
R311 G.n704 G.t153 132.208
R312 G.n702 G.t541 132.208
R313 G.n700 G.t345 132.208
R314 G.n698 G.t29 132.208
R315 G.n696 G.t713 132.208
R316 G.n694 G.t402 132.208
R317 G.n348 G.t1079 132.208
R318 G.n305 G.t766 132.208
R319 G.n262 G.t349 132.208
R320 G.n219 G.t34 132.208
R321 G.n1100 G.t714 132.208
R322 G.n1102 G.t405 132.208
R323 G.n1104 G.t1080 132.208
R324 G.n1106 G.t397 132.208
R325 G.n1108 G.t352 132.208
R326 G.n1110 G.t761 132.208
R327 G.n1112 G.t716 132.208
R328 G.n1114 G.t28 132.208
R329 G.n1116 G.t1084 132.208
R330 G.n1118 G.t818 132.208
R331 G.n1120 G.t389 132.208
R332 G.n1157 G.t115 132.208
R333 G.n1155 G.t521 132.208
R334 G.n1153 G.t811 132.208
R335 G.n1151 G.t862 132.208
R336 G.n1149 G.t443 132.208
R337 G.n1147 G.t493 132.208
R338 G.n1145 G.t71 132.208
R339 G.n1143 G.t124 132.208
R340 G.n1141 G.t808 132.208
R341 G.n1139 G.t130 132.208
R342 G.n1137 G.t442 132.208
R343 G.n1135 G.t867 132.208
R344 G.n259 G.t68 132.208
R345 G.n302 G.t496 132.208
R346 G.n345 G.t804 132.208
R347 G.n716 G.t127 132.208
R348 G.n718 G.t438 132.208
R349 G.n720 G.t865 132.208
R350 G.n722 G.t65 132.208
R351 G.n724 G.t252 132.208
R352 G.n726 G.t934 132.208
R353 G.n728 G.t989 132.208
R354 G.n752 G.t904 132.208
R355 G.n750 G.t883 132.208
R356 G.n748 G.t167 132.208
R357 G.n746 G.t1068 132.208
R358 G.n744 G.t746 132.208
R359 G.n742 G.t336 132.208
R360 G.n740 G.t12 132.208
R361 G.n738 G.t704 132.208
R362 G.n1525 G.t385 132.208
R363 G.n1171 G.t1070 132.208
R364 G.n1173 G.t751 132.208
R365 G.n1175 G.t338 132.208
R366 G.n1177 G.t15 132.208
R367 G.n1179 G.t705 132.208
R368 G.n1181 G.t8 132.208
R369 G.n1183 G.t1072 132.208
R370 G.n1185 G.t382 132.208
R371 G.n1187 G.t340 132.208
R372 G.n1189 G.t745 132.208
R373 G.n1191 G.t707 132.208
R374 G.n1193 G.t434 132.208
R375 G.n1195 G.t1 132.208
R376 G.n1228 G.t842 132.208
R377 G.n1226 G.t144 132.208
R378 G.n1224 G.t426 132.208
R379 G.n1222 G.t483 132.208
R380 G.n1220 G.t55 132.208
R381 G.n1218 G.t107 132.208
R382 G.n1216 G.t788 132.208
R383 G.n1214 G.t848 132.208
R384 G.n1212 G.t423 132.208
R385 G.n1210 G.t857 132.208
R386 G.n1208 G.t50 132.208
R387 G.n1474 G.t488 132.208
R388 G.n1499 G.t784 132.208
R389 G.n1524 G.t111 132.208
R390 G.n1551 G.t419 132.208
R391 G.n761 G.t853 132.208
R392 G.n763 G.t46 132.208
R393 G.n765 G.t484 132.208
R394 G.n767 G.t778 132.208
R395 G.n769 G.t974 132.208
R396 G.n771 G.t553 132.208
R397 G.n773 G.t597 132.208
R398 G.n791 G.t533 132.208
R399 G.n789 G.t512 132.208
R400 G.n787 G.t898 132.208
R401 G.n785 G.t690 132.208
R402 G.n783 G.t373 132.208
R403 G.n781 G.t1058 132.208
R404 G.n1580 G.t736 132.208
R405 G.n1556 G.t328 132.208
R406 G.n1530 G.t0 132.208
R407 G.n1503 G.t693 132.208
R408 G.n1478 G.t375 132.208
R409 G.n1453 G.t1060 132.208
R410 G.n1240 G.t739 132.208
R411 G.n1242 G.t330 132.208
R412 G.n1244 G.t732 132.208
R413 G.n1246 G.t695 132.208
R414 G.n1248 G.t1099 132.208
R415 G.n1250 G.t1064 132.208
R416 G.n1252 G.t372 132.208
R417 G.n1254 G.t332 132.208
R418 G.n1256 G.t45 132.208
R419 G.n1258 G.t725 132.208
R420 G.n1282 G.t456 132.208
R421 G.n1280 G.t875 132.208
R422 G.n1278 G.t38 132.208
R423 G.n1276 G.t98 132.208
R424 G.n1274 G.t774 132.208
R425 G.n1272 G.t834 132.208
R426 G.n1270 G.t407 132.208
R427 G.n1268 G.t468 132.208
R428 G.n1414 G.t36 132.208
R429 G.n1432 G.t475 132.208
R430 G.n1451 G.t768 132.208
R431 G.n1473 G.t101 132.208
R432 G.n1498 G.t404 132.208
R433 G.n1523 G.t839 132.208
R434 G.n1550 G.t33 132.208
R435 G.n1576 G.t473 132.208
R436 G.n1600 G.t765 132.208
R437 G.n798 G.t99 132.208
R438 G.n800 G.t400 132.208
R439 G.n802 G.t587 132.208
R440 G.n804 G.t180 132.208
R441 G.n806 G.t220 132.208
R442 G.n818 G.t157 132.208
R443 G.n816 G.t135 132.208
R444 G.n814 G.t527 132.208
R445 G.n812 G.t313 132.208
R446 G.n1624 G.t1091 132.208
R447 G.n1606 G.t677 132.208
R448 G.n1585 G.t361 132.208
R449 G.n1561 G.t1048 132.208
R450 G.n1535 G.t724 132.208
R451 G.n1508 G.t316 132.208
R452 G.n1483 G.t1093 132.208
R453 G.n1458 G.t680 132.208
R454 G.n1436 G.t363 132.208
R455 G.n1417 G.t1049 132.208
R456 G.n1399 G.t357 132.208
R457 G.n1291 G.t317 132.208
R458 G.n1293 G.t720 132.208
R459 G.n1295 G.t682 132.208
R460 G.n1297 G.t1089 132.208
R461 G.n1299 G.t1052 132.208
R462 G.n1301 G.t764 132.208
R463 G.n1303 G.t350 132.208
R464 G.n1317 G.t85 132.208
R465 G.n1314 G.t409 132.208
R466 G.n1311 G.t542 132.208
R467 G.n1308 G.t179 132.208
R468 G.n1306 G.t449 132.208
R469 G.n1372 G.t86 132.208
R470 G.n1384 G.t307 132.208
R471 G.n1397 G.t1045 132.208
R472 G.n1413 G.t173 132.208
R473 G.n1431 G.t814 132.208
R474 G.n1450 G.t70 132.208
R475 G.n1472 G.t669 132.208
R476 G.n1497 G.t1037 132.208
R477 G.n1522 G.t539 132.208
R478 G.n1549 G.t903 132.208
R479 G.n1575 G.t437 132.208
R480 G.n1599 G.t797 132.208
R481 G.n1620 G.t300 132.208
R482 G.n1638 G.t659 132.208
R483 G.n823 G.t388 132.208
R484 G.n825 G.t614 132.208
R485 G.n827 G.t256 132.208
R486 G.n834 G.t170 132.208
R487 G.n831 G.t537 132.208
R488 G.n1655 G.t305 132.208
R489 G.n1637 G.t557 132.208
R490 G.n1619 G.t198 132.208
R491 G.n1598 G.t702 132.208
R492 G.n1574 G.t337 132.208
R493 G.n1548 G.t856 132.208
R494 G.n1521 G.t490 132.208
R495 G.n1496 G.t933 132.208
R496 G.n1471 G.t567 132.208
R497 G.n1449 G.t1073 132.208
R498 G.n1430 G.t710 132.208
R499 G.n1412 G.t123 132.208
R500 G.n1396 G.t945 132.208
R501 G.n1383 G.t210 132.208
R502 G.n1371 G.t1083 132.208
R503 G.n1361 G.t348 132.208
R504 G.n1322 G.t134 132.208
R505 G.n1324 G.t500 132.208
R506 G.n1327 G.t319 132.208
R507 G.n1329 G.t1082 132.208
R508 G.n1674 G.t937 132.208
R509 G.n1669 G.t201 132.208
R510 G.n1660 G.t1077 132.208
R511 G.n1648 G.t240 132.208
R512 G.n1633 G.t982 132.208
R513 G.n1615 G.t377 132.208
R514 G.n1594 G.t6 132.208
R515 G.n1570 G.t518 132.208
R516 G.n1544 G.t149 132.208
R517 G.n1517 G.t613 132.208
R518 G.n1492 G.t255 132.208
R519 G.n1467 G.t743 132.208
R520 G.n1445 G.t387 132.208
R521 G.n1426 G.t886 132.208
R522 G.n1408 G.t629 132.208
R523 G.n1392 G.t996 132.208
R524 G.n1379 G.t760 132.208
R525 G.n1367 G.t20 132.208
R526 G.n1357 G.t894 132.208
R527 G.n1350 G.t155 132.208
R528 G.n1344 G.t1090 132.208
R529 G.n1339 G.t759 132.208
R530 G.n1336 G.t806 132.208
R531 G.n1334 G.t21 132.208
R532 G.n1347 G.t169 132.208
R533 G.n1353 G.t907 132.208
R534 G.n1360 G.t64 132.208
R535 G.n1370 G.t807 132.208
R536 G.n1382 G.t1030 132.208
R537 G.n1395 G.t666 132.208
R538 G.n1411 G.t901 132.208
R539 G.n1429 G.t430 132.208
R540 G.n1448 G.t792 132.208
R541 G.n1470 G.t296 132.208
R542 G.n1495 G.t655 132.208
R543 G.n1520 G.t164 132.208
R544 G.n1547 G.t534 132.208
R545 G.n1573 G.t49 132.208
R546 G.n1597 G.t414 132.208
R547 G.n1618 G.t1020 132.208
R548 G.n1636 G.t283 132.208
R549 G.n1651 G.t4 132.208
R550 G.n1663 G.t231 132.208
R551 G.n838 G.t977 132.208
R552 G.n837 G.t260 120.189
R553 G.n1333 G.t547 120.189
R554 G.n1342 G.t263 120.189
R555 G.n1343 G.t896 120.189
R556 G.n1346 G.t580 120.189
R557 G.n1349 G.t322 120.189
R558 G.n1352 G.t25 120.189
R559 G.n1356 G.t681 120.189
R560 G.n1359 G.t392 120.189
R561 G.n1366 G.t181 120.189
R562 G.n1369 G.t999 120.189
R563 G.n1378 G.t545 120.189
R564 G.n1381 G.t259 120.189
R565 G.n1391 G.t89 120.189
R566 G.n1394 G.t887 120.189
R567 G.n1407 G.t455 120.189
R568 G.n1410 G.t150 120.189
R569 G.n1425 G.t1047 120.189
R570 G.n1428 G.t749 120.189
R571 G.n1444 G.t310 120.189
R572 G.n1447 G.t7 120.189
R573 G.n1466 G.t910 120.189
R574 G.n1469 G.t617 120.189
R575 G.n1491 G.t73 120.189
R576 G.n1494 G.t882 120.189
R577 G.n1516 G.t813 120.189
R578 G.n1519 G.t520 120.189
R579 G.n1543 G.t1038 120.189
R580 G.n1546 G.t738 120.189
R581 G.n1569 G.t668 120.189
R582 G.n1572 G.t379 120.189
R583 G.n1593 G.t905 120.189
R584 G.n1596 G.t600 120.189
R585 G.n1614 G.t538 120.189
R586 G.n1617 G.t245 120.189
R587 G.n1632 G.t800 120.189
R588 G.n1635 G.t515 120.189
R589 G.n1647 G.t436 120.189
R590 G.n1650 G.t146 120.189
R591 G.n1659 G.t888 120.189
R592 G.n1662 G.t563 120.189
R593 G.n1668 G.t393 120.189
R594 G.n1671 G.t117 120.189
R595 G.n1673 G.t750 120.189
R596 G.n1676 G.t487 120.189
R597 G.n1330 G.t643 120.189
R598 G.n1321 G.t964 120.189
R599 G.n1325 G.t412 120.189
R600 G.n1354 G.t772 120.189
R601 G.n1364 G.t279 120.189
R602 G.n1376 G.t638 120.189
R603 G.n1389 G.t158 120.189
R604 G.n1405 G.t526 120.189
R605 G.n1423 G.t31 120.189
R606 G.n1442 G.t396 120.189
R607 G.n1464 G.t1006 120.189
R608 G.n1489 G.t152 120.189
R609 G.n1514 G.t890 120.189
R610 G.n1541 G.t14 120.189
R611 G.n1567 G.t755 120.189
R612 G.n1591 G.t992 120.189
R613 G.n1612 G.t623 120.189
R614 G.n1630 G.t885 120.189
R615 G.n1645 G.t523 120.189
R616 G.n1657 G.t944 120.189
R617 G.n1666 G.t499 120.189
R618 G.n832 G.t864 120.189
R619 G.n830 G.t347 120.189
R620 G.n821 G.t639 120.189
R621 G.n822 G.t32 120.189
R622 G.n1664 G.t773 120.189
R623 G.n1654 G.t159 120.189
R624 G.n1643 G.t825 120.189
R625 G.n1628 G.t79 120.189
R626 G.n1610 G.t911 120.189
R627 G.n1589 G.t177 120.189
R628 G.n1565 G.t1051 120.189
R629 G.n1539 G.t315 120.189
R630 G.n1512 G.t94 120.189
R631 G.n1487 G.t464 120.189
R632 G.n1462 G.t183 120.189
R633 G.n1440 G.t687 120.189
R634 G.n1421 G.t327 120.189
R635 G.n1403 G.t838 120.189
R636 G.n1387 G.t478 120.189
R637 G.n1374 G.t916 120.189
R638 G.n1362 G.t554 120.189
R639 G.n1309 G.t1063 120.189
R640 G.n1312 G.t698 120.189
R641 G.n1315 G.t166 120.189
R642 G.n1318 G.t921 120.189
R643 G.n1285 G.t1071 120.189
R644 G.n1286 G.t257 120.189
R645 G.n1287 G.t275 120.189
R646 G.n1288 G.t573 120.189
R647 G.n1289 G.t1007 120.189
R648 G.n1290 G.t211 120.189
R649 G.n1385 G.t632 120.189
R650 G.n1401 G.t941 120.189
R651 G.n1419 G.t270 120.189
R652 G.n1438 G.t568 120.189
R653 G.n1460 G.t1003 120.189
R654 G.n1485 G.t577 120.189
R655 G.n1510 G.t630 120.189
R656 G.n1537 G.t213 120.189
R657 G.n1563 G.t266 120.189
R658 G.n1587 G.t946 120.189
R659 G.n1608 G.t1000 120.189
R660 G.n1626 G.t574 120.189
R661 G.n1641 G.t626 120.189
R662 G.n1652 G.t11 120.189
R663 G.n811 G.t450 120.189
R664 G.n810 G.t744 120.189
R665 G.n809 G.t80 120.189
R666 G.n794 G.t428 120.189
R667 G.n795 G.t1097 120.189
R668 G.n796 G.t794 120.189
R669 G.n797 G.t369 120.189
R670 G.n1639 G.t978 120.189
R671 G.n1623 G.t924 120.189
R672 G.n1605 G.t241 120.189
R673 G.n1584 G.t191 120.189
R674 G.n1560 G.t602 120.189
R675 G.n1534 G.t558 120.189
R676 G.n1507 G.t980 120.189
R677 G.n1482 G.t926 120.189
R678 G.n1457 G.t246 120.189
R679 G.n1435 G.t922 120.189
R680 G.n1416 G.t606 120.189
R681 G.n1398 G.t189 120.189
R682 G.n1267 G.t983 120.189
R683 G.n1266 G.t555 120.189
R684 G.n1265 G.t248 120.189
R685 G.n1264 G.t923 120.189
R686 G.n1263 G.t609 120.189
R687 G.n1262 G.t592 120.189
R688 G.n1261 G.t323 120.189
R689 G.n1231 G.t351 120.189
R690 G.n1232 G.t636 120.189
R691 G.n1233 G.t652 120.189
R692 G.n1234 G.t954 120.189
R693 G.n1235 G.t290 120.189
R694 G.n1236 G.t588 120.189
R695 G.n1237 G.t1021 120.189
R696 G.n1238 G.t221 120.189
R697 G.n1239 G.t649 120.189
R698 G.n1433 G.t955 120.189
R699 G.n1455 G.t287 120.189
R700 G.n1480 G.t961 120.189
R701 G.n1505 G.t1017 120.189
R702 G.n1532 G.t590 120.189
R703 G.n1558 G.t646 120.189
R704 G.n1582 G.t224 120.189
R705 G.n1603 G.t284 120.189
R706 G.n1621 G.t959 120.189
R707 G.n780 G.t1015 120.189
R708 G.n779 G.t401 120.189
R709 G.n778 G.t835 120.189
R710 G.n777 G.t27 120.189
R711 G.n776 G.t469 120.189
R712 G.n755 G.t810 120.189
R713 G.n756 G.t381 120.189
R714 G.n757 G.t74 120.189
R715 G.n758 G.t742 120.189
R716 G.n759 G.t258 120.189
R717 G.n760 G.t206 120.189
R718 G.n1601 G.t620 120.189
R719 G.n1579 G.t569 120.189
R720 G.n1555 G.t993 120.189
R721 G.n1529 G.t938 120.189
R722 G.n1502 G.t261 120.189
R723 G.n1477 G.t205 120.189
R724 G.n1452 G.t624 120.189
R725 G.n1207 G.t202 120.189
R726 G.n1206 G.t997 120.189
R727 G.n1205 G.t566 120.189
R728 G.n1204 G.t264 120.189
R729 G.n1203 G.t936 120.189
R730 G.n1202 G.t627 120.189
R731 G.n1201 G.t204 120.189
R732 G.n1200 G.t1001 120.189
R733 G.n1199 G.t984 120.189
R734 G.n1198 G.t699 120.189
R735 G.n1160 G.t726 120.189
R736 G.n1161 G.t1022 120.189
R737 G.n1162 G.t1034 120.189
R738 G.n1163 G.t236 120.189
R739 G.n1164 G.t663 120.189
R740 G.n1165 G.t975 120.189
R741 G.n1166 G.t301 120.189
R742 G.n1167 G.t598 120.189
R743 G.n1168 G.t1031 120.189
R744 G.n1169 G.t232 120.189
R745 G.n1170 G.t661 120.189
R746 G.n1475 G.t242 120.189
R747 G.n1500 G.t299 120.189
R748 G.n1527 G.t979 120.189
R749 G.n1553 G.t1029 120.189
R750 G.n1577 G.t601 120.189
R751 G.n737 G.t660 120.189
R752 G.n736 G.t237 120.189
R753 G.n735 G.t297 120.189
R754 G.n734 G.t785 120.189
R755 G.n733 G.t112 120.189
R756 G.n732 G.t420 120.189
R757 G.n731 G.t854 120.189
R758 G.n709 G.t90 120.189
R759 G.n710 G.t756 120.189
R760 G.n711 G.t465 120.189
R761 G.n712 G.t22 120.189
R762 G.n713 G.t637 120.189
R763 G.n714 G.t583 120.189
R764 G.n715 G.t1010 120.189
R765 G.n387 G.t953 120.189
R766 G.n344 G.t276 120.189
R767 G.n301 G.t218 120.189
R768 G.n258 G.t640 120.189
R769 G.n1134 G.t584 120.189
R770 G.n1133 G.t1012 120.189
R771 G.n1132 G.t578 120.189
R772 G.n1131 G.t278 120.189
R773 G.n1130 G.t950 120.189
R774 G.n1129 G.t642 120.189
R775 G.n1128 G.t214 120.189
R776 G.n1127 G.t1014 120.189
R777 G.n1126 G.t581 120.189
R778 G.n1125 G.t280 120.189
R779 G.n1124 G.t267 120.189
R780 G.n1123 G.t1075 120.189
R781 G.n1089 G.t2 120.189
R782 G.n1090 G.t302 120.189
R783 G.n1091 G.t311 120.189
R784 G.n1092 G.t618 120.189
R785 G.n1093 G.t1042 120.189
R786 G.n1094 G.t253 120.189
R787 G.n1095 G.t673 120.189
R788 G.n1096 G.t990 120.189
R789 G.n1097 G.t308 120.189
R790 G.n1098 G.t615 120.189
R791 G.n1099 G.t1040 120.189
R792 G.n218 G.t625 120.189
R793 G.n261 G.t671 120.189
R794 G.n304 G.t262 120.189
R795 G.n347 G.t306 120.189
R796 G.n389 G.t994 120.189
R797 G.n693 G.t1039 120.189
R798 G.n692 G.t621 120.189
R799 G.n691 G.t670 120.189
R800 G.n690 G.t66 120.189
R801 G.n689 G.t494 120.189
R802 G.n688 G.t802 120.189
R803 G.n687 G.t125 120.189
R804 G.n668 G.t479 120.189
R805 G.n669 G.t39 120.189
R806 G.n670 G.t845 120.189
R807 G.n671 G.t410 120.189
R808 G.n672 G.t1023 120.189
R809 G.n673 G.t966 120.189
R810 G.n428 G.t291 120.189
R811 G.n391 G.t229 120.189
R812 G.n350 G.t653 120.189
R813 G.n307 G.t595 120.189
R814 G.n264 G.t1025 120.189
R815 G.n221 G.t971 120.189
R816 G.n181 G.t293 120.189
R817 G.n1067 G.t962 120.189
R818 G.n1066 G.t656 120.189
R819 G.n1065 G.t226 120.189
R820 G.n1064 G.t1027 120.189
R821 G.n1063 G.t591 120.189
R822 G.n1062 G.t295 120.189
R823 G.n1061 G.t965 120.189
R824 G.n1060 G.t658 120.189
R825 G.n1059 G.t644 120.189
R826 G.n1058 G.t358 120.189
R827 G.n1030 G.t390 120.189
R828 G.n1031 G.t675 120.189
R829 G.n1032 G.t688 120.189
R830 G.n1033 G.t1008 120.189
R831 G.n1034 G.t324 120.189
R832 G.n1035 G.t634 120.189
R833 G.n1036 G.t1054 120.189
R834 G.n1037 G.t272 120.189
R835 G.n1038 G.t684 120.189
R836 G.n147 G.t1004 120.189
R837 G.n184 G.t320 120.189
R838 G.n224 G.t1013 120.189
R839 G.n267 G.t1053 120.189
R840 G.n310 G.t641 120.189
R841 G.n353 G.t683 120.189
R842 G.n394 G.t277 120.189
R843 G.n430 G.t318 120.189
R844 G.n654 G.t1011 120.189
R845 G.n653 G.t1050 120.189
R846 G.n652 G.t452 120.189
R847 G.n651 G.t876 120.189
R848 G.n650 G.t81 120.189
R849 G.n649 G.t507 120.189
R850 G.n633 G.t779 120.189
R851 G.n634 G.t360 120.189
R852 G.n635 G.t47 120.189
R853 G.n636 G.t723 120.189
R854 G.n637 G.t228 120.189
R855 G.n463 G.t186 120.189
R856 G.n432 G.t593 120.189
R857 G.n397 G.t551 120.189
R858 G.n356 G.t967 120.189
R859 G.n313 G.t917 120.189
R860 G.n270 G.t230 120.189
R861 G.n227 G.t188 120.189
R862 G.n187 G.t596 120.189
R863 G.n150 G.t182 120.189
R864 G.n116 G.t972 120.189
R865 G.n1012 G.t550 120.189
R866 G.n1011 G.t233 120.189
R867 G.n1010 G.t915 120.189
R868 G.n1009 G.t599 120.189
R869 G.n1008 G.t184 120.189
R870 G.n1007 G.t976 120.189
R871 G.n1006 G.t956 120.189
R872 G.n1005 G.t678 120.189
R873 G.n980 G.t770 120.189
R874 G.n981 G.t1057 120.189
R875 G.n982 G.t1067 120.189
R876 G.n983 G.t288 120.189
R877 G.n984 G.t700 120.189
R878 G.n985 G.t1018 120.189
R879 G.n986 G.t334 120.189
R880 G.n987 G.t647 120.189
R881 G.n119 G.t1066 120.189
R882 G.n153 G.t285 120.189
R883 G.n190 G.t697 120.189
R884 G.n230 G.t294 120.189
R885 G.n273 G.t333 120.189
R886 G.n316 G.t1026 120.189
R887 G.n359 G.t1065 120.189
R888 G.n400 G.t654 120.189
R889 G.n435 G.t696 120.189
R890 G.n465 G.t292 120.189
R891 G.n622 G.t331 120.189
R892 G.n621 G.t836 120.189
R893 G.n620 G.t145 120.189
R894 G.n619 G.t470 120.189
R895 G.n618 G.t880 120.189
R896 G.n605 G.t63 120.189
R897 G.n606 G.t735 120.189
R898 G.n607 G.t435 120.189
R899 G.n608 G.t1103 120.189
R900 G.n493 G.t608 120.189
R901 G.n468 G.t562 120.189
R902 G.n438 G.t986 120.189
R903 G.n403 G.t932 120.189
R904 G.n362 G.t249 120.189
R905 G.n319 G.t200 120.189
R906 G.n276 G.t610 120.189
R907 G.n233 G.t565 120.189
R908 G.n193 G.t987 120.189
R909 G.n156 G.t559 120.189
R910 G.n122 G.t251 120.189
R911 G.n91 G.t928 120.189
R912 G.n964 G.t616 120.189
R913 G.n963 G.t194 120.189
R914 G.n962 G.t991 120.189
R915 G.n961 G.t560 120.189
R916 G.n960 G.t254 120.189
R917 G.n959 G.t238 120.189
R918 G.n958 G.t1061 120.189
R919 G.n939 G.t54 120.189
R920 G.n940 G.t335 120.189
R921 G.n941 G.t346 120.189
R922 G.n942 G.t665 120.189
R923 G.n943 G.t1078 120.189
R924 G.n944 G.t303 120.189
R925 G.n69 G.t712 120.189
R926 G.n94 G.t1033 120.189
R927 G.n125 G.t344 120.189
R928 G.n159 G.t662 120.189
R929 G.n196 G.t1076 120.189
R930 G.n236 G.t667 120.189
R931 G.n279 G.t709 120.189
R932 G.n322 G.t304 120.189
R933 G.n365 G.t343 120.189
R934 G.n406 G.t1036 120.189
R935 G.n441 G.t1074 120.189
R936 G.n471 G.t664 120.189
R937 G.n495 G.t708 120.189
R938 G.n517 G.t110 120.189
R939 G.n597 G.t522 120.189
R940 G.n596 G.t852 120.189
R941 G.n595 G.t148 120.189
R942 G.n585 G.t448 120.189
R943 G.n586 G.t10 120.189
R944 G.n587 G.t820 120.189
R945 G.n519 G.t383 120.189
R946 G.n498 G.t998 120.189
R947 G.n474 G.t943 120.189
R948 G.n444 G.t265 120.189
R949 G.n409 G.t212 120.189
R950 G.n368 G.t628 120.189
R951 G.n325 G.t576 120.189
R952 G.n282 G.t1002 120.189
R953 G.n239 G.t949 120.189
R954 G.n199 G.t269 120.189
R955 G.n162 G.t940 120.189
R956 G.n128 G.t631 120.189
R957 G.n97 G.t208 120.189
R958 G.n72 G.t1005 120.189
R959 G.n50 G.t571 120.189
R960 G.n927 G.t274 120.189
R961 G.n926 G.t942 120.189
R962 G.n925 G.t635 120.189
R963 G.n924 G.t619 120.189
R964 G.n923 G.t339 120.189
R965 G.n910 G.t440 120.189
R966 G.n911 G.t711 120.189
R967 G.n912 G.t721 120.189
R968 G.n913 G.t1044 120.189
R969 G.n34 G.t359 120.189
R970 G.n53 G.t674 120.189
R971 G.n75 G.t1088 120.189
R972 G.n100 G.t309 120.189
R973 G.n131 G.t719 120.189
R974 G.n165 G.t1041 120.189
R975 G.n202 G.t356 120.189
R976 G.n242 G.t1046 120.189
R977 G.n285 G.t1086 120.189
R978 G.n328 G.t676 120.189
R979 G.n371 G.t718 120.189
R980 G.n412 G.t312 120.189
R981 G.n447 G.t355 120.189
R982 G.n477 G.t1043 120.189
R983 G.n501 G.t1085 120.189
R984 G.n521 G.t495 120.189
R985 G.n537 G.t893 120.189
R986 G.n579 G.t126 120.189
R987 G.n578 G.t525 120.189
R988 G.n571 G.t832 120.189
R989 G.n572 G.t399 120.189
R990 G.n539 G.t96 120.189
R991 G.n524 G.t762 120.189
R992 G.n504 G.t282 120.189
R993 G.n480 G.t222 120.189
R994 G.n450 G.t645 120.189
R995 G.n415 G.t589 120.189
R996 G.n374 G.t1016 120.189
R997 G.n331 G.t960 120.189
R998 G.n288 G.t286 120.189
R999 G.n245 G.t225 120.189
R1000 G.n205 G.t648 120.189
R1001 G.n168 G.t219 120.189
R1002 G.n134 G.t1019 120.189
R1003 G.n103 G.t585 120.189
R1004 G.n78 G.t289 120.189
R1005 G.n56 G.t957 120.189
R1006 G.n37 G.t651 120.189
R1007 G.n21 G.t223 120.189
R1008 G.n902 G.t1024 120.189
R1009 G.n901 G.t1009 120.189
R1010 G.n900 G.t715 120.189
R1011 G.n893 G.t822 120.189
R1012 G.n894 G.t1087 120.189
R1013 G.n11 G.t1101 120.189
R1014 G.n24 G.t325 120.189
R1015 G.n40 G.t734 120.189
R1016 G.n59 G.t1056 120.189
R1017 G.n81 G.t371 120.189
R1018 G.n106 G.t686 120.189
R1019 G.n137 G.t1098 120.189
R1020 G.n171 G.t321 120.189
R1021 G.n208 G.t731 120.189
R1022 G.n248 G.t329 120.189
R1023 G.n291 G.t368 120.189
R1024 G.n334 G.t1059 120.189
R1025 G.n377 G.t1096 120.189
R1026 G.n418 G.t692 120.189
R1027 G.n453 G.t729 120.189
R1028 G.n483 G.t326 120.189
R1029 G.n507 G.t366 120.189
R1030 G.n527 G.t877 120.189
R1031 G.n541 G.t162 120.189
R1032 G.n551 G.t508 120.189
R1033 G.n567 G.t897 120.189
R1034 G.n564 G.t354 120.189
R1035 G.n553 G.t119 120.189
R1036 G.n544 G.t931 120.189
R1037 G.n530 G.t694 120.189
R1038 G.n510 G.t747 120.189
R1039 G.n486 G.t203 120.189
R1040 G.n456 G.t234 120.189
R1041 G.n421 G.t843 120.189
R1042 G.n380 G.t871 120.189
R1043 G.n337 G.t314 120.189
R1044 G.n294 G.t341 120.189
R1045 G.n251 G.t902 120.189
R1046 G.n211 G.t919 120.189
R1047 G.n174 G.t679 120.189
R1048 G.n140 G.t453 120.189
R1049 G.n109 G.t168 120.189
R1050 G.n84 G.t1032 120.189
R1051 G.n62 G.t781 120.189
R1052 G.n43 G.t531 120.189
R1053 G.n27 G.t268 120.189
R1054 G.n14 G.t18 120.189
R1055 G.n4 G.t516 120.189
R1056 G.n889 G.t939 120.189
R1057 G.n3 G.t689 120.189
R1058 G.n0 G.t828 120.189
R1059 G.n10 G.t970 120.189
R1060 G.n7 G.t685 120.189
R1061 G.n20 G.t988 120.189
R1062 G.n17 G.t128 120.189
R1063 G.n33 G.t192 120.189
R1064 G.n30 G.t790 120.189
R1065 G.n49 G.t612 120.189
R1066 G.n46 G.t575 120.189
R1067 G.n68 G.t925 120.189
R1068 G.n65 G.t165 120.189
R1069 G.n90 G.t250 120.189
R1070 G.n87 G.t1081 120.189
R1071 G.n115 G.t556 120.189
R1072 G.n112 G.t657 120.189
R1073 G.n146 G.t985 120.189
R1074 G.n143 G.t502 120.189
R1075 G.n180 G.t190 120.189
R1076 G.n177 G.t56 120.189
R1077 G.n217 G.t607 120.189
R1078 G.n214 G.t948 120.189
R1079 G.n257 G.t199 120.189
R1080 G.n254 G.t849 120.189
R1081 G.n300 G.t247 120.189
R1082 G.n297 G.t353 120.189
R1083 G.n343 G.t930 120.189
R1084 G.n340 G.t195 120.189
R1085 G.n386 G.t981 120.189
R1086 G.n383 G.t868 120.189
R1087 G.n427 G.t561 120.189
R1088 G.n424 G.t701 120.189
R1089 G.n462 G.t604 120.189
R1090 G.n459 G.t217 120.189
R1091 G.n492 G.t196 120.189
R1092 G.n489 G.t108 120.189
R1093 G.n516 G.t243 120.189
R1094 G.n513 G.t717 120.189
R1095 G.n536 G.t733 120.189
R1096 G.n533 G.t672 120.189
R1097 G.n550 G.t59 120.189
R1098 G.n547 G.t513 120.189
R1099 G.n559 G.t370 120.189
R1100 G.n556 G.t76 120.189
R1101 G.n562 G.t795 120.189
R1102 G.n560 G.t968 120.189
R1103 G.n1678 G.t1069 120.189
R1104 G.n827 G.n826 0.686
R1105 G.n825 G.n824 0.686
R1106 G.n1642 G.n1638 0.686
R1107 G.n1627 G.n1620 0.686
R1108 G.n1609 G.n1599 0.686
R1109 G.n1588 G.n1575 0.686
R1110 G.n1564 G.n1549 0.686
R1111 G.n1538 G.n1522 0.686
R1112 G.n1511 G.n1497 0.686
R1113 G.n1486 G.n1472 0.686
R1114 G.n1461 G.n1450 0.686
R1115 G.n1439 G.n1431 0.686
R1116 G.n1420 G.n1413 0.686
R1117 G.n1402 G.n1397 0.686
R1118 G.n1386 G.n1384 0.686
R1119 G.n1373 G.n1372 0.686
R1120 G.n1307 G.n1306 0.686
R1121 G.n1310 G.n1308 0.686
R1122 G.n1313 G.n1311 0.686
R1123 G.n1316 G.n1314 0.686
R1124 G.n1319 G.n1317 0.686
R1125 G.n819 G.n818 0.686
R1126 G.n817 G.n816 0.686
R1127 G.n815 G.n814 0.686
R1128 G.n813 G.n812 0.686
R1129 G.n1293 G.n1292 0.686
R1130 G.n1295 G.n1294 0.686
R1131 G.n1297 G.n1296 0.686
R1132 G.n1299 G.n1298 0.686
R1133 G.n1301 G.n1300 0.686
R1134 G.n1303 G.n1302 0.686
R1135 G.n806 G.n805 0.686
R1136 G.n804 G.n803 0.686
R1137 G.n802 G.n801 0.686
R1138 G.n800 G.n799 0.686
R1139 G.n1604 G.n1600 0.686
R1140 G.n1583 G.n1576 0.686
R1141 G.n1559 G.n1550 0.686
R1142 G.n1533 G.n1523 0.686
R1143 G.n1506 G.n1498 0.686
R1144 G.n1481 G.n1473 0.686
R1145 G.n1456 G.n1451 0.686
R1146 G.n1434 G.n1432 0.686
R1147 G.n1415 G.n1414 0.686
R1148 G.n1269 G.n1268 0.686
R1149 G.n1271 G.n1270 0.686
R1150 G.n1273 G.n1272 0.686
R1151 G.n1275 G.n1274 0.686
R1152 G.n1277 G.n1276 0.686
R1153 G.n1279 G.n1278 0.686
R1154 G.n1281 G.n1280 0.686
R1155 G.n1283 G.n1282 0.686
R1156 G.n792 G.n791 0.686
R1157 G.n790 G.n789 0.686
R1158 G.n788 G.n787 0.686
R1159 G.n786 G.n785 0.686
R1160 G.n784 G.n783 0.686
R1161 G.n782 G.n781 0.686
R1162 G.n1242 G.n1241 0.686
R1163 G.n1244 G.n1243 0.686
R1164 G.n1246 G.n1245 0.686
R1165 G.n1248 G.n1247 0.686
R1166 G.n1250 G.n1249 0.686
R1167 G.n1252 G.n1251 0.686
R1168 G.n1254 G.n1253 0.686
R1169 G.n1256 G.n1255 0.686
R1170 G.n1258 G.n1257 0.686
R1171 G.n773 G.n772 0.686
R1172 G.n771 G.n770 0.686
R1173 G.n769 G.n768 0.686
R1174 G.n767 G.n766 0.686
R1175 G.n765 G.n764 0.686
R1176 G.n763 G.n762 0.686
R1177 G.n1554 G.n1551 0.686
R1178 G.n1528 G.n1524 0.686
R1179 G.n1501 G.n1499 0.686
R1180 G.n1476 G.n1474 0.686
R1181 G.n1209 G.n1208 0.686
R1182 G.n1211 G.n1210 0.686
R1183 G.n1213 G.n1212 0.686
R1184 G.n1215 G.n1214 0.686
R1185 G.n1217 G.n1216 0.686
R1186 G.n1219 G.n1218 0.686
R1187 G.n1221 G.n1220 0.686
R1188 G.n1223 G.n1222 0.686
R1189 G.n1225 G.n1224 0.686
R1190 G.n1227 G.n1226 0.686
R1191 G.n1229 G.n1228 0.686
R1192 G.n753 G.n752 0.686
R1193 G.n751 G.n750 0.686
R1194 G.n749 G.n748 0.686
R1195 G.n747 G.n746 0.686
R1196 G.n745 G.n744 0.686
R1197 G.n743 G.n742 0.686
R1198 G.n741 G.n740 0.686
R1199 G.n739 G.n738 0.686
R1200 G.n1173 G.n1172 0.686
R1201 G.n1175 G.n1174 0.686
R1202 G.n1177 G.n1176 0.686
R1203 G.n1179 G.n1178 0.686
R1204 G.n1181 G.n1180 0.686
R1205 G.n1183 G.n1182 0.686
R1206 G.n1185 G.n1184 0.686
R1207 G.n1187 G.n1186 0.686
R1208 G.n1189 G.n1188 0.686
R1209 G.n1191 G.n1190 0.686
R1210 G.n1193 G.n1192 0.686
R1211 G.n1195 G.n1194 0.686
R1212 G.n728 G.n727 0.686
R1213 G.n726 G.n725 0.686
R1214 G.n724 G.n723 0.686
R1215 G.n722 G.n721 0.686
R1216 G.n720 G.n719 0.686
R1217 G.n718 G.n717 0.686
R1218 G.n346 G.n345 0.686
R1219 G.n303 G.n302 0.686
R1220 G.n260 G.n259 0.686
R1221 G.n1136 G.n1135 0.686
R1222 G.n1138 G.n1137 0.686
R1223 G.n1140 G.n1139 0.686
R1224 G.n1142 G.n1141 0.686
R1225 G.n1144 G.n1143 0.686
R1226 G.n1146 G.n1145 0.686
R1227 G.n1148 G.n1147 0.686
R1228 G.n1150 G.n1149 0.686
R1229 G.n1152 G.n1151 0.686
R1230 G.n1154 G.n1153 0.686
R1231 G.n1156 G.n1155 0.686
R1232 G.n1158 G.n1157 0.686
R1233 G.n707 G.n706 0.686
R1234 G.n705 G.n704 0.686
R1235 G.n703 G.n702 0.686
R1236 G.n701 G.n700 0.686
R1237 G.n699 G.n698 0.686
R1238 G.n697 G.n696 0.686
R1239 G.n695 G.n694 0.686
R1240 G.n1102 G.n1101 0.686
R1241 G.n1104 G.n1103 0.686
R1242 G.n1106 G.n1105 0.686
R1243 G.n1108 G.n1107 0.686
R1244 G.n1110 G.n1109 0.686
R1245 G.n1112 G.n1111 0.686
R1246 G.n1114 G.n1113 0.686
R1247 G.n1116 G.n1115 0.686
R1248 G.n1118 G.n1117 0.686
R1249 G.n1120 G.n1119 0.686
R1250 G.n684 G.n683 0.686
R1251 G.n682 G.n681 0.686
R1252 G.n680 G.n679 0.686
R1253 G.n678 G.n677 0.686
R1254 G.n676 G.n675 0.686
R1255 G.n393 G.n392 0.686
R1256 G.n352 G.n351 0.686
R1257 G.n309 G.n308 0.686
R1258 G.n266 G.n265 0.686
R1259 G.n223 G.n222 0.686
R1260 G.n183 G.n182 0.686
R1261 G.n1069 G.n1068 0.686
R1262 G.n1071 G.n1070 0.686
R1263 G.n1073 G.n1072 0.686
R1264 G.n1075 G.n1074 0.686
R1265 G.n1077 G.n1076 0.686
R1266 G.n1079 G.n1078 0.686
R1267 G.n1081 G.n1080 0.686
R1268 G.n1083 G.n1082 0.686
R1269 G.n1085 G.n1084 0.686
R1270 G.n1087 G.n1086 0.686
R1271 G.n666 G.n665 0.686
R1272 G.n664 G.n663 0.686
R1273 G.n662 G.n661 0.686
R1274 G.n660 G.n659 0.686
R1275 G.n658 G.n657 0.686
R1276 G.n656 G.n655 0.686
R1277 G.n1041 G.n1040 0.686
R1278 G.n1043 G.n1042 0.686
R1279 G.n1045 G.n1044 0.686
R1280 G.n1047 G.n1046 0.686
R1281 G.n1049 G.n1048 0.686
R1282 G.n1051 G.n1050 0.686
R1283 G.n1053 G.n1052 0.686
R1284 G.n1055 G.n1054 0.686
R1285 G.n646 G.n645 0.686
R1286 G.n644 G.n643 0.686
R1287 G.n642 G.n641 0.686
R1288 G.n640 G.n639 0.686
R1289 G.n434 G.n433 0.686
R1290 G.n399 G.n398 0.686
R1291 G.n358 G.n357 0.686
R1292 G.n315 G.n314 0.686
R1293 G.n272 G.n271 0.686
R1294 G.n229 G.n228 0.686
R1295 G.n189 G.n188 0.686
R1296 G.n152 G.n151 0.686
R1297 G.n118 G.n117 0.686
R1298 G.n1014 G.n1013 0.686
R1299 G.n1016 G.n1015 0.686
R1300 G.n1018 G.n1017 0.686
R1301 G.n1020 G.n1019 0.686
R1302 G.n1022 G.n1021 0.686
R1303 G.n1024 G.n1023 0.686
R1304 G.n1026 G.n1025 0.686
R1305 G.n1028 G.n1027 0.686
R1306 G.n631 G.n630 0.686
R1307 G.n629 G.n628 0.686
R1308 G.n627 G.n626 0.686
R1309 G.n625 G.n624 0.686
R1310 G.n990 G.n989 0.686
R1311 G.n992 G.n991 0.686
R1312 G.n994 G.n993 0.686
R1313 G.n996 G.n995 0.686
R1314 G.n998 G.n997 0.686
R1315 G.n1000 G.n999 0.686
R1316 G.n1002 G.n1001 0.686
R1317 G.n615 G.n614 0.686
R1318 G.n613 G.n612 0.686
R1319 G.n611 G.n610 0.686
R1320 G.n470 G.n469 0.686
R1321 G.n440 G.n439 0.686
R1322 G.n405 G.n404 0.686
R1323 G.n364 G.n363 0.686
R1324 G.n321 G.n320 0.686
R1325 G.n278 G.n277 0.686
R1326 G.n235 G.n234 0.686
R1327 G.n195 G.n194 0.686
R1328 G.n158 G.n157 0.686
R1329 G.n124 G.n123 0.686
R1330 G.n93 G.n92 0.686
R1331 G.n966 G.n965 0.686
R1332 G.n968 G.n967 0.686
R1333 G.n970 G.n969 0.686
R1334 G.n972 G.n971 0.686
R1335 G.n974 G.n973 0.686
R1336 G.n976 G.n975 0.686
R1337 G.n978 G.n977 0.686
R1338 G.n603 G.n602 0.686
R1339 G.n601 G.n600 0.686
R1340 G.n599 G.n598 0.686
R1341 G.n947 G.n946 0.686
R1342 G.n949 G.n948 0.686
R1343 G.n951 G.n950 0.686
R1344 G.n953 G.n952 0.686
R1345 G.n955 G.n954 0.686
R1346 G.n592 G.n591 0.686
R1347 G.n590 G.n589 0.686
R1348 G.n500 G.n499 0.686
R1349 G.n476 G.n475 0.686
R1350 G.n446 G.n445 0.686
R1351 G.n411 G.n410 0.686
R1352 G.n370 G.n369 0.686
R1353 G.n327 G.n326 0.686
R1354 G.n284 G.n283 0.686
R1355 G.n241 G.n240 0.686
R1356 G.n201 G.n200 0.686
R1357 G.n164 G.n163 0.686
R1358 G.n130 G.n129 0.686
R1359 G.n99 G.n98 0.686
R1360 G.n74 G.n73 0.686
R1361 G.n52 G.n51 0.686
R1362 G.n929 G.n928 0.686
R1363 G.n931 G.n930 0.686
R1364 G.n933 G.n932 0.686
R1365 G.n935 G.n934 0.686
R1366 G.n937 G.n936 0.686
R1367 G.n583 G.n582 0.686
R1368 G.n581 G.n580 0.686
R1369 G.n916 G.n915 0.686
R1370 G.n918 G.n917 0.686
R1371 G.n920 G.n919 0.686
R1372 G.n575 G.n574 0.686
R1373 G.n526 G.n525 0.686
R1374 G.n506 G.n505 0.686
R1375 G.n482 G.n481 0.686
R1376 G.n452 G.n451 0.686
R1377 G.n417 G.n416 0.686
R1378 G.n376 G.n375 0.686
R1379 G.n333 G.n332 0.686
R1380 G.n290 G.n289 0.686
R1381 G.n247 G.n246 0.686
R1382 G.n207 G.n206 0.686
R1383 G.n170 G.n169 0.686
R1384 G.n136 G.n135 0.686
R1385 G.n105 G.n104 0.686
R1386 G.n80 G.n79 0.686
R1387 G.n58 G.n57 0.686
R1388 G.n39 G.n38 0.686
R1389 G.n23 G.n22 0.686
R1390 G.n904 G.n903 0.686
R1391 G.n906 G.n905 0.686
R1392 G.n908 G.n907 0.686
R1393 G.n569 G.n568 0.686
R1394 G.n897 G.n896 0.686
R1395 G.n555 G.n554 0.686
R1396 G.n546 G.n545 0.686
R1397 G.n532 G.n531 0.686
R1398 G.n512 G.n511 0.686
R1399 G.n488 G.n487 0.686
R1400 G.n458 G.n457 0.686
R1401 G.n423 G.n422 0.686
R1402 G.n382 G.n381 0.686
R1403 G.n339 G.n338 0.686
R1404 G.n296 G.n295 0.686
R1405 G.n253 G.n252 0.686
R1406 G.n213 G.n212 0.686
R1407 G.n176 G.n175 0.686
R1408 G.n142 G.n141 0.686
R1409 G.n111 G.n110 0.686
R1410 G.n86 G.n85 0.686
R1411 G.n64 G.n63 0.686
R1412 G.n45 G.n44 0.686
R1413 G.n29 G.n28 0.686
R1414 G.n16 G.n15 0.686
R1415 G.n6 G.n5 0.686
R1416 G.n891 G.n890 0.686
R1417 G.n558 G.n557 0.686
R1418 G.n549 G.n548 0.686
R1419 G.n535 G.n534 0.686
R1420 G.n515 G.n514 0.686
R1421 G.n491 G.n490 0.686
R1422 G.n461 G.n460 0.686
R1423 G.n426 G.n425 0.686
R1424 G.n385 G.n384 0.686
R1425 G.n342 G.n341 0.686
R1426 G.n299 G.n298 0.686
R1427 G.n256 G.n255 0.686
R1428 G.n216 G.n215 0.686
R1429 G.n179 G.n178 0.686
R1430 G.n145 G.n144 0.686
R1431 G.n114 G.n113 0.686
R1432 G.n89 G.n88 0.686
R1433 G.n67 G.n66 0.686
R1434 G.n48 G.n47 0.686
R1435 G.n32 G.n31 0.686
R1436 G.n19 G.n18 0.686
R1437 G.n9 G.n8 0.686
R1438 G.n2 G.n1 0.686
R1439 G.n543 G.n542 0.686
R1440 G.n529 G.n528 0.686
R1441 G.n509 G.n508 0.686
R1442 G.n485 G.n484 0.686
R1443 G.n455 G.n454 0.686
R1444 G.n420 G.n419 0.686
R1445 G.n379 G.n378 0.686
R1446 G.n336 G.n335 0.686
R1447 G.n293 G.n292 0.686
R1448 G.n250 G.n249 0.686
R1449 G.n210 G.n209 0.686
R1450 G.n173 G.n172 0.686
R1451 G.n139 G.n138 0.686
R1452 G.n108 G.n107 0.686
R1453 G.n83 G.n82 0.686
R1454 G.n61 G.n60 0.686
R1455 G.n42 G.n41 0.686
R1456 G.n26 G.n25 0.686
R1457 G.n13 G.n12 0.686
R1458 G.n896 G.n895 0.686
R1459 G.n898 G.n897 0.686
R1460 G.n907 G.n906 0.686
R1461 G.n905 G.n904 0.686
R1462 G.n574 G.n573 0.686
R1463 G.n576 G.n575 0.686
R1464 G.n582 G.n581 0.686
R1465 G.n523 G.n522 0.686
R1466 G.n503 G.n502 0.686
R1467 G.n479 G.n478 0.686
R1468 G.n449 G.n448 0.686
R1469 G.n414 G.n413 0.686
R1470 G.n373 G.n372 0.686
R1471 G.n330 G.n329 0.686
R1472 G.n287 G.n286 0.686
R1473 G.n244 G.n243 0.686
R1474 G.n204 G.n203 0.686
R1475 G.n167 G.n166 0.686
R1476 G.n133 G.n132 0.686
R1477 G.n102 G.n101 0.686
R1478 G.n77 G.n76 0.686
R1479 G.n55 G.n54 0.686
R1480 G.n36 G.n35 0.686
R1481 G.n915 G.n914 0.686
R1482 G.n917 G.n916 0.686
R1483 G.n919 G.n918 0.686
R1484 G.n921 G.n920 0.686
R1485 G.n936 G.n935 0.686
R1486 G.n934 G.n933 0.686
R1487 G.n932 G.n931 0.686
R1488 G.n930 G.n929 0.686
R1489 G.n589 G.n588 0.686
R1490 G.n591 G.n590 0.686
R1491 G.n593 G.n592 0.686
R1492 G.n602 G.n601 0.686
R1493 G.n600 G.n599 0.686
R1494 G.n497 G.n496 0.686
R1495 G.n473 G.n472 0.686
R1496 G.n443 G.n442 0.686
R1497 G.n408 G.n407 0.686
R1498 G.n367 G.n366 0.686
R1499 G.n324 G.n323 0.686
R1500 G.n281 G.n280 0.686
R1501 G.n238 G.n237 0.686
R1502 G.n198 G.n197 0.686
R1503 G.n161 G.n160 0.686
R1504 G.n127 G.n126 0.686
R1505 G.n96 G.n95 0.686
R1506 G.n71 G.n70 0.686
R1507 G.n946 G.n945 0.686
R1508 G.n948 G.n947 0.686
R1509 G.n950 G.n949 0.686
R1510 G.n952 G.n951 0.686
R1511 G.n954 G.n953 0.686
R1512 G.n956 G.n955 0.686
R1513 G.n977 G.n976 0.686
R1514 G.n975 G.n974 0.686
R1515 G.n973 G.n972 0.686
R1516 G.n971 G.n970 0.686
R1517 G.n969 G.n968 0.686
R1518 G.n967 G.n966 0.686
R1519 G.n610 G.n609 0.686
R1520 G.n612 G.n611 0.686
R1521 G.n614 G.n613 0.686
R1522 G.n616 G.n615 0.686
R1523 G.n630 G.n629 0.686
R1524 G.n628 G.n627 0.686
R1525 G.n626 G.n625 0.686
R1526 G.n624 G.n623 0.686
R1527 G.n467 G.n466 0.686
R1528 G.n437 G.n436 0.686
R1529 G.n402 G.n401 0.686
R1530 G.n361 G.n360 0.686
R1531 G.n318 G.n317 0.686
R1532 G.n275 G.n274 0.686
R1533 G.n232 G.n231 0.686
R1534 G.n192 G.n191 0.686
R1535 G.n155 G.n154 0.686
R1536 G.n121 G.n120 0.686
R1537 G.n989 G.n988 0.686
R1538 G.n991 G.n990 0.686
R1539 G.n993 G.n992 0.686
R1540 G.n995 G.n994 0.686
R1541 G.n997 G.n996 0.686
R1542 G.n999 G.n998 0.686
R1543 G.n1001 G.n1000 0.686
R1544 G.n1003 G.n1002 0.686
R1545 G.n1027 G.n1026 0.686
R1546 G.n1025 G.n1024 0.686
R1547 G.n1023 G.n1022 0.686
R1548 G.n1021 G.n1020 0.686
R1549 G.n1019 G.n1018 0.686
R1550 G.n1017 G.n1016 0.686
R1551 G.n1015 G.n1014 0.686
R1552 G.n639 G.n638 0.686
R1553 G.n641 G.n640 0.686
R1554 G.n643 G.n642 0.686
R1555 G.n645 G.n644 0.686
R1556 G.n647 G.n646 0.686
R1557 G.n665 G.n664 0.686
R1558 G.n663 G.n662 0.686
R1559 G.n661 G.n660 0.686
R1560 G.n659 G.n658 0.686
R1561 G.n657 G.n656 0.686
R1562 G.n396 G.n395 0.686
R1563 G.n355 G.n354 0.686
R1564 G.n312 G.n311 0.686
R1565 G.n269 G.n268 0.686
R1566 G.n226 G.n225 0.686
R1567 G.n186 G.n185 0.686
R1568 G.n149 G.n148 0.686
R1569 G.n1040 G.n1039 0.686
R1570 G.n1042 G.n1041 0.686
R1571 G.n1044 G.n1043 0.686
R1572 G.n1046 G.n1045 0.686
R1573 G.n1048 G.n1047 0.686
R1574 G.n1050 G.n1049 0.686
R1575 G.n1052 G.n1051 0.686
R1576 G.n1054 G.n1053 0.686
R1577 G.n1056 G.n1055 0.686
R1578 G.n1086 G.n1085 0.686
R1579 G.n1084 G.n1083 0.686
R1580 G.n1082 G.n1081 0.686
R1581 G.n1080 G.n1079 0.686
R1582 G.n1078 G.n1077 0.686
R1583 G.n1076 G.n1075 0.686
R1584 G.n1074 G.n1073 0.686
R1585 G.n1072 G.n1071 0.686
R1586 G.n1070 G.n1069 0.686
R1587 G.n675 G.n674 0.686
R1588 G.n677 G.n676 0.686
R1589 G.n679 G.n678 0.686
R1590 G.n681 G.n680 0.686
R1591 G.n683 G.n682 0.686
R1592 G.n685 G.n684 0.686
R1593 G.n706 G.n705 0.686
R1594 G.n704 G.n703 0.686
R1595 G.n702 G.n701 0.686
R1596 G.n700 G.n699 0.686
R1597 G.n698 G.n697 0.686
R1598 G.n696 G.n695 0.686
R1599 G.n349 G.n348 0.686
R1600 G.n306 G.n305 0.686
R1601 G.n263 G.n262 0.686
R1602 G.n220 G.n219 0.686
R1603 G.n1101 G.n1100 0.686
R1604 G.n1103 G.n1102 0.686
R1605 G.n1105 G.n1104 0.686
R1606 G.n1107 G.n1106 0.686
R1607 G.n1109 G.n1108 0.686
R1608 G.n1111 G.n1110 0.686
R1609 G.n1113 G.n1112 0.686
R1610 G.n1115 G.n1114 0.686
R1611 G.n1117 G.n1116 0.686
R1612 G.n1119 G.n1118 0.686
R1613 G.n1121 G.n1120 0.686
R1614 G.n1157 G.n1156 0.686
R1615 G.n1155 G.n1154 0.686
R1616 G.n1153 G.n1152 0.686
R1617 G.n1151 G.n1150 0.686
R1618 G.n1149 G.n1148 0.686
R1619 G.n1147 G.n1146 0.686
R1620 G.n1145 G.n1144 0.686
R1621 G.n1143 G.n1142 0.686
R1622 G.n1141 G.n1140 0.686
R1623 G.n1139 G.n1138 0.686
R1624 G.n1137 G.n1136 0.686
R1625 G.n717 G.n716 0.686
R1626 G.n719 G.n718 0.686
R1627 G.n721 G.n720 0.686
R1628 G.n723 G.n722 0.686
R1629 G.n725 G.n724 0.686
R1630 G.n727 G.n726 0.686
R1631 G.n729 G.n728 0.686
R1632 G.n752 G.n751 0.686
R1633 G.n750 G.n749 0.686
R1634 G.n748 G.n747 0.686
R1635 G.n746 G.n745 0.686
R1636 G.n744 G.n743 0.686
R1637 G.n742 G.n741 0.686
R1638 G.n740 G.n739 0.686
R1639 G.n1526 G.n1525 0.686
R1640 G.n1172 G.n1171 0.686
R1641 G.n1174 G.n1173 0.686
R1642 G.n1176 G.n1175 0.686
R1643 G.n1178 G.n1177 0.686
R1644 G.n1180 G.n1179 0.686
R1645 G.n1182 G.n1181 0.686
R1646 G.n1184 G.n1183 0.686
R1647 G.n1186 G.n1185 0.686
R1648 G.n1188 G.n1187 0.686
R1649 G.n1190 G.n1189 0.686
R1650 G.n1192 G.n1191 0.686
R1651 G.n1194 G.n1193 0.686
R1652 G.n1196 G.n1195 0.686
R1653 G.n1228 G.n1227 0.686
R1654 G.n1226 G.n1225 0.686
R1655 G.n1224 G.n1223 0.686
R1656 G.n1222 G.n1221 0.686
R1657 G.n1220 G.n1219 0.686
R1658 G.n1218 G.n1217 0.686
R1659 G.n1216 G.n1215 0.686
R1660 G.n1214 G.n1213 0.686
R1661 G.n1212 G.n1211 0.686
R1662 G.n1210 G.n1209 0.686
R1663 G.n762 G.n761 0.686
R1664 G.n764 G.n763 0.686
R1665 G.n766 G.n765 0.686
R1666 G.n768 G.n767 0.686
R1667 G.n770 G.n769 0.686
R1668 G.n772 G.n771 0.686
R1669 G.n774 G.n773 0.686
R1670 G.n791 G.n790 0.686
R1671 G.n789 G.n788 0.686
R1672 G.n787 G.n786 0.686
R1673 G.n785 G.n784 0.686
R1674 G.n783 G.n782 0.686
R1675 G.n1581 G.n1580 0.686
R1676 G.n1557 G.n1556 0.686
R1677 G.n1531 G.n1530 0.686
R1678 G.n1504 G.n1503 0.686
R1679 G.n1479 G.n1478 0.686
R1680 G.n1454 G.n1453 0.686
R1681 G.n1241 G.n1240 0.686
R1682 G.n1243 G.n1242 0.686
R1683 G.n1245 G.n1244 0.686
R1684 G.n1247 G.n1246 0.686
R1685 G.n1249 G.n1248 0.686
R1686 G.n1251 G.n1250 0.686
R1687 G.n1253 G.n1252 0.686
R1688 G.n1255 G.n1254 0.686
R1689 G.n1257 G.n1256 0.686
R1690 G.n1259 G.n1258 0.686
R1691 G.n1282 G.n1281 0.686
R1692 G.n1280 G.n1279 0.686
R1693 G.n1278 G.n1277 0.686
R1694 G.n1276 G.n1275 0.686
R1695 G.n1274 G.n1273 0.686
R1696 G.n1272 G.n1271 0.686
R1697 G.n1270 G.n1269 0.686
R1698 G.n799 G.n798 0.686
R1699 G.n801 G.n800 0.686
R1700 G.n803 G.n802 0.686
R1701 G.n805 G.n804 0.686
R1702 G.n807 G.n806 0.686
R1703 G.n818 G.n817 0.686
R1704 G.n816 G.n815 0.686
R1705 G.n814 G.n813 0.686
R1706 G.n1625 G.n1624 0.686
R1707 G.n1607 G.n1606 0.686
R1708 G.n1586 G.n1585 0.686
R1709 G.n1562 G.n1561 0.686
R1710 G.n1536 G.n1535 0.686
R1711 G.n1509 G.n1508 0.686
R1712 G.n1484 G.n1483 0.686
R1713 G.n1459 G.n1458 0.686
R1714 G.n1437 G.n1436 0.686
R1715 G.n1418 G.n1417 0.686
R1716 G.n1400 G.n1399 0.686
R1717 G.n1292 G.n1291 0.686
R1718 G.n1294 G.n1293 0.686
R1719 G.n1296 G.n1295 0.686
R1720 G.n1298 G.n1297 0.686
R1721 G.n1300 G.n1299 0.686
R1722 G.n1302 G.n1301 0.686
R1723 G.n1304 G.n1303 0.686
R1724 G.n1317 G.n1316 0.686
R1725 G.n1314 G.n1313 0.686
R1726 G.n1311 G.n1310 0.686
R1727 G.n1308 G.n1307 0.686
R1728 G.n824 G.n823 0.686
R1729 G.n826 G.n825 0.686
R1730 G.n828 G.n827 0.686
R1731 G.n834 G.n833 0.686
R1732 G.n833 G.n831 0.686
R1733 G.n1644 G.n1637 0.686
R1734 G.n1629 G.n1619 0.686
R1735 G.n1611 G.n1598 0.686
R1736 G.n1590 G.n1574 0.686
R1737 G.n1566 G.n1548 0.686
R1738 G.n1540 G.n1521 0.686
R1739 G.n1513 G.n1496 0.686
R1740 G.n1488 G.n1471 0.686
R1741 G.n1463 G.n1449 0.686
R1742 G.n1441 G.n1430 0.686
R1743 G.n1422 G.n1412 0.686
R1744 G.n1404 G.n1396 0.686
R1745 G.n1388 G.n1383 0.686
R1746 G.n1375 G.n1371 0.686
R1747 G.n1363 G.n1361 0.686
R1748 G.n1323 G.n1322 0.686
R1749 G.n1326 G.n1324 0.686
R1750 G.n1327 G.n1326 0.686
R1751 G.n1331 G.n1329 0.686
R1752 G.n835 G.n834 0.686
R1753 G.n1656 G.n1655 0.686
R1754 G.n1324 G.n1323 0.686
R1755 G.n1328 G.n1327 0.686
R1756 G.n1329 G.n1328 0.686
R1757 G.n1667 G.n1663 0.686
R1758 G.n1658 G.n1651 0.686
R1759 G.n1646 G.n1636 0.686
R1760 G.n1631 G.n1618 0.686
R1761 G.n1613 G.n1597 0.686
R1762 G.n1592 G.n1573 0.686
R1763 G.n1568 G.n1547 0.686
R1764 G.n1542 G.n1520 0.686
R1765 G.n1515 G.n1495 0.686
R1766 G.n1490 G.n1470 0.686
R1767 G.n1465 G.n1448 0.686
R1768 G.n1443 G.n1429 0.686
R1769 G.n1424 G.n1411 0.686
R1770 G.n1406 G.n1395 0.686
R1771 G.n1390 G.n1382 0.686
R1772 G.n1377 G.n1370 0.686
R1773 G.n1365 G.n1360 0.686
R1774 G.n1355 G.n1353 0.686
R1775 G.n1348 G.n1347 0.686
R1776 G.n1335 G.n1334 0.686
R1777 G.n1337 G.n1336 0.686
R1778 G.n1675 G.n1674 0.686
R1779 G.n1670 G.n1669 0.686
R1780 G.n1661 G.n1660 0.686
R1781 G.n1649 G.n1648 0.686
R1782 G.n1634 G.n1633 0.686
R1783 G.n1616 G.n1615 0.686
R1784 G.n1595 G.n1594 0.686
R1785 G.n1571 G.n1570 0.686
R1786 G.n1545 G.n1544 0.686
R1787 G.n1518 G.n1517 0.686
R1788 G.n1493 G.n1492 0.686
R1789 G.n1468 G.n1467 0.686
R1790 G.n1446 G.n1445 0.686
R1791 G.n1427 G.n1426 0.686
R1792 G.n1409 G.n1408 0.686
R1793 G.n1393 G.n1392 0.686
R1794 G.n1380 G.n1379 0.686
R1795 G.n1368 G.n1367 0.686
R1796 G.n1358 G.n1357 0.686
R1797 G.n1351 G.n1350 0.686
R1798 G.n1345 G.n1344 0.686
R1799 G.n1340 G.n1339 0.686
R1800 G.n1336 G.n1335 0.686
R1801 G.n839 G.n838 0.686
R1802 G.n829 G.n828 0.655
R1803 G.n1320 G.n1319 0.655
R1804 G.n846 G.n820 0.655
R1805 G.n1305 G.n1304 0.655
R1806 G.n808 G.n807 0.655
R1807 G.n1284 G.n1283 0.655
R1808 G.n848 G.n793 0.655
R1809 G.n1260 G.n1259 0.655
R1810 G.n775 G.n774 0.655
R1811 G.n1230 G.n1229 0.655
R1812 G.n850 G.n754 0.655
R1813 G.n1197 G.n1196 0.655
R1814 G.n730 G.n729 0.655
R1815 G.n1159 G.n1158 0.655
R1816 G.n852 G.n708 0.655
R1817 G.n1122 G.n1121 0.655
R1818 G.n686 G.n685 0.655
R1819 G.n1088 G.n1087 0.655
R1820 G.n854 G.n667 0.655
R1821 G.n1057 G.n1056 0.655
R1822 G.n648 G.n647 0.655
R1823 G.n1029 G.n1028 0.655
R1824 G.n856 G.n632 0.655
R1825 G.n1004 G.n1003 0.655
R1826 G.n617 G.n616 0.655
R1827 G.n979 G.n978 0.655
R1828 G.n858 G.n604 0.655
R1829 G.n957 G.n956 0.655
R1830 G.n594 G.n593 0.655
R1831 G.n938 G.n937 0.655
R1832 G.n860 G.n584 0.655
R1833 G.n922 G.n921 0.655
R1834 G.n577 G.n576 0.655
R1835 G.n909 G.n908 0.655
R1836 G.n862 G.n570 0.655
R1837 G.n899 G.n898 0.655
R1838 G.n566 G.n565 0.655
R1839 G.n892 G.n891 0.655
R1840 G.n864 G.n563 0.655
R1841 G.n1724 G.n888 0.655
R1842 G.n1723 G.n892 0.655
R1843 G.n863 G.n566 0.655
R1844 G.n570 G.n569 0.655
R1845 G.n1722 G.n899 0.655
R1846 G.n1721 G.n909 0.655
R1847 G.n861 G.n577 0.655
R1848 G.n584 G.n583 0.655
R1849 G.n1720 G.n922 0.655
R1850 G.n1719 G.n938 0.655
R1851 G.n859 G.n594 0.655
R1852 G.n604 G.n603 0.655
R1853 G.n1718 G.n957 0.655
R1854 G.n1717 G.n979 0.655
R1855 G.n857 G.n617 0.655
R1856 G.n632 G.n631 0.655
R1857 G.n1716 G.n1004 0.655
R1858 G.n1715 G.n1029 0.655
R1859 G.n855 G.n648 0.655
R1860 G.n667 G.n666 0.655
R1861 G.n1714 G.n1057 0.655
R1862 G.n1713 G.n1088 0.655
R1863 G.n853 G.n686 0.655
R1864 G.n708 G.n707 0.655
R1865 G.n1712 G.n1122 0.655
R1866 G.n1711 G.n1159 0.655
R1867 G.n851 G.n730 0.655
R1868 G.n754 G.n753 0.655
R1869 G.n1710 G.n1197 0.655
R1870 G.n1709 G.n1230 0.655
R1871 G.n849 G.n775 0.655
R1872 G.n793 G.n792 0.655
R1873 G.n1708 G.n1260 0.655
R1874 G.n1707 G.n1284 0.655
R1875 G.n847 G.n808 0.655
R1876 G.n820 G.n819 0.655
R1877 G.n1706 G.n1305 0.655
R1878 G.n1332 G.n1331 0.655
R1879 G.n1705 G.n1320 0.655
R1880 G.n845 G.n829 0.655
R1881 G.n836 G.n835 0.655
R1882 G.n844 G.n836 0.655
R1883 G.n1704 G.n1332 0.655
R1884 G.n840 G.n839 0.655
R1885 G.n1338 G.n1337 0.655
R1886 G.n842 G.n841 0.655
R1887 G.n1341 G.n1340 0.655
R1888 G.n1702 G.n1341 0.655
R1889 G.n1703 G.n1338 0.655
R1890 G.n843 G.n840 0.655
R1891 G.n1702 G.n1701 0.645
R1892 G.n865 G.n864 0.644
R1893 G.n839 G.n837 0.624
R1894 G.n1337 G.n1333 0.624
R1895 G.n1701 G.n1342 0.624
R1896 G.n1700 G.n1346 0.624
R1897 G.n1349 G.n1348 0.624
R1898 G.n1699 G.n1352 0.624
R1899 G.n1356 G.n1355 0.624
R1900 G.n1698 G.n1359 0.624
R1901 G.n1366 G.n1365 0.624
R1902 G.n1697 G.n1369 0.624
R1903 G.n1378 G.n1377 0.624
R1904 G.n1696 G.n1381 0.624
R1905 G.n1391 G.n1390 0.624
R1906 G.n1695 G.n1394 0.624
R1907 G.n1407 G.n1406 0.624
R1908 G.n1694 G.n1410 0.624
R1909 G.n1425 G.n1424 0.624
R1910 G.n1693 G.n1428 0.624
R1911 G.n1444 G.n1443 0.624
R1912 G.n1692 G.n1447 0.624
R1913 G.n1466 G.n1465 0.624
R1914 G.n1691 G.n1469 0.624
R1915 G.n1491 G.n1490 0.624
R1916 G.n1690 G.n1494 0.624
R1917 G.n1516 G.n1515 0.624
R1918 G.n1689 G.n1519 0.624
R1919 G.n1543 G.n1542 0.624
R1920 G.n1688 G.n1546 0.624
R1921 G.n1569 G.n1568 0.624
R1922 G.n1687 G.n1572 0.624
R1923 G.n1593 G.n1592 0.624
R1924 G.n1686 G.n1596 0.624
R1925 G.n1614 G.n1613 0.624
R1926 G.n1685 G.n1617 0.624
R1927 G.n1632 G.n1631 0.624
R1928 G.n1684 G.n1635 0.624
R1929 G.n1647 G.n1646 0.624
R1930 G.n1683 G.n1650 0.624
R1931 G.n1659 G.n1658 0.624
R1932 G.n1682 G.n1662 0.624
R1933 G.n1668 G.n1667 0.624
R1934 G.n1681 G.n1671 0.624
R1935 G.n1673 G.n1672 0.624
R1936 G.n1680 G.n1676 0.624
R1937 G.n1676 G.n1675 0.624
R1938 G.n1678 G.n1677 0.624
R1939 G.n1671 G.n1670 0.624
R1940 G.n1662 G.n1661 0.624
R1941 G.n1650 G.n1649 0.624
R1942 G.n1635 G.n1634 0.624
R1943 G.n1617 G.n1616 0.624
R1944 G.n1596 G.n1595 0.624
R1945 G.n1572 G.n1571 0.624
R1946 G.n1546 G.n1545 0.624
R1947 G.n1519 G.n1518 0.624
R1948 G.n1494 G.n1493 0.624
R1949 G.n1469 G.n1468 0.624
R1950 G.n1447 G.n1446 0.624
R1951 G.n1428 G.n1427 0.624
R1952 G.n1410 G.n1409 0.624
R1953 G.n1394 G.n1393 0.624
R1954 G.n1381 G.n1380 0.624
R1955 G.n1369 G.n1368 0.624
R1956 G.n1359 G.n1358 0.624
R1957 G.n1352 G.n1351 0.624
R1958 G.n1346 G.n1345 0.624
R1959 G.n1675 G.n1673 0.624
R1960 G.n1670 G.n1668 0.624
R1961 G.n1661 G.n1659 0.624
R1962 G.n1649 G.n1647 0.624
R1963 G.n1634 G.n1632 0.624
R1964 G.n1616 G.n1614 0.624
R1965 G.n1595 G.n1593 0.624
R1966 G.n1571 G.n1569 0.624
R1967 G.n1545 G.n1543 0.624
R1968 G.n1518 G.n1516 0.624
R1969 G.n1493 G.n1491 0.624
R1970 G.n1468 G.n1466 0.624
R1971 G.n1446 G.n1444 0.624
R1972 G.n1427 G.n1425 0.624
R1973 G.n1409 G.n1407 0.624
R1974 G.n1393 G.n1391 0.624
R1975 G.n1380 G.n1378 0.624
R1976 G.n1368 G.n1366 0.624
R1977 G.n1358 G.n1356 0.624
R1978 G.n1351 G.n1349 0.624
R1979 G.n1658 G.n1657 0.624
R1980 G.n1646 G.n1645 0.624
R1981 G.n1631 G.n1630 0.624
R1982 G.n1613 G.n1612 0.624
R1983 G.n1592 G.n1591 0.624
R1984 G.n1568 G.n1567 0.624
R1985 G.n1542 G.n1541 0.624
R1986 G.n1515 G.n1514 0.624
R1987 G.n1490 G.n1489 0.624
R1988 G.n1465 G.n1464 0.624
R1989 G.n1443 G.n1442 0.624
R1990 G.n1424 G.n1423 0.624
R1991 G.n1406 G.n1405 0.624
R1992 G.n1390 G.n1389 0.624
R1993 G.n1377 G.n1376 0.624
R1994 G.n1365 G.n1364 0.624
R1995 G.n1355 G.n1354 0.624
R1996 G.n1667 G.n1666 0.624
R1997 G.n1331 G.n1330 0.624
R1998 G.n1328 G.n1321 0.624
R1999 G.n1326 G.n1325 0.624
R2000 G.n1364 G.n1363 0.624
R2001 G.n1376 G.n1375 0.624
R2002 G.n1389 G.n1388 0.624
R2003 G.n1405 G.n1404 0.624
R2004 G.n1423 G.n1422 0.624
R2005 G.n1442 G.n1441 0.624
R2006 G.n1464 G.n1463 0.624
R2007 G.n1489 G.n1488 0.624
R2008 G.n1514 G.n1513 0.624
R2009 G.n1541 G.n1540 0.624
R2010 G.n1567 G.n1566 0.624
R2011 G.n1591 G.n1590 0.624
R2012 G.n1612 G.n1611 0.624
R2013 G.n1630 G.n1629 0.624
R2014 G.n1645 G.n1644 0.624
R2015 G.n1657 G.n1656 0.624
R2016 G.n1666 G.n1665 0.624
R2017 G.n833 G.n832 0.624
R2018 G.n835 G.n830 0.624
R2019 G.n1665 G.n1664 0.624
R2020 G.n1656 G.n1654 0.624
R2021 G.n1644 G.n1643 0.624
R2022 G.n1629 G.n1628 0.624
R2023 G.n1611 G.n1610 0.624
R2024 G.n1590 G.n1589 0.624
R2025 G.n1566 G.n1565 0.624
R2026 G.n1540 G.n1539 0.624
R2027 G.n1513 G.n1512 0.624
R2028 G.n1488 G.n1487 0.624
R2029 G.n1463 G.n1462 0.624
R2030 G.n1441 G.n1440 0.624
R2031 G.n1422 G.n1421 0.624
R2032 G.n1404 G.n1403 0.624
R2033 G.n1388 G.n1387 0.624
R2034 G.n1375 G.n1374 0.624
R2035 G.n1363 G.n1362 0.624
R2036 G.n1304 G.n1285 0.624
R2037 G.n1302 G.n1286 0.624
R2038 G.n1300 G.n1287 0.624
R2039 G.n1298 G.n1288 0.624
R2040 G.n1296 G.n1289 0.624
R2041 G.n1294 G.n1290 0.624
R2042 G.n1401 G.n1400 0.624
R2043 G.n1419 G.n1418 0.624
R2044 G.n1438 G.n1437 0.624
R2045 G.n1460 G.n1459 0.624
R2046 G.n1485 G.n1484 0.624
R2047 G.n1510 G.n1509 0.624
R2048 G.n1537 G.n1536 0.624
R2049 G.n1563 G.n1562 0.624
R2050 G.n1587 G.n1586 0.624
R2051 G.n1608 G.n1607 0.624
R2052 G.n1626 G.n1625 0.624
R2053 G.n1641 G.n1640 0.624
R2054 G.n815 G.n811 0.624
R2055 G.n817 G.n810 0.624
R2056 G.n819 G.n809 0.624
R2057 G.n807 G.n794 0.624
R2058 G.n805 G.n795 0.624
R2059 G.n803 G.n796 0.624
R2060 G.n801 G.n797 0.624
R2061 G.n1623 G.n1622 0.624
R2062 G.n1605 G.n1604 0.624
R2063 G.n1584 G.n1583 0.624
R2064 G.n1560 G.n1559 0.624
R2065 G.n1534 G.n1533 0.624
R2066 G.n1507 G.n1506 0.624
R2067 G.n1482 G.n1481 0.624
R2068 G.n1457 G.n1456 0.624
R2069 G.n1435 G.n1434 0.624
R2070 G.n1416 G.n1415 0.624
R2071 G.n1271 G.n1267 0.624
R2072 G.n1273 G.n1266 0.624
R2073 G.n1275 G.n1265 0.624
R2074 G.n1277 G.n1264 0.624
R2075 G.n1279 G.n1263 0.624
R2076 G.n1281 G.n1262 0.624
R2077 G.n1283 G.n1261 0.624
R2078 G.n1259 G.n1231 0.624
R2079 G.n1257 G.n1232 0.624
R2080 G.n1255 G.n1233 0.624
R2081 G.n1253 G.n1234 0.624
R2082 G.n1251 G.n1235 0.624
R2083 G.n1249 G.n1236 0.624
R2084 G.n1247 G.n1237 0.624
R2085 G.n1245 G.n1238 0.624
R2086 G.n1243 G.n1239 0.624
R2087 G.n1455 G.n1454 0.624
R2088 G.n1480 G.n1479 0.624
R2089 G.n1505 G.n1504 0.624
R2090 G.n1532 G.n1531 0.624
R2091 G.n1558 G.n1557 0.624
R2092 G.n1582 G.n1581 0.624
R2093 G.n1603 G.n1602 0.624
R2094 G.n784 G.n780 0.624
R2095 G.n786 G.n779 0.624
R2096 G.n788 G.n778 0.624
R2097 G.n790 G.n777 0.624
R2098 G.n792 G.n776 0.624
R2099 G.n774 G.n755 0.624
R2100 G.n772 G.n756 0.624
R2101 G.n770 G.n757 0.624
R2102 G.n768 G.n758 0.624
R2103 G.n766 G.n759 0.624
R2104 G.n764 G.n760 0.624
R2105 G.n1579 G.n1578 0.624
R2106 G.n1555 G.n1554 0.624
R2107 G.n1529 G.n1528 0.624
R2108 G.n1502 G.n1501 0.624
R2109 G.n1477 G.n1476 0.624
R2110 G.n1211 G.n1207 0.624
R2111 G.n1213 G.n1206 0.624
R2112 G.n1215 G.n1205 0.624
R2113 G.n1217 G.n1204 0.624
R2114 G.n1219 G.n1203 0.624
R2115 G.n1221 G.n1202 0.624
R2116 G.n1223 G.n1201 0.624
R2117 G.n1225 G.n1200 0.624
R2118 G.n1227 G.n1199 0.624
R2119 G.n1229 G.n1198 0.624
R2120 G.n1196 G.n1160 0.624
R2121 G.n1194 G.n1161 0.624
R2122 G.n1192 G.n1162 0.624
R2123 G.n1190 G.n1163 0.624
R2124 G.n1188 G.n1164 0.624
R2125 G.n1186 G.n1165 0.624
R2126 G.n1184 G.n1166 0.624
R2127 G.n1182 G.n1167 0.624
R2128 G.n1180 G.n1168 0.624
R2129 G.n1178 G.n1169 0.624
R2130 G.n1176 G.n1170 0.624
R2131 G.n1527 G.n1526 0.624
R2132 G.n1553 G.n1552 0.624
R2133 G.n741 G.n737 0.624
R2134 G.n743 G.n736 0.624
R2135 G.n745 G.n735 0.624
R2136 G.n747 G.n734 0.624
R2137 G.n749 G.n733 0.624
R2138 G.n751 G.n732 0.624
R2139 G.n753 G.n731 0.624
R2140 G.n729 G.n709 0.624
R2141 G.n727 G.n710 0.624
R2142 G.n725 G.n711 0.624
R2143 G.n723 G.n712 0.624
R2144 G.n721 G.n713 0.624
R2145 G.n719 G.n714 0.624
R2146 G.n717 G.n715 0.624
R2147 G.n388 G.n387 0.624
R2148 G.n346 G.n344 0.624
R2149 G.n303 G.n301 0.624
R2150 G.n260 G.n258 0.624
R2151 G.n1136 G.n1134 0.624
R2152 G.n1138 G.n1133 0.624
R2153 G.n1140 G.n1132 0.624
R2154 G.n1142 G.n1131 0.624
R2155 G.n1144 G.n1130 0.624
R2156 G.n1146 G.n1129 0.624
R2157 G.n1148 G.n1128 0.624
R2158 G.n1150 G.n1127 0.624
R2159 G.n1152 G.n1126 0.624
R2160 G.n1154 G.n1125 0.624
R2161 G.n1156 G.n1124 0.624
R2162 G.n1158 G.n1123 0.624
R2163 G.n1121 G.n1089 0.624
R2164 G.n1119 G.n1090 0.624
R2165 G.n1117 G.n1091 0.624
R2166 G.n1115 G.n1092 0.624
R2167 G.n1113 G.n1093 0.624
R2168 G.n1111 G.n1094 0.624
R2169 G.n1109 G.n1095 0.624
R2170 G.n1107 G.n1096 0.624
R2171 G.n1105 G.n1097 0.624
R2172 G.n1103 G.n1098 0.624
R2173 G.n1101 G.n1099 0.624
R2174 G.n220 G.n218 0.624
R2175 G.n263 G.n261 0.624
R2176 G.n306 G.n304 0.624
R2177 G.n349 G.n347 0.624
R2178 G.n390 G.n389 0.624
R2179 G.n695 G.n693 0.624
R2180 G.n697 G.n692 0.624
R2181 G.n699 G.n691 0.624
R2182 G.n701 G.n690 0.624
R2183 G.n703 G.n689 0.624
R2184 G.n705 G.n688 0.624
R2185 G.n707 G.n687 0.624
R2186 G.n685 G.n668 0.624
R2187 G.n683 G.n669 0.624
R2188 G.n681 G.n670 0.624
R2189 G.n679 G.n671 0.624
R2190 G.n677 G.n672 0.624
R2191 G.n675 G.n673 0.624
R2192 G.n429 G.n428 0.624
R2193 G.n393 G.n391 0.624
R2194 G.n352 G.n350 0.624
R2195 G.n309 G.n307 0.624
R2196 G.n266 G.n264 0.624
R2197 G.n223 G.n221 0.624
R2198 G.n183 G.n181 0.624
R2199 G.n1069 G.n1067 0.624
R2200 G.n1071 G.n1066 0.624
R2201 G.n1073 G.n1065 0.624
R2202 G.n1075 G.n1064 0.624
R2203 G.n1077 G.n1063 0.624
R2204 G.n1079 G.n1062 0.624
R2205 G.n1081 G.n1061 0.624
R2206 G.n1083 G.n1060 0.624
R2207 G.n1085 G.n1059 0.624
R2208 G.n1087 G.n1058 0.624
R2209 G.n1056 G.n1030 0.624
R2210 G.n1054 G.n1031 0.624
R2211 G.n1052 G.n1032 0.624
R2212 G.n1050 G.n1033 0.624
R2213 G.n1048 G.n1034 0.624
R2214 G.n1046 G.n1035 0.624
R2215 G.n1044 G.n1036 0.624
R2216 G.n1042 G.n1037 0.624
R2217 G.n1040 G.n1038 0.624
R2218 G.n149 G.n147 0.624
R2219 G.n186 G.n184 0.624
R2220 G.n226 G.n224 0.624
R2221 G.n269 G.n267 0.624
R2222 G.n312 G.n310 0.624
R2223 G.n355 G.n353 0.624
R2224 G.n396 G.n394 0.624
R2225 G.n431 G.n430 0.624
R2226 G.n656 G.n654 0.624
R2227 G.n658 G.n653 0.624
R2228 G.n660 G.n652 0.624
R2229 G.n662 G.n651 0.624
R2230 G.n664 G.n650 0.624
R2231 G.n666 G.n649 0.624
R2232 G.n647 G.n633 0.624
R2233 G.n645 G.n634 0.624
R2234 G.n643 G.n635 0.624
R2235 G.n641 G.n636 0.624
R2236 G.n639 G.n637 0.624
R2237 G.n464 G.n463 0.624
R2238 G.n434 G.n432 0.624
R2239 G.n399 G.n397 0.624
R2240 G.n358 G.n356 0.624
R2241 G.n315 G.n313 0.624
R2242 G.n272 G.n270 0.624
R2243 G.n229 G.n227 0.624
R2244 G.n189 G.n187 0.624
R2245 G.n152 G.n150 0.624
R2246 G.n118 G.n116 0.624
R2247 G.n1014 G.n1012 0.624
R2248 G.n1016 G.n1011 0.624
R2249 G.n1018 G.n1010 0.624
R2250 G.n1020 G.n1009 0.624
R2251 G.n1022 G.n1008 0.624
R2252 G.n1024 G.n1007 0.624
R2253 G.n1026 G.n1006 0.624
R2254 G.n1028 G.n1005 0.624
R2255 G.n1003 G.n980 0.624
R2256 G.n1001 G.n981 0.624
R2257 G.n999 G.n982 0.624
R2258 G.n997 G.n983 0.624
R2259 G.n995 G.n984 0.624
R2260 G.n993 G.n985 0.624
R2261 G.n991 G.n986 0.624
R2262 G.n989 G.n987 0.624
R2263 G.n121 G.n119 0.624
R2264 G.n155 G.n153 0.624
R2265 G.n192 G.n190 0.624
R2266 G.n232 G.n230 0.624
R2267 G.n275 G.n273 0.624
R2268 G.n318 G.n316 0.624
R2269 G.n361 G.n359 0.624
R2270 G.n402 G.n400 0.624
R2271 G.n437 G.n435 0.624
R2272 G.n467 G.n465 0.624
R2273 G.n623 G.n622 0.624
R2274 G.n625 G.n621 0.624
R2275 G.n627 G.n620 0.624
R2276 G.n629 G.n619 0.624
R2277 G.n631 G.n618 0.624
R2278 G.n616 G.n605 0.624
R2279 G.n614 G.n606 0.624
R2280 G.n612 G.n607 0.624
R2281 G.n610 G.n608 0.624
R2282 G.n494 G.n493 0.624
R2283 G.n470 G.n468 0.624
R2284 G.n440 G.n438 0.624
R2285 G.n405 G.n403 0.624
R2286 G.n364 G.n362 0.624
R2287 G.n321 G.n319 0.624
R2288 G.n278 G.n276 0.624
R2289 G.n235 G.n233 0.624
R2290 G.n195 G.n193 0.624
R2291 G.n158 G.n156 0.624
R2292 G.n124 G.n122 0.624
R2293 G.n93 G.n91 0.624
R2294 G.n966 G.n964 0.624
R2295 G.n968 G.n963 0.624
R2296 G.n970 G.n962 0.624
R2297 G.n972 G.n961 0.624
R2298 G.n974 G.n960 0.624
R2299 G.n976 G.n959 0.624
R2300 G.n978 G.n958 0.624
R2301 G.n956 G.n939 0.624
R2302 G.n954 G.n940 0.624
R2303 G.n952 G.n941 0.624
R2304 G.n950 G.n942 0.624
R2305 G.n948 G.n943 0.624
R2306 G.n946 G.n944 0.624
R2307 G.n71 G.n69 0.624
R2308 G.n96 G.n94 0.624
R2309 G.n127 G.n125 0.624
R2310 G.n161 G.n159 0.624
R2311 G.n198 G.n196 0.624
R2312 G.n238 G.n236 0.624
R2313 G.n281 G.n279 0.624
R2314 G.n324 G.n322 0.624
R2315 G.n367 G.n365 0.624
R2316 G.n408 G.n406 0.624
R2317 G.n443 G.n441 0.624
R2318 G.n473 G.n471 0.624
R2319 G.n497 G.n495 0.624
R2320 G.n518 G.n517 0.624
R2321 G.n599 G.n597 0.624
R2322 G.n601 G.n596 0.624
R2323 G.n603 G.n595 0.624
R2324 G.n593 G.n585 0.624
R2325 G.n591 G.n586 0.624
R2326 G.n589 G.n587 0.624
R2327 G.n520 G.n519 0.624
R2328 G.n500 G.n498 0.624
R2329 G.n476 G.n474 0.624
R2330 G.n446 G.n444 0.624
R2331 G.n411 G.n409 0.624
R2332 G.n370 G.n368 0.624
R2333 G.n327 G.n325 0.624
R2334 G.n284 G.n282 0.624
R2335 G.n241 G.n239 0.624
R2336 G.n201 G.n199 0.624
R2337 G.n164 G.n162 0.624
R2338 G.n130 G.n128 0.624
R2339 G.n99 G.n97 0.624
R2340 G.n74 G.n72 0.624
R2341 G.n52 G.n50 0.624
R2342 G.n929 G.n927 0.624
R2343 G.n931 G.n926 0.624
R2344 G.n933 G.n925 0.624
R2345 G.n935 G.n924 0.624
R2346 G.n937 G.n923 0.624
R2347 G.n921 G.n910 0.624
R2348 G.n919 G.n911 0.624
R2349 G.n917 G.n912 0.624
R2350 G.n915 G.n913 0.624
R2351 G.n36 G.n34 0.624
R2352 G.n55 G.n53 0.624
R2353 G.n77 G.n75 0.624
R2354 G.n102 G.n100 0.624
R2355 G.n133 G.n131 0.624
R2356 G.n167 G.n165 0.624
R2357 G.n204 G.n202 0.624
R2358 G.n244 G.n242 0.624
R2359 G.n287 G.n285 0.624
R2360 G.n330 G.n328 0.624
R2361 G.n373 G.n371 0.624
R2362 G.n414 G.n412 0.624
R2363 G.n449 G.n447 0.624
R2364 G.n479 G.n477 0.624
R2365 G.n503 G.n501 0.624
R2366 G.n523 G.n521 0.624
R2367 G.n538 G.n537 0.624
R2368 G.n581 G.n579 0.624
R2369 G.n583 G.n578 0.624
R2370 G.n576 G.n571 0.624
R2371 G.n574 G.n572 0.624
R2372 G.n540 G.n539 0.624
R2373 G.n526 G.n524 0.624
R2374 G.n506 G.n504 0.624
R2375 G.n482 G.n480 0.624
R2376 G.n452 G.n450 0.624
R2377 G.n417 G.n415 0.624
R2378 G.n376 G.n374 0.624
R2379 G.n333 G.n331 0.624
R2380 G.n290 G.n288 0.624
R2381 G.n247 G.n245 0.624
R2382 G.n207 G.n205 0.624
R2383 G.n170 G.n168 0.624
R2384 G.n136 G.n134 0.624
R2385 G.n105 G.n103 0.624
R2386 G.n80 G.n78 0.624
R2387 G.n58 G.n56 0.624
R2388 G.n39 G.n37 0.624
R2389 G.n23 G.n21 0.624
R2390 G.n904 G.n902 0.624
R2391 G.n906 G.n901 0.624
R2392 G.n908 G.n900 0.624
R2393 G.n898 G.n893 0.624
R2394 G.n896 G.n894 0.624
R2395 G.n13 G.n11 0.624
R2396 G.n26 G.n24 0.624
R2397 G.n42 G.n40 0.624
R2398 G.n61 G.n59 0.624
R2399 G.n83 G.n81 0.624
R2400 G.n108 G.n106 0.624
R2401 G.n139 G.n137 0.624
R2402 G.n173 G.n171 0.624
R2403 G.n210 G.n208 0.624
R2404 G.n250 G.n248 0.624
R2405 G.n293 G.n291 0.624
R2406 G.n336 G.n334 0.624
R2407 G.n379 G.n377 0.624
R2408 G.n420 G.n418 0.624
R2409 G.n455 G.n453 0.624
R2410 G.n485 G.n483 0.624
R2411 G.n509 G.n507 0.624
R2412 G.n529 G.n527 0.624
R2413 G.n543 G.n541 0.624
R2414 G.n552 G.n551 0.624
R2415 G.n569 G.n567 0.624
R2416 G.n565 G.n564 0.624
R2417 G.n555 G.n553 0.624
R2418 G.n546 G.n544 0.624
R2419 G.n532 G.n530 0.624
R2420 G.n512 G.n510 0.624
R2421 G.n488 G.n486 0.624
R2422 G.n458 G.n456 0.624
R2423 G.n423 G.n421 0.624
R2424 G.n382 G.n380 0.624
R2425 G.n339 G.n337 0.624
R2426 G.n296 G.n294 0.624
R2427 G.n253 G.n251 0.624
R2428 G.n213 G.n211 0.624
R2429 G.n176 G.n174 0.624
R2430 G.n142 G.n140 0.624
R2431 G.n111 G.n109 0.624
R2432 G.n86 G.n84 0.624
R2433 G.n64 G.n62 0.624
R2434 G.n45 G.n43 0.624
R2435 G.n29 G.n27 0.624
R2436 G.n16 G.n14 0.624
R2437 G.n6 G.n4 0.624
R2438 G.n891 G.n889 0.624
R2439 G.n3 G.n2 0.624
R2440 G.n2 G.n0 0.624
R2441 G.n10 G.n9 0.624
R2442 G.n9 G.n7 0.624
R2443 G.n20 G.n19 0.624
R2444 G.n19 G.n17 0.624
R2445 G.n33 G.n32 0.624
R2446 G.n32 G.n30 0.624
R2447 G.n49 G.n48 0.624
R2448 G.n48 G.n46 0.624
R2449 G.n68 G.n67 0.624
R2450 G.n67 G.n65 0.624
R2451 G.n90 G.n89 0.624
R2452 G.n89 G.n87 0.624
R2453 G.n115 G.n114 0.624
R2454 G.n114 G.n112 0.624
R2455 G.n146 G.n145 0.624
R2456 G.n145 G.n143 0.624
R2457 G.n180 G.n179 0.624
R2458 G.n179 G.n177 0.624
R2459 G.n217 G.n216 0.624
R2460 G.n216 G.n214 0.624
R2461 G.n257 G.n256 0.624
R2462 G.n256 G.n254 0.624
R2463 G.n300 G.n299 0.624
R2464 G.n299 G.n297 0.624
R2465 G.n343 G.n342 0.624
R2466 G.n342 G.n340 0.624
R2467 G.n386 G.n385 0.624
R2468 G.n385 G.n383 0.624
R2469 G.n427 G.n426 0.624
R2470 G.n426 G.n424 0.624
R2471 G.n462 G.n461 0.624
R2472 G.n461 G.n459 0.624
R2473 G.n492 G.n491 0.624
R2474 G.n491 G.n489 0.624
R2475 G.n516 G.n515 0.624
R2476 G.n515 G.n513 0.624
R2477 G.n536 G.n535 0.624
R2478 G.n535 G.n533 0.624
R2479 G.n550 G.n549 0.624
R2480 G.n549 G.n547 0.624
R2481 G.n559 G.n558 0.624
R2482 G.n558 G.n556 0.624
R2483 G.n562 G.n561 0.624
R2484 G.n561 G.n560 0.624
R2485 G.n865 G.n562 0.624
R2486 G.n866 G.n559 0.624
R2487 G.n867 G.n550 0.624
R2488 G.n868 G.n536 0.624
R2489 G.n869 G.n516 0.624
R2490 G.n870 G.n492 0.624
R2491 G.n871 G.n462 0.624
R2492 G.n872 G.n427 0.624
R2493 G.n873 G.n386 0.624
R2494 G.n874 G.n343 0.624
R2495 G.n875 G.n300 0.624
R2496 G.n876 G.n257 0.624
R2497 G.n877 G.n217 0.624
R2498 G.n878 G.n180 0.624
R2499 G.n879 G.n146 0.624
R2500 G.n880 G.n115 0.624
R2501 G.n881 G.n90 0.624
R2502 G.n882 G.n68 0.624
R2503 G.n883 G.n49 0.624
R2504 G.n884 G.n33 0.624
R2505 G.n885 G.n20 0.624
R2506 G.n886 G.n10 0.624
R2507 G.n556 G.n555 0.624
R2508 G.n547 G.n546 0.624
R2509 G.n533 G.n532 0.624
R2510 G.n513 G.n512 0.624
R2511 G.n489 G.n488 0.624
R2512 G.n459 G.n458 0.624
R2513 G.n424 G.n423 0.624
R2514 G.n383 G.n382 0.624
R2515 G.n340 G.n339 0.624
R2516 G.n297 G.n296 0.624
R2517 G.n254 G.n253 0.624
R2518 G.n214 G.n213 0.624
R2519 G.n177 G.n176 0.624
R2520 G.n143 G.n142 0.624
R2521 G.n112 G.n111 0.624
R2522 G.n87 G.n86 0.624
R2523 G.n65 G.n64 0.624
R2524 G.n46 G.n45 0.624
R2525 G.n30 G.n29 0.624
R2526 G.n17 G.n16 0.624
R2527 G.n544 G.n543 0.624
R2528 G.n530 G.n529 0.624
R2529 G.n510 G.n509 0.624
R2530 G.n486 G.n485 0.624
R2531 G.n456 G.n455 0.624
R2532 G.n421 G.n420 0.624
R2533 G.n380 G.n379 0.624
R2534 G.n337 G.n336 0.624
R2535 G.n294 G.n293 0.624
R2536 G.n251 G.n250 0.624
R2537 G.n211 G.n210 0.624
R2538 G.n174 G.n173 0.624
R2539 G.n140 G.n139 0.624
R2540 G.n109 G.n108 0.624
R2541 G.n84 G.n83 0.624
R2542 G.n62 G.n61 0.624
R2543 G.n43 G.n42 0.624
R2544 G.n27 G.n26 0.624
R2545 G.n14 G.n13 0.624
R2546 G.n527 G.n526 0.624
R2547 G.n507 G.n506 0.624
R2548 G.n483 G.n482 0.624
R2549 G.n453 G.n452 0.624
R2550 G.n418 G.n417 0.624
R2551 G.n377 G.n376 0.624
R2552 G.n334 G.n333 0.624
R2553 G.n291 G.n290 0.624
R2554 G.n248 G.n247 0.624
R2555 G.n208 G.n207 0.624
R2556 G.n171 G.n170 0.624
R2557 G.n137 G.n136 0.624
R2558 G.n106 G.n105 0.624
R2559 G.n81 G.n80 0.624
R2560 G.n59 G.n58 0.624
R2561 G.n40 G.n39 0.624
R2562 G.n24 G.n23 0.624
R2563 G.n524 G.n523 0.624
R2564 G.n480 G.n479 0.624
R2565 G.n450 G.n449 0.624
R2566 G.n415 G.n414 0.624
R2567 G.n374 G.n373 0.624
R2568 G.n331 G.n330 0.624
R2569 G.n288 G.n287 0.624
R2570 G.n245 G.n244 0.624
R2571 G.n205 G.n204 0.624
R2572 G.n168 G.n167 0.624
R2573 G.n134 G.n133 0.624
R2574 G.n103 G.n102 0.624
R2575 G.n78 G.n77 0.624
R2576 G.n56 G.n55 0.624
R2577 G.n37 G.n36 0.624
R2578 G.n504 G.n503 0.624
R2579 G.n521 G.n520 0.624
R2580 G.n447 G.n446 0.624
R2581 G.n412 G.n411 0.624
R2582 G.n371 G.n370 0.624
R2583 G.n328 G.n327 0.624
R2584 G.n285 G.n284 0.624
R2585 G.n242 G.n241 0.624
R2586 G.n202 G.n201 0.624
R2587 G.n165 G.n164 0.624
R2588 G.n131 G.n130 0.624
R2589 G.n100 G.n99 0.624
R2590 G.n75 G.n74 0.624
R2591 G.n53 G.n52 0.624
R2592 G.n477 G.n476 0.624
R2593 G.n501 G.n500 0.624
R2594 G.n519 G.n518 0.624
R2595 G.n444 G.n443 0.624
R2596 G.n368 G.n367 0.624
R2597 G.n325 G.n324 0.624
R2598 G.n282 G.n281 0.624
R2599 G.n239 G.n238 0.624
R2600 G.n199 G.n198 0.624
R2601 G.n162 G.n161 0.624
R2602 G.n128 G.n127 0.624
R2603 G.n97 G.n96 0.624
R2604 G.n72 G.n71 0.624
R2605 G.n409 G.n408 0.624
R2606 G.n474 G.n473 0.624
R2607 G.n498 G.n497 0.624
R2608 G.n441 G.n440 0.624
R2609 G.n322 G.n321 0.624
R2610 G.n279 G.n278 0.624
R2611 G.n236 G.n235 0.624
R2612 G.n196 G.n195 0.624
R2613 G.n159 G.n158 0.624
R2614 G.n125 G.n124 0.624
R2615 G.n94 G.n93 0.624
R2616 G.n365 G.n364 0.624
R2617 G.n406 G.n405 0.624
R2618 G.n471 G.n470 0.624
R2619 G.n495 G.n494 0.624
R2620 G.n438 G.n437 0.624
R2621 G.n319 G.n318 0.624
R2622 G.n233 G.n232 0.624
R2623 G.n193 G.n192 0.624
R2624 G.n156 G.n155 0.624
R2625 G.n122 G.n121 0.624
R2626 G.n276 G.n275 0.624
R2627 G.n362 G.n361 0.624
R2628 G.n403 G.n402 0.624
R2629 G.n468 G.n467 0.624
R2630 G.n435 G.n434 0.624
R2631 G.n316 G.n315 0.624
R2632 G.n190 G.n189 0.624
R2633 G.n153 G.n152 0.624
R2634 G.n119 G.n118 0.624
R2635 G.n230 G.n229 0.624
R2636 G.n273 G.n272 0.624
R2637 G.n359 G.n358 0.624
R2638 G.n400 G.n399 0.624
R2639 G.n465 G.n464 0.624
R2640 G.n432 G.n431 0.624
R2641 G.n313 G.n312 0.624
R2642 G.n187 G.n186 0.624
R2643 G.n150 G.n149 0.624
R2644 G.n227 G.n226 0.624
R2645 G.n270 G.n269 0.624
R2646 G.n356 G.n355 0.624
R2647 G.n397 G.n396 0.624
R2648 G.n430 G.n429 0.624
R2649 G.n310 G.n309 0.624
R2650 G.n184 G.n183 0.624
R2651 G.n224 G.n223 0.624
R2652 G.n267 G.n266 0.624
R2653 G.n353 G.n352 0.624
R2654 G.n394 G.n393 0.624
R2655 G.n307 G.n306 0.624
R2656 G.n221 G.n220 0.624
R2657 G.n264 G.n263 0.624
R2658 G.n350 G.n349 0.624
R2659 G.n391 G.n390 0.624
R2660 G.n304 G.n303 0.624
R2661 G.n261 G.n260 0.624
R2662 G.n347 G.n346 0.624
R2663 G.n389 G.n388 0.624
R2664 G.n1528 G.n1527 0.624
R2665 G.n1501 G.n1500 0.624
R2666 G.n1476 G.n1475 0.624
R2667 G.n1554 G.n1553 0.624
R2668 G.n1578 G.n1577 0.624
R2669 G.n1602 G.n1601 0.624
R2670 G.n1531 G.n1529 0.624
R2671 G.n1504 G.n1502 0.624
R2672 G.n1479 G.n1477 0.624
R2673 G.n1454 G.n1452 0.624
R2674 G.n1557 G.n1555 0.624
R2675 G.n1581 G.n1579 0.624
R2676 G.n1604 G.n1603 0.624
R2677 G.n1583 G.n1582 0.624
R2678 G.n1559 G.n1558 0.624
R2679 G.n1533 G.n1532 0.624
R2680 G.n1506 G.n1505 0.624
R2681 G.n1481 G.n1480 0.624
R2682 G.n1456 G.n1455 0.624
R2683 G.n1434 G.n1433 0.624
R2684 G.n1622 G.n1621 0.624
R2685 G.n1607 G.n1605 0.624
R2686 G.n1586 G.n1584 0.624
R2687 G.n1562 G.n1560 0.624
R2688 G.n1536 G.n1534 0.624
R2689 G.n1509 G.n1507 0.624
R2690 G.n1484 G.n1482 0.624
R2691 G.n1459 G.n1457 0.624
R2692 G.n1437 G.n1435 0.624
R2693 G.n1418 G.n1416 0.624
R2694 G.n1400 G.n1398 0.624
R2695 G.n1625 G.n1623 0.624
R2696 G.n1640 G.n1639 0.624
R2697 G.n826 G.n822 0.624
R2698 G.n828 G.n821 0.624
R2699 G.n1654 G.n1653 0.624
R2700 G.n1653 G.n1652 0.624
R2701 G.n1643 G.n1642 0.624
R2702 G.n1642 G.n1641 0.624
R2703 G.n1628 G.n1627 0.624
R2704 G.n1627 G.n1626 0.624
R2705 G.n1610 G.n1609 0.624
R2706 G.n1609 G.n1608 0.624
R2707 G.n1589 G.n1588 0.624
R2708 G.n1588 G.n1587 0.624
R2709 G.n1565 G.n1564 0.624
R2710 G.n1564 G.n1563 0.624
R2711 G.n1539 G.n1538 0.624
R2712 G.n1538 G.n1537 0.624
R2713 G.n1512 G.n1511 0.624
R2714 G.n1511 G.n1510 0.624
R2715 G.n1487 G.n1486 0.624
R2716 G.n1486 G.n1485 0.624
R2717 G.n1462 G.n1461 0.624
R2718 G.n1461 G.n1460 0.624
R2719 G.n1440 G.n1439 0.624
R2720 G.n1439 G.n1438 0.624
R2721 G.n1421 G.n1420 0.624
R2722 G.n1420 G.n1419 0.624
R2723 G.n1403 G.n1402 0.624
R2724 G.n1402 G.n1401 0.624
R2725 G.n1387 G.n1386 0.624
R2726 G.n1386 G.n1385 0.624
R2727 G.n1374 G.n1373 0.624
R2728 G.n1310 G.n1309 0.624
R2729 G.n1313 G.n1312 0.624
R2730 G.n1316 G.n1315 0.624
R2731 G.n1319 G.n1318 0.624
R2732 G.n539 G.n538 0.624
R2733 G.n541 G.n540 0.624
R2734 G.n553 G.n552 0.624
R2735 G.n7 G.n6 0.624
R2736 G.n887 G.n3 0.624
R2737 G.n1345 G.n1343 0.624
R2738 G.n1679 G.n1678 0.624
R2739 G G.n887 0.339
R2740 G.n1680 G.n1679 0.305
R2741 G.n1681 G.n1680 0.305
R2742 G.n1682 G.n1681 0.305
R2743 G.n1683 G.n1682 0.305
R2744 G.n1684 G.n1683 0.305
R2745 G.n1685 G.n1684 0.305
R2746 G.n1686 G.n1685 0.305
R2747 G.n1687 G.n1686 0.305
R2748 G.n1688 G.n1687 0.305
R2749 G.n1689 G.n1688 0.305
R2750 G.n1690 G.n1689 0.305
R2751 G.n1691 G.n1690 0.305
R2752 G.n1692 G.n1691 0.305
R2753 G.n1693 G.n1692 0.305
R2754 G.n1694 G.n1693 0.305
R2755 G.n1695 G.n1694 0.305
R2756 G.n1696 G.n1695 0.305
R2757 G.n1697 G.n1696 0.305
R2758 G.n1698 G.n1697 0.305
R2759 G.n1699 G.n1698 0.305
R2760 G.n1700 G.n1699 0.305
R2761 G.n1701 G.n1700 0.305
R2762 G.n866 G.n865 0.305
R2763 G.n867 G.n866 0.305
R2764 G.n868 G.n867 0.305
R2765 G.n869 G.n868 0.305
R2766 G.n870 G.n869 0.305
R2767 G.n871 G.n870 0.305
R2768 G.n872 G.n871 0.305
R2769 G.n873 G.n872 0.305
R2770 G.n874 G.n873 0.305
R2771 G.n875 G.n874 0.305
R2772 G.n876 G.n875 0.305
R2773 G.n877 G.n876 0.305
R2774 G.n878 G.n877 0.305
R2775 G.n879 G.n878 0.305
R2776 G.n880 G.n879 0.305
R2777 G.n881 G.n880 0.305
R2778 G.n882 G.n881 0.305
R2779 G.n883 G.n882 0.305
R2780 G.n884 G.n883 0.305
R2781 G.n885 G.n884 0.305
R2782 G.n886 G.n885 0.305
R2783 G.n887 G.n886 0.305
R2784 G.n843 G.n842 0.305
R2785 G.n844 G.n843 0.305
R2786 G.n845 G.n844 0.305
R2787 G.n846 G.n845 0.305
R2788 G.n847 G.n846 0.305
R2789 G.n848 G.n847 0.305
R2790 G.n849 G.n848 0.305
R2791 G.n850 G.n849 0.305
R2792 G.n851 G.n850 0.305
R2793 G.n852 G.n851 0.305
R2794 G.n853 G.n852 0.305
R2795 G.n854 G.n853 0.305
R2796 G.n855 G.n854 0.305
R2797 G.n856 G.n855 0.305
R2798 G.n857 G.n856 0.305
R2799 G.n858 G.n857 0.305
R2800 G.n859 G.n858 0.305
R2801 G.n860 G.n859 0.305
R2802 G.n861 G.n860 0.305
R2803 G.n862 G.n861 0.305
R2804 G.n863 G.n862 0.305
R2805 G.n864 G.n863 0.305
R2806 G.n1703 G.n1702 0.305
R2807 G.n1704 G.n1703 0.305
R2808 G.n1705 G.n1704 0.305
R2809 G.n1706 G.n1705 0.305
R2810 G.n1707 G.n1706 0.305
R2811 G.n1708 G.n1707 0.305
R2812 G.n1709 G.n1708 0.305
R2813 G.n1710 G.n1709 0.305
R2814 G.n1711 G.n1710 0.305
R2815 G.n1712 G.n1711 0.305
R2816 G.n1713 G.n1712 0.305
R2817 G.n1714 G.n1713 0.305
R2818 G.n1715 G.n1714 0.305
R2819 G.n1716 G.n1715 0.305
R2820 G.n1717 G.n1716 0.305
R2821 G.n1718 G.n1717 0.305
R2822 G.n1719 G.n1718 0.305
R2823 G.n1720 G.n1719 0.305
R2824 G.n1721 G.n1720 0.305
R2825 G.n1722 G.n1721 0.305
R2826 G.n1723 G.n1722 0.305
R2827 G.n1724 G.n1723 0.305
R2828 G G.n1724 0.305
R2829 S.n5401 S.n5400 153.554
R2830 S.n3032 S.n3031 153.554
R2831 S.n3544 S.n3543 153.554
R2832 S.n4043 S.n4042 153.554
R2833 S.n4488 S.n4487 153.554
R2834 S.n4961 S.n4960 153.554
R2835 S.n1952 S.n1951 153.554
R2836 S.n2496 S.n2495 153.554
R2837 S.n779 S.n778 153.554
R2838 S.n1338 S.n1337 153.554
R2839 S.n132 S.n131 153.554
R2840 S.n4372 S.n4371 153.118
R2841 S.n4803 S.n4802 153.118
R2842 S.n3904 S.n3903 153.118
R2843 S.n3419 S.n3418 153.118
R2844 S.n2923 S.n2922 153.118
R2845 S.n2400 S.n2399 153.118
R2846 S.n1872 S.n1871 153.118
R2847 S.n1309 S.n1308 153.118
R2848 S.n5691 S.n5690 153.118
R2849 S.n465 S.n464 153.118
R2850 S.n5260 S.n5259 153.118
R2851 S.n719 S.n718 146.135
R2852 S.n622 S.n621 146.135
R2853 S.n716 S.n715 146.135
R2854 S.n637 S.n636 146.135
R2855 S.n684 S.n683 146.135
R2856 S.n701 S.n700 146.135
R2857 S.n610 S.n609 146.135
R2858 S.n712 S.n711 146.135
R2859 S.n598 S.n597 146.135
R2860 S.n708 S.n707 146.135
R2861 S.n704 S.n703 146.135
R2862 S.n5791 S.n5790 145.699
R2863 S.n5798 S.n5797 145.699
R2864 S.n5784 S.n5783 145.699
R2865 S.n5777 S.n5776 145.699
R2866 S.n5770 S.n5769 145.699
R2867 S.n5763 S.n5762 145.699
R2868 S.n5756 S.n5755 145.699
R2869 S.n5747 S.n5746 145.699
R2870 S.n5733 S.n5732 145.699
R2871 S.n5738 S.n5737 145.699
R2872 S.n5829 S.n5828 145.699
R2873 S.n119 S.n118 101.08
R2874 S.n768 S.n767 101.08
R2875 S.n1328 S.n1327 101.08
R2876 S.n1941 S.n1940 101.08
R2877 S.n2486 S.n2485 101.08
R2878 S.n3021 S.n3020 101.08
R2879 S.n3534 S.n3533 101.08
R2880 S.n4032 S.n4031 101.08
R2881 S.n4478 S.n4477 101.08
R2882 S.n4950 S.n4949 101.08
R2883 S.n5386 S.n5385 101.08
R2884 S.n450 S.n449 98.123
R2885 S.n5711 S.n5710 88.439
R2886 S.n121 S.n120 68.042
R2887 S.n1550 S.n1549 68.042
R2888 S.n1883 S.n1882 68.042
R2889 S.n2411 S.n2410 68.042
R2890 S.n2933 S.n2932 68.042
R2891 S.n3429 S.n3428 68.042
R2892 S.n3914 S.n3913 68.042
R2893 S.n4820 S.n4819 68.042
R2894 S.n4838 S.n4837 68.042
R2895 S.n5704 S.n5703 68.042
R2896 S.n5388 S.n5387 65.312
R2897 S.n5695 S.n5694 62.872
R2898 S.n4841 S.n4840 62.872
R2899 S.n4823 S.n4822 62.872
R2900 S.n3917 S.n3916 62.872
R2901 S.n3432 S.n3431 62.872
R2902 S.n2936 S.n2935 62.872
R2903 S.n2414 S.n2413 62.872
R2904 S.n1886 S.n1885 62.872
R2905 S.n1553 S.n1552 62.872
R2906 S.n744 S.n743 62.872
R2907 S.n453 S.n452 62.872
R2908 S.t191 S.t12 18.142
R2909 S.n458 S.t24 15.833
R2910 S.n122 S.t180 15.833
R2911 S.n749 S.t0 15.833
R2912 S.n769 S.t8 15.833
R2913 S.n1558 S.t95 15.833
R2914 S.n1329 S.t62 15.833
R2915 S.n1891 S.t103 15.833
R2916 S.n1942 S.t2 15.833
R2917 S.n2419 S.t81 15.833
R2918 S.n2487 S.t42 15.833
R2919 S.n2941 S.t10 15.833
R2920 S.n3022 S.t47 15.833
R2921 S.n3437 S.t99 15.833
R2922 S.n3535 S.t22 15.833
R2923 S.n3922 S.t112 15.833
R2924 S.n4033 S.t38 15.833
R2925 S.n4828 S.t85 15.833
R2926 S.n4479 S.t50 15.833
R2927 S.n4846 S.t75 15.833
R2928 S.n4951 S.t16 15.833
R2929 S.n5700 S.t40 15.833
R2930 S.n5390 S.t60 15.833
R2931 S.t151 S.n408 15.305
R2932 S.t213 S.n280 15.305
R2933 S.t58 S.n1032 15.305
R2934 S.t14 S.n961 15.305
R2935 S.t18 S.n1627 15.305
R2936 S.t32 S.n1502 15.305
R2937 S.t290 S.n2191 15.305
R2938 S.t56 S.n2093 15.305
R2939 S.t256 S.n2740 15.305
R2940 S.t68 S.n2620 15.305
R2941 S.t30 S.n3268 15.305
R2942 S.t27 S.n3137 15.305
R2943 S.t200 S.n3783 15.305
R2944 S.t6 S.n3631 15.305
R2945 S.t77 S.n4279 15.305
R2946 S.t65 S.n4113 15.305
R2947 S.t20 S.n4439 15.305
R2948 S.t4 S.n4532 15.305
R2949 S.t36 S.n4886 15.305
R2950 S.t45 S.n4997 15.305
R2951 S.t34 S.n5665 15.305
R2952 S.t52 S.n5449 15.305
R2953 S.t240 S.n5735 15.305
R2954 S.n5712 S.n5711 10.138
R2955 S.n5831 S.t686 6.541
R2956 S.n5723 S.t461 6.541
R2957 S.n4372 S.t78 6.541
R2958 S.n4211 S.n4210 6.541
R2959 S.n4219 S.t971 6.541
R2960 S.n4222 S.t499 6.541
R2961 S.n4214 S.n4213 6.541
R2962 S.n4793 S.n4792 6.541
R2963 S.n4797 S.t668 6.541
R2964 S.n4800 S.t114 6.541
R2965 S.n4790 S.n4789 6.541
R2966 S.n5791 S.t79 6.541
R2967 S.n5789 S.t1003 6.541
R2968 S.n5554 S.n5553 6.541
R2969 S.n5559 S.t1058 6.541
R2970 S.n5562 S.t823 6.541
R2971 S.n5551 S.n5550 6.541
R2972 S.n5298 S.n5297 6.541
R2973 S.n5305 S.t297 6.541
R2974 S.n5302 S.t516 6.541
R2975 S.n5295 S.n5294 6.541
R2976 S.n5084 S.n5083 6.541
R2977 S.n5089 S.t1097 6.541
R2978 S.n5092 S.t94 6.541
R2979 S.n5081 S.n5080 6.541
R2980 S.n5230 S.n5229 6.541
R2981 S.n5234 S.t674 6.541
R2982 S.n5237 S.t462 6.541
R2983 S.n5227 S.n5226 6.541
R2984 S.n4633 S.n4632 6.541
R2985 S.n4638 S.t1073 6.541
R2986 S.n4641 S.t86 6.541
R2987 S.n4630 S.n4629 6.541
R2988 S.n4803 S.t625 6.541
R2989 S.n4805 S.t898 6.541
R2990 S.n5798 S.t820 6.541
R2991 S.n5796 S.t629 6.541
R2992 S.n5567 S.n5566 6.541
R2993 S.n5575 S.t678 6.541
R2994 S.n5578 S.t441 6.541
R2995 S.n5570 S.n5569 6.541
R2996 S.n5279 S.n5278 6.541
R2997 S.n5290 S.t1012 6.541
R2998 S.n5287 S.t122 6.541
R2999 S.n5282 S.n5281 6.541
R3000 S.n5102 S.n5101 6.541
R3001 S.n5110 S.t705 6.541
R3002 S.n5113 S.t833 6.541
R3003 S.n5105 S.n5104 6.541
R3004 S.n5245 S.n5244 6.541
R3005 S.n5254 S.t304 6.541
R3006 S.n5257 S.t633 6.541
R3007 S.n5248 S.n5247 6.541
R3008 S.n4651 S.n4650 6.541
R3009 S.n4662 S.t334 6.541
R3010 S.n4665 S.t986 6.541
R3011 S.n4654 S.n4653 6.541
R3012 S.n4376 S.t165 6.541
R3013 S.n3904 S.t976 6.541
R3014 S.n3713 S.n3712 6.541
R3015 S.n3721 S.t445 6.541
R3016 S.n3724 S.t1083 6.541
R3017 S.n3716 S.n3715 6.541
R3018 S.n3937 S.n3936 6.541
R3019 S.n3944 S.t1049 6.541
R3020 S.n3941 S.t700 6.541
R3021 S.n3934 S.n3933 6.541
R3022 S.n5784 S.t472 6.541
R3023 S.n5782 S.t280 6.541
R3024 S.n5538 S.n5537 6.541
R3025 S.n5543 S.t346 6.541
R3026 S.n5546 S.t84 6.541
R3027 S.n5535 S.n5534 6.541
R3028 S.n5313 S.n5312 6.541
R3029 S.n5320 S.t664 6.541
R3030 S.n5317 S.t902 6.541
R3031 S.n5310 S.n5309 6.541
R3032 S.n5068 S.n5067 6.541
R3033 S.n5073 S.t373 6.541
R3034 S.n5076 S.t492 6.541
R3035 S.n5065 S.n5064 6.541
R3036 S.n5215 S.n5214 6.541
R3037 S.n5219 S.t1072 6.541
R3038 S.n5222 S.t879 6.541
R3039 S.n5212 S.n5211 6.541
R3040 S.n4617 S.n4616 6.541
R3041 S.n4622 S.t351 6.541
R3042 S.n4625 S.t481 6.541
R3043 S.n4614 S.n4613 6.541
R3044 S.n4777 S.n4776 6.541
R3045 S.n4781 S.t1054 6.541
R3046 S.n4784 S.t807 6.541
R3047 S.n4774 S.n4773 6.541
R3048 S.n4198 S.n4197 6.541
R3049 S.n4203 S.t345 6.541
R3050 S.n4206 S.t473 6.541
R3051 S.n4195 S.n4194 6.541
R3052 S.n3908 S.t541 6.541
R3053 S.n3419 S.t459 6.541
R3054 S.n3203 S.n3202 6.541
R3055 S.n3211 S.t1025 6.541
R3056 S.n3214 S.t306 6.541
R3057 S.n3206 S.n3205 6.541
R3058 S.n3452 S.n3451 6.541
R3059 S.n3459 S.t1041 6.541
R3060 S.n3456 S.t230 6.541
R3061 S.n3449 S.n3448 6.541
R3062 S.n5777 S.t751 6.541
R3063 S.n5775 S.t656 6.541
R3064 S.n5522 S.n5521 6.541
R3065 S.n5527 S.t646 6.541
R3066 S.n5530 S.t469 6.541
R3067 S.n5519 S.n5518 6.541
R3068 S.n5328 S.n5327 6.541
R3069 S.n5335 S.t1056 6.541
R3070 S.n5332 S.t150 6.541
R3071 S.n5325 S.n5324 6.541
R3072 S.n5052 S.n5051 6.541
R3073 S.n5057 S.t760 6.541
R3074 S.n5060 S.t862 6.541
R3075 S.n5049 S.n5048 6.541
R3076 S.n5200 S.n5199 6.541
R3077 S.n5204 S.t362 6.541
R3078 S.n5207 S.t159 6.541
R3079 S.n5197 S.n5196 6.541
R3080 S.n4601 S.n4600 6.541
R3081 S.n4606 S.t734 6.541
R3082 S.n4609 S.t811 6.541
R3083 S.n4598 S.n4597 6.541
R3084 S.n4762 S.n4761 6.541
R3085 S.n4766 S.t332 6.541
R3086 S.n4769 S.t139 6.541
R3087 S.n4759 S.n4758 6.541
R3088 S.n4182 S.n4181 6.541
R3089 S.n4187 S.t721 6.541
R3090 S.n4190 S.t812 6.541
R3091 S.n4179 S.n4178 6.541
R3092 S.n3952 S.n3951 6.541
R3093 S.n3959 S.t321 6.541
R3094 S.n3956 S.t125 6.541
R3095 S.n3949 S.n3948 6.541
R3096 S.n3700 S.n3699 6.541
R3097 S.n3705 S.t711 6.541
R3098 S.n3708 S.t837 6.541
R3099 S.n3697 S.n3696 6.541
R3100 S.n3423 S.t907 6.541
R3101 S.n2923 S.t1034 6.541
R3102 S.n2670 S.n2669 6.541
R3103 S.n2678 S.t558 6.541
R3104 S.n2681 S.t958 6.541
R3105 S.n2673 S.n2672 6.541
R3106 S.n2956 S.n2955 6.541
R3107 S.n2963 S.t300 6.541
R3108 S.n2960 S.t815 6.541
R3109 S.n2953 S.n2952 6.541
R3110 S.n5770 S.t61 6.541
R3111 S.n5768 S.t1036 6.541
R3112 S.n5506 S.n5505 6.541
R3113 S.n5511 S.t1039 6.541
R3114 S.n5514 S.t850 6.541
R3115 S.n5503 S.n5502 6.541
R3116 S.n5343 S.n5342 6.541
R3117 S.n5350 S.t333 6.541
R3118 S.n5347 S.t497 6.541
R3119 S.n5340 S.n5339 6.541
R3120 S.n5036 S.n5035 6.541
R3121 S.n5041 S.t1060 6.541
R3122 S.n5044 S.t128 6.541
R3123 S.n5033 S.n5032 6.541
R3124 S.n5185 S.n5184 6.541
R3125 S.n5189 S.t729 6.541
R3126 S.n5192 S.t563 6.541
R3127 S.n5182 S.n5181 6.541
R3128 S.n4585 S.n4584 6.541
R3129 S.n4590 S.t1128 6.541
R3130 S.n4593 S.t126 6.541
R3131 S.n4582 S.n4581 6.541
R3132 S.n4747 S.n4746 6.541
R3133 S.n4751 S.t722 6.541
R3134 S.n4754 S.t544 6.541
R3135 S.n4744 S.n4743 6.541
R3136 S.n4166 S.n4165 6.541
R3137 S.n4171 S.t1113 6.541
R3138 S.n4174 S.t113 6.541
R3139 S.n4163 S.n4162 6.541
R3140 S.n3967 S.n3966 6.541
R3141 S.n3974 S.t712 6.541
R3142 S.n3971 S.t519 6.541
R3143 S.n3964 S.n3963 6.541
R3144 S.n3684 S.n3683 6.541
R3145 S.n3689 S.t1095 6.541
R3146 S.n3692 S.t100 6.541
R3147 S.n3681 S.n3680 6.541
R3148 S.n3467 S.n3466 6.541
R3149 S.n3474 S.t262 6.541
R3150 S.n3471 S.t504 6.541
R3151 S.n3464 S.n3463 6.541
R3152 S.n3190 S.n3189 6.541
R3153 S.n3195 S.t1078 6.541
R3154 S.n3198 S.t809 6.541
R3155 S.n3187 S.n3186 6.541
R3156 S.n2927 S.t155 6.541
R3157 S.n2400 S.t552 6.541
R3158 S.n2127 S.n2126 6.541
R3159 S.n2135 S.t1141 6.541
R3160 S.n2138 S.t450 6.541
R3161 S.n2130 S.n2129 6.541
R3162 S.n2434 S.n2433 6.541
R3163 S.n2441 S.t665 6.541
R3164 S.n2438 S.t281 6.541
R3165 S.n2431 S.n2430 6.541
R3166 S.n5763 S.t451 6.541
R3167 S.n5761 S.t312 6.541
R3168 S.n5490 S.n5489 6.541
R3169 S.n5495 S.t310 6.541
R3170 S.n5498 S.t123 6.541
R3171 S.n5487 S.n5486 6.541
R3172 S.n5358 S.n5357 6.541
R3173 S.n5365 S.t720 6.541
R3174 S.n5362 S.t867 6.541
R3175 S.n5355 S.n5354 6.541
R3176 S.n5020 S.n5019 6.541
R3177 S.n5025 S.t349 6.541
R3178 S.n5028 S.t537 6.541
R3179 S.n5017 S.n5016 6.541
R3180 S.n5170 S.n5169 6.541
R3181 S.n5174 S.t1126 6.541
R3182 S.n5177 S.t857 6.541
R3183 S.n5167 S.n5166 6.541
R3184 S.n4569 S.n4568 6.541
R3185 S.n4574 S.t316 6.541
R3186 S.n4577 S.t465 6.541
R3187 S.n4566 S.n4565 6.541
R3188 S.n4732 S.n4731 6.541
R3189 S.n4736 S.t1114 6.541
R3190 S.n4739 S.t920 6.541
R3191 S.n4729 S.n4728 6.541
R3192 S.n4150 S.n4149 6.541
R3193 S.n4155 S.t392 6.541
R3194 S.n4158 S.t505 6.541
R3195 S.n4147 S.n4146 6.541
R3196 S.n3982 S.n3981 6.541
R3197 S.n3989 S.t1086 6.541
R3198 S.n3986 S.t905 6.541
R3199 S.n3979 S.n3978 6.541
R3200 S.n3668 S.n3667 6.541
R3201 S.n3673 S.t379 6.541
R3202 S.n3676 S.t487 6.541
R3203 S.n3665 S.n3664 6.541
R3204 S.n3482 S.n3481 6.541
R3205 S.n3489 S.t698 6.541
R3206 S.n3486 S.t886 6.541
R3207 S.n3479 S.n3478 6.541
R3208 S.n3174 S.n3173 6.541
R3209 S.n3179 S.t364 6.541
R3210 S.n3182 S.t11 6.541
R3211 S.n3171 S.n3170 6.541
R3212 S.n2971 S.n2970 6.541
R3213 S.n2978 S.t677 6.541
R3214 S.n2975 S.t864 6.541
R3215 S.n2968 S.n2967 6.541
R3216 S.n2657 S.n2656 6.541
R3217 S.n2662 S.t348 6.541
R3218 S.n2665 S.t82 6.541
R3219 S.n2654 S.n2653 6.541
R3220 S.n2404 S.t555 6.541
R3221 S.n1872 S.t19 6.541
R3222 S.n1319 S.n1318 6.541
R3223 S.n1536 S.t636 6.541
R3224 S.n1539 S.t1046 6.541
R3225 S.n1542 S.n1541 6.541
R3226 S.n1906 S.n1905 6.541
R3227 S.n1914 S.t1045 6.541
R3228 S.n1911 S.t919 6.541
R3229 S.n1903 S.n1902 6.541
R3230 S.n5756 S.t835 6.541
R3231 S.n5754 S.t697 6.541
R3232 S.n5587 S.n5586 6.541
R3233 S.n5584 S.t691 6.541
R3234 S.n5581 S.t515 6.541
R3235 S.n5378 S.n5377 6.541
R3236 S.n5373 S.n5372 6.541
R3237 S.n5597 S.t1112 6.541
R3238 S.n5594 S.t143 6.541
R3239 S.n5370 S.n5369 6.541
R3240 S.n5153 S.n5152 6.541
R3241 S.n5150 S.t725 6.541
R3242 S.n5147 S.t876 6.541
R3243 S.n5144 S.n5143 6.541
R3244 S.n5139 S.n5138 6.541
R3245 S.n5159 S.t402 6.541
R3246 S.n5162 S.t131 6.541
R3247 S.n5136 S.n5135 6.541
R3248 S.n4554 S.n4553 6.541
R3249 S.n4558 S.t707 6.541
R3250 S.n4561 S.t903 6.541
R3251 S.n4551 S.n4550 6.541
R3252 S.n4716 S.n4715 6.541
R3253 S.n4721 S.t385 6.541
R3254 S.n4724 S.t120 6.541
R3255 S.n4713 S.n4712 6.541
R3256 S.n4135 S.n4134 6.541
R3257 S.n4139 S.t696 6.541
R3258 S.n4142 S.t883 6.541
R3259 S.n4132 S.n4131 6.541
R3260 S.n3997 S.n3996 6.541
R3261 S.n4005 S.t329 6.541
R3262 S.n4002 S.t173 6.541
R3263 S.n3994 S.n3993 6.541
R3264 S.n3653 S.n3652 6.541
R3265 S.n3657 S.t765 6.541
R3266 S.n3660 S.t865 6.541
R3267 S.n3650 S.n3649 6.541
R3268 S.n3497 S.n3496 6.541
R3269 S.n3505 S.t1081 6.541
R3270 S.n3502 S.t163 6.541
R3271 S.n3494 S.n3493 6.541
R3272 S.n3159 S.n3158 6.541
R3273 S.n3163 S.t737 6.541
R3274 S.n3166 S.t490 6.541
R3275 S.n3156 S.n3155 6.541
R3276 S.n2986 S.n2985 6.541
R3277 S.n2994 S.t1066 6.541
R3278 S.n2991 S.t142 6.541
R3279 S.n2983 S.n2982 6.541
R3280 S.n2642 S.n2641 6.541
R3281 S.n2646 S.t670 6.541
R3282 S.n2649 S.t468 6.541
R3283 S.n2639 S.n2638 6.541
R3284 S.n2449 S.n2448 6.541
R3285 S.n2457 S.t1014 6.541
R3286 S.n2454 S.t129 6.541
R3287 S.n2446 S.n2445 6.541
R3288 S.n2115 S.n2114 6.541
R3289 S.n2119 S.t710 6.541
R3290 S.n2122 S.t453 6.541
R3291 S.n2112 S.n2111 6.541
R3292 S.n1876 S.t911 6.541
R3293 S.n1309 S.t653 6.541
R3294 S.n965 S.n964 6.541
R3295 S.n973 S.t119 6.541
R3296 S.n976 S.t483 6.541
R3297 S.n968 S.n967 6.541
R3298 S.n1573 S.n1572 6.541
R3299 S.n1580 S.t305 6.541
R3300 S.n1577 S.t396 6.541
R3301 S.n1570 S.n1569 6.541
R3302 S.n5747 S.t228 6.541
R3303 S.n5745 S.t449 6.541
R3304 S.n5473 S.n5472 6.541
R3305 S.n5479 S.t1065 6.541
R3306 S.n5482 S.t899 6.541
R3307 S.n5470 S.n5469 6.541
R3308 S.n5605 S.n5604 6.541
R3309 S.n5616 S.t389 6.541
R3310 S.n5613 S.t554 6.541
R3311 S.n5602 S.n5601 6.541
R3312 S.n5122 S.n5121 6.541
R3313 S.n5119 S.t1118 6.541
R3314 S.n5116 S.t179 6.541
R3315 S.n4941 S.n4940 6.541
R3316 S.n4936 S.n4935 6.541
R3317 S.n5128 S.t741 6.541
R3318 S.n5131 S.t526 6.541
R3319 S.n4933 S.n4932 6.541
R3320 S.n4539 S.n4538 6.541
R3321 S.n4543 S.t1101 6.541
R3322 S.n4546 S.t168 6.541
R3323 S.n4536 S.n4535 6.541
R3324 S.n4700 S.n4699 6.541
R3325 S.n4705 S.t778 6.541
R3326 S.n4708 S.t510 6.541
R3327 S.n4697 S.n4696 6.541
R3328 S.n4120 S.n4119 6.541
R3329 S.n4124 S.t1076 6.541
R3330 S.n4127 S.t160 6.541
R3331 S.n4117 S.n4116 6.541
R3332 S.n4013 S.n4012 6.541
R3333 S.n4021 S.t762 6.541
R3334 S.n4018 S.t500 6.541
R3335 S.n4010 S.n4009 6.541
R3336 S.n3638 S.n3637 6.541
R3337 S.n3642 S.t1064 6.541
R3338 S.n3645 S.t140 6.541
R3339 S.n3635 S.n3634 6.541
R3340 S.n3513 S.n3512 6.541
R3341 S.n3521 S.t331 6.541
R3342 S.n3518 S.t566 6.541
R3343 S.n3510 S.n3509 6.541
R3344 S.n3144 S.n3143 6.541
R3345 S.n3148 S.t1131 6.541
R3346 S.n3151 S.t858 6.541
R3347 S.n3141 S.n3140 6.541
R3348 S.n3002 S.n3001 6.541
R3349 S.n3010 S.t359 6.541
R3350 S.n3007 S.t534 6.541
R3351 S.n2999 S.n2998 6.541
R3352 S.n2627 S.n2626 6.541
R3353 S.n2631 S.t1116 6.541
R3354 S.n2634 S.t847 6.541
R3355 S.n2624 S.n2623 6.541
R3356 S.n2465 S.n2464 6.541
R3357 S.n2473 S.t337 6.541
R3358 S.n2470 S.t525 6.541
R3359 S.n2462 S.n2461 6.541
R3360 S.n2100 S.n2099 6.541
R3361 S.n2104 S.t1100 6.541
R3362 S.n2107 S.t844 6.541
R3363 S.n2097 S.n2096 6.541
R3364 S.n1922 S.n1921 6.541
R3365 S.n1930 S.t313 6.541
R3366 S.n1927 S.t507 6.541
R3367 S.n1919 S.n1918 6.541
R3368 S.n1525 S.n1524 6.541
R3369 S.n1530 S.t1075 6.541
R3370 S.n1533 S.t832 6.541
R3371 S.n1522 S.n1521 6.541
R3372 S.n1313 S.t1099 6.541
R3373 S.n5734 S.t988 6.541
R3374 S.n5733 S.t208 6.541
R3375 S.n5691 S.t870 6.541
R3376 S.n5637 S.t162 6.541
R3377 S.n382 S.n381 6.541
R3378 S.n406 S.t172 6.541
R3379 S.n403 S.t796 6.541
R3380 S.n385 S.n384 6.541
R3381 S.n1048 S.n1047 6.541
R3382 S.n1058 S.t189 6.541
R3383 S.n1061 S.t1055 6.541
R3384 S.n1045 S.n1044 6.541
R3385 S.n5402 S.t540 6.541
R3386 S.n5645 S.n5644 6.541
R3387 S.n5663 S.t35 6.541
R3388 S.n5660 S.t836 6.541
R3389 S.n5642 S.n5641 6.541
R3390 S.n4970 S.n4969 6.541
R3391 S.n4981 S.t983 6.541
R3392 S.n4978 S.t325 6.541
R3393 S.n4967 S.n4966 6.541
R3394 S.n4869 S.n4868 6.541
R3395 S.n4884 S.t1023 6.541
R3396 S.n4881 S.t592 6.541
R3397 S.n4866 S.n4865 6.541
R3398 S.n4519 S.n4518 6.541
R3399 S.n4530 S.t704 6.541
R3400 S.n4527 S.t941 6.541
R3401 S.n4516 S.n4515 6.541
R3402 S.n4422 S.n4421 6.541
R3403 S.n4437 S.t413 6.541
R3404 S.n4434 S.t157 6.541
R3405 S.n4419 S.n4418 6.541
R3406 S.n4100 S.n4099 6.541
R3407 S.n4111 S.t753 6.541
R3408 S.n4108 S.t931 6.541
R3409 S.n4097 S.n4096 6.541
R3410 S.n4295 S.n4294 6.541
R3411 S.n4307 S.t419 6.541
R3412 S.n4310 S.t108 6.541
R3413 S.n4292 S.n4291 6.541
R3414 S.n3618 S.n3617 6.541
R3415 S.n3629 S.t727 6.541
R3416 S.n3626 S.t921 6.541
R3417 S.n3615 S.n3614 6.541
R3418 S.n3799 S.n3798 6.541
R3419 S.n3811 S.t1088 6.541
R3420 S.n3814 S.t136 6.541
R3421 S.n3796 S.n3795 6.541
R3422 S.n3124 S.n3123 6.541
R3423 S.n3135 S.t713 6.541
R3424 S.n3132 S.t524 6.541
R3425 S.n3121 S.n3120 6.541
R3426 S.n3284 S.n3283 6.541
R3427 S.n3296 S.t1094 6.541
R3428 S.n3299 S.t121 6.541
R3429 S.n3281 S.n3280 6.541
R3430 S.n2607 S.n2606 6.541
R3431 S.n2618 S.t692 6.541
R3432 S.n2615 S.t511 6.541
R3433 S.n2604 S.n2603 6.541
R3434 S.n2756 S.n2755 6.541
R3435 S.n2768 S.t1105 6.541
R3436 S.n2771 S.t176 6.541
R3437 S.n2753 S.n2752 6.541
R3438 S.n2080 S.n2079 6.541
R3439 S.n2091 S.t767 6.541
R3440 S.n2088 S.t501 6.541
R3441 S.n2077 S.n2076 6.541
R3442 S.n2207 S.n2206 6.541
R3443 S.n2218 S.t1084 6.541
R3444 S.n2221 S.t164 6.541
R3445 S.n2204 S.n2203 6.541
R3446 S.n1488 S.n1487 6.541
R3447 S.n1500 S.t748 6.541
R3448 S.n1497 S.t488 6.541
R3449 S.n1485 S.n1484 6.541
R3450 S.n1643 S.n1642 6.541
R3451 S.n1655 S.t1068 6.541
R3452 S.n1658 S.t145 6.541
R3453 S.n1640 S.n1639 6.541
R3454 S.n948 S.n947 6.541
R3455 S.n959 S.t708 6.541
R3456 S.n956 S.t614 6.541
R3457 S.n945 S.n944 6.541
R3458 S.n360 S.n359 6.541
R3459 S.n363 S.t583 6.541
R3460 S.n366 S.t649 6.541
R3461 S.n369 S.n368 6.541
R3462 S.n284 S.n283 6.541
R3463 S.n295 S.t1008 6.541
R3464 S.n298 S.t1077 6.541
R3465 S.n287 S.n286 6.541
R3466 S.n465 S.t170 6.541
R3467 S.n440 S.t365 6.541
R3468 S.n5738 S.t622 6.541
R3469 S.n5736 S.t780 6.541
R3470 S.n5454 S.n5453 6.541
R3471 S.n5462 S.t358 6.541
R3472 S.n5465 S.t183 6.541
R3473 S.n5457 S.n5456 6.541
R3474 S.n5624 S.n5623 6.541
R3475 S.n5635 S.t831 6.541
R3476 S.n5632 S.t452 6.541
R3477 S.n5627 S.n5626 6.541
R3478 S.n5001 S.n5000 6.541
R3479 S.n5009 S.t612 6.541
R3480 S.n5012 S.t580 6.541
R3481 S.n5004 S.n5003 6.541
R3482 S.n4917 S.n4916 6.541
R3483 S.n4925 S.t37 6.541
R3484 S.n4928 S.t897 6.541
R3485 S.n4920 S.n4919 6.541
R3486 S.n4467 S.n4466 6.541
R3487 S.n4668 S.t327 6.541
R3488 S.n4671 S.t571 6.541
R3489 S.n4674 S.n4673 6.541
R3490 S.n4681 S.n4680 6.541
R3491 S.n4689 S.t21 6.541
R3492 S.n4692 S.t889 6.541
R3493 S.n4684 S.n4683 6.541
R3494 S.n4025 S.n4024 6.541
R3495 S.n4225 S.t368 6.541
R3496 S.n4228 S.t564 6.541
R3497 S.n4231 S.n4230 6.541
R3498 S.n4238 S.n4237 6.541
R3499 S.n4249 S.t1142 6.541
R3500 S.n4246 S.t872 6.541
R3501 S.n4241 S.n4240 6.541
R3502 S.n3525 S.n3524 6.541
R3503 S.n3727 S.t356 6.541
R3504 S.n3730 S.t545 6.541
R3505 S.n3733 S.n3732 6.541
R3506 S.n3740 S.n3739 6.541
R3507 S.n3751 S.t738 6.541
R3508 S.n3748 S.t808 6.541
R3509 S.n3743 S.n3742 6.541
R3510 S.n3014 S.n3013 6.541
R3511 S.n3217 S.t335 6.541
R3512 S.n3220 S.t132 6.541
R3513 S.n3223 S.n3222 6.541
R3514 S.n3230 S.n3229 6.541
R3515 S.n3241 S.t726 6.541
R3516 S.n3238 S.t923 6.541
R3517 S.n3233 S.n3232 6.541
R3518 S.n2477 S.n2476 6.541
R3519 S.n2684 S.t403 6.541
R3520 S.n2687 S.t115 6.541
R3521 S.n2690 S.n2689 6.541
R3522 S.n2697 S.n2696 6.541
R3523 S.n2708 S.t715 6.541
R3524 S.n2705 S.t906 6.541
R3525 S.n2700 S.n2699 6.541
R3526 S.n1934 S.n1933 6.541
R3527 S.n2141 S.t328 6.541
R3528 S.n2144 S.t104 6.541
R3529 S.n2147 S.n2146 6.541
R3530 S.n2154 S.n2153 6.541
R3531 S.n2165 S.t689 6.541
R3532 S.n2162 S.t891 6.541
R3533 S.n2157 S.n2156 6.541
R3534 S.n1506 S.n1505 6.541
R3535 S.n1514 S.t341 6.541
R3536 S.n1517 S.t96 6.541
R3537 S.n1509 S.n1508 6.541
R3538 S.n1584 S.n1583 6.541
R3539 S.n1595 S.t684 6.541
R3540 S.n1592 S.t869 6.541
R3541 S.n1587 S.n1586 6.541
R3542 S.n761 S.n760 6.541
R3543 S.n979 S.t354 6.541
R3544 S.n982 S.t283 6.541
R3545 S.n985 S.n984 6.541
R3546 S.n992 S.n991 6.541
R3547 S.n1007 S.t877 6.541
R3548 S.n1004 S.t181 6.541
R3549 S.n995 S.n994 6.541
R3550 S.n616 S.t192 6.541
R3551 S.n97 S.n96 6.541
R3552 S.n108 S.t977 6.541
R3553 S.n105 S.t679 6.541
R3554 S.n100 S.n99 6.541
R3555 S.n1201 S.n1200 6.541
R3556 S.n1211 S.t984 6.541
R3557 S.n1214 S.t688 6.541
R3558 S.n1198 S.n1197 6.541
R3559 S.n3033 S.t277 6.541
R3560 S.n3249 S.n3248 6.541
R3561 S.n3266 S.t901 6.541
R3562 S.n3263 S.t330 6.541
R3563 S.n3246 S.n3245 6.541
R3564 S.n2505 S.n2504 6.541
R3565 S.n2516 S.t498 6.541
R3566 S.n2513 S.t1137 6.541
R3567 S.n2502 S.n2501 6.541
R3568 S.n2905 S.n2904 6.541
R3569 S.n2917 S.t660 6.541
R3570 S.n2920 S.t90 6.541
R3571 S.n2902 S.n2901 6.541
R3572 S.n1980 S.n1979 6.541
R3573 S.n1991 S.t248 6.541
R3574 S.n1988 S.t202 6.541
R3575 S.n1977 S.n1976 6.541
R3576 S.n2350 S.n2349 6.541
R3577 S.n2361 S.t743 6.541
R3578 S.n2364 S.t881 6.541
R3579 S.n2347 S.n2346 6.541
R3580 S.n1386 S.n1385 6.541
R3581 S.n1398 S.t388 6.541
R3582 S.n1395 S.t188 6.541
R3583 S.n1383 S.n1382 6.541
R3584 S.n1789 S.n1788 6.541
R3585 S.n1801 S.t782 6.541
R3586 S.n1804 S.t896 6.541
R3587 S.n1786 S.n1785 6.541
R3588 S.n843 S.n842 6.541
R3589 S.n854 S.t378 6.541
R3590 S.n851 S.t371 6.541
R3591 S.n840 S.n839 6.541
R3592 S.n714 S.t978 6.541
R3593 S.n12 S.n11 6.541
R3594 S.n468 S.t620 6.541
R3595 S.n471 S.t377 6.541
R3596 S.n474 S.n473 6.541
R3597 S.n3545 S.t1144 6.541
R3598 S.n3763 S.n3762 6.541
R3599 S.n3781 S.t773 6.541
R3600 S.n3778 S.t221 6.541
R3601 S.n3766 S.n3765 6.541
R3602 S.n3041 S.n3040 6.541
R3603 S.n3052 S.t367 6.541
R3604 S.n3049 S.t998 6.541
R3605 S.n3044 S.n3043 6.541
R3606 S.n3396 S.n3395 6.541
R3607 S.n3413 S.t586 6.541
R3608 S.n3416 S.t1057 6.541
R3609 S.n3399 S.n3398 6.541
R3610 S.n2524 S.n2523 6.541
R3611 S.n2535 S.t105 6.541
R3612 S.n2532 S.t939 6.541
R3613 S.n2527 S.n2526 6.541
R3614 S.n2868 S.n2867 6.541
R3615 S.n2885 S.t434 6.541
R3616 S.n2888 S.t560 6.541
R3617 S.n2871 S.n2870 6.541
R3618 S.n1997 S.n1996 6.541
R3619 S.n2008 S.t1122 6.541
R3620 S.n2005 S.t915 6.541
R3621 S.n2000 S.n1999 6.541
R3622 S.n2313 S.n2312 6.541
R3623 S.n2330 S.t424 6.541
R3624 S.n2333 S.t530 6.541
R3625 S.n2316 S.n2315 6.541
R3626 S.n1404 S.n1403 6.541
R3627 S.n1415 S.t1110 6.541
R3628 S.n1412 S.t918 6.541
R3629 S.n1407 S.n1406 6.541
R3630 S.n1752 S.n1751 6.541
R3631 S.n1769 S.t411 6.541
R3632 S.n1772 S.t514 6.541
R3633 S.n1755 S.n1754 6.541
R3634 S.n860 S.n859 6.541
R3635 S.n873 S.t1092 6.541
R3636 S.n870 S.t1085 6.541
R3637 S.n863 S.n862 6.541
R3638 S.n881 S.n880 6.541
R3639 S.n895 S.t702 6.541
R3640 S.n892 S.t701 6.541
R3641 S.n884 S.n883 6.541
R3642 S.n1132 S.n1131 6.541
R3643 S.n1153 S.t232 6.541
R3644 S.n1156 S.t1109 6.541
R3645 S.n1135 S.n1134 6.541
R3646 S.n112 S.n111 6.541
R3647 S.n301 S.t610 6.541
R3648 S.n304 S.t676 6.541
R3649 S.n307 S.n306 6.541
R3650 S.n315 S.n314 6.541
R3651 S.n330 S.t220 6.541
R3652 S.n327 S.t1096 6.541
R3653 S.n318 S.n317 6.541
R3654 S.n630 S.t621 6.541
R3655 S.n1728 S.n1727 6.541
R3656 S.n1740 S.t1125 6.541
R3657 S.n1743 S.t110 6.541
R3658 S.n1725 S.n1724 6.541
R3659 S.n2290 S.n2289 6.541
R3660 S.n2301 S.t1138 6.541
R3661 S.n2304 S.t138 6.541
R3662 S.n2287 S.n2286 6.541
R3663 S.n2840 S.n2839 6.541
R3664 S.n2852 S.t1150 6.541
R3665 S.n2855 S.t149 6.541
R3666 S.n2837 S.n2836 6.541
R3667 S.n3368 S.n3367 6.541
R3668 S.n3380 S.t31 6.541
R3669 S.n3383 S.t167 6.541
R3670 S.n3365 S.n3364 6.541
R3671 S.n3886 S.n3885 6.541
R3672 S.n3898 S.t442 6.541
R3673 S.n3901 S.t973 6.541
R3674 S.n3883 S.n3882 6.541
R3675 S.n4260 S.n4259 6.541
R3676 S.n4277 S.t521 6.541
R3677 S.n4274 S.t91 6.541
R3678 S.n4257 S.n4256 6.541
R3679 S.n4044 S.t1000 6.541
R3680 S.n3553 S.n3552 6.541
R3681 S.n3564 S.t246 6.541
R3682 S.n3561 S.t763 6.541
R3683 S.n3550 S.n3549 6.541
R3684 S.n3060 S.n3059 6.541
R3685 S.n3071 S.t1074 6.541
R3686 S.n3068 S.t576 6.541
R3687 S.n3057 S.n3056 6.541
R3688 S.n2543 S.n2542 6.541
R3689 S.n2554 S.t755 6.541
R3690 S.n2551 S.t569 6.541
R3691 S.n2540 S.n2539 6.541
R3692 S.n2016 S.n2015 6.541
R3693 S.n2027 S.t732 6.541
R3694 S.n2024 S.t561 6.541
R3695 S.n2013 S.n2012 6.541
R3696 S.n1423 S.n1422 6.541
R3697 S.n1435 S.t716 6.541
R3698 S.n1432 S.t529 6.541
R3699 S.n1420 S.n1419 6.541
R3700 S.n1104 S.n1103 6.541
R3701 S.n1119 S.t959 6.541
R3702 S.n1122 S.t719 6.541
R3703 S.n1107 S.n1106 6.541
R3704 S.n240 S.n239 6.541
R3705 S.n259 S.t236 6.541
R3706 S.n256 S.t303 6.541
R3707 S.n243 S.n242 6.541
R3708 S.n646 S.n645 6.541
R3709 S.n649 S.t938 6.541
R3710 S.n652 S.t671 6.541
R3711 S.n655 S.n654 6.541
R3712 S.n641 S.t218 6.541
R3713 S.n4489 S.t895 6.541
R3714 S.n4452 S.n4451 6.541
R3715 S.n4460 S.t384 6.541
R3716 S.n4463 S.t1062 6.541
R3717 S.n4449 S.n4448 6.541
R3718 S.n4061 S.n4060 6.541
R3719 S.n4070 S.t117 6.541
R3720 S.n4067 S.t630 6.541
R3721 S.n4058 S.n4057 6.541
R3722 S.n4348 S.n4347 6.541
R3723 S.n4366 S.t203 6.541
R3724 S.n4369 S.t829 6.541
R3725 S.n4345 S.n4344 6.541
R3726 S.n3581 S.n3580 6.541
R3727 S.n3590 S.t979 6.541
R3728 S.n3587 S.t584 6.541
R3729 S.n3578 S.n3577 6.541
R3730 S.n3848 S.n3847 6.541
R3731 S.n3866 S.t791 6.541
R3732 S.n3869 S.t908 6.541
R3733 S.n3845 S.n3844 6.541
R3734 S.n3088 S.n3087 6.541
R3735 S.n3096 S.t382 6.541
R3736 S.n3093 S.t186 6.541
R3737 S.n3085 S.n3084 6.541
R3738 S.n3333 S.n3332 6.541
R3739 S.n3348 S.t746 6.541
R3740 S.n3351 S.t894 6.541
R3741 S.n3330 S.n3329 6.541
R3742 S.n2571 S.n2570 6.541
R3743 S.n2579 S.t372 6.541
R3744 S.n2576 S.t154 6.541
R3745 S.n2568 S.n2567 6.541
R3746 S.n2805 S.n2804 6.541
R3747 S.n2820 S.t774 6.541
R3748 S.n2823 S.t874 6.541
R3749 S.n2802 S.n2801 6.541
R3750 S.n2044 S.n2043 6.541
R3751 S.n2052 S.t360 6.541
R3752 S.n2049 S.t146 6.541
R3753 S.n2041 S.n2040 6.541
R3754 S.n2255 S.n2254 6.541
R3755 S.n2270 S.t757 6.541
R3756 S.n2273 S.t860 6.541
R3757 S.n2252 S.n2251 6.541
R3758 S.n1452 S.n1451 6.541
R3759 S.n1460 S.t343 6.541
R3760 S.n1457 S.t137 6.541
R3761 S.n1449 S.n1448 6.541
R3762 S.n1692 S.n1691 6.541
R3763 S.n1707 S.t730 6.541
R3764 S.n1710 S.t925 6.541
R3765 S.n1689 S.n1688 6.541
R3766 S.n911 S.n910 6.541
R3767 S.n919 S.t407 6.541
R3768 S.n916 S.t314 6.541
R3769 S.n908 S.n907 6.541
R3770 S.n1070 S.n1069 6.541
R3771 S.n1086 S.t581 6.541
R3772 S.n1089 S.t344 6.541
R3773 S.n1073 S.n1072 6.541
R3774 S.n264 S.n263 6.541
R3775 S.n278 S.t957 6.541
R3776 S.n275 S.t1028 6.541
R3777 S.n267 S.n266 6.541
R3778 S.n931 S.n930 6.541
R3779 S.n940 S.t1115 6.541
R3780 S.n937 S.t1044 6.541
R3781 S.n928 S.n927 6.541
R3782 S.n1667 S.n1666 6.541
R3783 S.n1675 S.t361 6.541
R3784 S.n1678 S.t550 6.541
R3785 S.n1670 S.n1669 6.541
R3786 S.n1466 S.n1465 6.541
R3787 S.n1480 S.t1091 6.541
R3788 S.n1477 S.t859 6.541
R3789 S.n1469 S.n1468 6.541
R3790 S.n2230 S.n2229 6.541
R3791 S.n2238 S.t370 6.541
R3792 S.n2241 S.t567 6.541
R3793 S.n2233 S.n2232 6.541
R3794 S.n2058 S.n2057 6.541
R3795 S.n2072 S.t1067 6.541
R3796 S.n2069 S.t873 6.541
R3797 S.n2061 S.n2060 6.541
R3798 S.n2780 S.n2779 6.541
R3799 S.n2788 S.t386 6.541
R3800 S.n2791 S.t470 6.541
R3801 S.n2783 S.n2782 6.541
R3802 S.n2585 S.n2584 6.541
R3803 S.n2599 S.t1082 6.541
R3804 S.n2596 S.t892 6.541
R3805 S.n2588 S.n2587 6.541
R3806 S.n3308 S.n3307 6.541
R3807 S.n3316 S.t409 6.541
R3808 S.n3319 S.t512 6.541
R3809 S.n3311 S.n3310 6.541
R3810 S.n3102 S.n3101 6.541
R3811 S.n3116 S.t1106 6.541
R3812 S.n3113 S.t912 6.541
R3813 S.n3105 S.n3104 6.541
R3814 S.n3823 S.n3822 6.541
R3815 S.n3831 S.t421 6.541
R3816 S.n3834 S.t522 6.541
R3817 S.n3826 S.n3825 6.541
R3818 S.n3596 S.n3595 6.541
R3819 S.n3610 S.t1120 6.541
R3820 S.n3607 S.t195 6.541
R3821 S.n3599 S.n3598 6.541
R3822 S.n4323 S.n4322 6.541
R3823 S.n4331 S.t740 6.541
R3824 S.n4334 S.t543 6.541
R3825 S.n4326 S.n4325 6.541
R3826 S.n4078 S.n4077 6.541
R3827 S.n4092 S.t818 6.541
R3828 S.n4089 S.t207 6.541
R3829 S.n4081 S.n4080 6.541
R3830 S.n4394 S.n4393 6.541
R3831 S.n4405 S.t49 6.541
R3832 S.n4402 S.t680 6.541
R3833 S.n4397 S.n4396 6.541
R3834 S.n4497 S.n4496 6.541
R3835 S.n4511 S.t1093 6.541
R3836 S.n4508 S.t466 6.541
R3837 S.n4500 S.n4499 6.541
R3838 S.n4898 S.n4897 6.541
R3839 S.n4906 S.t254 6.541
R3840 S.n4909 S.t967 6.541
R3841 S.n4901 S.n4900 6.541
R3842 S.n4962 S.t769 6.541
R3843 S.n689 S.t943 6.541
R3844 S.n339 S.n338 6.541
R3845 S.n356 S.t553 6.541
R3846 S.n353 S.t318 6.541
R3847 S.n342 S.n341 6.541
R3848 S.n1165 S.n1164 6.541
R3849 S.n1181 S.t611 6.541
R3850 S.n1184 S.t268 6.541
R3851 S.n1168 S.n1167 6.541
R3852 S.n224 S.n223 6.541
R3853 S.n235 S.t935 6.541
R3854 S.n232 S.t1069 6.541
R3855 S.n227 S.n226 6.541
R3856 S.n207 S.n206 6.541
R3857 S.n218 S.t214 6.541
R3858 S.n215 S.t355 6.541
R3859 S.n210 S.n209 6.541
R3860 S.n604 S.t969 6.541
R3861 S.n65 S.n64 6.541
R3862 S.n76 S.t631 6.541
R3863 S.n73 S.t350 6.541
R3864 S.n68 S.n67 6.541
R3865 S.n1260 S.n1259 6.541
R3866 S.n1270 S.t637 6.541
R3867 S.n1273 S.t366 6.541
R3868 S.n1257 S.n1256 6.541
R3869 S.n1953 S.t562 6.541
R3870 S.n2173 S.n2172 6.541
R3871 S.n2189 S.t1145 6.541
R3872 S.n2186 S.t607 6.541
R3873 S.n2170 S.n2169 6.541
R3874 S.n1347 S.n1346 6.541
R3875 S.n1359 S.t736 6.541
R3876 S.n1356 S.t255 6.541
R3877 S.n1344 S.n1343 6.541
R3878 S.n1854 S.n1853 6.541
R3879 S.n1866 S.t955 6.541
R3880 S.n1869 S.t336 6.541
R3881 S.n1851 S.n1850 6.541
R3882 S.n807 S.n806 6.541
R3883 S.n818 S.t496 6.541
R3884 S.n815 S.t1139 6.541
R3885 S.n804 S.n803 6.541
R3886 S.n710 S.t587 6.541
R3887 S.n506 S.n505 6.541
R3888 S.n509 S.t247 6.541
R3889 S.n512 S.t1061 6.541
R3890 S.n515 S.n514 6.541
R3891 S.n2497 S.t422 6.541
R3892 S.n2720 S.n2719 6.541
R3893 S.n2738 S.t1001 6.541
R3894 S.n2735 S.t489 6.541
R3895 S.n2723 S.n2722 6.541
R3896 S.n1961 S.n1960 6.541
R3897 S.n1972 S.t627 6.541
R3898 S.n1969 S.t158 6.541
R3899 S.n1964 S.n1963 6.541
R3900 S.n2377 S.n2376 6.541
R3901 S.n2394 S.t822 6.541
R3902 S.n2397 S.t237 6.541
R3903 S.n2380 S.n2379 6.541
R3904 S.n1367 S.n1366 6.541
R3905 S.n1378 S.t363 6.541
R3906 S.n1375 S.t579 6.541
R3907 S.n1370 S.n1369 6.541
R3908 S.n1817 S.n1816 6.541
R3909 S.n1834 S.t29 6.541
R3910 S.n1837 S.t153 6.541
R3911 S.n1820 S.n1819 6.541
R3912 S.n824 S.n823 6.541
R3913 S.n835 S.t759 6.541
R3914 S.n832 S.t758 6.541
R3915 S.n827 S.n826 6.541
R3916 S.n1223 S.n1222 6.541
R3917 S.n1240 S.t250 6.541
R3918 S.n1243 S.t1079 6.541
R3919 S.n1226 S.n1225 6.541
R3920 S.n189 S.n188 6.541
R3921 S.n200 S.t597 6.541
R3922 S.n197 S.t731 6.541
R3923 S.n192 S.n191 6.541
R3924 S.n172 S.n171 6.541
R3925 S.n183 S.t965 6.541
R3926 S.n180 S.t1127 6.541
R3927 S.n175 S.n174 6.541
R3928 S.n591 S.t642 6.541
R3929 S.n33 S.n32 6.541
R3930 S.n44 S.t981 6.541
R3931 S.n41 S.t513 6.541
R3932 S.n36 S.n35 6.541
R3933 S.n1015 S.n1014 6.541
R3934 S.n1030 S.t59 6.541
R3935 S.n1027 S.t768 6.541
R3936 S.n1012 S.n1011 6.541
R3937 S.n780 S.t532 6.541
R3938 S.n706 S.t222 6.541
R3939 S.n544 S.n543 6.541
R3940 S.n547 S.t994 6.541
R3941 S.n550 S.t724 6.541
R3942 S.n553 S.n552 6.541
R3943 S.n1339 S.t601 6.541
R3944 S.n1607 S.n1606 6.541
R3945 S.n1625 S.t156 6.541
R3946 S.n1622 S.t718 6.541
R3947 S.n1610 S.n1609 6.541
R3948 S.n788 S.n787 6.541
R3949 S.n799 S.t868 6.541
R3950 S.n796 S.t204 6.541
R3951 S.n791 S.n790 6.541
R3952 S.n1286 S.n1285 6.541
R3953 S.n1303 S.t848 6.541
R3954 S.n1306 S.t326 6.541
R3955 S.n1289 S.n1288 6.541
R3956 S.n154 S.n153 6.541
R3957 S.n165 S.t546 6.541
R3958 S.n162 S.t401 6.541
R3959 S.n157 S.n156 6.541
R3960 S.n138 S.n137 6.541
R3961 S.n149 S.t922 6.541
R3962 S.n146 S.t296 6.541
R3963 S.n141 S.n140 6.541
R3964 S.n702 S.t1009 6.541
R3965 S.n421 S.n420 6.541
R3966 S.n410 S.t210 6.541
R3967 S.n434 S.t893 6.541
R3968 S.n424 S.n423 6.541
R3969 S.n133 S.t663 6.541
R3970 S.n728 S.t535 6.541
R3971 S.n5418 S.n5417 6.541
R3972 S.n5421 S.t270 6.541
R3973 S.n5260 S.t1098 6.541
R3974 S.n5262 S.t551 6.541
R3975 S.n5829 S.t437 6.541
R3976 S.n5827 S.t253 6.541
R3977 S.n5677 S.n5676 6.541
R3978 S.n5685 S.t644 6.541
R3979 S.n5688 S.t1136 6.541
R3980 S.n5680 S.n5679 6.541
R3981 S.n4984 S.n4983 6.541
R3982 S.n4995 S.t854 6.541
R3983 S.n4992 S.t339 6.541
R3984 S.n4987 S.n4986 6.541
R3985 S.n5411 S.n5410 6.541
R3986 S.n5414 S.t41 6.541
R3987 S.n5444 S.n5443 6.541
R3988 S.n5447 S.t238 6.541
R3989 S.n5439 S.n5438 6.541
R3990 S.n5424 S.t474 6.541
R3991 S.n4211 S.t632 6.105
R3992 S.n4219 S.n4218 6.105
R3993 S.n4222 S.n4221 6.105
R3994 S.n4214 S.t54 6.105
R3995 S.n4793 S.t934 6.105
R3996 S.n4797 S.n4796 6.105
R3997 S.n4800 S.n4799 6.105
R3998 S.n4790 S.t375 6.105
R3999 S.n5792 S.t990 6.105
R4000 S.n5554 S.t669 6.105
R4001 S.n5559 S.n5558 6.105
R4002 S.n5562 S.n5561 6.105
R4003 S.n5551 S.t1102 6.105
R4004 S.n5298 S.t278 6.105
R4005 S.n5305 S.n5304 6.105
R4006 S.n5302 S.n5301 6.105
R4007 S.n5295 S.t536 6.105
R4008 S.n5084 S.t752 6.105
R4009 S.n5089 S.n5088 6.105
R4010 S.n5092 S.n5091 6.105
R4011 S.n5081 S.t412 6.105
R4012 S.n5230 S.t647 6.105
R4013 S.n5234 S.n5233 6.105
R4014 S.n5237 S.n5236 6.105
R4015 S.n5227 S.t929 6.105
R4016 S.n4633 S.t706 6.105
R4017 S.n4638 S.n4637 6.105
R4018 S.n4641 S.n4640 6.105
R4019 S.n4630 S.t426 6.105
R4020 S.n4807 S.t225 6.105
R4021 S.n5799 S.t605 6.105
R4022 S.n5567 S.t338 6.105
R4023 S.n5575 S.n5574 6.105
R4024 S.n5578 S.n5577 6.105
R4025 S.n5570 S.t714 6.105
R4026 S.n5279 S.t1002 6.105
R4027 S.n5290 S.n5289 6.105
R4028 S.n5287 S.n5286 6.105
R4029 S.n5282 S.t135 6.105
R4030 S.n5102 S.t340 6.105
R4031 S.n5110 S.n5109 6.105
R4032 S.n5113 S.n5112 6.105
R4033 S.n5105 S.t17 6.105
R4034 S.n5245 S.t299 6.105
R4035 S.n5254 S.n5253 6.105
R4036 S.n5257 S.n5256 6.105
R4037 S.n5248 S.t887 6.105
R4038 S.n4651 S.t1130 6.105
R4039 S.n4662 S.n4661 6.105
R4040 S.n4665 S.n4664 6.105
R4041 S.n4654 S.t578 6.105
R4042 S.n4374 S.t594 6.105
R4043 S.n3713 S.t106 6.105
R4044 S.n3721 S.n3720 6.105
R4045 S.n3724 S.n3723 6.105
R4046 S.n3716 S.t655 6.105
R4047 S.n3937 S.t428 6.105
R4048 S.n3944 S.n3943 6.105
R4049 S.n3941 S.n3940 6.105
R4050 S.n3934 S.t945 6.105
R4051 S.n5785 S.t273 6.105
R4052 S.n5538 S.t1104 6.105
R4053 S.n5543 S.n5542 6.105
R4054 S.n5546 S.n5545 6.105
R4055 S.n5535 S.t381 6.105
R4056 S.n5313 S.t645 6.105
R4057 S.n5320 S.n5319 6.105
R4058 S.n5317 S.n5316 6.105
R4059 S.n5310 S.t917 6.105
R4060 S.n5068 S.t1135 6.105
R4061 S.n5073 S.n5072 6.105
R4062 S.n5076 S.n5075 6.105
R4063 S.n5065 S.t804 6.105
R4064 S.n5215 S.t1038 6.105
R4065 S.n5219 S.n5218 6.105
R4066 S.n5222 S.n5221 6.105
R4067 S.n5212 S.t206 6.105
R4068 S.n4617 S.t1119 6.105
R4069 S.n4622 S.n4621 6.105
R4070 S.n4625 S.n4624 6.105
R4071 S.n4614 S.t793 6.105
R4072 S.n4777 S.t1018 6.105
R4073 S.n4781 S.n4780 6.105
R4074 S.n4784 S.n4783 6.105
R4075 S.n4774 S.t182 6.105
R4076 S.n4198 S.t1103 6.105
R4077 S.n4203 S.n4202 6.105
R4078 S.n4206 S.n4205 6.105
R4079 S.n4195 S.t783 6.105
R4080 S.n3906 S.t962 6.105
R4081 S.n3203 S.t699 6.105
R4082 S.n3211 S.n3210 6.105
R4083 S.n3214 S.n3213 6.105
R4084 S.n3206 S.t198 6.105
R4085 S.n3452 S.t201 6.105
R4086 S.n3459 S.n3458 6.105
R4087 S.n3456 S.n3455 6.105
R4088 S.n3449 S.t480 6.105
R4089 S.n5778 S.t615 6.105
R4090 S.n5522 S.t324 6.105
R4091 S.n5527 S.n5526 6.105
R4092 S.n5530 S.n5529 6.105
R4093 S.n5519 S.t771 6.105
R4094 S.n5328 S.t1026 6.105
R4095 S.n5335 S.n5334 6.105
R4096 S.n5332 S.n5331 6.105
R4097 S.n5325 S.t190 6.105
R4098 S.n5052 S.t417 6.105
R4099 S.n5057 S.n5056 6.105
R4100 S.n5060 S.n5059 6.105
R4101 S.n5049 S.t72 6.105
R4102 S.n5200 S.t267 6.105
R4103 S.n5204 S.n5203 6.105
R4104 S.n5207 S.n5206 6.105
R4105 S.n5197 S.t590 6.105
R4106 S.n4601 S.t406 6.105
R4107 S.n4606 S.n4605 6.105
R4108 S.n4609 S.n4608 6.105
R4109 S.n4598 S.t51 6.105
R4110 S.n4762 S.t269 6.105
R4111 S.n4766 S.n4765 6.105
R4112 S.n4769 S.n4768 6.105
R4113 S.n4759 S.t582 6.105
R4114 S.n4182 S.t380 6.105
R4115 S.n4187 S.n4186 6.105
R4116 S.n4190 S.n4189 6.105
R4117 S.n4179 S.t39 6.105
R4118 S.n3952 S.t294 6.105
R4119 S.n3959 S.n3958 6.105
R4120 S.n3956 S.n3955 6.105
R4121 S.n3949 S.t549 6.105
R4122 S.n3700 S.t369 6.105
R4123 S.n3705 S.n3704 6.105
R4124 S.n3708 S.n3707 6.105
R4125 S.n3697 S.t23 6.105
R4126 S.n3421 S.t954 6.105
R4127 S.n2670 S.t231 6.105
R4128 S.n2678 S.n2677 6.105
R4129 S.n2681 S.n2680 6.105
R4130 S.n2673 S.t797 6.105
R4131 S.n2956 S.t789 6.105
R4132 S.n2963 S.n2962 6.105
R4133 S.n2960 S.n2959 6.105
R4134 S.n2953 S.t249 6.105
R4135 S.n5771 S.t980 6.105
R4136 S.n5506 S.t772 6.105
R4137 S.n5511 S.n5510 6.105
R4138 S.n5514 S.n5513 6.105
R4139 S.n5503 S.t1143 6.105
R4140 S.n5343 S.t261 6.105
R4141 S.n5350 S.n5349 6.105
R4142 S.n5347 S.n5346 6.105
R4143 S.n5340 S.t508 6.105
R4144 S.n5036 S.t787 6.105
R4145 S.n5041 S.n5040 6.105
R4146 S.n5044 S.n5043 6.105
R4147 S.n5033 S.t463 6.105
R4148 S.n5185 S.t695 6.105
R4149 S.n5189 S.n5188 6.105
R4150 S.n5192 S.n5191 6.105
R4151 S.n5182 S.t972 6.105
R4152 S.n4585 S.t745 6.105
R4153 S.n4590 S.n4589 6.105
R4154 S.n4593 S.n4592 6.105
R4155 S.n4582 S.t448 6.105
R4156 S.n4747 S.t681 6.105
R4157 S.n4751 S.n4750 6.105
R4158 S.n4754 S.n4753 6.105
R4159 S.n4744 S.t947 6.105
R4160 S.n4166 S.t770 6.105
R4161 S.n4171 S.n4170 6.105
R4162 S.n4174 S.n4173 6.105
R4163 S.n4163 S.t440 6.105
R4164 S.n3967 S.t661 6.105
R4165 S.n3974 S.n3973 6.105
R4166 S.n3971 S.n3970 6.105
R4167 S.n3964 S.t942 6.105
R4168 S.n3684 S.t754 6.105
R4169 S.n3689 S.n3688 6.105
R4170 S.n3692 S.n3691 6.105
R4171 S.n3681 S.t393 6.105
R4172 S.n3467 S.t288 6.105
R4173 S.n3474 S.n3473 6.105
R4174 S.n3471 S.n3470 6.105
R4175 S.n3464 S.t932 6.105
R4176 S.n3190 S.t728 6.105
R4177 S.n3195 S.n3194 6.105
R4178 S.n3198 S.n3197 6.105
R4179 S.n3187 S.t427 6.105
R4180 S.n2925 S.t217 6.105
R4181 S.n2127 S.t814 6.105
R4182 S.n2135 S.n2134 6.105
R4183 S.n2138 S.n2137 6.105
R4184 S.n2130 S.t292 6.105
R4185 S.n2434 S.t257 6.105
R4186 S.n2441 S.n2440 6.105
R4187 S.n2438 S.n2437 6.105
R4188 S.n2431 S.t842 6.105
R4189 S.n5764 S.t244 6.105
R4190 S.n5490 S.t1149 6.105
R4191 S.n5495 S.n5494 6.105
R4192 S.n5498 S.n5497 6.105
R4193 S.n5487 S.t432 6.105
R4194 S.n5358 S.t640 6.105
R4195 S.n5365 S.n5364 6.105
R4196 S.n5362 S.n5361 6.105
R4197 S.n5355 S.t880 6.105
R4198 S.n5020 S.t46 6.105
R4199 S.n5025 S.n5024 6.105
R4200 S.n5028 S.n5027 6.105
R4201 S.n5017 S.t845 6.105
R4202 S.n5170 S.t1019 6.105
R4203 S.n5174 S.n5173 6.105
R4204 S.n5177 S.n5176 6.105
R4205 S.n5167 S.t178 6.105
R4206 S.n4569 S.t5 6.105
R4207 S.n4574 S.n4573 6.105
R4208 S.n4577 S.n4576 6.105
R4209 S.n4566 S.t834 6.105
R4210 S.n4732 S.t1063 6.105
R4211 S.n4736 S.n4735 6.105
R4212 S.n4739 S.n4738 6.105
R4213 S.n4729 S.t235 6.105
R4214 S.n4150 S.t1146 6.105
R4215 S.n4155 S.n4154 6.105
R4216 S.n4158 S.n4157 6.105
R4217 S.n4147 S.t824 6.105
R4218 S.n3982 S.t1021 6.105
R4219 S.n3989 S.n3988 6.105
R4220 S.n3986 S.n3985 6.105
R4221 S.n3979 S.t219 6.105
R4222 S.n3668 S.t1087 6.105
R4223 S.n3673 S.n3672 6.105
R4224 S.n3676 S.n3675 6.105
R4225 S.n3665 S.t806 6.105
R4226 S.n3482 S.t658 6.105
R4227 S.n3489 S.n3488 6.105
R4228 S.n3486 S.n3485 6.105
R4229 S.n3479 S.t199 6.105
R4230 S.n3174 S.t1121 6.105
R4231 S.n3179 S.n3178 6.105
R4232 S.n3182 S.n3181 6.105
R4233 S.n3171 S.t794 6.105
R4234 S.n2971 S.t652 6.105
R4235 S.n2978 S.n2977 6.105
R4236 S.n2975 S.n2974 6.105
R4237 S.n2968 S.t928 6.105
R4238 S.n2657 S.t1108 6.105
R4239 S.n2662 S.n2661 6.105
R4240 S.n2665 S.n2664 6.105
R4241 S.n2654 S.t786 6.105
R4242 S.n2402 S.t589 6.105
R4243 S.n1319 S.t286 6.105
R4244 S.n1536 S.n1535 6.105
R4245 S.n1539 S.n1538 6.105
R4246 S.n1542 S.t933 6.105
R4247 S.n1906 S.t882 6.105
R4248 S.n1914 S.n1913 6.105
R4249 S.n1911 S.n1910 6.105
R4250 S.n1903 S.t265 6.105
R4251 S.n5757 S.t635 6.105
R4252 S.n5587 S.t433 6.105
R4253 S.n5584 S.n5583 6.105
R4254 S.n5581 S.n5580 6.105
R4255 S.n5378 S.t801 6.105
R4256 S.n5373 S.t1007 6.105
R4257 S.n5597 S.n5596 6.105
R4258 S.n5594 S.n5593 6.105
R4259 S.n5370 S.t166 6.105
R4260 S.n5153 S.t395 6.105
R4261 S.n5150 S.n5149 6.105
R4262 S.n5147 S.n5146 6.105
R4263 S.n5144 S.t107 6.105
R4264 S.n5139 S.t271 6.105
R4265 S.n5159 S.n5158 6.105
R4266 S.n5162 S.n5161 6.105
R4267 S.n5136 S.t538 6.105
R4268 S.n4554 S.t436 6.105
R4269 S.n4558 S.n4557 6.105
R4270 S.n4561 S.n4560 6.105
R4271 S.n4551 S.t98 6.105
R4272 S.n4716 S.t287 6.105
R4273 S.n4721 S.n4720 6.105
R4274 S.n4724 S.n4723 6.105
R4275 S.n4713 S.t568 6.105
R4276 S.n4135 S.t430 6.105
R4277 S.n4139 S.n4138 6.105
R4278 S.n4142 S.n4141 6.105
R4279 S.n4132 S.t88 6.105
R4280 S.n3997 S.t323 6.105
R4281 S.n4005 S.n4004 6.105
R4282 S.n4002 S.n4001 6.105
R4283 S.n3994 S.t616 6.105
R4284 S.n3653 S.t418 6.105
R4285 S.n3657 S.n3656 6.105
R4286 S.n3660 S.n3659 6.105
R4287 S.n3650 S.t73 6.105
R4288 S.n3497 S.t1048 6.105
R4289 S.n3505 S.n3504 6.105
R4290 S.n3502 S.n3501 6.105
R4291 S.n3494 S.t591 6.105
R4292 S.n3159 S.t408 6.105
R4293 S.n3163 S.n3162 6.105
R4294 S.n3166 S.n3165 6.105
R4295 S.n3156 S.t48 6.105
R4296 S.n2986 S.t1032 6.105
R4297 S.n2994 S.n2993 6.105
R4298 S.n2991 S.n2990 6.105
R4299 S.n2983 S.t197 6.105
R4300 S.n2642 S.t383 6.105
R4301 S.n2646 S.n2645 6.105
R4302 S.n2649 S.n2648 6.105
R4303 S.n2639 S.t43 6.105
R4304 S.n2449 S.t1024 6.105
R4305 S.n2457 S.n2456 6.105
R4306 S.n2454 S.n2453 6.105
R4307 S.n2446 S.t187 6.105
R4308 S.n2115 S.t374 6.105
R4309 S.n2119 S.n2118 6.105
R4310 S.n2122 S.n2121 6.105
R4311 S.n2112 S.t26 6.105
R4312 S.n1874 S.t956 6.105
R4313 S.n965 S.t916 6.105
R4314 S.n973 S.n972 6.105
R4315 S.n976 S.n975 6.105
R4316 S.n968 S.t435 6.105
R4317 S.n1573 S.t376 6.105
R4318 S.n1580 S.n1579 6.105
R4319 S.n1577 S.n1576 6.105
R4320 S.n1570 S.t950 6.105
R4321 S.n5748 S.t353 6.105
R4322 S.n5473 S.t802 6.105
R4323 S.n5479 S.n5478 6.105
R4324 S.n5482 S.n5481 6.105
R4325 S.n5470 S.t67 6.105
R4326 S.n5605 S.t285 6.105
R4327 S.n5616 S.n5615 6.105
R4328 S.n5613 S.n5612 6.105
R4329 S.n5602 S.t557 6.105
R4330 S.n5122 S.t810 6.105
R4331 S.n5119 S.n5118 6.105
R4332 S.n5116 S.n5115 6.105
R4333 S.n4941 S.t467 6.105
R4334 S.n4936 S.t667 6.105
R4335 S.n5128 S.n5127 6.105
R4336 S.n5131 S.n5130 6.105
R4337 S.n4933 S.t949 6.105
R4338 S.n4539 S.t816 6.105
R4339 S.n4543 S.n4542 6.105
R4340 S.n4546 S.n4545 6.105
R4341 S.n4536 S.t493 6.105
R4342 S.n4700 S.t609 6.105
R4343 S.n4705 S.n4704 6.105
R4344 S.n4708 S.n4707 6.105
R4345 S.n4697 S.t936 6.105
R4346 S.n4120 S.t800 6.105
R4347 S.n4124 S.n4123 6.105
R4348 S.n4127 S.n4126 6.105
R4349 S.n4117 S.t482 6.105
R4350 S.n4013 S.t651 6.105
R4351 S.n4021 S.n4020 6.105
R4352 S.n4018 S.n4017 6.105
R4353 S.n4010 S.t927 6.105
R4354 S.n3638 S.t790 6.105
R4355 S.n3642 S.n3641 6.105
R4356 S.n3645 S.n3644 6.105
R4357 S.n3635 S.t475 6.105
R4358 S.n3513 S.t315 6.105
R4359 S.n3521 S.n3520 6.105
R4360 S.n3518 S.n3517 6.105
R4361 S.n3510 S.t974 6.105
R4362 S.n3144 S.t781 6.105
R4363 S.n3148 S.n3147 6.105
R4364 S.n3151 S.n3150 6.105
R4365 S.n3141 S.t454 6.105
R4366 S.n3002 S.t308 6.105
R4367 S.n3010 S.n3009 6.105
R4368 S.n3007 S.n3006 6.105
R4369 S.n2999 S.t585 6.105
R4370 S.n2627 S.t775 6.105
R4371 S.n2631 S.n2630 6.105
R4372 S.n2634 S.n2633 6.105
R4373 S.n2624 S.t443 6.105
R4374 S.n2465 S.t298 6.105
R4375 S.n2473 S.n2472 6.105
R4376 S.n2470 S.n2469 6.105
R4377 S.n2462 S.t577 6.105
R4378 S.n2100 S.t756 6.105
R4379 S.n2104 S.n2103 6.105
R4380 S.n2107 S.n2106 6.105
R4381 S.n2097 S.t397 6.105
R4382 S.n1922 S.t291 6.105
R4383 S.n1930 S.n1929 6.105
R4384 S.n1927 S.n1926 6.105
R4385 S.n1919 S.t570 6.105
R4386 S.n1525 S.t735 6.105
R4387 S.n1530 S.n1529 6.105
R4388 S.n1533 S.n1532 6.105
R4389 S.n1522 S.t429 6.105
R4390 S.n1311 S.t420 6.105
R4391 S.n5731 S.t1013 6.105
R4392 S.n5272 S.t171 6.105
R4393 S.n719 S.t175 6.105
R4394 S.n585 S.t1040 6.105
R4395 S.n575 S.t13 6.105
R4396 S.n382 S.t502 6.105
R4397 S.n406 S.n405 6.105
R4398 S.n403 S.n402 6.105
R4399 S.n385 S.t1035 6.105
R4400 S.n1048 S.t148 6.105
R4401 S.n1058 S.n1057 6.105
R4402 S.n1061 S.n1060 6.105
R4403 S.n1045 S.t387 6.105
R4404 S.n5401 S.t391 6.105
R4405 S.n5380 S.t890 6.105
R4406 S.n5645 S.t1133 6.105
R4407 S.n5663 S.n5662 6.105
R4408 S.n5660 S.n5659 6.105
R4409 S.n5642 S.t252 6.105
R4410 S.n4970 S.t657 6.105
R4411 S.n4981 S.n4980 6.105
R4412 S.n4978 S.n4977 6.105
R4413 S.n4967 S.t747 6.105
R4414 S.n4869 S.t966 6.105
R4415 S.n4884 S.n4883 6.105
R4416 S.n4881 S.n4880 6.105
R4417 S.n4866 S.t76 6.105
R4418 S.n4519 S.t477 6.105
R4419 S.n4530 S.n4529 6.105
R4420 S.n4527 S.n4526 6.105
R4421 S.n4516 S.t134 6.105
R4422 S.n4422 S.t320 6.105
R4423 S.n4437 S.n4436 6.105
R4424 S.n4434 S.n4433 6.105
R4425 S.n4419 S.t593 6.105
R4426 S.n4100 S.t456 6.105
R4427 S.n4111 S.n4110 6.105
R4428 S.n4108 S.n4107 6.105
R4429 S.n4097 S.t124 6.105
R4430 S.n4295 S.t307 6.105
R4431 S.n4307 S.n4306 6.105
R4432 S.n4310 S.n4309 6.105
R4433 S.n4292 S.t533 6.105
R4434 S.n3618 S.t447 6.105
R4435 S.n3629 S.n3628 6.105
R4436 S.n3626 S.n3625 6.105
R4437 S.n3615 S.t116 6.105
R4438 S.n3799 S.t1027 6.105
R4439 S.n3811 S.n3810 6.105
R4440 S.n3814 S.n3813 6.105
R4441 S.n3796 S.t575 6.105
R4442 S.n3124 S.t438 6.105
R4443 S.n3135 S.n3134 6.105
R4444 S.n3132 S.n3131 6.105
R4445 S.n3121 S.t101 6.105
R4446 S.n3284 S.t1005 6.105
R4447 S.n3296 S.n3295 6.105
R4448 S.n3299 S.n3298 6.105
R4449 S.n3281 S.t174 6.105
R4450 S.n2607 S.t431 6.105
R4451 S.n2618 S.n2617 6.105
R4452 S.n2615 S.n2614 6.105
R4453 S.n2604 S.t89 6.105
R4454 S.n2756 S.t1059 6.105
R4455 S.n2768 S.n2767 6.105
R4456 S.n2771 S.n2770 6.105
R4457 S.n2753 S.t233 6.105
R4458 S.n2080 S.t423 6.105
R4459 S.n2091 S.n2090 6.105
R4460 S.n2088 S.n2087 6.105
R4461 S.n2077 S.t3 6.105
R4462 S.n2207 S.t1050 6.105
R4463 S.n2218 S.n2217 6.105
R4464 S.n2221 S.n2220 6.105
R4465 S.n2204 S.t216 6.105
R4466 S.n1488 S.t400 6.105
R4467 S.n1500 S.n1499 6.105
R4468 S.n1497 S.n1496 6.105
R4469 S.n1485 S.t63 6.105
R4470 S.n1643 S.t1033 6.105
R4471 S.n1655 S.n1654 6.105
R4472 S.n1658 S.n1657 6.105
R4473 S.n1640 S.t205 6.105
R4474 S.n948 S.t390 6.105
R4475 S.n959 S.n958 6.105
R4476 S.n956 S.n955 6.105
R4477 S.n945 S.t44 6.105
R4478 S.n360 S.t229 6.105
R4479 S.n363 S.n362 6.105
R4480 S.n366 S.n365 6.105
R4481 S.n369 S.t989 6.105
R4482 S.n284 S.t682 6.105
R4483 S.n295 S.n294 6.105
R4484 S.n298 S.n297 6.105
R4485 S.n287 S.t604 6.105
R4486 S.n442 S.t784 6.105
R4487 S.n5739 S.t733 6.105
R4488 S.n5454 S.t53 6.105
R4489 S.n5462 S.n5461 6.105
R4490 S.n5465 S.n5464 6.105
R4491 S.n5457 S.t509 6.105
R4492 S.n5624 S.t750 6.105
R4493 S.n5635 S.n5634 6.105
R4494 S.n5632 S.n5631 6.105
R4495 S.n5627 S.t985 6.105
R4496 S.n5001 S.t71 6.105
R4497 S.n5009 S.n5008 6.105
R4498 S.n5012 S.n5011 6.105
R4499 S.n5004 S.t875 6.105
R4500 S.n4917 S.t1053 6.105
R4501 S.n4925 S.n4924 6.105
R4502 S.n4928 S.n4927 6.105
R4503 S.n4920 S.t226 6.105
R4504 S.n4467 S.t74 6.105
R4505 S.n4668 S.n4667 6.105
R4506 S.n4671 S.n4670 6.105
R4507 S.n4674 S.t861 6.105
R4508 S.n4681 S.t1047 6.105
R4509 S.n4689 S.n4688 6.105
R4510 S.n4692 S.n4691 6.105
R4511 S.n4684 S.t211 6.105
R4512 S.n4025 S.t66 6.105
R4513 S.n4225 S.n4224 6.105
R4514 S.n4228 S.n4227 6.105
R4515 S.n4231 S.t851 6.105
R4516 S.n4238 S.t1029 6.105
R4517 S.n4249 S.n4248 6.105
R4518 S.n4246 S.n4245 6.105
R4519 S.n4241 S.t196 6.105
R4520 S.n3525 S.t55 6.105
R4521 S.n3727 S.n3726 6.105
R4522 S.n3730 S.n3729 6.105
R4523 S.n3733 S.t846 6.105
R4524 S.n3740 S.t602 6.105
R4525 S.n3751 S.n3750 6.105
R4526 S.n3748 S.n3747 6.105
R4527 S.n3743 S.t185 6.105
R4528 S.n3014 S.t28 6.105
R4529 S.n3217 S.n3216 6.105
R4530 S.n3220 S.n3219 6.105
R4531 S.n3223 S.t838 6.105
R4532 S.n3230 S.t687 6.105
R4533 S.n3241 S.n3240 6.105
R4534 S.n3238 S.n3237 6.105
R4535 S.n3233 S.t968 6.105
R4536 S.n2477 S.t1148 6.105
R4537 S.n2684 S.n2683 6.105
R4538 S.n2687 S.n2686 6.105
R4539 S.n2690 S.t825 6.105
R4540 S.n2697 S.t672 6.105
R4541 S.n2708 S.n2707 6.105
R4542 S.n2705 S.n2704 6.105
R4543 S.n2700 S.t953 6.105
R4544 S.n1934 S.t1140 6.105
R4545 S.n2141 S.n2140 6.105
R4546 S.n2144 S.n2143 6.105
R4547 S.n2147 S.t813 6.105
R4548 S.n2154 S.t659 6.105
R4549 S.n2165 S.n2164 6.105
R4550 S.n2162 S.n2161 6.105
R4551 S.n2157 S.t940 6.105
R4552 S.n1506 S.t1089 6.105
R4553 S.n1514 S.n1513 6.105
R4554 S.n1517 S.n1516 6.105
R4555 S.n1509 S.t795 6.105
R4556 S.n1584 S.t654 6.105
R4557 S.n1595 S.n1594 6.105
R4558 S.n1592 S.n1591 6.105
R4559 S.n1587 S.t930 6.105
R4560 S.n761 S.t1111 6.105
R4561 S.n979 S.n978 6.105
R4562 S.n982 S.n981 6.105
R4563 S.n985 S.t788 6.105
R4564 S.n992 S.t995 6.105
R4565 S.n1007 S.n1006 6.105
R4566 S.n1004 S.n1003 6.105
R4567 S.n995 S.t457 6.105
R4568 S.n622 S.t650 6.105
R4569 S.n615 S.t991 6.105
R4570 S.n97 S.t884 6.105
R4571 S.n108 S.n107 6.105
R4572 S.n105 S.n104 6.105
R4573 S.n100 S.t1117 6.105
R4574 S.n1201 S.t904 6.105
R4575 S.n1211 S.n1210 6.105
R4576 S.n1214 S.n1213 6.105
R4577 S.n1198 S.t1132 6.105
R4578 S.n3032 S.t415 6.105
R4579 S.n3016 S.t542 6.105
R4580 S.n3249 S.t856 6.105
R4581 S.n3266 S.n3265 6.105
R4582 S.n3263 S.n3262 6.105
R4583 S.n3246 S.t1080 6.105
R4584 S.n2505 S.t215 6.105
R4585 S.n2516 S.n2515 6.105
R4586 S.n2513 S.n2512 6.105
R4587 S.n2502 S.t274 6.105
R4588 S.n2905 S.t608 6.105
R4589 S.n2917 S.n2916 6.105
R4590 S.n2920 S.n2919 6.105
R4591 S.n2902 S.t841 6.105
R4592 S.n1980 S.t92 6.105
R4593 S.n1991 S.n1990 6.105
R4594 S.n1988 S.n1987 6.105
R4595 S.n1977 S.t888 6.105
R4596 S.n2350 S.t675 6.105
R4597 S.n2361 S.n2360 6.105
R4598 S.n2364 S.n2363 6.105
R4599 S.n2347 S.t961 6.105
R4600 S.n1386 S.t83 6.105
R4601 S.n1398 S.n1397 6.105
R4602 S.n1395 S.n1394 6.105
R4603 S.n1383 S.t866 6.105
R4604 S.n1789 S.t666 6.105
R4605 S.n1801 S.n1800 6.105
R4606 S.n1804 S.n1803 6.105
R4607 S.n1786 S.t944 6.105
R4608 S.n843 S.t70 6.105
R4609 S.n854 S.n853 6.105
R4610 S.n851 S.n850 6.105
R4611 S.n840 S.t855 6.105
R4612 S.n716 S.t279 6.105
R4613 S.n717 S.t626 6.105
R4614 S.n12 S.t574 6.105
R4615 S.n468 S.n467 6.105
R4616 S.n471 S.n470 6.105
R4617 S.n474 S.t739 6.105
R4618 S.n3544 S.t264 6.105
R4619 S.n3527 S.t399 6.105
R4620 S.n3763 S.t723 6.105
R4621 S.n3781 S.n3780 6.105
R4622 S.n3778 S.n3777 6.105
R4623 S.n3766 S.t819 6.105
R4624 S.n3041 S.t64 6.105
R4625 S.n3052 S.n3051 6.105
R4626 S.n3049 S.n3048 6.105
R4627 S.n3044 S.t133 6.105
R4628 S.n3396 S.t486 6.105
R4629 S.n3413 S.n3412 6.105
R4630 S.n3416 S.n3415 6.105
R4631 S.n3399 S.t693 6.105
R4632 S.n2524 S.t830 6.105
R4633 S.n2535 S.n2534 6.105
R4634 S.n2532 S.n2531 6.105
R4635 S.n2527 S.t520 6.105
R4636 S.n2868 S.t311 6.105
R4637 S.n2885 S.n2884 6.105
R4638 S.n2888 S.n2887 6.105
R4639 S.n2871 S.t595 6.105
R4640 S.n1997 S.t828 6.105
R4641 S.n2008 S.n2007 6.105
R4642 S.n2005 S.n2004 6.105
R4643 S.n2000 S.t506 6.105
R4644 S.n2313 S.t302 6.105
R4645 S.n2330 S.n2329 6.105
R4646 S.n2333 S.n2332 6.105
R4647 S.n2316 S.t539 6.105
R4648 S.n1404 S.t817 6.105
R4649 S.n1415 S.n1414 6.105
R4650 S.n1412 S.n1411 6.105
R4651 S.n1407 S.t495 6.105
R4652 S.n1752 S.t295 6.105
R4653 S.n1769 S.n1768 6.105
R4654 S.n1772 S.n1771 6.105
R4655 S.n1755 S.t573 6.105
R4656 S.n860 S.t805 6.105
R4657 S.n873 S.n872 6.105
R4658 S.n870 S.n869 6.105
R4659 S.n863 S.t485 6.105
R4660 S.n881 S.t414 6.105
R4661 S.n895 S.n894 6.105
R4662 S.n892 S.n891 6.105
R4663 S.n884 S.t9 6.105
R4664 S.n1132 S.t193 6.105
R4665 S.n1153 S.n1152 6.105
R4666 S.n1156 S.n1155 6.105
R4667 S.n1135 S.t398 6.105
R4668 S.n112 S.t245 6.105
R4669 S.n301 S.n300 6.105
R4670 S.n304 S.n303 6.105
R4671 S.n307 S.t1006 6.105
R4672 S.n315 S.t184 6.105
R4673 S.n330 S.n329 6.105
R4674 S.n327 S.n326 6.105
R4675 S.n318 S.t425 6.105
R4676 S.n637 S.t999 6.105
R4677 S.n629 S.t242 6.105
R4678 S.n1728 S.t1011 6.105
R4679 S.n1740 S.n1739 6.105
R4680 S.n1743 S.n1742 6.105
R4681 S.n1725 S.t177 6.105
R4682 S.n2290 S.t1017 6.105
R4683 S.n2301 S.n2300 6.105
R4684 S.n2304 S.n2303 6.105
R4685 S.n2287 S.t194 6.105
R4686 S.n2840 S.t1043 6.105
R4687 S.n2852 S.n2851 6.105
R4688 S.n2855 S.n2854 6.105
R4689 S.n2837 S.t209 6.105
R4690 S.n3368 S.t1052 6.105
R4691 S.n3380 S.n3379 6.105
R4692 S.n3383 S.n3382 6.105
R4693 S.n3365 S.t224 6.105
R4694 S.n3886 S.t347 6.105
R4695 S.n3898 S.n3897 6.105
R4696 S.n3901 S.n3900 6.105
R4697 S.n3883 S.t464 6.105
R4698 S.n4260 S.t491 6.105
R4699 S.n4277 S.n4276 6.105
R4700 S.n4274 S.n4273 6.105
R4701 S.n4257 S.t690 6.105
R4702 S.n4043 S.t147 6.105
R4703 S.n4027 S.t258 6.105
R4704 S.n3553 S.t1030 6.105
R4705 S.n3564 S.n3563 6.105
R4706 S.n3561 S.n3560 6.105
R4707 S.n3550 S.t1124 6.105
R4708 S.n3060 S.t478 6.105
R4709 S.n3071 S.n3070 6.105
R4710 S.n3068 S.n3067 6.105
R4711 S.n3057 S.t141 6.105
R4712 S.n2543 S.t458 6.105
R4713 S.n2554 S.n2553 6.105
R4714 S.n2551 S.n2550 6.105
R4715 S.n2540 S.t127 6.105
R4716 S.n2016 S.t446 6.105
R4717 S.n2027 S.n2026 6.105
R4718 S.n2024 S.n2023 6.105
R4719 S.n2013 S.t118 6.105
R4720 S.n1423 S.t439 6.105
R4721 S.n1435 S.n1434 6.105
R4722 S.n1432 S.n1431 6.105
R4723 S.n1420 S.t97 6.105
R4724 S.n1104 S.t926 6.105
R4725 S.n1119 S.n1118 6.105
R4726 S.n1122 S.n1121 6.105
R4727 S.n1107 S.t1 6.105
R4728 S.n240 S.t946 6.105
R4729 S.n259 S.n258 6.105
R4730 S.n256 S.n255 6.105
R4731 S.n243 S.t639 6.105
R4732 S.n646 S.t910 6.105
R4733 S.n649 S.n648 6.105
R4734 S.n652 S.n651 6.105
R4735 S.n655 S.t1090 6.105
R4736 S.n684 S.t638 6.105
R4737 S.n640 S.t964 6.105
R4738 S.n4488 S.t1134 6.105
R4739 S.n4469 S.t144 6.105
R4740 S.n4452 S.t357 6.105
R4741 S.n4460 S.n4459 6.105
R4742 S.n4463 S.n4462 6.105
R4743 S.n4449 S.t624 6.105
R4744 S.n4061 S.t937 6.105
R4745 S.n4070 S.n4069 6.105
R4746 S.n4067 S.n4066 6.105
R4747 S.n4058 S.t993 6.105
R4748 S.n4348 S.t93 6.105
R4749 S.n4366 S.n4365 6.105
R4750 S.n4369 S.n4368 6.105
R4751 S.n4345 S.t263 6.105
R4752 S.n3581 S.t7 6.105
R4753 S.n3590 S.n3589 6.105
R4754 S.n3587 S.n3586 6.105
R4755 S.n3578 S.t885 6.105
R4756 S.n3848 S.t683 6.105
R4757 S.n3866 S.n3865 6.105
R4758 S.n3869 S.n3868 6.105
R4759 S.n3845 S.t227 6.105
R4760 S.n3088 S.t80 6.105
R4761 S.n3096 S.n3095 6.105
R4762 S.n3093 S.n3092 6.105
R4763 S.n3085 S.t863 6.105
R4764 S.n3333 S.t662 6.105
R4765 S.n3348 S.n3347 6.105
R4766 S.n3351 S.n3350 6.105
R4767 S.n3330 S.t948 6.105
R4768 S.n2571 S.t69 6.105
R4769 S.n2579 S.n2578 6.105
R4770 S.n2576 S.n2575 6.105
R4771 S.n2568 S.t853 6.105
R4772 S.n2805 S.t618 6.105
R4773 S.n2820 S.n2819 6.105
R4774 S.n2823 S.n2822 6.105
R4775 S.n2802 S.t878 6.105
R4776 S.n2044 S.t57 6.105
R4777 S.n2052 S.n2051 6.105
R4778 S.n2049 S.n2048 6.105
R4779 S.n2041 S.t849 6.105
R4780 S.n2255 S.t648 6.105
R4781 S.n2270 S.n2269 6.105
R4782 S.n2273 S.n2272 6.105
R4783 S.n2252 S.t924 6.105
R4784 S.n1452 S.t33 6.105
R4785 S.n1460 S.n1459 6.105
R4786 S.n1457 S.n1456 6.105
R4787 S.n1449 S.t839 6.105
R4788 S.n1692 S.t694 6.105
R4789 S.n1707 S.n1706 6.105
R4790 S.n1710 S.n1709 6.105
R4791 S.n1689 S.t970 6.105
R4792 S.n911 S.t15 6.105
R4793 S.n919 S.n918 6.105
R4794 S.n916 S.n915 6.105
R4795 S.n908 S.t826 6.105
R4796 S.n1070 S.t531 6.105
R4797 S.n1086 S.n1085 6.105
R4798 S.n1089 S.n1088 6.105
R4799 S.n1073 S.t777 6.105
R4800 S.n264 S.t623 6.105
R4801 S.n278 S.n277 6.105
R4802 S.n275 S.n274 6.105
R4803 S.n267 S.t260 6.105
R4804 S.n931 S.t776 6.105
R4805 S.n940 S.n939 6.105
R4806 S.n937 S.n936 6.105
R4807 S.n928 S.t444 6.105
R4808 S.n1667 S.t309 6.105
R4809 S.n1675 S.n1674 6.105
R4810 S.n1678 S.n1677 6.105
R4811 S.n1670 S.t588 6.105
R4812 S.n1466 S.t742 6.105
R4813 S.n1480 S.n1479 6.105
R4814 S.n1477 S.n1476 6.105
R4815 S.n1469 S.t455 6.105
R4816 S.n2230 S.t317 6.105
R4817 S.n2238 S.n2237 6.105
R4818 S.n2241 S.n2240 6.105
R4819 S.n2233 S.t599 6.105
R4820 S.n2058 S.t792 6.105
R4821 S.n2072 S.n2071 6.105
R4822 S.n2069 S.n2068 6.105
R4823 S.n2061 S.t476 6.105
R4824 S.n2780 S.t282 6.105
R4825 S.n2788 S.n2787 6.105
R4826 S.n2791 S.n2790 6.105
R4827 S.n2783 S.t559 6.105
R4828 S.n2585 S.t799 6.105
R4829 S.n2599 S.n2598 6.105
R4830 S.n2596 S.n2595 6.105
R4831 S.n2588 S.t484 6.105
R4832 S.n3308 S.t293 6.105
R4833 S.n3316 S.n3315 6.105
R4834 S.n3319 S.n3318 6.105
R4835 S.n3311 S.t548 6.105
R4836 S.n3102 S.t821 6.105
R4837 S.n3116 S.n3115 6.105
R4838 S.n3113 S.n3112 6.105
R4839 S.n3105 S.t494 6.105
R4840 S.n3823 S.t259 6.105
R4841 S.n3831 S.n3830 6.105
R4842 S.n3834 S.n3833 6.105
R4843 S.n3826 S.t951 6.105
R4844 S.n3596 S.t827 6.105
R4845 S.n3610 S.n3609 6.105
R4846 S.n3607 S.n3606 6.105
R4847 S.n3599 S.t503 6.105
R4848 S.n4323 S.t673 6.105
R4849 S.n4331 S.n4330 6.105
R4850 S.n4334 S.n4333 6.105
R4851 S.n4326 S.t963 6.105
R4852 S.n4078 S.t840 6.105
R4853 S.n4092 S.n4091 6.105
R4854 S.n4089 S.n4088 6.105
R4855 S.n4081 S.t518 6.105
R4856 S.n4394 S.t1020 6.105
R4857 S.n4405 S.n4404 6.105
R4858 S.n4402 S.n4401 6.105
R4859 S.n4397 S.t234 6.105
R4860 S.n4497 S.t803 6.105
R4861 S.n4511 S.n4510 6.105
R4862 S.n4508 S.n4507 6.105
R4863 S.n4500 S.t871 6.105
R4864 S.n4898 S.t239 6.105
R4865 S.n4906 S.n4905 6.105
R4866 S.n4909 S.n4908 6.105
R4867 S.n4901 S.t479 6.105
R4868 S.n4961 S.t982 6.105
R4869 S.n4943 S.t1129 6.105
R4870 S.n701 S.t251 6.105
R4871 S.n688 S.t598 6.105
R4872 S.n339 S.t528 6.105
R4873 S.n356 S.n355 6.105
R4874 S.n353 S.n352 6.105
R4875 S.n342 S.t761 6.105
R4876 S.n1165 S.t517 6.105
R4877 S.n1181 S.n1180 6.105
R4878 S.n1184 S.n1183 6.105
R4879 S.n1168 S.t749 6.105
R4880 S.n224 S.t634 6.105
R4881 S.n235 S.n234 6.105
R4882 S.n232 S.n231 6.105
R4883 S.n227 S.t284 6.105
R4884 S.n207 S.t997 6.105
R4885 S.n218 S.n217 6.105
R4886 S.n215 S.n214 6.105
R4887 S.n210 S.t613 6.105
R4888 S.n610 S.t301 6.105
R4889 S.n603 S.t619 6.105
R4890 S.n65 S.t565 6.105
R4891 S.n76 S.n75 6.105
R4892 S.n73 S.n72 6.105
R4893 S.n68 S.t779 6.105
R4894 S.n1260 S.t572 6.105
R4895 S.n1270 S.n1269 6.105
R4896 S.n1273 S.n1272 6.105
R4897 S.n1257 S.t785 6.105
R4898 S.n1952 S.t643 6.105
R4899 S.n1936 S.t766 6.105
R4900 S.n2173 S.t1107 6.105
R4901 S.n2189 S.n2188 6.105
R4902 S.n2186 S.n2185 6.105
R4903 S.n2170 S.t243 6.105
R4904 S.n1347 S.t394 6.105
R4905 S.n1359 S.n1358 6.105
R4906 S.n1356 S.n1355 6.105
R4907 S.n1344 S.t523 6.105
R4908 S.n1854 S.t852 6.105
R4909 S.n1866 S.n1865 6.105
R4910 S.n1869 S.n1868 6.105
R4911 S.n1851 S.t1071 6.105
R4912 S.n807 S.t843 6.105
R4913 S.n818 S.n817 6.105
R4914 S.n815 S.n814 6.105
R4915 S.n804 S.t527 6.105
R4916 S.n712 S.t1031 6.105
R4917 S.n713 S.t275 6.105
R4918 S.n506 S.t161 6.105
R4919 S.n509 S.n508 6.105
R4920 S.n512 S.n511 6.105
R4921 S.n515 S.t404 6.105
R4922 S.n2496 S.t547 6.105
R4923 S.n2479 S.t641 6.105
R4924 S.n2720 S.t987 6.105
R4925 S.n2738 S.n2737 6.105
R4926 S.n2735 S.n2734 6.105
R4927 S.n2723 S.t102 6.105
R4928 S.n1961 S.t266 6.105
R4929 S.n1972 S.n1971 6.105
R4930 S.n1969 S.n1968 6.105
R4931 S.n1964 S.t405 6.105
R4932 S.n2377 S.t717 6.105
R4933 S.n2394 S.n2393 6.105
R4934 S.n2397 S.n2396 6.105
R4935 S.n2380 S.t975 6.105
R4936 S.n1367 S.t471 6.105
R4937 S.n1378 S.n1377 6.105
R4938 S.n1375 S.n1374 6.105
R4939 S.n1370 S.t109 6.105
R4940 S.n1817 S.t1015 6.105
R4941 S.n1834 S.n1833 6.105
R4942 S.n1837 S.n1836 6.105
R4943 S.n1820 S.t223 6.105
R4944 S.n824 S.t460 6.105
R4945 S.n835 S.n834 6.105
R4946 S.n832 S.n831 6.105
R4947 S.n827 S.t130 6.105
R4948 S.n1223 S.t169 6.105
R4949 S.n1240 S.n1239 6.105
R4950 S.n1243 S.n1242 6.105
R4951 S.n1226 S.t416 6.105
R4952 S.n189 S.t276 6.105
R4953 S.n200 S.n199 6.105
R4954 S.n197 S.n196 6.105
R4955 S.n192 S.t1042 6.105
R4956 S.n172 S.t603 6.105
R4957 S.n183 S.n182 6.105
R4958 S.n180 S.n179 6.105
R4959 S.n175 S.t319 6.105
R4960 S.n598 S.t1070 6.105
R4961 S.n590 S.t289 6.105
R4962 S.n33 S.t900 6.105
R4963 S.n44 S.n43 6.105
R4964 S.n41 S.n40 6.105
R4965 S.n36 S.t1123 6.105
R4966 S.n1015 S.t1147 6.105
R4967 S.n1030 S.n1029 6.105
R4968 S.n1027 S.n1026 6.105
R4969 S.n1012 S.t272 6.105
R4970 S.n779 S.t913 6.105
R4971 S.n763 S.t1004 6.105
R4972 S.n708 S.t685 6.105
R4973 S.n709 S.t1010 6.105
R4974 S.n544 S.t914 6.105
R4975 S.n547 S.n546 6.105
R4976 S.n550 S.n549 6.105
R4977 S.n553 S.t25 6.105
R4978 S.n1338 S.t744 6.105
R4979 S.n1321 S.t909 6.105
R4980 S.n1607 S.t111 6.105
R4981 S.n1625 S.n1624 6.105
R4982 S.n1622 S.n1621 6.105
R4983 S.n1610 S.t352 6.105
R4984 S.n788 S.t596 6.105
R4985 S.n799 S.n798 6.105
R4986 S.n796 S.n795 6.105
R4987 S.n791 S.t628 6.105
R4988 S.n1286 S.t764 6.105
R4989 S.n1303 S.n1302 6.105
R4990 S.n1306 S.n1305 6.105
R4991 S.n1289 S.t992 6.105
R4992 S.n154 S.t1022 6.105
R4993 S.n165 S.n164 6.105
R4994 S.n162 S.n161 6.105
R4995 S.n157 S.t703 6.105
R4996 S.n138 S.t606 6.105
R4997 S.n149 S.n148 6.105
R4998 S.n146 S.n145 6.105
R4999 S.n141 S.t617 6.105
R5000 S.n704 S.t798 6.105
R5001 S.n705 S.t709 6.105
R5002 S.n421 S.t152 6.105
R5003 S.n410 S.n409 6.105
R5004 S.n434 S.n433 6.105
R5005 S.n424 S.t410 6.105
R5006 S.n132 S.t952 6.105
R5007 S.n114 S.t1037 6.105
R5008 S.n726 S.t212 6.105
R5009 S.n5418 S.t1051 6.105
R5010 S.n5421 S.n5420 6.105
R5011 S.n5264 S.t960 6.105
R5012 S.n5830 S.t241 6.105
R5013 S.n5677 S.t87 6.105
R5014 S.n5685 S.n5684 6.105
R5015 S.n5688 S.n5687 6.105
R5016 S.n5680 S.t600 6.105
R5017 S.n4984 S.t556 6.105
R5018 S.n4995 S.n4994 6.105
R5019 S.n4992 S.n4991 6.105
R5020 S.n4987 S.t1016 6.105
R5021 S.n5411 S.t342 6.105
R5022 S.n5414 S.n5413 6.105
R5023 S.n5444 S.t996 6.105
R5024 S.n5447 S.n5446 6.105
R5025 S.n5439 S.t322 6.105
R5026 S.n5424 S.n5423 6.105
R5027 S.n5390 S.n5388 4.263
R5028 S.n454 S.n453 3.857
R5029 S.n745 S.n744 3.857
R5030 S.n1554 S.n1553 3.857
R5031 S.n1887 S.n1886 3.857
R5032 S.n2415 S.n2414 3.857
R5033 S.n2937 S.n2936 3.857
R5034 S.n3433 S.n3432 3.857
R5035 S.n3918 S.n3917 3.857
R5036 S.n4824 S.n4823 3.857
R5037 S.n4842 S.n4841 3.857
R5038 S.n5696 S.n5695 3.857
R5039 S.n5720 S.n5717 0.178
R5040 S.n580 S.n577 0.164
R5041 S.n5845 S.n5844 0.144
R5042 S.n451 S.n450 0.136
R5043 S.n739 S.n731 0.123
R5044 S.n558 S.n530 0.123
R5045 S.n593 S.n592 0.123
R5046 S.n570 S.n568 0.123
R5047 S.n456 S.n455 0.117
R5048 S.n747 S.n746 0.117
R5049 S.n1556 S.n1555 0.117
R5050 S.n1889 S.n1888 0.117
R5051 S.n2417 S.n2416 0.117
R5052 S.n2939 S.n2938 0.117
R5053 S.n3435 S.n3434 0.117
R5054 S.n3920 S.n3919 0.117
R5055 S.n4826 S.n4825 0.117
R5056 S.n4844 S.n4843 0.117
R5057 S.n5698 S.n5697 0.117
R5058 S.n5854 S.n1316 0.116
R5059 S.n5852 S.n2407 0.114
R5060 S.n5853 S.n1879 0.114
R5061 S.n5845 S.n5709 0.11
R5062 S.n5847 S.n4834 0.11
R5063 S.n5848 S.n4378 0.11
R5064 S.n5849 S.n3910 0.11
R5065 S.n5850 S.n3425 0.11
R5066 S.n5851 S.n2929 0.11
R5067 S.n5846 S.n5270 0.11
R5068 S.n5730 S.n5729 0.109
R5069 S.n4505 S.n4503 0.109
R5070 S.n4086 S.n4084 0.109
R5071 S.n3604 S.n3602 0.109
R5072 S.n3110 S.n3108 0.109
R5073 S.n2593 S.n2591 0.109
R5074 S.n2066 S.n2064 0.109
R5075 S.n1474 S.n1472 0.109
R5076 S.n924 S.n922 0.109
R5077 S.n85 S.n80 0.104
R5078 S.n53 S.n48 0.104
R5079 S.n21 S.n16 0.104
R5080 S.n1551 S.n1550 0.103
R5081 S.n1884 S.n1883 0.103
R5082 S.n2412 S.n2411 0.103
R5083 S.n2934 S.n2933 0.103
R5084 S.n3430 S.n3429 0.103
R5085 S.n3915 S.n3914 0.103
R5086 S.n4821 S.n4820 0.103
R5087 S.n4839 S.n4838 0.103
R5088 S.n5705 S.n5704 0.103
R5089 S.n1000 S.n999 0.097
R5090 S.n1080 S.n1079 0.097
R5091 S.n84 S.n81 0.097
R5092 S.n52 S.n49 0.097
R5093 S.n20 S.n17 0.097
R5094 S.n5667 S.n5666 0.096
R5095 S.n5384 S.n5383 0.093
R5096 S.n4946 S.n4945 0.093
R5097 S.n4493 S.n4492 0.093
R5098 S.n4074 S.n4073 0.093
R5099 S.n3037 S.n3035 0.093
R5100 S.n2520 S.n2518 0.093
R5101 S.n1957 S.n1955 0.093
R5102 S.n1363 S.n1361 0.093
R5103 S.n784 S.n782 0.093
R5104 S.n397 S.n393 0.092
R5105 S.n5428 S.n5427 0.092
R5106 S.n4064 S.n4063 0.091
R5107 S.n3584 S.n3583 0.091
R5108 S S.n5855 0.09
R5109 S.n1148 S.n1147 0.087
R5110 S.n461 S.n460 0.082
R5111 S.n752 S.n751 0.082
R5112 S.n1561 S.n1560 0.082
R5113 S.n1894 S.n1893 0.082
R5114 S.n2422 S.n2421 0.082
R5115 S.n2944 S.n2943 0.082
R5116 S.n3440 S.n3439 0.082
R5117 S.n3925 S.n3924 0.082
R5118 S.n4831 S.n4830 0.082
R5119 S.n4849 S.n4848 0.082
R5120 S.n5707 S.n5702 0.082
R5121 S.n1082 S.n1081 0.08
R5122 S.n5722 S.n5721 0.079
R5123 S.n292 S.n291 0.077
R5124 S.n901 S.n900 0.077
R5125 S.n1441 S.n1440 0.077
R5126 S.n2033 S.n2032 0.077
R5127 S.n2560 S.n2559 0.077
R5128 S.n3077 S.n3076 0.077
R5129 S.n3570 S.n3569 0.077
R5130 S.n4050 S.n4049 0.077
R5131 S.n253 S.n252 0.077
R5132 S.n272 S.n271 0.077
R5133 S.n4484 S.n4483 0.076
R5134 S.n5397 S.n5396 0.074
R5135 S.n4038 S.n4037 0.074
R5136 S.n4956 S.n4955 0.074
R5137 S.n3540 S.n3539 0.074
R5138 S.n3027 S.n3026 0.074
R5139 S.n2492 S.n2491 0.074
R5140 S.n1947 S.n1946 0.074
R5141 S.n774 S.n773 0.074
R5142 S.n1334 S.n1333 0.074
R5143 S.n127 S.n126 0.074
R5144 S.n5787 S.n5786 0.073
R5145 S.n5795 S.n5794 0.073
R5146 S.n5780 S.n5779 0.073
R5147 S.n5773 S.n5772 0.073
R5148 S.n5766 S.n5765 0.073
R5149 S.n5759 S.n5758 0.073
R5150 S.n5750 S.n5749 0.073
R5151 S.n5741 S.n5740 0.073
R5152 S.n5801 S.n5800 0.071
R5153 S.n5803 S.n5802 0.071
R5154 S.n1076 S.n1075 0.071
R5155 S.t240 S.n5753 0.068
R5156 S.t240 S.n5744 0.068
R5157 S.t240 S.n5726 0.068
R5158 S.n4831 S.n4818 0.067
R5159 S.n4831 S.n4817 0.067
R5160 S.n3925 S.n3912 0.067
R5161 S.n3925 S.n3911 0.067
R5162 S.n3440 S.n3427 0.067
R5163 S.n3440 S.n3426 0.067
R5164 S.n2944 S.n2931 0.067
R5165 S.n2944 S.n2930 0.067
R5166 S.n2422 S.n2409 0.067
R5167 S.n2422 S.n2408 0.067
R5168 S.n1894 S.n1881 0.067
R5169 S.n1894 S.n1880 0.067
R5170 S.n1561 S.n1548 0.067
R5171 S.n1561 S.n1547 0.067
R5172 S.n461 S.n448 0.067
R5173 S.n461 S.n446 0.067
R5174 S.n723 S.n722 0.067
R5175 S.n626 S.n624 0.067
R5176 S.n626 S.n625 0.067
R5177 S.n664 S.n663 0.067
R5178 S.n664 S.n662 0.067
R5179 S.n698 S.n696 0.067
R5180 S.n698 S.n697 0.067
R5181 S.n492 S.n481 0.067
R5182 S.n492 S.n480 0.067
R5183 S.n613 S.n611 0.067
R5184 S.n613 S.n612 0.067
R5185 S.n523 S.n522 0.067
R5186 S.n523 S.n521 0.067
R5187 S.n601 S.n599 0.067
R5188 S.n601 S.n600 0.067
R5189 S.n588 S.n586 0.067
R5190 S.n561 S.n560 0.067
R5191 S.n561 S.n559 0.067
R5192 S.n588 S.n587 0.067
R5193 S.n573 S.n572 0.067
R5194 S.n573 S.n571 0.067
R5195 S.n723 S.n721 0.067
R5196 S.n4849 S.n4836 0.067
R5197 S.n4849 S.n4835 0.067
R5198 S.n5707 S.n5706 0.067
R5199 S.n5707 S.n5693 0.067
R5200 S.n462 S.n444 0.064
R5201 S.n4658 S.n4657 0.064
R5202 S.n4852 S.n4849 0.063
R5203 S.n1056 S.n1055 0.063
R5204 S.n954 S.n953 0.063
R5205 S.n1653 S.n1652 0.063
R5206 S.n1495 S.n1494 0.063
R5207 S.n2216 S.n2215 0.063
R5208 S.n2086 S.n2085 0.063
R5209 S.n2766 S.n2765 0.063
R5210 S.n2613 S.n2612 0.063
R5211 S.n3294 S.n3293 0.063
R5212 S.n3130 S.n3129 0.063
R5213 S.n3809 S.n3808 0.063
R5214 S.n3624 S.n3623 0.063
R5215 S.n4305 S.n4304 0.063
R5216 S.n4106 S.n4105 0.063
R5217 S.n4525 S.n4524 0.063
R5218 S.n4976 S.n4975 0.063
R5219 S.n1151 S.n1127 0.063
R5220 S.n890 S.n876 0.063
R5221 S.n1738 S.n1737 0.063
R5222 S.n1430 S.n1429 0.063
R5223 S.n2299 S.n2298 0.063
R5224 S.n2022 S.n2021 0.063
R5225 S.n2850 S.n2849 0.063
R5226 S.n2549 S.n2548 0.063
R5227 S.n3066 S.n3065 0.063
R5228 S.n3559 S.n3558 0.063
R5229 S.n659 S.n658 0.063
R5230 S.n1084 S.n1064 0.063
R5231 S.n1673 S.n1661 0.063
R5232 S.n2236 S.n2224 0.063
R5233 S.n2786 S.n2774 0.063
R5234 S.n3314 S.n3302 0.063
R5235 S.n3829 S.n3817 0.063
R5236 S.n351 S.n335 0.063
R5237 S.n2328 S.n2307 0.063
R5238 S.n1767 S.n1746 0.063
R5239 S.n1179 S.n1160 0.063
R5240 S.n477 S.n8 0.063
R5241 S.n1209 S.n1208 0.063
R5242 S.n849 S.n848 0.063
R5243 S.n1799 S.n1798 0.063
R5244 S.n1393 S.n1392 0.063
R5245 S.n1986 S.n1985 0.063
R5246 S.n2511 S.n2510 0.063
R5247 S.n1238 S.n1218 0.063
R5248 S.n518 S.n500 0.063
R5249 S.n813 S.n812 0.063
R5250 S.n1354 S.n1353 0.063
R5251 S.n556 S.n532 0.063
R5252 S.n432 S.n431 0.063
R5253 S.n5608 S.n5607 0.062
R5254 S.n5610 S.n5609 0.062
R5255 S.n5621 S.n5618 0.062
R5256 S.n5620 S.n5619 0.062
R5257 S.n4914 S.n4911 0.062
R5258 S.n4913 S.n4912 0.062
R5259 S.n724 S.n723 0.062
R5260 S.n614 S.n613 0.062
R5261 S.n602 S.n601 0.062
R5262 S.n589 S.n588 0.062
R5263 S.n675 S.n664 0.061
R5264 S.n493 S.n492 0.06
R5265 S.n524 S.n523 0.06
R5266 S.n562 S.n561 0.06
R5267 S.n574 S.n573 0.06
R5268 S.n5654 S.n5653 0.059
R5269 S.n4888 S.n4887 0.059
R5270 S.n4384 S.n4383 0.059
R5271 S.n4313 S.n4312 0.059
R5272 S.n3388 S.n3387 0.059
R5273 S.n2860 S.n2859 0.059
R5274 S.n2369 S.n2368 0.059
R5275 S.n1809 S.n1808 0.059
R5276 S.n1278 S.n1277 0.059
R5277 S.n1723 S.n1713 0.059
R5278 S.n627 S.n626 0.059
R5279 S.n1895 S.n1894 0.058
R5280 S.n1562 S.n1561 0.058
R5281 S.n462 S.n461 0.058
R5282 S.n5708 S.n5707 0.058
R5283 S.n3926 S.n3925 0.058
R5284 S.n3441 S.n3440 0.058
R5285 S.n2945 S.n2944 0.058
R5286 S.n2423 S.n2422 0.058
R5287 S.n2 S.n1 0.056
R5288 S.n693 S.n692 0.056
R5289 S.n496 S.n495 0.056
R5290 S.n527 S.n526 0.056
R5291 S.n565 S.n564 0.056
R5292 S.n584 S.n575 0.055
R5293 S.n4806 S.n4805 0.055
R5294 S.n4377 S.n4376 0.055
R5295 S.n3909 S.n3908 0.055
R5296 S.n3424 S.n3423 0.055
R5297 S.n2928 S.n2927 0.055
R5298 S.n2405 S.n2404 0.055
R5299 S.n1877 S.n1876 0.055
R5300 S.n1314 S.n1313 0.055
R5301 S.n441 S.n440 0.055
R5302 S.n5263 S.n5262 0.055
R5303 S.n5692 S.n5272 0.054
R5304 S.n5399 S.n5380 0.054
R5305 S.n3030 S.n3016 0.054
R5306 S.n3542 S.n3527 0.054
R5307 S.n4041 S.n4027 0.054
R5308 S.n4486 S.n4469 0.054
R5309 S.n4959 S.n4943 0.054
R5310 S.n1950 S.n1936 0.054
R5311 S.n2494 S.n2479 0.054
R5312 S.n777 S.n763 0.054
R5313 S.n1336 S.n1321 0.054
R5314 S.n130 S.n114 0.054
R5315 S.n905 S.n904 0.054
R5316 S.n1446 S.n1445 0.054
R5317 S.n2038 S.n2037 0.054
R5318 S.n2565 S.n2564 0.054
R5319 S.n3082 S.n3081 0.054
R5320 S.n3575 S.n3574 0.054
R5321 S.n4055 S.n4054 0.054
R5322 S.n249 S.n248 0.054
R5323 S.n5722 S.n5720 0.054
R5324 S.n492 S.n491 0.054
R5325 S.n4223 S.n4222 0.054
R5326 S.n4801 S.n4800 0.054
R5327 S.n5563 S.n5562 0.054
R5328 S.n5303 S.n5302 0.054
R5329 S.n5093 S.n5092 0.054
R5330 S.n5238 S.n5237 0.054
R5331 S.n4642 S.n4641 0.054
R5332 S.n5579 S.n5578 0.054
R5333 S.n5288 S.n5287 0.054
R5334 S.n5114 S.n5113 0.054
R5335 S.n5258 S.n5257 0.054
R5336 S.n4666 S.n4665 0.054
R5337 S.n3725 S.n3724 0.054
R5338 S.n3942 S.n3941 0.054
R5339 S.n5547 S.n5546 0.054
R5340 S.n5318 S.n5317 0.054
R5341 S.n5077 S.n5076 0.054
R5342 S.n5223 S.n5222 0.054
R5343 S.n4626 S.n4625 0.054
R5344 S.n4785 S.n4784 0.054
R5345 S.n4207 S.n4206 0.054
R5346 S.n3215 S.n3214 0.054
R5347 S.n3457 S.n3456 0.054
R5348 S.n5531 S.n5530 0.054
R5349 S.n5333 S.n5332 0.054
R5350 S.n5061 S.n5060 0.054
R5351 S.n5208 S.n5207 0.054
R5352 S.n4610 S.n4609 0.054
R5353 S.n4770 S.n4769 0.054
R5354 S.n4191 S.n4190 0.054
R5355 S.n3957 S.n3956 0.054
R5356 S.n3709 S.n3708 0.054
R5357 S.n2682 S.n2681 0.054
R5358 S.n2961 S.n2960 0.054
R5359 S.n5515 S.n5514 0.054
R5360 S.n5348 S.n5347 0.054
R5361 S.n5045 S.n5044 0.054
R5362 S.n5193 S.n5192 0.054
R5363 S.n4594 S.n4593 0.054
R5364 S.n4755 S.n4754 0.054
R5365 S.n4175 S.n4174 0.054
R5366 S.n3972 S.n3971 0.054
R5367 S.n3693 S.n3692 0.054
R5368 S.n3472 S.n3471 0.054
R5369 S.n3199 S.n3198 0.054
R5370 S.n2139 S.n2138 0.054
R5371 S.n2439 S.n2438 0.054
R5372 S.n5499 S.n5498 0.054
R5373 S.n5363 S.n5362 0.054
R5374 S.n5029 S.n5028 0.054
R5375 S.n5178 S.n5177 0.054
R5376 S.n4578 S.n4577 0.054
R5377 S.n4740 S.n4739 0.054
R5378 S.n4159 S.n4158 0.054
R5379 S.n3987 S.n3986 0.054
R5380 S.n3677 S.n3676 0.054
R5381 S.n3487 S.n3486 0.054
R5382 S.n3183 S.n3182 0.054
R5383 S.n2976 S.n2975 0.054
R5384 S.n2666 S.n2665 0.054
R5385 S.n1540 S.n1539 0.054
R5386 S.n1912 S.n1911 0.054
R5387 S.n5582 S.n5581 0.054
R5388 S.n5595 S.n5594 0.054
R5389 S.n5148 S.n5147 0.054
R5390 S.n5163 S.n5162 0.054
R5391 S.n4562 S.n4561 0.054
R5392 S.n4725 S.n4724 0.054
R5393 S.n4143 S.n4142 0.054
R5394 S.n4003 S.n4002 0.054
R5395 S.n3661 S.n3660 0.054
R5396 S.n3503 S.n3502 0.054
R5397 S.n3167 S.n3166 0.054
R5398 S.n2992 S.n2991 0.054
R5399 S.n2650 S.n2649 0.054
R5400 S.n2455 S.n2454 0.054
R5401 S.n2123 S.n2122 0.054
R5402 S.n977 S.n976 0.054
R5403 S.n1578 S.n1577 0.054
R5404 S.n5483 S.n5482 0.054
R5405 S.n5614 S.n5613 0.054
R5406 S.n5117 S.n5116 0.054
R5407 S.n5132 S.n5131 0.054
R5408 S.n4547 S.n4546 0.054
R5409 S.n4709 S.n4708 0.054
R5410 S.n4128 S.n4127 0.054
R5411 S.n4019 S.n4018 0.054
R5412 S.n3646 S.n3645 0.054
R5413 S.n3519 S.n3518 0.054
R5414 S.n3152 S.n3151 0.054
R5415 S.n3008 S.n3007 0.054
R5416 S.n2635 S.n2634 0.054
R5417 S.n2471 S.n2470 0.054
R5418 S.n2108 S.n2107 0.054
R5419 S.n1928 S.n1927 0.054
R5420 S.n1534 S.n1533 0.054
R5421 S.n404 S.n403 0.054
R5422 S.n1062 S.n1061 0.054
R5423 S.n5661 S.n5660 0.054
R5424 S.n4979 S.n4978 0.054
R5425 S.n4882 S.n4881 0.054
R5426 S.n4528 S.n4527 0.054
R5427 S.n4435 S.n4434 0.054
R5428 S.n4109 S.n4108 0.054
R5429 S.n4311 S.n4310 0.054
R5430 S.n3627 S.n3626 0.054
R5431 S.n3815 S.n3814 0.054
R5432 S.n3133 S.n3132 0.054
R5433 S.n3300 S.n3299 0.054
R5434 S.n2616 S.n2615 0.054
R5435 S.n2772 S.n2771 0.054
R5436 S.n2089 S.n2088 0.054
R5437 S.n2222 S.n2221 0.054
R5438 S.n1498 S.n1497 0.054
R5439 S.n1659 S.n1658 0.054
R5440 S.n957 S.n956 0.054
R5441 S.n367 S.n366 0.054
R5442 S.n299 S.n298 0.054
R5443 S.n5466 S.n5465 0.054
R5444 S.n5633 S.n5632 0.054
R5445 S.n5013 S.n5012 0.054
R5446 S.n4929 S.n4928 0.054
R5447 S.n4672 S.n4671 0.054
R5448 S.n4693 S.n4692 0.054
R5449 S.n4229 S.n4228 0.054
R5450 S.n4247 S.n4246 0.054
R5451 S.n3731 S.n3730 0.054
R5452 S.n3749 S.n3748 0.054
R5453 S.n3221 S.n3220 0.054
R5454 S.n3239 S.n3238 0.054
R5455 S.n2688 S.n2687 0.054
R5456 S.n2706 S.n2705 0.054
R5457 S.n2145 S.n2144 0.054
R5458 S.n2163 S.n2162 0.054
R5459 S.n1518 S.n1517 0.054
R5460 S.n1593 S.n1592 0.054
R5461 S.n983 S.n982 0.054
R5462 S.n1005 S.n1004 0.054
R5463 S.n106 S.n105 0.054
R5464 S.n1215 S.n1214 0.054
R5465 S.n3264 S.n3263 0.054
R5466 S.n2514 S.n2513 0.054
R5467 S.n2921 S.n2920 0.054
R5468 S.n1989 S.n1988 0.054
R5469 S.n2365 S.n2364 0.054
R5470 S.n1396 S.n1395 0.054
R5471 S.n1805 S.n1804 0.054
R5472 S.n852 S.n851 0.054
R5473 S.n472 S.n471 0.054
R5474 S.n3779 S.n3778 0.054
R5475 S.n3050 S.n3049 0.054
R5476 S.n3417 S.n3416 0.054
R5477 S.n2533 S.n2532 0.054
R5478 S.n2889 S.n2888 0.054
R5479 S.n2006 S.n2005 0.054
R5480 S.n2334 S.n2333 0.054
R5481 S.n1413 S.n1412 0.054
R5482 S.n1773 S.n1772 0.054
R5483 S.n871 S.n870 0.054
R5484 S.n893 S.n892 0.054
R5485 S.n1157 S.n1156 0.054
R5486 S.n305 S.n304 0.054
R5487 S.n328 S.n327 0.054
R5488 S.n1744 S.n1743 0.054
R5489 S.n2305 S.n2304 0.054
R5490 S.n2856 S.n2855 0.054
R5491 S.n3384 S.n3383 0.054
R5492 S.n3902 S.n3901 0.054
R5493 S.n4275 S.n4274 0.054
R5494 S.n3562 S.n3561 0.054
R5495 S.n3069 S.n3068 0.054
R5496 S.n2552 S.n2551 0.054
R5497 S.n2025 S.n2024 0.054
R5498 S.n1433 S.n1432 0.054
R5499 S.n1123 S.n1122 0.054
R5500 S.n257 S.n256 0.054
R5501 S.n653 S.n652 0.054
R5502 S.n4464 S.n4463 0.054
R5503 S.n4068 S.n4067 0.054
R5504 S.n4370 S.n4369 0.054
R5505 S.n3588 S.n3587 0.054
R5506 S.n3870 S.n3869 0.054
R5507 S.n3094 S.n3093 0.054
R5508 S.n3352 S.n3351 0.054
R5509 S.n2577 S.n2576 0.054
R5510 S.n2824 S.n2823 0.054
R5511 S.n2050 S.n2049 0.054
R5512 S.n2274 S.n2273 0.054
R5513 S.n1458 S.n1457 0.054
R5514 S.n1711 S.n1710 0.054
R5515 S.n917 S.n916 0.054
R5516 S.n1090 S.n1089 0.054
R5517 S.n276 S.n275 0.054
R5518 S.n938 S.n937 0.054
R5519 S.n1679 S.n1678 0.054
R5520 S.n1478 S.n1477 0.054
R5521 S.n2242 S.n2241 0.054
R5522 S.n2070 S.n2069 0.054
R5523 S.n2792 S.n2791 0.054
R5524 S.n2597 S.n2596 0.054
R5525 S.n3320 S.n3319 0.054
R5526 S.n3114 S.n3113 0.054
R5527 S.n3835 S.n3834 0.054
R5528 S.n3608 S.n3607 0.054
R5529 S.n4335 S.n4334 0.054
R5530 S.n4090 S.n4089 0.054
R5531 S.n4403 S.n4402 0.054
R5532 S.n4509 S.n4508 0.054
R5533 S.n4910 S.n4909 0.054
R5534 S.n354 S.n353 0.054
R5535 S.n1185 S.n1184 0.054
R5536 S.n233 S.n232 0.054
R5537 S.n216 S.n215 0.054
R5538 S.n74 S.n73 0.054
R5539 S.n1274 S.n1273 0.054
R5540 S.n2187 S.n2186 0.054
R5541 S.n1357 S.n1356 0.054
R5542 S.n1870 S.n1869 0.054
R5543 S.n816 S.n815 0.054
R5544 S.n513 S.n512 0.054
R5545 S.n2736 S.n2735 0.054
R5546 S.n1970 S.n1969 0.054
R5547 S.n2398 S.n2397 0.054
R5548 S.n1376 S.n1375 0.054
R5549 S.n1838 S.n1837 0.054
R5550 S.n833 S.n832 0.054
R5551 S.n1244 S.n1243 0.054
R5552 S.n198 S.n197 0.054
R5553 S.n181 S.n180 0.054
R5554 S.n42 S.n41 0.054
R5555 S.n1028 S.n1027 0.054
R5556 S.n551 S.n550 0.054
R5557 S.n1623 S.n1622 0.054
R5558 S.n797 S.n796 0.054
R5559 S.n1307 S.n1306 0.054
R5560 S.n163 S.n162 0.054
R5561 S.n147 S.n146 0.054
R5562 S.n435 S.n434 0.054
R5563 S.n5689 S.n5688 0.054
R5564 S.n4993 S.n4992 0.054
R5565 S.n699 S.n698 0.053
R5566 S.n5815 S.n5814 0.053
R5567 S.n5842 S.n5723 0.053
R5568 S.n5395 S.n5393 0.052
R5569 S.n125 S.n124 0.052
R5570 S.n772 S.n771 0.052
R5571 S.n1332 S.n1331 0.052
R5572 S.n1945 S.n1944 0.052
R5573 S.n2490 S.n2489 0.052
R5574 S.n3025 S.n3024 0.052
R5575 S.n3538 S.n3537 0.052
R5576 S.n4036 S.n4035 0.052
R5577 S.n4482 S.n4481 0.052
R5578 S.n4954 S.n4953 0.052
R5579 S.n1565 S.n1564 0.052
R5580 S.n757 S.n756 0.052
R5581 S.n396 S.n394 0.051
R5582 S.n4270 S.n4268 0.051
R5583 S.n3755 S.n3754 0.051
R5584 S.n3259 S.n3257 0.051
R5585 S.n2712 S.n2711 0.051
R5586 S.n2182 S.n2180 0.051
R5587 S.n1023 S.n1021 0.051
R5588 S.n1599 S.n1598 0.051
R5589 S.n415 S.n413 0.051
R5590 S.n5821 S.n5820 0.051
R5591 S.n5823 S.n5822 0.051
R5592 S.n446 S.n445 0.051
R5593 S.n5837 S.n5836 0.051
R5594 S.n5839 S.n5838 0.051
R5595 S.n448 S.n447 0.051
R5596 S.n900 S.n899 0.051
R5597 S.n1440 S.n1439 0.051
R5598 S.n2032 S.n2031 0.051
R5599 S.n2559 S.n2558 0.051
R5600 S.n3076 S.n3075 0.051
R5601 S.n3569 S.n3568 0.051
R5602 S.n4049 S.n4048 0.051
R5603 S.n252 S.n251 0.051
R5604 S.n4432 S.n4431 0.05
R5605 S.n4879 S.n4878 0.05
R5606 S.n5658 S.n5657 0.05
R5607 S.n3378 S.n3377 0.05
R5608 S.n3896 S.n3895 0.05
R5609 S.n4272 S.n4271 0.05
R5610 S.n4329 S.n4316 0.05
R5611 S.n4400 S.n4387 0.05
R5612 S.n4904 S.n4891 0.05
R5613 S.n345 S.n344 0.05
R5614 S.n3773 S.n3770 0.05
R5615 S.n3776 S.n3757 0.05
R5616 S.n3411 S.n3389 0.05
R5617 S.n2883 S.n2861 0.05
R5618 S.n2359 S.n2358 0.05
R5619 S.n2915 S.n2914 0.05
R5620 S.n3261 S.n3260 0.05
R5621 S.n2728 S.n2727 0.05
R5622 S.n2733 S.n2714 0.05
R5623 S.n2392 S.n2370 0.05
R5624 S.n1832 S.n1810 0.05
R5625 S.n1268 S.n1267 0.05
R5626 S.n1864 S.n1863 0.05
R5627 S.n2184 S.n2183 0.05
R5628 S.n1025 S.n1024 0.05
R5629 S.n1615 S.n1614 0.05
R5630 S.n1620 S.n1601 0.05
R5631 S.n1301 S.n1279 0.05
R5632 S.n432 S.n416 0.05
R5633 S.n312 S.n311 0.05
R5634 S.n5441 S.n5440 0.05
R5635 S.n4852 S.n4851 0.05
R5636 S.n379 S.n378 0.049
R5637 S.n290 S.n289 0.049
R5638 S.n906 S.n905 0.049
R5639 S.n1447 S.n1446 0.049
R5640 S.n2039 S.n2038 0.049
R5641 S.n2566 S.n2565 0.049
R5642 S.n3083 S.n3082 0.049
R5643 S.n3576 S.n3575 0.049
R5644 S.n4056 S.n4055 0.049
R5645 S.n250 S.n249 0.049
R5646 S.n270 S.n269 0.049
R5647 S.n5674 S.n5669 0.049
R5648 S.n4832 S.n4831 0.048
R5649 S.n753 S.n752 0.048
R5650 S.n5270 S.n4853 0.048
R5651 S.n1145 S.n1140 0.048
R5652 S.n3880 S.n3879 0.048
R5653 S.n3362 S.n3361 0.048
R5654 S.n2834 S.n2833 0.048
R5655 S.n2284 S.n2283 0.048
R5656 S.n1722 S.n1721 0.048
R5657 S.n4217 S.n4215 0.047
R5658 S.n4795 S.n4791 0.047
R5659 S.n5557 S.n5552 0.047
R5660 S.n5300 S.n5296 0.047
R5661 S.n5087 S.n5082 0.047
R5662 S.n5232 S.n5228 0.047
R5663 S.n4636 S.n4631 0.047
R5664 S.n4834 S.n4808 0.047
R5665 S.n5573 S.n5571 0.047
R5666 S.n5285 S.n5283 0.047
R5667 S.n5108 S.n5106 0.047
R5668 S.n5252 S.n5249 0.047
R5669 S.n4660 S.n4655 0.047
R5670 S.n4378 S.n4375 0.047
R5671 S.n3719 S.n3717 0.047
R5672 S.n3939 S.n3935 0.047
R5673 S.n5541 S.n5536 0.047
R5674 S.n5315 S.n5311 0.047
R5675 S.n5071 S.n5066 0.047
R5676 S.n5217 S.n5213 0.047
R5677 S.n4620 S.n4615 0.047
R5678 S.n4779 S.n4775 0.047
R5679 S.n4201 S.n4196 0.047
R5680 S.n3910 S.n3907 0.047
R5681 S.n3209 S.n3207 0.047
R5682 S.n3454 S.n3450 0.047
R5683 S.n5525 S.n5520 0.047
R5684 S.n5330 S.n5326 0.047
R5685 S.n5055 S.n5050 0.047
R5686 S.n5202 S.n5198 0.047
R5687 S.n4604 S.n4599 0.047
R5688 S.n4764 S.n4760 0.047
R5689 S.n4185 S.n4180 0.047
R5690 S.n3954 S.n3950 0.047
R5691 S.n3703 S.n3698 0.047
R5692 S.n3425 S.n3422 0.047
R5693 S.n2676 S.n2674 0.047
R5694 S.n2958 S.n2954 0.047
R5695 S.n5509 S.n5504 0.047
R5696 S.n5345 S.n5341 0.047
R5697 S.n5039 S.n5034 0.047
R5698 S.n5187 S.n5183 0.047
R5699 S.n4588 S.n4583 0.047
R5700 S.n4749 S.n4745 0.047
R5701 S.n4169 S.n4164 0.047
R5702 S.n3969 S.n3965 0.047
R5703 S.n3687 S.n3682 0.047
R5704 S.n3469 S.n3465 0.047
R5705 S.n3193 S.n3188 0.047
R5706 S.n2929 S.n2926 0.047
R5707 S.n2133 S.n2131 0.047
R5708 S.n2436 S.n2432 0.047
R5709 S.n5493 S.n5488 0.047
R5710 S.n5360 S.n5356 0.047
R5711 S.n5023 S.n5018 0.047
R5712 S.n5172 S.n5168 0.047
R5713 S.n4572 S.n4567 0.047
R5714 S.n4734 S.n4730 0.047
R5715 S.n4153 S.n4148 0.047
R5716 S.n3984 S.n3980 0.047
R5717 S.n3671 S.n3666 0.047
R5718 S.n3484 S.n3480 0.047
R5719 S.n3177 S.n3172 0.047
R5720 S.n2973 S.n2969 0.047
R5721 S.n2660 S.n2655 0.047
R5722 S.n2406 S.n2403 0.047
R5723 S.n1545 S.n1543 0.047
R5724 S.n1909 S.n1904 0.047
R5725 S.n5589 S.n5379 0.047
R5726 S.n5592 S.n5371 0.047
R5727 S.n5155 S.n5145 0.047
R5728 S.n5157 S.n5137 0.047
R5729 S.n4556 S.n4552 0.047
R5730 S.n4719 S.n4714 0.047
R5731 S.n4137 S.n4133 0.047
R5732 S.n4000 S.n3995 0.047
R5733 S.n3655 S.n3651 0.047
R5734 S.n3500 S.n3495 0.047
R5735 S.n3161 S.n3157 0.047
R5736 S.n2989 S.n2984 0.047
R5737 S.n2644 S.n2640 0.047
R5738 S.n2452 S.n2447 0.047
R5739 S.n2117 S.n2113 0.047
R5740 S.n1878 S.n1875 0.047
R5741 S.n971 S.n969 0.047
R5742 S.n1575 S.n1571 0.047
R5743 S.n5477 S.n5471 0.047
R5744 S.n5611 S.n5603 0.047
R5745 S.n5124 S.n4942 0.047
R5746 S.n5126 S.n4934 0.047
R5747 S.n4541 S.n4537 0.047
R5748 S.n4703 S.n4698 0.047
R5749 S.n4122 S.n4118 0.047
R5750 S.n4016 S.n4011 0.047
R5751 S.n3640 S.n3636 0.047
R5752 S.n3516 S.n3511 0.047
R5753 S.n3146 S.n3142 0.047
R5754 S.n3005 S.n3000 0.047
R5755 S.n2629 S.n2625 0.047
R5756 S.n2468 S.n2463 0.047
R5757 S.n2102 S.n2098 0.047
R5758 S.n1925 S.n1920 0.047
R5759 S.n1528 S.n1523 0.047
R5760 S.n1315 S.n1312 0.047
R5761 S.n401 S.n386 0.047
R5762 S.n1056 S.n1046 0.047
R5763 S.n5658 S.n5643 0.047
R5764 S.n4976 S.n4968 0.047
R5765 S.n4879 S.n4867 0.047
R5766 S.n4525 S.n4517 0.047
R5767 S.n4432 S.n4420 0.047
R5768 S.n4106 S.n4098 0.047
R5769 S.n4305 S.n4293 0.047
R5770 S.n3624 S.n3616 0.047
R5771 S.n3809 S.n3797 0.047
R5772 S.n3130 S.n3122 0.047
R5773 S.n3294 S.n3282 0.047
R5774 S.n2613 S.n2605 0.047
R5775 S.n2766 S.n2754 0.047
R5776 S.n2086 S.n2078 0.047
R5777 S.n2216 S.n2205 0.047
R5778 S.n1495 S.n1486 0.047
R5779 S.n1653 S.n1641 0.047
R5780 S.n954 S.n946 0.047
R5781 S.n377 S.n370 0.047
R5782 S.n293 S.n288 0.047
R5783 S.n463 S.n443 0.047
R5784 S.n5460 S.n5458 0.047
R5785 S.n5630 S.n5628 0.047
R5786 S.n5007 S.n5005 0.047
R5787 S.n4923 S.n4921 0.047
R5788 S.n4677 S.n4675 0.047
R5789 S.n4687 S.n4685 0.047
R5790 S.n4234 S.n4232 0.047
R5791 S.n4244 S.n4242 0.047
R5792 S.n3736 S.n3734 0.047
R5793 S.n3746 S.n3744 0.047
R5794 S.n3226 S.n3224 0.047
R5795 S.n3236 S.n3234 0.047
R5796 S.n2693 S.n2691 0.047
R5797 S.n2703 S.n2701 0.047
R5798 S.n2150 S.n2148 0.047
R5799 S.n2160 S.n2158 0.047
R5800 S.n1512 S.n1510 0.047
R5801 S.n1590 S.n1588 0.047
R5802 S.n988 S.n986 0.047
R5803 S.n1002 S.n996 0.047
R5804 S.n103 S.n101 0.047
R5805 S.n1209 S.n1199 0.047
R5806 S.n3261 S.n3247 0.047
R5807 S.n2511 S.n2503 0.047
R5808 S.n2915 S.n2903 0.047
R5809 S.n1986 S.n1978 0.047
R5810 S.n2359 S.n2348 0.047
R5811 S.n1393 S.n1384 0.047
R5812 S.n1799 S.n1787 0.047
R5813 S.n849 S.n841 0.047
R5814 S.n477 S.n475 0.047
R5815 S.n3776 S.n3767 0.047
R5816 S.n3047 S.n3045 0.047
R5817 S.n3411 S.n3400 0.047
R5818 S.n2530 S.n2528 0.047
R5819 S.n2883 S.n2872 0.047
R5820 S.n2003 S.n2001 0.047
R5821 S.n2328 S.n2317 0.047
R5822 S.n1410 S.n1408 0.047
R5823 S.n1767 S.n1756 0.047
R5824 S.n868 S.n864 0.047
R5825 S.n890 S.n885 0.047
R5826 S.n1151 S.n1136 0.047
R5827 S.n310 S.n308 0.047
R5828 S.n325 S.n319 0.047
R5829 S.n1738 S.n1726 0.047
R5830 S.n2299 S.n2288 0.047
R5831 S.n2850 S.n2838 0.047
R5832 S.n3378 S.n3366 0.047
R5833 S.n3896 S.n3884 0.047
R5834 S.n4272 S.n4258 0.047
R5835 S.n3559 S.n3551 0.047
R5836 S.n3066 S.n3058 0.047
R5837 S.n2549 S.n2541 0.047
R5838 S.n2022 S.n2014 0.047
R5839 S.n1430 S.n1421 0.047
R5840 S.n1117 S.n1108 0.047
R5841 S.n254 S.n244 0.047
R5842 S.n659 S.n656 0.047
R5843 S.n4458 S.n4450 0.047
R5844 S.n4065 S.n4059 0.047
R5845 S.n4364 S.n4346 0.047
R5846 S.n3585 S.n3579 0.047
R5847 S.n3864 S.n3846 0.047
R5848 S.n3091 S.n3086 0.047
R5849 S.n3346 S.n3331 0.047
R5850 S.n2574 S.n2569 0.047
R5851 S.n2818 S.n2803 0.047
R5852 S.n2047 S.n2042 0.047
R5853 S.n2268 S.n2253 0.047
R5854 S.n1455 S.n1450 0.047
R5855 S.n1705 S.n1690 0.047
R5856 S.n914 S.n909 0.047
R5857 S.n1084 S.n1074 0.047
R5858 S.n273 S.n268 0.047
R5859 S.n935 S.n929 0.047
R5860 S.n1673 S.n1671 0.047
R5861 S.n1475 S.n1470 0.047
R5862 S.n2236 S.n2234 0.047
R5863 S.n2067 S.n2062 0.047
R5864 S.n2786 S.n2784 0.047
R5865 S.n2594 S.n2589 0.047
R5866 S.n3314 S.n3312 0.047
R5867 S.n3111 S.n3106 0.047
R5868 S.n3829 S.n3827 0.047
R5869 S.n3605 S.n3600 0.047
R5870 S.n4329 S.n4327 0.047
R5871 S.n4087 S.n4082 0.047
R5872 S.n4400 S.n4398 0.047
R5873 S.n4506 S.n4501 0.047
R5874 S.n4904 S.n4902 0.047
R5875 S.n351 S.n343 0.047
R5876 S.n1179 S.n1169 0.047
R5877 S.n230 S.n228 0.047
R5878 S.n213 S.n211 0.047
R5879 S.n71 S.n69 0.047
R5880 S.n1268 S.n1258 0.047
R5881 S.n2184 S.n2171 0.047
R5882 S.n1354 S.n1345 0.047
R5883 S.n1864 S.n1852 0.047
R5884 S.n813 S.n805 0.047
R5885 S.n518 S.n516 0.047
R5886 S.n2733 S.n2724 0.047
R5887 S.n1967 S.n1965 0.047
R5888 S.n2392 S.n2381 0.047
R5889 S.n1373 S.n1371 0.047
R5890 S.n1832 S.n1821 0.047
R5891 S.n830 S.n828 0.047
R5892 S.n1238 S.n1227 0.047
R5893 S.n195 S.n193 0.047
R5894 S.n178 S.n176 0.047
R5895 S.n39 S.n37 0.047
R5896 S.n1025 S.n1013 0.047
R5897 S.n556 S.n554 0.047
R5898 S.n1620 S.n1611 0.047
R5899 S.n794 S.n792 0.047
R5900 S.n1301 S.n1290 0.047
R5901 S.n160 S.n158 0.047
R5902 S.n144 S.n142 0.047
R5903 S.n432 S.n425 0.047
R5904 S.n5270 S.n5265 0.047
R5905 S.n5683 S.n5681 0.047
R5906 S.n4990 S.n4988 0.047
R5907 S.n5416 S.n5412 0.047
R5908 S.n687 S.n686 0.046
R5909 S.t191 S.n628 0.046
R5910 S.t191 S.n618 0.046
R5911 S.t191 S.n606 0.046
R5912 S.t191 S.n594 0.046
R5913 S.n5251 S.n5250 0.046
R5914 S.n635 S.n633 0.045
R5915 S.n5833 S.n5832 0.045
R5916 S.n372 S.n371 0.045
R5917 S.n643 S.n642 0.045
R5918 S.n1099 S.n1091 0.045
R5919 S.n1702 S.n1694 0.045
R5920 S.n2265 S.n2257 0.045
R5921 S.n2815 S.n2807 0.045
R5922 S.n3343 S.n3335 0.045
R5923 S.n3852 S.n3851 0.045
R5924 S.n4352 S.n4351 0.045
R5925 S.n5818 S.n5817 0.045
R5926 S.n1264 S.n1263 0.045
R5927 S.n675 S.n674 0.044
R5928 S.n1909 S.n1908 0.044
R5929 S.n2452 S.n2451 0.044
R5930 S.n2989 S.n2988 0.044
R5931 S.n3500 S.n3499 0.044
R5932 S.n4000 S.n3999 0.044
R5933 S.n4719 S.n4718 0.044
R5934 S.n5157 S.n5156 0.044
R5935 S.n5592 S.n5591 0.044
R5936 S.n1925 S.n1924 0.044
R5937 S.n2468 S.n2467 0.044
R5938 S.n3005 S.n3004 0.044
R5939 S.n3516 S.n3515 0.044
R5940 S.n4016 S.n4015 0.044
R5941 S.n4703 S.n4702 0.044
R5942 S.n5126 S.n5125 0.044
R5943 S.n5816 S.n5815 0.044
R5944 S.n5725 S.n5724 0.044
R5945 S.n4687 S.n4678 0.043
R5946 S.n4244 S.n4235 0.043
R5947 S.n3746 S.n3737 0.043
R5948 S.n3236 S.n3227 0.043
R5949 S.n2703 S.n2694 0.043
R5950 S.n2160 S.n2151 0.043
R5951 S.n1002 S.n989 0.043
R5952 S.n122 S.n121 0.043
R5953 S.n5657 S.n5656 0.043
R5954 S.n322 S.n321 0.043
R5955 S.n4316 S.n4315 0.043
R5956 S.n4387 S.n4386 0.043
R5957 S.n4891 S.n4890 0.043
R5958 S.n3389 S.n3386 0.043
R5959 S.n2861 S.n2858 0.043
R5960 S.n93 S.n92 0.043
R5961 S.n2370 S.n2367 0.043
R5962 S.n1810 S.n1807 0.043
R5963 S.n1279 S.n1276 0.043
R5964 S.n4875 S.n4872 0.043
R5965 S.n4428 S.n4425 0.043
R5966 S.n2911 S.n2908 0.043
R5967 S.n2355 S.n2353 0.043
R5968 S.n3892 S.n3889 0.043
R5969 S.n3374 S.n3371 0.043
R5970 S.n1860 S.n1857 0.043
R5971 S.n570 S.n569 0.043
R5972 S.n691 S.n690 0.043
R5973 S.n1350 S.n1349 0.042
R5974 S.n1162 S.n1161 0.042
R5975 S.n1748 S.n1747 0.042
R5976 S.n2309 S.n2308 0.042
R5977 S.n1220 S.n1219 0.042
R5978 S.n428 S.n427 0.042
R5979 S.n4301 S.n4298 0.042
R5980 S.n3805 S.n3802 0.042
R5981 S.n3290 S.n3287 0.042
R5982 S.n2762 S.n2759 0.042
R5983 S.n2212 S.n2210 0.042
R5984 S.n1491 S.n1490 0.042
R5985 S.n1649 S.n1646 0.042
R5986 S.n1389 S.n1388 0.042
R5987 S.n1795 S.n1792 0.042
R5988 S.n2846 S.n2843 0.042
R5989 S.n2295 S.n2293 0.042
R5990 S.n1426 S.n1425 0.042
R5991 S.n1734 S.n1731 0.042
R5992 S.n479 S.n478 0.042
R5993 S.n661 S.n660 0.042
R5994 S.n520 S.n519 0.042
R5995 S.n558 S.n557 0.042
R5996 S.n3819 S.n3818 0.042
R5997 S.n3304 S.n3303 0.042
R5998 S.n2776 S.n2775 0.042
R5999 S.n2226 S.n2225 0.042
R6000 S.n1663 S.n1662 0.042
R6001 S.n1066 S.n1065 0.042
R6002 S.n4255 S.n4254 0.041
R6003 S.n695 S.n694 0.041
R6004 S.n4 S.n3 0.041
R6005 S.n498 S.n497 0.041
R6006 S.n529 S.n528 0.041
R6007 S.n567 S.n566 0.041
R6008 S.n582 S.n580 0.041
R6009 S.n439 S.n438 0.041
R6010 S.n678 S.n677 0.04
R6011 S.n503 S.n502 0.04
R6012 S.n125 S.n116 0.04
R6013 S.n772 S.n765 0.04
R6014 S.n1332 S.n1325 0.04
R6015 S.n1945 S.n1938 0.04
R6016 S.n2490 S.n2483 0.04
R6017 S.n3025 S.n3018 0.04
R6018 S.n3538 S.n3531 0.04
R6019 S.n4036 S.n4029 0.04
R6020 S.n4482 S.n4475 0.04
R6021 S.n4954 S.n4947 0.04
R6022 S.n5395 S.n5394 0.04
R6023 S.n579 S.n578 0.039
R6024 S.n124 S.n117 0.039
R6025 S.n771 S.n766 0.039
R6026 S.n1331 S.n1326 0.039
R6027 S.n1944 S.n1939 0.039
R6028 S.n2489 S.n2484 0.039
R6029 S.n3024 S.n3019 0.039
R6030 S.n3537 S.n3532 0.039
R6031 S.n4035 S.n4030 0.039
R6032 S.n4481 S.n4476 0.039
R6033 S.n4953 S.n4948 0.039
R6034 S.n5393 S.n5392 0.039
R6035 S.n5814 S.n5801 0.039
R6036 S.n5804 S.n5803 0.039
R6037 S.n5384 S.n5382 0.038
R6038 S.n4074 S.n4072 0.038
R6039 S.n4493 S.n4491 0.038
R6040 S.n4946 S.n4944 0.038
R6041 S.n3037 S.n3036 0.038
R6042 S.n2520 S.n2519 0.038
R6043 S.n1957 S.n1956 0.038
R6044 S.n1363 S.n1362 0.038
R6045 S.n784 S.n783 0.038
R6046 S.n4863 S.n4862 0.038
R6047 S.n4416 S.n4415 0.038
R6048 S.n4289 S.n4288 0.038
R6049 S.n3793 S.n3792 0.038
R6050 S.n3278 S.n3277 0.038
R6051 S.n2750 S.n2749 0.038
R6052 S.n2201 S.n2200 0.038
R6053 S.n1637 S.n1636 0.038
R6054 S.n1042 S.n1041 0.038
R6055 S.n2899 S.n2898 0.038
R6056 S.n2344 S.n2343 0.038
R6057 S.n1783 S.n1782 0.038
R6058 S.n1195 S.n1194 0.038
R6059 S.n3409 S.n3404 0.038
R6060 S.n2881 S.n2876 0.038
R6061 S.n2326 S.n2321 0.038
R6062 S.n1765 S.n1760 0.038
R6063 S.n1177 S.n1173 0.038
R6064 S.n1848 S.n1847 0.038
R6065 S.n1254 S.n1253 0.038
R6066 S.n2390 S.n2385 0.038
R6067 S.n1830 S.n1825 0.038
R6068 S.n1236 S.n1231 0.038
R6069 S.n1299 S.n1294 0.038
R6070 S.n1705 S.n1687 0.038
R6071 S.n2268 S.n2250 0.038
R6072 S.n2818 S.n2800 0.038
R6073 S.n3346 S.n3328 0.038
R6074 S.n3864 S.n3843 0.038
R6075 S.n4364 S.n4343 0.038
R6076 S.n4458 S.n4447 0.038
R6077 S.n1117 S.n1112 0.038
R6078 S.n4457 S.n4455 0.037
R6079 S.n1084 S.n1076 0.037
R6080 S.n1879 S.n1546 0.037
R6081 S.n5276 S.n5275 0.037
R6082 S.n5242 S.n5241 0.037
R6083 S.n729 S.n728 0.036
R6084 S.n463 S.n439 0.036
R6085 S.n934 S.n933 0.036
R6086 S.n1463 S.n1462 0.036
R6087 S.n2055 S.n2054 0.036
R6088 S.n2582 S.n2581 0.036
R6089 S.n3099 S.n3098 0.036
R6090 S.n3593 S.n3592 0.036
R6091 S.n5674 S.n5673 0.036
R6092 S.n1994 S.n1993 0.035
R6093 S.n1401 S.n1400 0.035
R6094 S.n857 S.n856 0.035
R6095 S.n821 S.n820 0.035
R6096 S.n5752 S.n5751 0.035
R6097 S.n5743 S.n5742 0.035
R6098 S.n5638 S.n5637 0.035
R6099 S.n5403 S.n5402 0.035
R6100 S.n3034 S.n3033 0.035
R6101 S.n3546 S.n3545 0.035
R6102 S.n4045 S.n4044 0.035
R6103 S.n4490 S.n4489 0.035
R6104 S.n4963 S.n4962 0.035
R6105 S.n1954 S.n1953 0.035
R6106 S.n2498 S.n2497 0.035
R6107 S.n781 S.n780 0.035
R6108 S.n1340 S.n1339 0.035
R6109 S.n134 S.n133 0.035
R6110 S.n4863 S.n4858 0.035
R6111 S.n4416 S.n4411 0.035
R6112 S.n4289 S.n4284 0.035
R6113 S.n3793 S.n3788 0.035
R6114 S.n3278 S.n3273 0.035
R6115 S.n2750 S.n2745 0.035
R6116 S.n2201 S.n2196 0.035
R6117 S.n1637 S.n1632 0.035
R6118 S.n1042 S.n1037 0.035
R6119 S.n2899 S.n2894 0.035
R6120 S.n2344 S.n2339 0.035
R6121 S.n1783 S.n1778 0.035
R6122 S.n1195 S.n1190 0.035
R6123 S.n4272 S.n4255 0.035
R6124 S.n4361 S.n4360 0.035
R6125 S.n3861 S.n3860 0.035
R6126 S.n1177 S.n1176 0.035
R6127 S.n1765 S.n1764 0.035
R6128 S.n2326 S.n2325 0.035
R6129 S.n2881 S.n2880 0.035
R6130 S.n3409 S.n3408 0.035
R6131 S.n1848 S.n1843 0.035
R6132 S.n1254 S.n1249 0.035
R6133 S.n1236 S.n1235 0.035
R6134 S.n1830 S.n1829 0.035
R6135 S.n2390 S.n2389 0.035
R6136 S.n1299 S.n1298 0.035
R6137 S.t240 S.n5789 0.035
R6138 S.t240 S.n5796 0.035
R6139 S.t240 S.n5782 0.035
R6140 S.t240 S.n5775 0.035
R6141 S.t240 S.n5768 0.035
R6142 S.t240 S.n5761 0.035
R6143 S.t240 S.n5754 0.035
R6144 S.t240 S.n5745 0.035
R6145 S.t240 S.n5734 0.035
R6146 S.t240 S.n5736 0.035
R6147 S.t191 S.n616 0.035
R6148 S.t191 S.n714 0.035
R6149 S.t191 S.n630 0.035
R6150 S.t191 S.n641 0.035
R6151 S.t191 S.n689 0.035
R6152 S.t191 S.n604 0.035
R6153 S.t191 S.n710 0.035
R6154 S.t191 S.n591 0.035
R6155 S.t191 S.n706 0.035
R6156 S.t191 S.n702 0.035
R6157 S.t240 S.n5827 0.035
R6158 S.n5728 S.n5727 0.035
R6159 S.n627 S.n623 0.034
R6160 S.n620 S.n619 0.034
R6161 S.n608 S.n607 0.034
R6162 S.n596 S.n595 0.034
R6163 S.n1878 S.n1566 0.034
R6164 S.n1315 S.n758 0.034
R6165 S.n397 S.n396 0.034
R6166 S.n4038 S.n4028 0.034
R6167 S.n3540 S.n3530 0.034
R6168 S.n3027 S.n3017 0.034
R6169 S.n2492 S.n2482 0.034
R6170 S.n1947 S.n1937 0.034
R6171 S.n774 S.n764 0.034
R6172 S.n1334 S.n1324 0.034
R6173 S.n127 S.n115 0.034
R6174 S.t240 S.n5792 0.034
R6175 S.t240 S.n5799 0.034
R6176 S.t240 S.n5785 0.034
R6177 S.t240 S.n5778 0.034
R6178 S.t240 S.n5771 0.034
R6179 S.t240 S.n5764 0.034
R6180 S.t240 S.n5757 0.034
R6181 S.t240 S.n5748 0.034
R6182 S.t240 S.n5731 0.034
R6183 S.t240 S.n5739 0.034
R6184 S.t191 S.n615 0.034
R6185 S.t191 S.n717 0.034
R6186 S.t191 S.n629 0.034
R6187 S.t191 S.n640 0.034
R6188 S.t191 S.n688 0.034
R6189 S.t191 S.n603 0.034
R6190 S.t191 S.n713 0.034
R6191 S.t191 S.n590 0.034
R6192 S.t191 S.n709 0.034
R6193 S.t191 S.n705 0.034
R6194 S.t240 S.n5830 0.034
R6195 S.n889 S.n888 0.033
R6196 S.n5415 S.n5414 0.033
R6197 S.n582 S.n581 0.032
R6198 S.n5397 S.n5384 0.032
R6199 S.n4075 S.n4074 0.032
R6200 S.n4494 S.n4493 0.032
R6201 S.n4956 S.n4946 0.032
R6202 S.n1018 S.n1017 0.031
R6203 S.n3038 S.n3037 0.031
R6204 S.n2521 S.n2520 0.031
R6205 S.n1958 S.n1957 0.031
R6206 S.n1364 S.n1363 0.031
R6207 S.n785 S.n784 0.031
R6208 S.t34 S.n5638 0.031
R6209 S.t52 S.n5403 0.031
R6210 S.t27 S.n3034 0.031
R6211 S.t6 S.n3546 0.031
R6212 S.t65 S.n4045 0.031
R6213 S.t4 S.n4490 0.031
R6214 S.t45 S.n4963 0.031
R6215 S.t56 S.n1954 0.031
R6216 S.t68 S.n2498 0.031
R6217 S.t14 S.n781 0.031
R6218 S.t32 S.n1340 0.031
R6219 S.t213 S.n134 0.031
R6220 S.n4858 S.n4857 0.031
R6221 S.n4411 S.n4410 0.031
R6222 S.n4284 S.n4283 0.031
R6223 S.n3788 S.n3787 0.031
R6224 S.n3273 S.n3272 0.031
R6225 S.n2745 S.n2744 0.031
R6226 S.n2196 S.n2195 0.031
R6227 S.n1632 S.n1631 0.031
R6228 S.n1037 S.n1036 0.031
R6229 S.n437 S.n436 0.031
R6230 S.n2894 S.n2893 0.031
R6231 S.n2339 S.n2338 0.031
R6232 S.n1778 S.n1777 0.031
R6233 S.n1190 S.n1189 0.031
R6234 S.n1176 S.n1175 0.031
R6235 S.n1764 S.n1763 0.031
R6236 S.n2325 S.n2324 0.031
R6237 S.n2880 S.n2879 0.031
R6238 S.n3408 S.n3407 0.031
R6239 S.n1843 S.n1842 0.031
R6240 S.n1249 S.n1248 0.031
R6241 S.n1235 S.n1234 0.031
R6242 S.n1829 S.n1828 0.031
R6243 S.n2389 S.n2388 0.031
R6244 S.n1298 S.n1297 0.031
R6245 S.n5442 S.n5426 0.031
R6246 S.n5855 S.n5854 0.031
R6247 S.n5854 S.n5853 0.031
R6248 S.n5853 S.n5852 0.031
R6249 S.n5852 S.n5851 0.031
R6250 S.n5851 S.n5850 0.031
R6251 S.n5850 S.n5849 0.031
R6252 S.n5849 S.n5848 0.031
R6253 S.n5848 S.n5847 0.031
R6254 S.n5847 S.n5846 0.031
R6255 S.n5846 S.n5845 0.031
R6256 S.n733 S.n732 0.031
R6257 S.n734 S.n733 0.031
R6258 S.n735 S.n734 0.031
R6259 S.n736 S.n735 0.031
R6260 S.n737 S.n736 0.031
R6261 S.n738 S.n737 0.031
R6262 S.n739 S.n738 0.031
R6263 S.n5426 S.n5425 0.031
R6264 S.n2731 S.n2730 0.031
R6265 S.n1618 S.n1617 0.031
R6266 S.n3759 S.n3758 0.03
R6267 S.n2716 S.n2715 0.03
R6268 S.n1603 S.n1602 0.03
R6269 S.n4356 S.n4355 0.03
R6270 S.n3856 S.n3855 0.03
R6271 S.n3340 S.n3339 0.03
R6272 S.n2812 S.n2811 0.03
R6273 S.n2262 S.n2261 0.03
R6274 S.n1699 S.n1698 0.03
R6275 S.n1096 S.n1095 0.03
R6276 S.n669 S.n668 0.03
R6277 S.n730 S.n727 0.029
R6278 S.n3254 S.n3251 0.029
R6279 S.n4265 S.n4262 0.029
R6280 S.n2177 S.n2175 0.029
R6281 S.n1649 S.n1648 0.029
R6282 S.n2212 S.n2211 0.029
R6283 S.n2762 S.n2761 0.029
R6284 S.n3290 S.n3289 0.029
R6285 S.n3805 S.n3804 0.029
R6286 S.n4301 S.n4300 0.029
R6287 S.n1734 S.n1733 0.029
R6288 S.n2295 S.n2294 0.029
R6289 S.n2846 S.n2845 0.029
R6290 S.n1795 S.n1794 0.029
R6291 S.n3339 S.n3338 0.029
R6292 S.n2811 S.n2810 0.029
R6293 S.n2261 S.n2260 0.029
R6294 S.n1698 S.n1697 0.029
R6295 S.n1095 S.n1094 0.029
R6296 S.n668 S.n667 0.029
R6297 S.n4788 S.n4787 0.029
R6298 S.n3881 S.n3880 0.028
R6299 S.n3363 S.n3362 0.028
R6300 S.n2835 S.n2834 0.028
R6301 S.n2285 S.n2284 0.028
R6302 S.n4858 S.n4855 0.028
R6303 S.n4411 S.n4408 0.028
R6304 S.n4284 S.n4281 0.028
R6305 S.n3788 S.n3785 0.028
R6306 S.n3273 S.n3270 0.028
R6307 S.n2745 S.n2742 0.028
R6308 S.n2196 S.n2193 0.028
R6309 S.n1632 S.n1629 0.028
R6310 S.n1037 S.n1034 0.028
R6311 S.n2894 S.n2891 0.028
R6312 S.n2339 S.n2336 0.028
R6313 S.n1778 S.n1775 0.028
R6314 S.n1190 S.n1187 0.028
R6315 S.n1764 S.n1761 0.028
R6316 S.n2325 S.n2322 0.028
R6317 S.n2880 S.n2877 0.028
R6318 S.n3408 S.n3405 0.028
R6319 S.n1843 S.n1840 0.028
R6320 S.n1249 S.n1246 0.028
R6321 S.n1235 S.n1232 0.028
R6322 S.n1829 S.n1826 0.028
R6323 S.n2389 S.n2386 0.028
R6324 S.n1298 S.n1295 0.028
R6325 S.n998 S.n997 0.028
R6326 S.n1000 S.n998 0.028
R6327 S.n1111 S.n1110 0.028
R6328 S.n904 S.n903 0.028
R6329 S.n1686 S.n1685 0.028
R6330 S.n1445 S.n1444 0.028
R6331 S.n2249 S.n2248 0.028
R6332 S.n2037 S.n2036 0.028
R6333 S.n2799 S.n2798 0.028
R6334 S.n2564 S.n2563 0.028
R6335 S.n3327 S.n3326 0.028
R6336 S.n3081 S.n3080 0.028
R6337 S.n3842 S.n3841 0.028
R6338 S.n3574 S.n3573 0.028
R6339 S.n4342 S.n4341 0.028
R6340 S.n4054 S.n4053 0.028
R6341 S.n4446 S.n4445 0.028
R6342 S.n248 S.n247 0.028
R6343 S.n1078 S.n1077 0.028
R6344 S.n1080 S.n1078 0.028
R6345 S.n4428 S.n4427 0.028
R6346 S.n4875 S.n4874 0.028
R6347 S.n5651 S.n5650 0.028
R6348 S.n3374 S.n3373 0.028
R6349 S.n3892 S.n3891 0.028
R6350 S.n4265 S.n4264 0.028
R6351 S.n2355 S.n2354 0.028
R6352 S.n2911 S.n2910 0.028
R6353 S.n3254 S.n3253 0.028
R6354 S.n1860 S.n1859 0.028
R6355 S.n2177 S.n2176 0.028
R6356 S.n903 S.n902 0.028
R6357 S.n1444 S.n1443 0.028
R6358 S.n2036 S.n2035 0.028
R6359 S.n2563 S.n2562 0.028
R6360 S.n3080 S.n3079 0.028
R6361 S.n3573 S.n3572 0.028
R6362 S.n4053 S.n4052 0.028
R6363 S.n247 S.n246 0.028
R6364 S.n5276 S.n5274 0.027
R6365 S.n5242 S.n5240 0.027
R6366 S.n5591 S.n5590 0.027
R6367 S.n5476 S.n5475 0.027
R6368 S.n5451 S.n5450 0.027
R6369 S.n1723 S.n1722 0.027
R6370 S.n1315 S.n741 0.027
R6371 S.n347 S.n346 0.027
R6372 S.n3772 S.n3771 0.027
R6373 S.n2730 S.n2729 0.027
R6374 S.n1617 S.n1616 0.027
R6375 S.n5270 S.n5269 0.027
R6376 S.n866 S.n865 0.027
R6377 S.n4834 S.n4380 0.026
R6378 S.n4378 S.n3930 0.026
R6379 S.n3910 S.n3445 0.026
R6380 S.n3425 S.n2949 0.026
R6381 S.n2929 S.n2427 0.026
R6382 S.n2406 S.n1899 0.026
R6383 S.n1056 S.n1051 0.026
R6384 S.n954 S.n951 0.026
R6385 S.n1653 S.n1650 0.026
R6386 S.n1495 S.n1492 0.026
R6387 S.n2216 S.n2213 0.026
R6388 S.n2086 S.n2083 0.026
R6389 S.n2766 S.n2763 0.026
R6390 S.n2613 S.n2610 0.026
R6391 S.n3294 S.n3291 0.026
R6392 S.n3130 S.n3127 0.026
R6393 S.n3809 S.n3806 0.026
R6394 S.n3624 S.n3621 0.026
R6395 S.n4305 S.n4302 0.026
R6396 S.n4106 S.n4103 0.026
R6397 S.n4432 S.n4429 0.026
R6398 S.n4525 S.n4522 0.026
R6399 S.n4879 S.n4876 0.026
R6400 S.n4976 S.n4973 0.026
R6401 S.n5658 S.n5652 0.026
R6402 S.n1151 S.n1129 0.026
R6403 S.n890 S.n878 0.026
R6404 S.n1738 S.n1735 0.026
R6405 S.n1430 S.n1427 0.026
R6406 S.n2299 S.n2296 0.026
R6407 S.n2022 S.n2019 0.026
R6408 S.n2850 S.n2847 0.026
R6409 S.n2549 S.n2546 0.026
R6410 S.n3378 S.n3375 0.026
R6411 S.n3066 S.n3063 0.026
R6412 S.n3896 S.n3893 0.026
R6413 S.n3559 S.n3556 0.026
R6414 S.n4272 S.n4266 0.026
R6415 S.n901 S.n898 0.026
R6416 S.n1441 S.n1438 0.026
R6417 S.n2033 S.n2030 0.026
R6418 S.n2560 S.n2557 0.026
R6419 S.n3077 S.n3074 0.026
R6420 S.n3570 S.n3567 0.026
R6421 S.n4050 S.n4047 0.026
R6422 S.n4505 S.n4504 0.026
R6423 S.n4086 S.n4085 0.026
R6424 S.n3604 S.n3603 0.026
R6425 S.n3110 S.n3109 0.026
R6426 S.n2593 S.n2592 0.026
R6427 S.n2066 S.n2065 0.026
R6428 S.n1474 S.n1473 0.026
R6429 S.n924 S.n923 0.026
R6430 S.n1084 S.n1067 0.026
R6431 S.n1673 S.n1664 0.026
R6432 S.n2236 S.n2227 0.026
R6433 S.n2786 S.n2777 0.026
R6434 S.n3314 S.n3305 0.026
R6435 S.n3829 S.n3820 0.026
R6436 S.n4329 S.n4320 0.026
R6437 S.n4400 S.n4391 0.026
R6438 S.n4904 S.n4895 0.026
R6439 S.n351 S.n337 0.026
R6440 S.n3776 S.n3760 0.026
R6441 S.n3411 S.n3393 0.026
R6442 S.n2883 S.n2865 0.026
R6443 S.n2328 S.n2310 0.026
R6444 S.n1767 S.n1749 0.026
R6445 S.n1179 S.n1163 0.026
R6446 S.n477 S.n10 0.026
R6447 S.n1209 S.n1204 0.026
R6448 S.n849 S.n846 0.026
R6449 S.n1799 S.n1796 0.026
R6450 S.n1393 S.n1390 0.026
R6451 S.n2359 S.n2356 0.026
R6452 S.n1986 S.n1983 0.026
R6453 S.n2915 S.n2912 0.026
R6454 S.n2511 S.n2508 0.026
R6455 S.n3261 S.n3255 0.026
R6456 S.n2733 S.n2717 0.026
R6457 S.n2392 S.n2374 0.026
R6458 S.n1832 S.n1814 0.026
R6459 S.n1238 S.n1221 0.026
R6460 S.n518 S.n504 0.026
R6461 S.n1268 S.n1265 0.026
R6462 S.n813 S.n810 0.026
R6463 S.n1864 S.n1861 0.026
R6464 S.n1354 S.n1351 0.026
R6465 S.n2184 S.n2178 0.026
R6466 S.n1025 S.n1019 0.026
R6467 S.n1620 S.n1604 0.026
R6468 S.n1301 S.n1283 0.026
R6469 S.n556 S.n542 0.026
R6470 S.n432 S.n419 0.026
R6471 S.n432 S.n429 0.026
R6472 S.n5434 S.n5433 0.026
R6473 S.n418 S.n417 0.026
R6474 S.n325 S.n324 0.026
R6475 S.n389 S.n388 0.026
R6476 S.n5669 S.n5668 0.025
R6477 S.n3880 S.n3875 0.025
R6478 S.n3362 S.n3357 0.025
R6479 S.n2834 S.n2829 0.025
R6480 S.n2284 S.n2279 0.025
R6481 S.n1722 S.n1717 0.025
R6482 S.n1705 S.n1683 0.025
R6483 S.n2268 S.n2246 0.025
R6484 S.n2818 S.n2796 0.025
R6485 S.n3346 S.n3324 0.025
R6486 S.n3864 S.n3839 0.025
R6487 S.n4364 S.n4339 0.025
R6488 S.n4458 S.n4443 0.025
R6489 S.n1117 S.n1116 0.025
R6490 S.n1145 S.n1144 0.025
R6491 S.n3930 S.n3929 0.025
R6492 S.n3445 S.n3444 0.025
R6493 S.n2949 S.n2948 0.025
R6494 S.n2427 S.n2426 0.025
R6495 S.n1899 S.n1898 0.025
R6496 S.t191 S.n4 0.025
R6497 S.t191 S.n695 0.025
R6498 S.t191 S.n498 0.025
R6499 S.t191 S.n529 0.025
R6500 S.t191 S.n567 0.025
R6501 S.n4380 S.n4379 0.024
R6502 S.n457 S.n454 0.024
R6503 S.n123 S.n119 0.024
R6504 S.n748 S.n745 0.024
R6505 S.n770 S.n768 0.024
R6506 S.n1557 S.n1554 0.024
R6507 S.n1330 S.n1328 0.024
R6508 S.n1890 S.n1887 0.024
R6509 S.n1943 S.n1941 0.024
R6510 S.n2418 S.n2415 0.024
R6511 S.n2488 S.n2486 0.024
R6512 S.n2940 S.n2937 0.024
R6513 S.n3023 S.n3021 0.024
R6514 S.n3436 S.n3433 0.024
R6515 S.n3536 S.n3534 0.024
R6516 S.n3921 S.n3918 0.024
R6517 S.n4034 S.n4032 0.024
R6518 S.n4827 S.n4824 0.024
R6519 S.n4480 S.n4478 0.024
R6520 S.n4845 S.n4842 0.024
R6521 S.n4952 S.n4950 0.024
R6522 S.n5699 S.n5696 0.024
R6523 S.n5391 S.n5386 0.024
R6524 S.n5714 S.n5712 0.024
R6525 S.n5269 S.n5268 0.024
R6526 S.n5719 S.n5718 0.024
R6527 S.n741 S.n740 0.024
R6528 S.n1084 S.n1083 0.024
R6529 S.n19 S.n18 0.024
R6530 S.n5841 S.n5833 0.023
R6531 S.n3928 S.n3927 0.023
R6532 S.n4813 S.n4811 0.023
R6533 S.n4659 S.n4658 0.023
R6534 S.n4382 S.n4381 0.023
R6535 S.n3443 S.n3442 0.023
R6536 S.n2947 S.n2946 0.023
R6537 S.n2425 S.n2424 0.023
R6538 S.n1897 S.n1896 0.023
R6539 S.n1565 S.n1563 0.023
R6540 S.n757 S.n755 0.023
R6541 S.n754 S.n753 0.023
R6542 S.n375 S.n372 0.023
R6543 S.n1002 S.n1000 0.023
R6544 S.n93 S.n91 0.023
R6545 S.n323 S.n320 0.023
R6546 S.n1116 S.n1115 0.023
R6547 S.n681 S.n679 0.023
R6548 S.t191 S.n682 0.023
R6549 S.n4471 S.n4470 0.023
R6550 S.n4443 S.n4442 0.023
R6551 S.n4339 S.n4338 0.023
R6552 S.n3839 S.n3838 0.023
R6553 S.n3324 S.n3323 0.023
R6554 S.n2796 S.n2795 0.023
R6555 S.n2246 S.n2245 0.023
R6556 S.n1683 S.n1682 0.023
R6557 S.n681 S.n680 0.023
R6558 S.n682 S.n681 0.023
R6559 S.n250 S.n245 0.023
R6560 S.n1083 S.n1082 0.023
R6561 S.n348 S.n347 0.023
R6562 S.n1084 S.n1080 0.023
R6563 S.n1117 S.n1113 0.023
R6564 S.n3773 S.n3772 0.023
R6565 S.n94 S.n89 0.023
R6566 S.n61 S.n60 0.023
R6567 S.n58 S.n57 0.023
R6568 S.n62 S.n58 0.023
R6569 S.n29 S.n28 0.023
R6570 S.n26 S.n25 0.023
R6571 S.n537 S.n534 0.023
R6572 S.n30 S.n26 0.023
R6573 S.n5826 S.n5818 0.023
R6574 S.n5267 S.n5266 0.023
R6575 S.n1150 S.n1149 0.023
R6576 S.n2864 S.n2863 0.022
R6577 S.n3392 S.n3391 0.022
R6578 S.n1813 S.n1812 0.022
R6579 S.n2373 S.n2372 0.022
R6580 S.n1282 S.n1281 0.022
R6581 S.n3875 S.n3873 0.022
R6582 S.n3357 S.n3355 0.022
R6583 S.n2829 S.n2827 0.022
R6584 S.n2279 S.n2277 0.022
R6585 S.n1717 S.n1715 0.022
R6586 S.n1144 S.n1142 0.022
R6587 S.n5656 S.n5655 0.022
R6588 S.n1149 S.n1148 0.022
R6589 S.n4357 S.n4354 0.022
R6590 S.n3857 S.n3854 0.022
R6591 S.n3341 S.n3337 0.022
R6592 S.n2813 S.n2809 0.022
R6593 S.n2263 S.n2259 0.022
R6594 S.n1700 S.n1696 0.022
R6595 S.n1097 S.n1093 0.022
R6596 S.n670 S.n666 0.022
R6597 S.n4315 S.n4314 0.022
R6598 S.n4386 S.n4385 0.022
R6599 S.n4890 S.n4889 0.022
R6600 S.n3386 S.n3385 0.022
R6601 S.n2858 S.n2857 0.022
R6602 S.n85 S.n84 0.022
R6603 S.n2367 S.n2366 0.022
R6604 S.n1807 S.n1806 0.022
R6605 S.n53 S.n52 0.022
R6606 S.n1276 S.n1275 0.022
R6607 S.n21 S.n20 0.022
R6608 S.n4270 S.n4269 0.022
R6609 S.n3755 S.n3753 0.022
R6610 S.n3259 S.n3258 0.022
R6611 S.n2712 S.n2710 0.022
R6612 S.n2182 S.n2181 0.022
R6613 S.n1023 S.n1022 0.022
R6614 S.n1599 S.n1597 0.022
R6615 S.n415 S.n414 0.022
R6616 S.n4894 S.n4893 0.022
R6617 S.n4390 S.n4389 0.022
R6618 S.n4319 S.n4318 0.022
R6619 S.n5651 S.n5648 0.021
R6620 S.n5416 S.n5415 0.021
R6621 S.n1054 S.n1053 0.021
R6622 S.n1648 S.n1647 0.021
R6623 S.n1646 S.n1645 0.021
R6624 S.n2210 S.n2209 0.021
R6625 S.n2761 S.n2760 0.021
R6626 S.n2759 S.n2758 0.021
R6627 S.n3289 S.n3288 0.021
R6628 S.n3287 S.n3286 0.021
R6629 S.n3804 S.n3803 0.021
R6630 S.n3802 S.n3801 0.021
R6631 S.n4300 S.n4299 0.021
R6632 S.n4298 S.n4297 0.021
R6633 S.n4427 S.n4426 0.021
R6634 S.n4874 S.n4873 0.021
R6635 S.n5650 S.n5649 0.021
R6636 S.n1126 S.n1125 0.021
R6637 S.n1733 S.n1732 0.021
R6638 S.n1731 S.n1730 0.021
R6639 S.n2293 S.n2292 0.021
R6640 S.n2845 S.n2844 0.021
R6641 S.n2843 S.n2842 0.021
R6642 S.n3373 S.n3372 0.021
R6643 S.n3891 S.n3890 0.021
R6644 S.n4264 S.n4263 0.021
R6645 S.n1207 S.n1206 0.021
R6646 S.n1794 S.n1793 0.021
R6647 S.n1792 S.n1791 0.021
R6648 S.n2910 S.n2909 0.021
R6649 S.n3253 S.n3252 0.021
R6650 S.n1859 S.n1858 0.021
R6651 S.n5610 S.n5608 0.021
R6652 S.n4857 S.n4856 0.021
R6653 S.n4410 S.n4409 0.021
R6654 S.n4283 S.n4282 0.021
R6655 S.n3787 S.n3786 0.021
R6656 S.n3272 S.n3271 0.021
R6657 S.n2744 S.n2743 0.021
R6658 S.n2195 S.n2194 0.021
R6659 S.n1631 S.n1630 0.021
R6660 S.n1036 S.n1035 0.021
R6661 S.n5621 S.n5620 0.021
R6662 S.n4914 S.n4913 0.021
R6663 S.n2893 S.n2892 0.021
R6664 S.n2338 S.n2337 0.021
R6665 S.n1777 S.n1776 0.021
R6666 S.n1189 S.n1188 0.021
R6667 S.n3875 S.n3874 0.021
R6668 S.n3357 S.n3356 0.021
R6669 S.n2829 S.n2828 0.021
R6670 S.n2279 S.n2278 0.021
R6671 S.n1717 S.n1716 0.021
R6672 S.n4271 S.n4270 0.021
R6673 S.n4457 S.n4456 0.021
R6674 S.n4363 S.n4362 0.021
R6675 S.n3863 S.n3862 0.021
R6676 S.n1144 S.n1143 0.021
R6677 S.n1175 S.n1174 0.021
R6678 S.n1763 S.n1762 0.021
R6679 S.n2324 S.n2323 0.021
R6680 S.n2879 S.n2878 0.021
R6681 S.n3407 S.n3406 0.021
R6682 S.n3757 S.n3755 0.021
R6683 S.n3260 S.n3259 0.021
R6684 S.n1842 S.n1841 0.021
R6685 S.n1248 S.n1247 0.021
R6686 S.n1234 S.n1233 0.021
R6687 S.n1828 S.n1827 0.021
R6688 S.n2388 S.n2387 0.021
R6689 S.n2714 S.n2712 0.021
R6690 S.n2183 S.n2182 0.021
R6691 S.n1024 S.n1023 0.021
R6692 S.n1297 S.n1296 0.021
R6693 S.n1601 S.n1599 0.021
R6694 S.n416 S.n415 0.021
R6695 S.n398 S.n392 0.021
R6696 S.n86 S.n79 0.021
R6697 S.n54 S.n47 0.021
R6698 S.n22 S.n15 0.021
R6699 S.n374 S.n373 0.02
R6700 S.n5825 S.n5824 0.02
R6701 S.n5840 S.n5834 0.02
R6702 S.n677 S.n676 0.02
R6703 S.n333 S.n332 0.02
R6704 S.n7 S.n6 0.02
R6705 S.n502 S.n501 0.02
R6706 S.n427 S.n426 0.02
R6707 S.n5673 S.n5672 0.02
R6708 S.n4431 S.n4430 0.02
R6709 S.n4878 S.n4877 0.02
R6710 S.n5657 S.n5654 0.02
R6711 S.n3377 S.n3376 0.02
R6712 S.n3895 S.n3894 0.02
R6713 S.n4271 S.n4267 0.02
R6714 S.n4316 S.n4313 0.02
R6715 S.n4387 S.n4384 0.02
R6716 S.n4891 S.n4888 0.02
R6717 S.n3757 S.n3756 0.02
R6718 S.n3389 S.n3388 0.02
R6719 S.n2861 S.n2860 0.02
R6720 S.n2358 S.n2357 0.02
R6721 S.n2914 S.n2913 0.02
R6722 S.n3260 S.n3256 0.02
R6723 S.n2714 S.n2713 0.02
R6724 S.n2370 S.n2369 0.02
R6725 S.n1810 S.n1809 0.02
R6726 S.n1267 S.n1266 0.02
R6727 S.n1863 S.n1862 0.02
R6728 S.n2183 S.n2179 0.02
R6729 S.n1024 S.n1020 0.02
R6730 S.n1601 S.n1600 0.02
R6731 S.n1279 S.n1278 0.02
R6732 S.n416 S.n412 0.02
R6733 S.n686 S.n685 0.02
R6734 S.n4474 S.n4473 0.019
R6735 S.n4815 S.n4814 0.019
R6736 S.t191 S.n635 0.019
R6737 S.n644 S.n643 0.019
R6738 S.n926 S.n925 0.019
R6739 S.n3345 S.n3344 0.019
R6740 S.n2817 S.n2816 0.019
R6741 S.n2267 S.n2266 0.019
R6742 S.n1704 S.n1703 0.019
R6743 S.n1101 S.n1100 0.019
R6744 S.n4425 S.n4424 0.019
R6745 S.n4872 S.n4871 0.019
R6746 S.n3371 S.n3370 0.019
R6747 S.n3889 S.n3888 0.019
R6748 S.n2353 S.n2352 0.019
R6749 S.n2908 S.n2907 0.019
R6750 S.n1263 S.n1262 0.019
R6751 S.n1857 S.n1856 0.019
R6752 S.n5099 S.n5098 0.018
R6753 S.n4648 S.n4647 0.018
R6754 S.n635 S.n634 0.018
R6755 S.n4442 S.n4441 0.018
R6756 S.n4447 S.n4446 0.018
R6757 S.n4338 S.n4337 0.018
R6758 S.n4343 S.n4342 0.018
R6759 S.n3838 S.n3837 0.018
R6760 S.n3843 S.n3842 0.018
R6761 S.n3323 S.n3322 0.018
R6762 S.n3328 S.n3327 0.018
R6763 S.n2795 S.n2794 0.018
R6764 S.n2800 S.n2799 0.018
R6765 S.n2245 S.n2244 0.018
R6766 S.n2250 S.n2249 0.018
R6767 S.n1682 S.n1681 0.018
R6768 S.n1687 S.n1686 0.018
R6769 S.n1115 S.n1114 0.018
R6770 S.n1112 S.n1111 0.018
R6771 S S.n739 0.018
R6772 S.n639 S.n638 0.018
R6773 S.n83 S.n82 0.018
R6774 S.n51 S.n50 0.018
R6775 S.n5096 S.n5095 0.017
R6776 S.n4645 S.n4644 0.017
R6777 S.n400 S.n399 0.017
R6778 S.n88 S.n87 0.017
R6779 S.n56 S.n55 0.017
R6780 S.n24 S.n23 0.017
R6781 S.n5409 S.n5408 0.017
R6782 S.n5431 S.n5430 0.017
R6783 S.n4660 S.n4656 0.017
R6784 S.n79 S.n78 0.017
R6785 S.n47 S.n46 0.017
R6786 S.n539 S.n538 0.017
R6787 S.n1447 S.n1442 0.016
R6788 S.n2039 S.n2034 0.016
R6789 S.n2566 S.n2561 0.016
R6790 S.n3083 S.n3078 0.016
R6791 S.n3576 S.n3571 0.016
R6792 S.n4056 S.n4051 0.016
R6793 S.n1151 S.n1150 0.016
R6794 S.n890 S.n886 0.016
R6795 S.n3776 S.n3768 0.016
R6796 S.n2733 S.n2725 0.016
R6797 S.n1620 S.n1612 0.016
R6798 S.n3873 S.n3872 0.016
R6799 S.n3355 S.n3354 0.016
R6800 S.n2827 S.n2826 0.016
R6801 S.n2277 S.n2276 0.016
R6802 S.n1715 S.n1714 0.016
R6803 S.n1142 S.n1141 0.016
R6804 S.n5274 S.n5273 0.015
R6805 S.n5240 S.n5239 0.015
R6806 S.n5098 S.n5097 0.015
R6807 S.n4647 S.n4646 0.015
R6808 S.n4834 S.n4832 0.015
R6809 S.t240 S.n5752 0.015
R6810 S.t240 S.n5743 0.015
R6811 S.n5648 S.n5647 0.015
R6812 S.t240 S.n5728 0.015
R6813 S.n2863 S.n2862 0.015
R6814 S.n3391 S.n3390 0.015
R6815 S.n4358 S.n4352 0.015
R6816 S.n4358 S.n4357 0.015
R6817 S.n4357 S.n4356 0.015
R6818 S.n3858 S.n3852 0.015
R6819 S.n3858 S.n3857 0.015
R6820 S.n3857 S.n3856 0.015
R6821 S.n3343 S.n3342 0.015
R6822 S.n3342 S.n3341 0.015
R6823 S.n3341 S.n3340 0.015
R6824 S.n2815 S.n2814 0.015
R6825 S.n2814 S.n2813 0.015
R6826 S.n2813 S.n2812 0.015
R6827 S.n2265 S.n2264 0.015
R6828 S.n2264 S.n2263 0.015
R6829 S.n2263 S.n2262 0.015
R6830 S.n1702 S.n1701 0.015
R6831 S.n1701 S.n1700 0.015
R6832 S.n1700 S.n1699 0.015
R6833 S.n1099 S.n1098 0.015
R6834 S.n1098 S.n1097 0.015
R6835 S.n1097 S.n1096 0.015
R6836 S.n671 S.n670 0.015
R6837 S.n670 S.n669 0.015
R6838 S.n4893 S.n4892 0.015
R6839 S.n4389 S.n4388 0.015
R6840 S.n4318 S.n4317 0.015
R6841 S.n350 S.n349 0.015
R6842 S.n1812 S.n1811 0.015
R6843 S.n2372 S.n2371 0.015
R6844 S.n1281 S.n1280 0.015
R6845 S.n1151 S.n1146 0.015
R6846 S.n4860 S.n4859 0.015
R6847 S.n4413 S.n4412 0.015
R6848 S.n4286 S.n4285 0.015
R6849 S.n3790 S.n3789 0.015
R6850 S.n3275 S.n3274 0.015
R6851 S.n2747 S.n2746 0.015
R6852 S.n2198 S.n2197 0.015
R6853 S.n1634 S.n1633 0.015
R6854 S.n1039 S.n1038 0.015
R6855 S.n2896 S.n2895 0.015
R6856 S.n2341 S.n2340 0.015
R6857 S.n1780 S.n1779 0.015
R6858 S.n1192 S.n1191 0.015
R6859 S.n3402 S.n3401 0.015
R6860 S.n2874 S.n2873 0.015
R6861 S.n2319 S.n2318 0.015
R6862 S.n1758 S.n1757 0.015
R6863 S.n1171 S.n1170 0.015
R6864 S.n1845 S.n1844 0.015
R6865 S.n1251 S.n1250 0.015
R6866 S.n2383 S.n2382 0.015
R6867 S.n1823 S.n1822 0.015
R6868 S.n1229 S.n1228 0.015
R6869 S.n1292 S.n1291 0.015
R6870 S.n674 S.n673 0.014
R6871 S.n537 S.n536 0.014
R6872 S.n1043 S.n1042 0.014
R6873 S.n1196 S.n1195 0.014
R6874 S.n1766 S.n1765 0.014
R6875 S.n2327 S.n2326 0.014
R6876 S.n2882 S.n2881 0.014
R6877 S.n3410 S.n3409 0.014
R6878 S.n1255 S.n1254 0.014
R6879 S.n1831 S.n1830 0.014
R6880 S.n2391 S.n2390 0.014
R6881 S.n1300 S.n1299 0.014
R6882 S.n5285 S.n5276 0.014
R6883 S.n5252 S.n5242 0.014
R6884 S.n867 S.n866 0.014
R6885 S.n1146 S.n1145 0.014
R6886 S.n4864 S.n4863 0.013
R6887 S.n4417 S.n4416 0.013
R6888 S.n4290 S.n4289 0.013
R6889 S.n3794 S.n3793 0.013
R6890 S.n3279 S.n3278 0.013
R6891 S.n2751 S.n2750 0.013
R6892 S.n2202 S.n2201 0.013
R6893 S.n1638 S.n1637 0.013
R6894 S.n2900 S.n2899 0.013
R6895 S.n2345 S.n2344 0.013
R6896 S.n1784 S.n1783 0.013
R6897 S.n1178 S.n1177 0.013
R6898 S.n1849 S.n1848 0.013
R6899 S.n1237 S.n1236 0.013
R6900 S.n4455 S.n4454 0.013
R6901 S.n4832 S.n4816 0.013
R6902 S.n1002 S.n1001 0.013
R6903 S.n392 S.n391 0.013
R6904 S.n205 S.n204 0.013
R6905 S.n170 S.n169 0.013
R6906 S.n15 S.n14 0.013
R6907 S.t191 S.n699 0.012
R6908 S.t191 S.n0 0.012
R6909 S.t191 S.n494 0.012
R6910 S.t191 S.n525 0.012
R6911 S.t191 S.n563 0.012
R6912 S.n4861 S.n4860 0.012
R6913 S.n4414 S.n4413 0.012
R6914 S.n4287 S.n4286 0.012
R6915 S.n3791 S.n3790 0.012
R6916 S.n3276 S.n3275 0.012
R6917 S.n2748 S.n2747 0.012
R6918 S.n2199 S.n2198 0.012
R6919 S.n1635 S.n1634 0.012
R6920 S.n1040 S.n1039 0.012
R6921 S.n396 S.n395 0.012
R6922 S.n2897 S.n2896 0.012
R6923 S.n2342 S.n2341 0.012
R6924 S.n1781 S.n1780 0.012
R6925 S.n1193 S.n1192 0.012
R6926 S.n3403 S.n3402 0.012
R6927 S.n2875 S.n2874 0.012
R6928 S.n2320 S.n2319 0.012
R6929 S.n1759 S.n1758 0.012
R6930 S.n1139 S.n1138 0.012
R6931 S.n3878 S.n3877 0.012
R6932 S.n3360 S.n3359 0.012
R6933 S.n2832 S.n2831 0.012
R6934 S.n2282 S.n2281 0.012
R6935 S.n1720 S.n1719 0.012
R6936 S.n1172 S.n1171 0.012
R6937 S.n84 S.n83 0.012
R6938 S.n1846 S.n1845 0.012
R6939 S.n1252 S.n1251 0.012
R6940 S.n2384 S.n2383 0.012
R6941 S.n1824 S.n1823 0.012
R6942 S.n1230 S.n1229 0.012
R6943 S.n52 S.n51 0.012
R6944 S.n1293 S.n1292 0.012
R6945 S.n5822 S.n5821 0.012
R6946 S.n5838 S.n5837 0.012
R6947 S.n376 S.n375 0.011
R6948 S.n401 S.n389 0.011
R6949 S.n540 S.n539 0.011
R6950 S.n5437 S.n5434 0.011
R6951 S.n4816 S.n4815 0.011
R6952 S.n4360 S.n4350 0.011
R6953 S.n3860 S.n3850 0.011
R6954 S.n541 S.n540 0.01
R6955 S.n5108 S.n5096 0.01
R6956 S.n4660 S.n4645 0.01
R6957 S.n221 S.n220 0.01
R6958 S.n186 S.n185 0.01
R6959 S.n4253 S.n4252 0.01
R6960 S.n4834 S.n4382 0.01
R6961 S.n4378 S.n3928 0.01
R6962 S.n3910 S.n3443 0.01
R6963 S.n3425 S.n2947 0.01
R6964 S.n2929 S.n2425 0.01
R6965 S.n2406 S.n1897 0.01
R6966 S.n1878 S.n1565 0.01
R6967 S.n1315 S.n754 0.01
R6968 S.n1315 S.n757 0.01
R6969 S.n293 S.n290 0.01
R6970 S.n401 S.n400 0.01
R6971 S.n325 S.n323 0.01
R6972 S.n914 S.n906 0.01
R6973 S.n1455 S.n1447 0.01
R6974 S.n2047 S.n2039 0.01
R6975 S.n2574 S.n2566 0.01
R6976 S.n3091 S.n3083 0.01
R6977 S.n3585 S.n3576 0.01
R6978 S.n4065 S.n4056 0.01
R6979 S.n254 S.n250 0.01
R6980 S.n4506 S.n4502 0.01
R6981 S.n4087 S.n4083 0.01
R6982 S.n3605 S.n3601 0.01
R6983 S.n3111 S.n3107 0.01
R6984 S.n2594 S.n2590 0.01
R6985 S.n2067 S.n2063 0.01
R6986 S.n1475 S.n1471 0.01
R6987 S.n935 S.n926 0.01
R6988 S.n273 S.n270 0.01
R6989 S.n103 S.n94 0.01
R6990 S.n103 S.n88 0.01
R6991 S.n71 S.n62 0.01
R6992 S.n71 S.n56 0.01
R6993 S.n39 S.n30 0.01
R6994 S.n39 S.n24 0.01
R6995 S.n5270 S.n5267 0.01
R6996 S.n5416 S.n5409 0.01
R6997 S.n5437 S.n5431 0.01
R6998 S.n889 S.n887 0.01
R6999 S.n4485 S.n4474 0.01
R7000 S.n3541 S.n3529 0.01
R7001 S.n2493 S.n2481 0.01
R7002 S.n1335 S.n1323 0.01
R7003 S.n5270 S.n4852 0.009
R7004 S.n5709 S.n5271 0.009
R7005 S.n536 S.n535 0.009
R7006 S.n5611 S.n5610 0.009
R7007 S.n5630 S.n5621 0.009
R7008 S.n4923 S.n4914 0.009
R7009 S.n4458 S.n4457 0.009
R7010 S.n4363 S.n4361 0.009
R7011 S.n4364 S.n4363 0.009
R7012 S.n3863 S.n3861 0.009
R7013 S.n3864 S.n3863 0.009
R7014 S.n204 S.n203 0.009
R7015 S.n169 S.n168 0.009
R7016 S.n399 S.n398 0.008
R7017 S.n87 S.n86 0.008
R7018 S.n55 S.n54 0.008
R7019 S.n23 S.n22 0.008
R7020 S.n5408 S.n5407 0.008
R7021 S.n5430 S.n5429 0.008
R7022 S.n5825 S.n5823 0.008
R7023 S.n5840 S.n5839 0.008
R7024 S.n4862 S.n4861 0.008
R7025 S.n4415 S.n4414 0.008
R7026 S.n4288 S.n4287 0.008
R7027 S.n3792 S.n3791 0.008
R7028 S.n3277 S.n3276 0.008
R7029 S.n2749 S.n2748 0.008
R7030 S.n2200 S.n2199 0.008
R7031 S.n1636 S.n1635 0.008
R7032 S.n1041 S.n1040 0.008
R7033 S.n2898 S.n2897 0.008
R7034 S.n2343 S.n2342 0.008
R7035 S.n1782 S.n1781 0.008
R7036 S.n1194 S.n1193 0.008
R7037 S.n3404 S.n3403 0.008
R7038 S.n2876 S.n2875 0.008
R7039 S.n2321 S.n2320 0.008
R7040 S.n1760 S.n1759 0.008
R7041 S.n1173 S.n1172 0.008
R7042 S.n1847 S.n1846 0.008
R7043 S.n1253 S.n1252 0.008
R7044 S.n2385 S.n2384 0.008
R7045 S.n1825 S.n1824 0.008
R7046 S.n1231 S.n1230 0.008
R7047 S.n1294 S.n1293 0.008
R7048 S.n4660 S.n4659 0.008
R7049 S.n1055 S.n1052 0.008
R7050 S.n953 S.n952 0.008
R7051 S.n1652 S.n1651 0.008
R7052 S.n1494 S.n1493 0.008
R7053 S.n2215 S.n2214 0.008
R7054 S.n2085 S.n2084 0.008
R7055 S.n2765 S.n2764 0.008
R7056 S.n2612 S.n2611 0.008
R7057 S.n3293 S.n3292 0.008
R7058 S.n3129 S.n3128 0.008
R7059 S.n3808 S.n3807 0.008
R7060 S.n3623 S.n3622 0.008
R7061 S.n4304 S.n4303 0.008
R7062 S.n4105 S.n4104 0.008
R7063 S.n4524 S.n4523 0.008
R7064 S.n4975 S.n4974 0.008
R7065 S.n463 S.n437 0.008
R7066 S.n293 S.n292 0.008
R7067 S.n1127 S.n1124 0.008
R7068 S.n876 S.n875 0.008
R7069 S.n1737 S.n1736 0.008
R7070 S.n1429 S.n1428 0.008
R7071 S.n2298 S.n2297 0.008
R7072 S.n2021 S.n2020 0.008
R7073 S.n2849 S.n2848 0.008
R7074 S.n2548 S.n2547 0.008
R7075 S.n3065 S.n3064 0.008
R7076 S.n3558 S.n3557 0.008
R7077 S.n914 S.n901 0.008
R7078 S.n1455 S.n1441 0.008
R7079 S.n2047 S.n2033 0.008
R7080 S.n2574 S.n2560 0.008
R7081 S.n3091 S.n3077 0.008
R7082 S.n3585 S.n3570 0.008
R7083 S.n4065 S.n4050 0.008
R7084 S.n658 S.n657 0.008
R7085 S.n254 S.n253 0.008
R7086 S.n4506 S.n4505 0.008
R7087 S.n4087 S.n4086 0.008
R7088 S.n3605 S.n3604 0.008
R7089 S.n3111 S.n3110 0.008
R7090 S.n2594 S.n2593 0.008
R7091 S.n2067 S.n2066 0.008
R7092 S.n1475 S.n1474 0.008
R7093 S.n935 S.n924 0.008
R7094 S.n1064 S.n1063 0.008
R7095 S.n1661 S.n1660 0.008
R7096 S.n2224 S.n2223 0.008
R7097 S.n2774 S.n2773 0.008
R7098 S.n3302 S.n3301 0.008
R7099 S.n3817 S.n3816 0.008
R7100 S.n335 S.n334 0.008
R7101 S.n349 S.n345 0.008
R7102 S.n349 S.n348 0.008
R7103 S.n273 S.n272 0.008
R7104 S.n3775 S.n3773 0.008
R7105 S.n2307 S.n2306 0.008
R7106 S.n1746 S.n1745 0.008
R7107 S.n1160 S.n1159 0.008
R7108 S.n8 S.n5 0.008
R7109 S.n1208 S.n1205 0.008
R7110 S.n848 S.n847 0.008
R7111 S.n1798 S.n1797 0.008
R7112 S.n1392 S.n1391 0.008
R7113 S.n1985 S.n1984 0.008
R7114 S.n2510 S.n2509 0.008
R7115 S.n2732 S.n2728 0.008
R7116 S.n1218 S.n1217 0.008
R7117 S.n500 S.n499 0.008
R7118 S.n812 S.n811 0.008
R7119 S.n1353 S.n1352 0.008
R7120 S.n1619 S.n1615 0.008
R7121 S.n532 S.n531 0.008
R7122 S.n431 S.n430 0.008
R7123 S.n5671 S.n5670 0.008
R7124 S.t191 S.n627 0.007
R7125 S.t191 S.n620 0.007
R7126 S.t191 S.n608 0.007
R7127 S.t191 S.n596 0.007
R7128 S.n5095 S.n5094 0.007
R7129 S.n4644 S.n4643 0.007
R7130 S.n4360 S.n4359 0.007
R7131 S.n3860 S.n3859 0.007
R7132 S.n673 S.n672 0.007
R7133 S.n419 S.n418 0.007
R7134 S.t240 S.n5793 0.006
R7135 S.t240 S.n5788 0.006
R7136 S.t240 S.n5781 0.006
R7137 S.t240 S.n5774 0.006
R7138 S.t240 S.n5767 0.006
R7139 S.t240 S.n5760 0.006
R7140 S.n20 S.n19 0.006
R7141 S.n1055 S.n1054 0.006
R7142 S.n1127 S.n1126 0.006
R7143 S.n335 S.n333 0.006
R7144 S.n8 S.n7 0.006
R7145 S.n1208 S.n1207 0.006
R7146 S.n5672 S.n5671 0.006
R7147 S.n375 S.n374 0.006
R7148 S.n5826 S.n5825 0.006
R7149 S.n5841 S.n5840 0.006
R7150 S.n401 S.n379 0.006
R7151 S.n325 S.n312 0.006
R7152 S.n1140 S.n1139 0.005
R7153 S.n3879 S.n3878 0.005
R7154 S.n3361 S.n3360 0.005
R7155 S.n2833 S.n2832 0.005
R7156 S.n2283 S.n2282 0.005
R7157 S.n1721 S.n1720 0.005
R7158 S.n391 S.n390 0.005
R7159 S.t191 S.n632 0.005
R7160 S.n3770 S.n3769 0.005
R7161 S.n2727 S.n2726 0.005
R7162 S.n1614 S.n1613 0.005
R7163 S.n5823 S.n5819 0.005
R7164 S.n5839 S.n5835 0.005
R7165 S.t191 S.n675 0.005
R7166 S.n4215 S.n4214 0.004
R7167 S.n4791 S.n4790 0.004
R7168 S.n5552 S.n5551 0.004
R7169 S.n5296 S.n5295 0.004
R7170 S.n5082 S.n5081 0.004
R7171 S.n5228 S.n5227 0.004
R7172 S.n4631 S.n4630 0.004
R7173 S.n4808 S.n4807 0.004
R7174 S.n5571 S.n5570 0.004
R7175 S.n5283 S.n5282 0.004
R7176 S.n5106 S.n5105 0.004
R7177 S.n5249 S.n5248 0.004
R7178 S.n4655 S.n4654 0.004
R7179 S.n4375 S.n4374 0.004
R7180 S.n3717 S.n3716 0.004
R7181 S.n3935 S.n3934 0.004
R7182 S.n5536 S.n5535 0.004
R7183 S.n5311 S.n5310 0.004
R7184 S.n5066 S.n5065 0.004
R7185 S.n5213 S.n5212 0.004
R7186 S.n4615 S.n4614 0.004
R7187 S.n4775 S.n4774 0.004
R7188 S.n4196 S.n4195 0.004
R7189 S.n3907 S.n3906 0.004
R7190 S.n3207 S.n3206 0.004
R7191 S.n3450 S.n3449 0.004
R7192 S.n5520 S.n5519 0.004
R7193 S.n5326 S.n5325 0.004
R7194 S.n5050 S.n5049 0.004
R7195 S.n5198 S.n5197 0.004
R7196 S.n4599 S.n4598 0.004
R7197 S.n4760 S.n4759 0.004
R7198 S.n4180 S.n4179 0.004
R7199 S.n3950 S.n3949 0.004
R7200 S.n3698 S.n3697 0.004
R7201 S.n3422 S.n3421 0.004
R7202 S.n2674 S.n2673 0.004
R7203 S.n2954 S.n2953 0.004
R7204 S.n5504 S.n5503 0.004
R7205 S.n5341 S.n5340 0.004
R7206 S.n5034 S.n5033 0.004
R7207 S.n5183 S.n5182 0.004
R7208 S.n4583 S.n4582 0.004
R7209 S.n4745 S.n4744 0.004
R7210 S.n4164 S.n4163 0.004
R7211 S.n3965 S.n3964 0.004
R7212 S.n3682 S.n3681 0.004
R7213 S.n3465 S.n3464 0.004
R7214 S.n3188 S.n3187 0.004
R7215 S.n2926 S.n2925 0.004
R7216 S.n2131 S.n2130 0.004
R7217 S.n2432 S.n2431 0.004
R7218 S.n5488 S.n5487 0.004
R7219 S.n5356 S.n5355 0.004
R7220 S.n5018 S.n5017 0.004
R7221 S.n5168 S.n5167 0.004
R7222 S.n4567 S.n4566 0.004
R7223 S.n4730 S.n4729 0.004
R7224 S.n4148 S.n4147 0.004
R7225 S.n3980 S.n3979 0.004
R7226 S.n3666 S.n3665 0.004
R7227 S.n3480 S.n3479 0.004
R7228 S.n3172 S.n3171 0.004
R7229 S.n2969 S.n2968 0.004
R7230 S.n2655 S.n2654 0.004
R7231 S.n2403 S.n2402 0.004
R7232 S.n1543 S.n1542 0.004
R7233 S.n1904 S.n1903 0.004
R7234 S.n5379 S.n5378 0.004
R7235 S.n5371 S.n5370 0.004
R7236 S.n5145 S.n5144 0.004
R7237 S.n5137 S.n5136 0.004
R7238 S.n4552 S.n4551 0.004
R7239 S.n4714 S.n4713 0.004
R7240 S.n4133 S.n4132 0.004
R7241 S.n3995 S.n3994 0.004
R7242 S.n3651 S.n3650 0.004
R7243 S.n3495 S.n3494 0.004
R7244 S.n3157 S.n3156 0.004
R7245 S.n2984 S.n2983 0.004
R7246 S.n2640 S.n2639 0.004
R7247 S.n2447 S.n2446 0.004
R7248 S.n2113 S.n2112 0.004
R7249 S.n1875 S.n1874 0.004
R7250 S.n969 S.n968 0.004
R7251 S.n1571 S.n1570 0.004
R7252 S.n5471 S.n5470 0.004
R7253 S.n5603 S.n5602 0.004
R7254 S.n4942 S.n4941 0.004
R7255 S.n4934 S.n4933 0.004
R7256 S.n4537 S.n4536 0.004
R7257 S.n4698 S.n4697 0.004
R7258 S.n4118 S.n4117 0.004
R7259 S.n4011 S.n4010 0.004
R7260 S.n3636 S.n3635 0.004
R7261 S.n3511 S.n3510 0.004
R7262 S.n3142 S.n3141 0.004
R7263 S.n3000 S.n2999 0.004
R7264 S.n2625 S.n2624 0.004
R7265 S.n2463 S.n2462 0.004
R7266 S.n2098 S.n2097 0.004
R7267 S.n1920 S.n1919 0.004
R7268 S.n1523 S.n1522 0.004
R7269 S.n1312 S.n1311 0.004
R7270 S.n386 S.n385 0.004
R7271 S.n1046 S.n1045 0.004
R7272 S.n5643 S.n5642 0.004
R7273 S.n4968 S.n4967 0.004
R7274 S.n4867 S.n4866 0.004
R7275 S.n4517 S.n4516 0.004
R7276 S.n4420 S.n4419 0.004
R7277 S.n4098 S.n4097 0.004
R7278 S.n4293 S.n4292 0.004
R7279 S.n3616 S.n3615 0.004
R7280 S.n3797 S.n3796 0.004
R7281 S.n3122 S.n3121 0.004
R7282 S.n3282 S.n3281 0.004
R7283 S.n2605 S.n2604 0.004
R7284 S.n2754 S.n2753 0.004
R7285 S.n2078 S.n2077 0.004
R7286 S.n2205 S.n2204 0.004
R7287 S.n1486 S.n1485 0.004
R7288 S.n1641 S.n1640 0.004
R7289 S.n946 S.n945 0.004
R7290 S.n370 S.n369 0.004
R7291 S.n288 S.n287 0.004
R7292 S.n443 S.n442 0.004
R7293 S.n5458 S.n5457 0.004
R7294 S.n5628 S.n5627 0.004
R7295 S.n5005 S.n5004 0.004
R7296 S.n4921 S.n4920 0.004
R7297 S.n4675 S.n4674 0.004
R7298 S.n4685 S.n4684 0.004
R7299 S.n4232 S.n4231 0.004
R7300 S.n4242 S.n4241 0.004
R7301 S.n3734 S.n3733 0.004
R7302 S.n3744 S.n3743 0.004
R7303 S.n3224 S.n3223 0.004
R7304 S.n3234 S.n3233 0.004
R7305 S.n2691 S.n2690 0.004
R7306 S.n2701 S.n2700 0.004
R7307 S.n2148 S.n2147 0.004
R7308 S.n2158 S.n2157 0.004
R7309 S.n1510 S.n1509 0.004
R7310 S.n1588 S.n1587 0.004
R7311 S.n986 S.n985 0.004
R7312 S.n996 S.n995 0.004
R7313 S.n101 S.n100 0.004
R7314 S.n1199 S.n1198 0.004
R7315 S.n3247 S.n3246 0.004
R7316 S.n2503 S.n2502 0.004
R7317 S.n2903 S.n2902 0.004
R7318 S.n1978 S.n1977 0.004
R7319 S.n2348 S.n2347 0.004
R7320 S.n1384 S.n1383 0.004
R7321 S.n1787 S.n1786 0.004
R7322 S.n841 S.n840 0.004
R7323 S.n475 S.n474 0.004
R7324 S.n3767 S.n3766 0.004
R7325 S.n3045 S.n3044 0.004
R7326 S.n3400 S.n3399 0.004
R7327 S.n2528 S.n2527 0.004
R7328 S.n2872 S.n2871 0.004
R7329 S.n2001 S.n2000 0.004
R7330 S.n2317 S.n2316 0.004
R7331 S.n1408 S.n1407 0.004
R7332 S.n1756 S.n1755 0.004
R7333 S.n864 S.n863 0.004
R7334 S.n885 S.n884 0.004
R7335 S.n1136 S.n1135 0.004
R7336 S.n308 S.n307 0.004
R7337 S.n319 S.n318 0.004
R7338 S.n1726 S.n1725 0.004
R7339 S.n2288 S.n2287 0.004
R7340 S.n2838 S.n2837 0.004
R7341 S.n3366 S.n3365 0.004
R7342 S.n3884 S.n3883 0.004
R7343 S.n4258 S.n4257 0.004
R7344 S.n3551 S.n3550 0.004
R7345 S.n3058 S.n3057 0.004
R7346 S.n2541 S.n2540 0.004
R7347 S.n2014 S.n2013 0.004
R7348 S.n1421 S.n1420 0.004
R7349 S.n1108 S.n1107 0.004
R7350 S.n244 S.n243 0.004
R7351 S.n656 S.n655 0.004
R7352 S.n4450 S.n4449 0.004
R7353 S.n4059 S.n4058 0.004
R7354 S.n4346 S.n4345 0.004
R7355 S.n3579 S.n3578 0.004
R7356 S.n3846 S.n3845 0.004
R7357 S.n3086 S.n3085 0.004
R7358 S.n3331 S.n3330 0.004
R7359 S.n2569 S.n2568 0.004
R7360 S.n2803 S.n2802 0.004
R7361 S.n2042 S.n2041 0.004
R7362 S.n2253 S.n2252 0.004
R7363 S.n1450 S.n1449 0.004
R7364 S.n1690 S.n1689 0.004
R7365 S.n909 S.n908 0.004
R7366 S.n1074 S.n1073 0.004
R7367 S.n268 S.n267 0.004
R7368 S.n929 S.n928 0.004
R7369 S.n1671 S.n1670 0.004
R7370 S.n1470 S.n1469 0.004
R7371 S.n2234 S.n2233 0.004
R7372 S.n2062 S.n2061 0.004
R7373 S.n2784 S.n2783 0.004
R7374 S.n2589 S.n2588 0.004
R7375 S.n3312 S.n3311 0.004
R7376 S.n3106 S.n3105 0.004
R7377 S.n3827 S.n3826 0.004
R7378 S.n3600 S.n3599 0.004
R7379 S.n4327 S.n4326 0.004
R7380 S.n4082 S.n4081 0.004
R7381 S.n4398 S.n4397 0.004
R7382 S.n4501 S.n4500 0.004
R7383 S.n4902 S.n4901 0.004
R7384 S.n343 S.n342 0.004
R7385 S.n1169 S.n1168 0.004
R7386 S.n228 S.n227 0.004
R7387 S.n211 S.n210 0.004
R7388 S.n69 S.n68 0.004
R7389 S.n1258 S.n1257 0.004
R7390 S.n2171 S.n2170 0.004
R7391 S.n1345 S.n1344 0.004
R7392 S.n1852 S.n1851 0.004
R7393 S.n805 S.n804 0.004
R7394 S.n516 S.n515 0.004
R7395 S.n2724 S.n2723 0.004
R7396 S.n1965 S.n1964 0.004
R7397 S.n2381 S.n2380 0.004
R7398 S.n1371 S.n1370 0.004
R7399 S.n1821 S.n1820 0.004
R7400 S.n828 S.n827 0.004
R7401 S.n1227 S.n1226 0.004
R7402 S.n193 S.n192 0.004
R7403 S.n176 S.n175 0.004
R7404 S.n37 S.n36 0.004
R7405 S.n1013 S.n1012 0.004
R7406 S.n554 S.n553 0.004
R7407 S.n1611 S.n1610 0.004
R7408 S.n792 S.n791 0.004
R7409 S.n1290 S.n1289 0.004
R7410 S.n158 S.n157 0.004
R7411 S.n142 S.n141 0.004
R7412 S.n425 S.n424 0.004
R7413 S.n727 S.n726 0.004
R7414 S.n5265 S.n5264 0.004
R7415 S.n5681 S.n5680 0.004
R7416 S.n4988 S.n4987 0.004
R7417 S.n5412 S.n5411 0.004
R7418 S.n5440 S.n5439 0.004
R7419 S.n5425 S.n5424 0.004
R7420 S.t191 S.n639 0.004
R7421 S.n477 S.n476 0.004
R7422 S.n103 S.n102 0.004
R7423 S.n518 S.n517 0.004
R7424 S.n71 S.n70 0.004
R7425 S.n556 S.n555 0.004
R7426 S.n39 S.n38 0.004
R7427 S.t191 S.n687 0.004
R7428 S.n4040 S.n4039 0.004
R7429 S.n129 S.n128 0.004
R7430 S.n4813 S.n4812 0.004
R7431 S.n4354 S.n4353 0.004
R7432 S.n3854 S.n3853 0.004
R7433 S.n3337 S.n3336 0.004
R7434 S.n2809 S.n2808 0.004
R7435 S.n2259 S.n2258 0.004
R7436 S.n1696 S.n1695 0.004
R7437 S.n1093 S.n1092 0.004
R7438 S.n666 S.n665 0.004
R7439 S.n5398 S.n5397 0.004
R7440 S.n4040 S.n4038 0.004
R7441 S.n273 S.n261 0.004
R7442 S.n935 S.n934 0.004
R7443 S.n1475 S.n1463 0.004
R7444 S.n2067 S.n2055 0.004
R7445 S.n2594 S.n2582 0.004
R7446 S.n3111 S.n3099 0.004
R7447 S.n3605 S.n3593 0.004
R7448 S.n4087 S.n4075 0.004
R7449 S.n4506 S.n4494 0.004
R7450 S.n4958 S.n4956 0.004
R7451 S.n3541 S.n3540 0.004
R7452 S.n230 S.n221 0.004
R7453 S.n3029 S.n3027 0.004
R7454 S.n2493 S.n2492 0.004
R7455 S.n195 S.n186 0.004
R7456 S.n1949 S.n1947 0.004
R7457 S.n776 S.n774 0.004
R7458 S.n1335 S.n1334 0.004
R7459 S.n129 S.n127 0.004
R7460 S.n5683 S.n5674 0.004
R7461 S.n4834 S.n4833 0.004
R7462 S.n1138 S.n1137 0.004
R7463 S.n3877 S.n3876 0.004
R7464 S.n3359 S.n3358 0.004
R7465 S.n2831 S.n2830 0.004
R7466 S.n2281 S.n2280 0.004
R7467 S.n1719 S.n1718 0.004
R7468 S.n4485 S.n4471 0.004
R7469 S.n3345 S.n3343 0.004
R7470 S.n2817 S.n2815 0.004
R7471 S.n2267 S.n2265 0.004
R7472 S.n1704 S.n1702 0.004
R7473 S.n1101 S.n1099 0.004
R7474 S.n890 S.n889 0.004
R7475 S.n3776 S.n3775 0.004
R7476 S.n3541 S.n3528 0.004
R7477 S.n2733 S.n2732 0.004
R7478 S.n2493 S.n2480 0.004
R7479 S.n1620 S.n1619 0.004
R7480 S.n1335 S.n1322 0.004
R7481 S.n160 S.n152 0.004
R7482 S.t240 S.n5787 0.004
R7483 S.t240 S.n5795 0.004
R7484 S.t240 S.n5780 0.004
R7485 S.t240 S.n5773 0.004
R7486 S.t240 S.n5766 0.004
R7487 S.t240 S.n5759 0.004
R7488 S.t240 S.n5750 0.004
R7489 S.t240 S.n5741 0.004
R7490 S.n5445 S.n5444 0.004
R7491 S.t191 S.n585 0.004
R7492 S.t52 S.n5401 0.004
R7493 S.t191 S.n622 0.004
R7494 S.t27 S.n3032 0.004
R7495 S.t191 S.n716 0.004
R7496 S.t6 S.n3544 0.004
R7497 S.t191 S.n637 0.004
R7498 S.t65 S.n4043 0.004
R7499 S.t191 S.n684 0.004
R7500 S.t4 S.n4488 0.004
R7501 S.t45 S.n4961 0.004
R7502 S.t191 S.n701 0.004
R7503 S.t191 S.n610 0.004
R7504 S.t56 S.n1952 0.004
R7505 S.t191 S.n712 0.004
R7506 S.t68 S.n2496 0.004
R7507 S.t191 S.n598 0.004
R7508 S.t14 S.n779 0.004
R7509 S.t191 S.n708 0.004
R7510 S.t32 S.n1338 0.004
R7511 S.t191 S.n704 0.004
R7512 S.t213 S.n132 0.004
R7513 S.t240 S.n5791 0.004
R7514 S.t240 S.n5798 0.004
R7515 S.t240 S.n5784 0.004
R7516 S.t240 S.n5777 0.004
R7517 S.t240 S.n5770 0.004
R7518 S.t240 S.n5763 0.004
R7519 S.t240 S.n5756 0.004
R7520 S.t240 S.n5747 0.004
R7521 S.t240 S.n5738 0.004
R7522 S.t240 S.n5829 0.004
R7523 S.t240 S.n5730 0.004
R7524 S.n730 S.n725 0.004
R7525 S.t34 S.n5691 0.004
R7526 S.t240 S.n5733 0.004
R7527 S.t191 S.n493 0.004
R7528 S.t191 S.n524 0.004
R7529 S.t191 S.n562 0.004
R7530 S.t191 S.n574 0.004
R7531 S.n310 S.n309 0.004
R7532 S.n730 S.n724 0.004
R7533 S.t191 S.n614 0.004
R7534 S.t191 S.n602 0.004
R7535 S.t191 S.n589 0.004
R7536 S.n4958 S.n4957 0.004
R7537 S.n3559 S.n3548 0.004
R7538 S.n3066 S.n3055 0.004
R7539 S.n2549 S.n2538 0.004
R7540 S.n2022 S.n2011 0.004
R7541 S.n1430 S.n1418 0.004
R7542 S.n720 S.n719 0.003
R7543 S.n5419 S.n5418 0.003
R7544 S.n4373 S.n4372 0.003
R7545 S.n4220 S.n4219 0.003
R7546 S.n4798 S.n4797 0.003
R7547 S.n5560 S.n5559 0.003
R7548 S.n5306 S.n5305 0.003
R7549 S.n5090 S.n5089 0.003
R7550 S.n5235 S.n5234 0.003
R7551 S.n4639 S.n4638 0.003
R7552 S.n4804 S.n4803 0.003
R7553 S.n5576 S.n5575 0.003
R7554 S.n5291 S.n5290 0.003
R7555 S.n5111 S.n5110 0.003
R7556 S.n5255 S.n5254 0.003
R7557 S.n4663 S.n4662 0.003
R7558 S.n3905 S.n3904 0.003
R7559 S.n3722 S.n3721 0.003
R7560 S.n3945 S.n3944 0.003
R7561 S.n5544 S.n5543 0.003
R7562 S.n5321 S.n5320 0.003
R7563 S.n5074 S.n5073 0.003
R7564 S.n5220 S.n5219 0.003
R7565 S.n4623 S.n4622 0.003
R7566 S.n4782 S.n4781 0.003
R7567 S.n4204 S.n4203 0.003
R7568 S.n3420 S.n3419 0.003
R7569 S.n3212 S.n3211 0.003
R7570 S.n3460 S.n3459 0.003
R7571 S.n5528 S.n5527 0.003
R7572 S.n5336 S.n5335 0.003
R7573 S.n5058 S.n5057 0.003
R7574 S.n5205 S.n5204 0.003
R7575 S.n4607 S.n4606 0.003
R7576 S.n4767 S.n4766 0.003
R7577 S.n4188 S.n4187 0.003
R7578 S.n3960 S.n3959 0.003
R7579 S.n3706 S.n3705 0.003
R7580 S.n2924 S.n2923 0.003
R7581 S.n2679 S.n2678 0.003
R7582 S.n2964 S.n2963 0.003
R7583 S.n5512 S.n5511 0.003
R7584 S.n5351 S.n5350 0.003
R7585 S.n5042 S.n5041 0.003
R7586 S.n5190 S.n5189 0.003
R7587 S.n4591 S.n4590 0.003
R7588 S.n4752 S.n4751 0.003
R7589 S.n4172 S.n4171 0.003
R7590 S.n3975 S.n3974 0.003
R7591 S.n3690 S.n3689 0.003
R7592 S.n3475 S.n3474 0.003
R7593 S.n3196 S.n3195 0.003
R7594 S.n2401 S.n2400 0.003
R7595 S.n2136 S.n2135 0.003
R7596 S.n2442 S.n2441 0.003
R7597 S.n5496 S.n5495 0.003
R7598 S.n5366 S.n5365 0.003
R7599 S.n5026 S.n5025 0.003
R7600 S.n5175 S.n5174 0.003
R7601 S.n4575 S.n4574 0.003
R7602 S.n4737 S.n4736 0.003
R7603 S.n4156 S.n4155 0.003
R7604 S.n3990 S.n3989 0.003
R7605 S.n3674 S.n3673 0.003
R7606 S.n3490 S.n3489 0.003
R7607 S.n3180 S.n3179 0.003
R7608 S.n2979 S.n2978 0.003
R7609 S.n2663 S.n2662 0.003
R7610 S.n1873 S.n1872 0.003
R7611 S.n1537 S.n1536 0.003
R7612 S.n1915 S.n1914 0.003
R7613 S.n5585 S.n5584 0.003
R7614 S.n5598 S.n5597 0.003
R7615 S.n5151 S.n5150 0.003
R7616 S.n5160 S.n5159 0.003
R7617 S.n4559 S.n4558 0.003
R7618 S.n4722 S.n4721 0.003
R7619 S.n4140 S.n4139 0.003
R7620 S.n4006 S.n4005 0.003
R7621 S.n3658 S.n3657 0.003
R7622 S.n3506 S.n3505 0.003
R7623 S.n3164 S.n3163 0.003
R7624 S.n2995 S.n2994 0.003
R7625 S.n2647 S.n2646 0.003
R7626 S.n2458 S.n2457 0.003
R7627 S.n2120 S.n2119 0.003
R7628 S.n1310 S.n1309 0.003
R7629 S.n974 S.n973 0.003
R7630 S.n1581 S.n1580 0.003
R7631 S.n5480 S.n5479 0.003
R7632 S.n5617 S.n5616 0.003
R7633 S.n5120 S.n5119 0.003
R7634 S.n5129 S.n5128 0.003
R7635 S.n4544 S.n4543 0.003
R7636 S.n4706 S.n4705 0.003
R7637 S.n4125 S.n4124 0.003
R7638 S.n4022 S.n4021 0.003
R7639 S.n3643 S.n3642 0.003
R7640 S.n3522 S.n3521 0.003
R7641 S.n3149 S.n3148 0.003
R7642 S.n3011 S.n3010 0.003
R7643 S.n2632 S.n2631 0.003
R7644 S.n2474 S.n2473 0.003
R7645 S.n2105 S.n2104 0.003
R7646 S.n1931 S.n1930 0.003
R7647 S.n1531 S.n1530 0.003
R7648 S.n407 S.n406 0.003
R7649 S.n1059 S.n1058 0.003
R7650 S.n5664 S.n5663 0.003
R7651 S.n4982 S.n4981 0.003
R7652 S.n4885 S.n4884 0.003
R7653 S.n4531 S.n4530 0.003
R7654 S.n4438 S.n4437 0.003
R7655 S.n4112 S.n4111 0.003
R7656 S.n4308 S.n4307 0.003
R7657 S.n3630 S.n3629 0.003
R7658 S.n3812 S.n3811 0.003
R7659 S.n3136 S.n3135 0.003
R7660 S.n3297 S.n3296 0.003
R7661 S.n2619 S.n2618 0.003
R7662 S.n2769 S.n2768 0.003
R7663 S.n2092 S.n2091 0.003
R7664 S.n2219 S.n2218 0.003
R7665 S.n1501 S.n1500 0.003
R7666 S.n1656 S.n1655 0.003
R7667 S.n960 S.n959 0.003
R7668 S.n364 S.n363 0.003
R7669 S.n296 S.n295 0.003
R7670 S.n466 S.n465 0.003
R7671 S.n5463 S.n5462 0.003
R7672 S.n5636 S.n5635 0.003
R7673 S.n5010 S.n5009 0.003
R7674 S.n4926 S.n4925 0.003
R7675 S.n4669 S.n4668 0.003
R7676 S.n4690 S.n4689 0.003
R7677 S.n4226 S.n4225 0.003
R7678 S.n4250 S.n4249 0.003
R7679 S.n3728 S.n3727 0.003
R7680 S.n3752 S.n3751 0.003
R7681 S.n3218 S.n3217 0.003
R7682 S.n3242 S.n3241 0.003
R7683 S.n2685 S.n2684 0.003
R7684 S.n2709 S.n2708 0.003
R7685 S.n2142 S.n2141 0.003
R7686 S.n2166 S.n2165 0.003
R7687 S.n1515 S.n1514 0.003
R7688 S.n1596 S.n1595 0.003
R7689 S.n980 S.n979 0.003
R7690 S.n1008 S.n1007 0.003
R7691 S.n109 S.n108 0.003
R7692 S.n1212 S.n1211 0.003
R7693 S.n3267 S.n3266 0.003
R7694 S.n2517 S.n2516 0.003
R7695 S.n2918 S.n2917 0.003
R7696 S.n1992 S.n1991 0.003
R7697 S.n2362 S.n2361 0.003
R7698 S.n1399 S.n1398 0.003
R7699 S.n1802 S.n1801 0.003
R7700 S.n855 S.n854 0.003
R7701 S.n469 S.n468 0.003
R7702 S.n3782 S.n3781 0.003
R7703 S.n3053 S.n3052 0.003
R7704 S.n3414 S.n3413 0.003
R7705 S.n2536 S.n2535 0.003
R7706 S.n2886 S.n2885 0.003
R7707 S.n2009 S.n2008 0.003
R7708 S.n2331 S.n2330 0.003
R7709 S.n1416 S.n1415 0.003
R7710 S.n1770 S.n1769 0.003
R7711 S.n874 S.n873 0.003
R7712 S.n896 S.n895 0.003
R7713 S.n1154 S.n1153 0.003
R7714 S.n302 S.n301 0.003
R7715 S.n331 S.n330 0.003
R7716 S.n1741 S.n1740 0.003
R7717 S.n2302 S.n2301 0.003
R7718 S.n2853 S.n2852 0.003
R7719 S.n3381 S.n3380 0.003
R7720 S.n3899 S.n3898 0.003
R7721 S.n4278 S.n4277 0.003
R7722 S.n3565 S.n3564 0.003
R7723 S.n3072 S.n3071 0.003
R7724 S.n2555 S.n2554 0.003
R7725 S.n2028 S.n2027 0.003
R7726 S.n1436 S.n1435 0.003
R7727 S.n1120 S.n1119 0.003
R7728 S.n260 S.n259 0.003
R7729 S.n650 S.n649 0.003
R7730 S.n4461 S.n4460 0.003
R7731 S.n4071 S.n4070 0.003
R7732 S.n4367 S.n4366 0.003
R7733 S.n3591 S.n3590 0.003
R7734 S.n3867 S.n3866 0.003
R7735 S.n3097 S.n3096 0.003
R7736 S.n3349 S.n3348 0.003
R7737 S.n2580 S.n2579 0.003
R7738 S.n2821 S.n2820 0.003
R7739 S.n2053 S.n2052 0.003
R7740 S.n2271 S.n2270 0.003
R7741 S.n1461 S.n1460 0.003
R7742 S.n1708 S.n1707 0.003
R7743 S.n920 S.n919 0.003
R7744 S.n1087 S.n1086 0.003
R7745 S.n279 S.n278 0.003
R7746 S.n941 S.n940 0.003
R7747 S.n1676 S.n1675 0.003
R7748 S.n1481 S.n1480 0.003
R7749 S.n2239 S.n2238 0.003
R7750 S.n2073 S.n2072 0.003
R7751 S.n2789 S.n2788 0.003
R7752 S.n2600 S.n2599 0.003
R7753 S.n3317 S.n3316 0.003
R7754 S.n3117 S.n3116 0.003
R7755 S.n3832 S.n3831 0.003
R7756 S.n3611 S.n3610 0.003
R7757 S.n4332 S.n4331 0.003
R7758 S.n4093 S.n4092 0.003
R7759 S.n4406 S.n4405 0.003
R7760 S.n4512 S.n4511 0.003
R7761 S.n4907 S.n4906 0.003
R7762 S.n357 S.n356 0.003
R7763 S.n1182 S.n1181 0.003
R7764 S.n236 S.n235 0.003
R7765 S.n219 S.n218 0.003
R7766 S.n77 S.n76 0.003
R7767 S.n1271 S.n1270 0.003
R7768 S.n2190 S.n2189 0.003
R7769 S.n1360 S.n1359 0.003
R7770 S.n1867 S.n1866 0.003
R7771 S.n819 S.n818 0.003
R7772 S.n510 S.n509 0.003
R7773 S.n2739 S.n2738 0.003
R7774 S.n1973 S.n1972 0.003
R7775 S.n2395 S.n2394 0.003
R7776 S.n1379 S.n1378 0.003
R7777 S.n1835 S.n1834 0.003
R7778 S.n836 S.n835 0.003
R7779 S.n1241 S.n1240 0.003
R7780 S.n201 S.n200 0.003
R7781 S.n184 S.n183 0.003
R7782 S.n45 S.n44 0.003
R7783 S.n1031 S.n1030 0.003
R7784 S.n548 S.n547 0.003
R7785 S.n1626 S.n1625 0.003
R7786 S.n800 S.n799 0.003
R7787 S.n1304 S.n1303 0.003
R7788 S.n166 S.n165 0.003
R7789 S.n150 S.n149 0.003
R7790 S.n411 S.n410 0.003
R7791 S.n5422 S.n5421 0.003
R7792 S.n5261 S.n5260 0.003
R7793 S.n5686 S.n5685 0.003
R7794 S.n4996 S.n4995 0.003
R7795 S.n5448 S.n5447 0.003
R7796 S.n868 S.n867 0.003
R7797 S.n4217 S.n4212 0.003
R7798 S.n4795 S.n4794 0.003
R7799 S.n5557 S.n5555 0.003
R7800 S.n5300 S.n5299 0.003
R7801 S.n5087 S.n5085 0.003
R7802 S.n5232 S.n5231 0.003
R7803 S.n4636 S.n4634 0.003
R7804 S.n5573 S.n5568 0.003
R7805 S.n5285 S.n5280 0.003
R7806 S.n5108 S.n5103 0.003
R7807 S.n5252 S.n5246 0.003
R7808 S.n4660 S.n4652 0.003
R7809 S.n3719 S.n3714 0.003
R7810 S.n3939 S.n3938 0.003
R7811 S.n5541 S.n5539 0.003
R7812 S.n5315 S.n5314 0.003
R7813 S.n5071 S.n5069 0.003
R7814 S.n5217 S.n5216 0.003
R7815 S.n4620 S.n4618 0.003
R7816 S.n4779 S.n4778 0.003
R7817 S.n4201 S.n4199 0.003
R7818 S.n3209 S.n3204 0.003
R7819 S.n3454 S.n3453 0.003
R7820 S.n5525 S.n5523 0.003
R7821 S.n5330 S.n5329 0.003
R7822 S.n5055 S.n5053 0.003
R7823 S.n5202 S.n5201 0.003
R7824 S.n4604 S.n4602 0.003
R7825 S.n4764 S.n4763 0.003
R7826 S.n4185 S.n4183 0.003
R7827 S.n3954 S.n3953 0.003
R7828 S.n3703 S.n3701 0.003
R7829 S.n2676 S.n2671 0.003
R7830 S.n2958 S.n2957 0.003
R7831 S.n5509 S.n5507 0.003
R7832 S.n5345 S.n5344 0.003
R7833 S.n5039 S.n5037 0.003
R7834 S.n5187 S.n5186 0.003
R7835 S.n4588 S.n4586 0.003
R7836 S.n4749 S.n4748 0.003
R7837 S.n4169 S.n4167 0.003
R7838 S.n3969 S.n3968 0.003
R7839 S.n3687 S.n3685 0.003
R7840 S.n3469 S.n3468 0.003
R7841 S.n3193 S.n3191 0.003
R7842 S.n2133 S.n2128 0.003
R7843 S.n2436 S.n2435 0.003
R7844 S.n5493 S.n5491 0.003
R7845 S.n5360 S.n5359 0.003
R7846 S.n5023 S.n5021 0.003
R7847 S.n5172 S.n5171 0.003
R7848 S.n4572 S.n4570 0.003
R7849 S.n4734 S.n4733 0.003
R7850 S.n4153 S.n4151 0.003
R7851 S.n3984 S.n3983 0.003
R7852 S.n3671 S.n3669 0.003
R7853 S.n3484 S.n3483 0.003
R7854 S.n3177 S.n3175 0.003
R7855 S.n2973 S.n2972 0.003
R7856 S.n2660 S.n2658 0.003
R7857 S.n1545 S.n1320 0.003
R7858 S.n1909 S.n1907 0.003
R7859 S.n5589 S.n5588 0.003
R7860 S.n5592 S.n5374 0.003
R7861 S.n5155 S.n5154 0.003
R7862 S.n5157 S.n5140 0.003
R7863 S.n4556 S.n4555 0.003
R7864 S.n4719 S.n4717 0.003
R7865 S.n4137 S.n4136 0.003
R7866 S.n4000 S.n3998 0.003
R7867 S.n3655 S.n3654 0.003
R7868 S.n3500 S.n3498 0.003
R7869 S.n3161 S.n3160 0.003
R7870 S.n2989 S.n2987 0.003
R7871 S.n2644 S.n2643 0.003
R7872 S.n2452 S.n2450 0.003
R7873 S.n2117 S.n2116 0.003
R7874 S.n971 S.n966 0.003
R7875 S.n1575 S.n1574 0.003
R7876 S.n5477 S.n5474 0.003
R7877 S.n5611 S.n5606 0.003
R7878 S.n5124 S.n5123 0.003
R7879 S.n5126 S.n4937 0.003
R7880 S.n4541 S.n4540 0.003
R7881 S.n4703 S.n4701 0.003
R7882 S.n4122 S.n4121 0.003
R7883 S.n4016 S.n4014 0.003
R7884 S.n3640 S.n3639 0.003
R7885 S.n3516 S.n3514 0.003
R7886 S.n3146 S.n3145 0.003
R7887 S.n3005 S.n3003 0.003
R7888 S.n2629 S.n2628 0.003
R7889 S.n2468 S.n2466 0.003
R7890 S.n2102 S.n2101 0.003
R7891 S.n1925 S.n1923 0.003
R7892 S.n1528 S.n1526 0.003
R7893 S.n401 S.n383 0.003
R7894 S.n1056 S.n1049 0.003
R7895 S.n5658 S.n5646 0.003
R7896 S.n4976 S.n4971 0.003
R7897 S.n4879 S.n4870 0.003
R7898 S.n4525 S.n4520 0.003
R7899 S.n4432 S.n4423 0.003
R7900 S.n4106 S.n4101 0.003
R7901 S.n4305 S.n4296 0.003
R7902 S.n3624 S.n3619 0.003
R7903 S.n3809 S.n3800 0.003
R7904 S.n3130 S.n3125 0.003
R7905 S.n3294 S.n3285 0.003
R7906 S.n2613 S.n2608 0.003
R7907 S.n2766 S.n2757 0.003
R7908 S.n2086 S.n2081 0.003
R7909 S.n2216 S.n2208 0.003
R7910 S.n1495 S.n1489 0.003
R7911 S.n1653 S.n1644 0.003
R7912 S.n954 S.n949 0.003
R7913 S.n377 S.n361 0.003
R7914 S.n293 S.n285 0.003
R7915 S.n5460 S.n5455 0.003
R7916 S.n5630 S.n5625 0.003
R7917 S.n5007 S.n5002 0.003
R7918 S.n4923 S.n4918 0.003
R7919 S.n4677 S.n4468 0.003
R7920 S.n4687 S.n4682 0.003
R7921 S.n4234 S.n4026 0.003
R7922 S.n4244 S.n4239 0.003
R7923 S.n3736 S.n3526 0.003
R7924 S.n3746 S.n3741 0.003
R7925 S.n3226 S.n3015 0.003
R7926 S.n3236 S.n3231 0.003
R7927 S.n2693 S.n2478 0.003
R7928 S.n2703 S.n2698 0.003
R7929 S.n2150 S.n1935 0.003
R7930 S.n2160 S.n2155 0.003
R7931 S.n1512 S.n1507 0.003
R7932 S.n1590 S.n1585 0.003
R7933 S.n988 S.n762 0.003
R7934 S.n1002 S.n993 0.003
R7935 S.n103 S.n98 0.003
R7936 S.n1209 S.n1202 0.003
R7937 S.n3261 S.n3250 0.003
R7938 S.n2511 S.n2506 0.003
R7939 S.n2915 S.n2906 0.003
R7940 S.n1986 S.n1981 0.003
R7941 S.n2359 S.n2351 0.003
R7942 S.n1393 S.n1387 0.003
R7943 S.n1799 S.n1790 0.003
R7944 S.n849 S.n844 0.003
R7945 S.n477 S.n13 0.003
R7946 S.n3776 S.n3764 0.003
R7947 S.n3047 S.n3042 0.003
R7948 S.n3411 S.n3397 0.003
R7949 S.n2530 S.n2525 0.003
R7950 S.n2883 S.n2869 0.003
R7951 S.n2003 S.n1998 0.003
R7952 S.n2328 S.n2314 0.003
R7953 S.n1410 S.n1405 0.003
R7954 S.n1767 S.n1753 0.003
R7955 S.n868 S.n861 0.003
R7956 S.n890 S.n882 0.003
R7957 S.n1151 S.n1133 0.003
R7958 S.n310 S.n113 0.003
R7959 S.n325 S.n316 0.003
R7960 S.n1738 S.n1729 0.003
R7961 S.n2299 S.n2291 0.003
R7962 S.n2850 S.n2841 0.003
R7963 S.n3378 S.n3369 0.003
R7964 S.n3896 S.n3887 0.003
R7965 S.n4272 S.n4261 0.003
R7966 S.n3559 S.n3554 0.003
R7967 S.n3066 S.n3061 0.003
R7968 S.n2549 S.n2544 0.003
R7969 S.n2022 S.n2017 0.003
R7970 S.n1430 S.n1424 0.003
R7971 S.n1117 S.n1105 0.003
R7972 S.n254 S.n241 0.003
R7973 S.n659 S.n647 0.003
R7974 S.n4458 S.n4453 0.003
R7975 S.n4065 S.n4062 0.003
R7976 S.n4364 S.n4349 0.003
R7977 S.n3585 S.n3582 0.003
R7978 S.n3864 S.n3849 0.003
R7979 S.n3091 S.n3089 0.003
R7980 S.n3346 S.n3334 0.003
R7981 S.n2574 S.n2572 0.003
R7982 S.n2818 S.n2806 0.003
R7983 S.n2047 S.n2045 0.003
R7984 S.n2268 S.n2256 0.003
R7985 S.n1455 S.n1453 0.003
R7986 S.n1705 S.n1693 0.003
R7987 S.n914 S.n912 0.003
R7988 S.n1084 S.n1071 0.003
R7989 S.n273 S.n265 0.003
R7990 S.n935 S.n932 0.003
R7991 S.n1673 S.n1668 0.003
R7992 S.n1475 S.n1467 0.003
R7993 S.n2236 S.n2231 0.003
R7994 S.n2067 S.n2059 0.003
R7995 S.n2786 S.n2781 0.003
R7996 S.n2594 S.n2586 0.003
R7997 S.n3314 S.n3309 0.003
R7998 S.n3111 S.n3103 0.003
R7999 S.n3829 S.n3824 0.003
R8000 S.n3605 S.n3597 0.003
R8001 S.n4329 S.n4324 0.003
R8002 S.n4087 S.n4079 0.003
R8003 S.n4400 S.n4395 0.003
R8004 S.n4506 S.n4498 0.003
R8005 S.n4904 S.n4899 0.003
R8006 S.n351 S.n340 0.003
R8007 S.n1179 S.n1166 0.003
R8008 S.n230 S.n225 0.003
R8009 S.n213 S.n208 0.003
R8010 S.n71 S.n66 0.003
R8011 S.n1268 S.n1261 0.003
R8012 S.n2184 S.n2174 0.003
R8013 S.n1354 S.n1348 0.003
R8014 S.n1864 S.n1855 0.003
R8015 S.n813 S.n808 0.003
R8016 S.n518 S.n507 0.003
R8017 S.n2733 S.n2721 0.003
R8018 S.n1967 S.n1962 0.003
R8019 S.n2392 S.n2378 0.003
R8020 S.n1373 S.n1368 0.003
R8021 S.n1832 S.n1818 0.003
R8022 S.n830 S.n825 0.003
R8023 S.n1238 S.n1224 0.003
R8024 S.n195 S.n190 0.003
R8025 S.n178 S.n173 0.003
R8026 S.n39 S.n34 0.003
R8027 S.n1025 S.n1016 0.003
R8028 S.n556 S.n545 0.003
R8029 S.n1620 S.n1608 0.003
R8030 S.n794 S.n789 0.003
R8031 S.n1301 S.n1287 0.003
R8032 S.n160 S.n155 0.003
R8033 S.n144 S.n139 0.003
R8034 S.n432 S.n422 0.003
R8035 S.n5683 S.n5678 0.003
R8036 S.n4990 S.n4985 0.003
R8037 S.n695 S.n693 0.003
R8038 S.n4 S.n2 0.003
R8039 S.n498 S.n496 0.003
R8040 S.n529 S.n527 0.003
R8041 S.n567 S.n565 0.003
R8042 S.n5844 S.n5843 0.003
R8043 S.n5844 S.n5722 0.003
R8044 S.n4485 S.n4484 0.003
R8045 S.n679 S.n678 0.003
R8046 S.n337 S.n336 0.003
R8047 S.n10 S.n9 0.003
R8048 S.n504 S.n503 0.003
R8049 S.n542 S.n541 0.003
R8050 S.n4814 S.n4809 0.003
R8051 S.n323 S.n322 0.003
R8052 S.n4473 S.n4472 0.003
R8053 S.n3346 S.n3345 0.003
R8054 S.n2818 S.n2817 0.003
R8055 S.n2268 S.n2267 0.003
R8056 S.n1705 S.n1704 0.003
R8057 S.n1117 S.n1101 0.003
R8058 S.n94 S.n93 0.003
R8059 S.n62 S.n61 0.003
R8060 S.n538 S.n533 0.003
R8061 S.n538 S.n537 0.003
R8062 S.n30 S.n29 0.003
R8063 S.n4378 S.n3926 0.003
R8064 S.n3910 S.n3441 0.003
R8065 S.n3425 S.n2945 0.003
R8066 S.n2929 S.n2423 0.003
R8067 S.t240 S.n5831 0.003
R8068 S.n463 S.n462 0.003
R8069 S.n5398 S.n5381 0.003
R8070 S.n3029 S.n3028 0.003
R8071 S.n1949 S.n1948 0.003
R8072 S.n776 S.n775 0.003
R8073 S.n4795 S.n4788 0.003
R8074 S.t240 S.n5725 0.003
R8075 S.t240 S.n5816 0.003
R8076 S.n4895 S.n4894 0.003
R8077 S.n4391 S.n4390 0.003
R8078 S.n4320 S.n4319 0.003
R8079 S.n2406 S.n1895 0.003
R8080 S.n1878 S.n1562 0.003
R8081 S.n3047 S.n3038 0.003
R8082 S.n2530 S.n2521 0.003
R8083 S.n2003 S.n1994 0.003
R8084 S.n1410 S.n1401 0.003
R8085 S.n868 S.n857 0.003
R8086 S.n1967 S.n1958 0.003
R8087 S.n1373 S.n1364 0.003
R8088 S.n830 S.n821 0.003
R8089 S.n794 S.n785 0.003
R8090 S.n5709 S.n5708 0.003
R8091 S.n377 S.n376 0.003
R8092 S.n1265 S.n1264 0.003
R8093 S.n1019 S.n1018 0.003
R8094 S.n4359 S.n4358 0.003
R8095 S.n3859 S.n3858 0.003
R8096 S.n672 S.n671 0.003
R8097 S.n4660 S.n4649 0.002
R8098 S.n5252 S.n5243 0.002
R8099 S.n5108 S.n5100 0.002
R8100 S.n5285 S.n5277 0.002
R8101 S.n5573 S.n5565 0.002
R8102 S.n5557 S.n5548 0.002
R8103 S.n5300 S.n5292 0.002
R8104 S.n5087 S.n5078 0.002
R8105 S.n5232 S.n5224 0.002
R8106 S.n4636 S.n4627 0.002
R8107 S.n4795 S.n4786 0.002
R8108 S.n4217 S.n4209 0.002
R8109 S.n5541 S.n5532 0.002
R8110 S.n5315 S.n5307 0.002
R8111 S.n5071 S.n5062 0.002
R8112 S.n5217 S.n5209 0.002
R8113 S.n4620 S.n4611 0.002
R8114 S.n4779 S.n4771 0.002
R8115 S.n4201 S.n4192 0.002
R8116 S.n3939 S.n3931 0.002
R8117 S.n3719 S.n3711 0.002
R8118 S.n5525 S.n5516 0.002
R8119 S.n5330 S.n5322 0.002
R8120 S.n5055 S.n5046 0.002
R8121 S.n5202 S.n5194 0.002
R8122 S.n4604 S.n4595 0.002
R8123 S.n4764 S.n4756 0.002
R8124 S.n4185 S.n4176 0.002
R8125 S.n3954 S.n3946 0.002
R8126 S.n3703 S.n3694 0.002
R8127 S.n3454 S.n3446 0.002
R8128 S.n3209 S.n3201 0.002
R8129 S.n5509 S.n5500 0.002
R8130 S.n5345 S.n5337 0.002
R8131 S.n5039 S.n5030 0.002
R8132 S.n5187 S.n5179 0.002
R8133 S.n4588 S.n4579 0.002
R8134 S.n4749 S.n4741 0.002
R8135 S.n4169 S.n4160 0.002
R8136 S.n3969 S.n3961 0.002
R8137 S.n3687 S.n3678 0.002
R8138 S.n3469 S.n3461 0.002
R8139 S.n3193 S.n3184 0.002
R8140 S.n2958 S.n2950 0.002
R8141 S.n2676 S.n2668 0.002
R8142 S.n5493 S.n5484 0.002
R8143 S.n5360 S.n5352 0.002
R8144 S.n5023 S.n5014 0.002
R8145 S.n5172 S.n5164 0.002
R8146 S.n4572 S.n4563 0.002
R8147 S.n4734 S.n4726 0.002
R8148 S.n4153 S.n4144 0.002
R8149 S.n3984 S.n3976 0.002
R8150 S.n3671 S.n3662 0.002
R8151 S.n3484 S.n3476 0.002
R8152 S.n3177 S.n3168 0.002
R8153 S.n2973 S.n2965 0.002
R8154 S.n2660 S.n2651 0.002
R8155 S.n2436 S.n2428 0.002
R8156 S.n2133 S.n2125 0.002
R8157 S.n5589 S.n5375 0.002
R8158 S.n5592 S.n5367 0.002
R8159 S.n5155 S.n5141 0.002
R8160 S.n5157 S.n5133 0.002
R8161 S.n4556 S.n4548 0.002
R8162 S.n4719 S.n4710 0.002
R8163 S.n4137 S.n4129 0.002
R8164 S.n4000 S.n3991 0.002
R8165 S.n3655 S.n3647 0.002
R8166 S.n3500 S.n3491 0.002
R8167 S.n3161 S.n3153 0.002
R8168 S.n2989 S.n2980 0.002
R8169 S.n2644 S.n2636 0.002
R8170 S.n2452 S.n2443 0.002
R8171 S.n2117 S.n2109 0.002
R8172 S.n1909 S.n1900 0.002
R8173 S.n5477 S.n5467 0.002
R8174 S.n5611 S.n5599 0.002
R8175 S.n5124 S.n4938 0.002
R8176 S.n5126 S.n4930 0.002
R8177 S.n4541 S.n4533 0.002
R8178 S.n4703 S.n4694 0.002
R8179 S.n4122 S.n4114 0.002
R8180 S.n4016 S.n4007 0.002
R8181 S.n3640 S.n3632 0.002
R8182 S.n3516 S.n3507 0.002
R8183 S.n3146 S.n3138 0.002
R8184 S.n3005 S.n2996 0.002
R8185 S.n2629 S.n2621 0.002
R8186 S.n2468 S.n2459 0.002
R8187 S.n2102 S.n2094 0.002
R8188 S.n1925 S.n1916 0.002
R8189 S.n1528 S.n1519 0.002
R8190 S.n1575 S.n1567 0.002
R8191 S.n1002 S.n990 0.002
R8192 S.n988 S.n759 0.002
R8193 S.n1590 S.n1582 0.002
R8194 S.n1512 S.n1504 0.002
R8195 S.n2160 S.n2152 0.002
R8196 S.n2150 S.n1932 0.002
R8197 S.n2703 S.n2695 0.002
R8198 S.n2693 S.n2475 0.002
R8199 S.n3236 S.n3228 0.002
R8200 S.n3226 S.n3012 0.002
R8201 S.n3746 S.n3738 0.002
R8202 S.n3736 S.n3523 0.002
R8203 S.n4244 S.n4236 0.002
R8204 S.n4234 S.n4023 0.002
R8205 S.n4687 S.n4679 0.002
R8206 S.n4677 S.n4465 0.002
R8207 S.n4923 S.n4915 0.002
R8208 S.n5007 S.n4999 0.002
R8209 S.n5630 S.n5622 0.002
R8210 S.n5460 S.n5452 0.002
R8211 S.n478 S.n477 0.002
R8212 S.n230 S.n222 0.002
R8213 S.n1179 S.n1158 0.002
R8214 S.n868 S.n858 0.002
R8215 S.n1767 S.n1750 0.002
R8216 S.n1410 S.n1402 0.002
R8217 S.n2328 S.n2311 0.002
R8218 S.n2003 S.n1995 0.002
R8219 S.n2883 S.n2866 0.002
R8220 S.n2530 S.n2522 0.002
R8221 S.n3411 S.n3394 0.002
R8222 S.n3047 S.n3039 0.002
R8223 S.n660 S.n659 0.002
R8224 S.n254 S.n238 0.002
R8225 S.n1117 S.n1102 0.002
R8226 S.n914 S.n897 0.002
R8227 S.n1705 S.n1680 0.002
R8228 S.n1455 S.n1437 0.002
R8229 S.n2268 S.n2243 0.002
R8230 S.n2047 S.n2029 0.002
R8231 S.n2818 S.n2793 0.002
R8232 S.n2574 S.n2556 0.002
R8233 S.n3346 S.n3321 0.002
R8234 S.n3091 S.n3073 0.002
R8235 S.n3864 S.n3836 0.002
R8236 S.n3585 S.n3566 0.002
R8237 S.n4364 S.n4336 0.002
R8238 S.n4065 S.n4046 0.002
R8239 S.n4506 S.n4495 0.002
R8240 S.n4400 S.n4392 0.002
R8241 S.n4087 S.n4076 0.002
R8242 S.n4329 S.n4321 0.002
R8243 S.n3605 S.n3594 0.002
R8244 S.n3829 S.n3821 0.002
R8245 S.n3111 S.n3100 0.002
R8246 S.n3314 S.n3306 0.002
R8247 S.n2594 S.n2583 0.002
R8248 S.n2786 S.n2778 0.002
R8249 S.n2067 S.n2056 0.002
R8250 S.n2236 S.n2228 0.002
R8251 S.n1475 S.n1464 0.002
R8252 S.n1673 S.n1665 0.002
R8253 S.n935 S.n921 0.002
R8254 S.n1084 S.n1068 0.002
R8255 S.n273 S.n262 0.002
R8256 S.n519 S.n518 0.002
R8257 S.n195 S.n187 0.002
R8258 S.n1238 S.n1216 0.002
R8259 S.n830 S.n822 0.002
R8260 S.n1832 S.n1815 0.002
R8261 S.n1373 S.n1365 0.002
R8262 S.n2392 S.n2375 0.002
R8263 S.n1967 S.n1959 0.002
R8264 S.n557 S.n556 0.002
R8265 S.n160 S.n151 0.002
R8266 S.n1301 S.n1284 0.002
R8267 S.n794 S.n786 0.002
R8268 S.n5683 S.n5675 0.002
R8269 S.n5416 S.n5405 0.002
R8270 S.n5812 S.n5811 0.002
R8271 S.n3776 S.n3761 0.002
R8272 S.n4458 S.n4440 0.002
R8273 S.n4904 S.n4896 0.002
R8274 S.n2733 S.n2718 0.002
R8275 S.n1620 S.n1605 0.002
R8276 S.n398 S.n397 0.002
R8277 S.n86 S.n85 0.002
R8278 S.n54 S.n53 0.002
R8279 S.n22 S.n21 0.002
R8280 S.n5407 S.n5406 0.002
R8281 S.n5429 S.n5428 0.002
R8282 S.n1110 S.n1109 0.002
R8283 S.n4429 S.n4428 0.002
R8284 S.n4876 S.n4875 0.002
R8285 S.n5652 S.n5651 0.002
R8286 S.n3375 S.n3374 0.002
R8287 S.n3893 S.n3892 0.002
R8288 S.n4266 S.n4265 0.002
R8289 S.n2356 S.n2355 0.002
R8290 S.n2912 S.n2911 0.002
R8291 S.n3255 S.n3254 0.002
R8292 S.n1861 S.n1860 0.002
R8293 S.n2178 S.n2177 0.002
R8294 S.n5252 S.n5251 0.002
R8295 S.n5108 S.n5107 0.002
R8296 S.n5285 S.n5284 0.002
R8297 S.n5573 S.n5572 0.002
R8298 S.n3939 S.n3932 0.002
R8299 S.n3454 S.n3447 0.002
R8300 S.n2958 S.n2951 0.002
R8301 S.n2436 S.n2429 0.002
R8302 S.n1909 S.n1901 0.002
R8303 S.n1575 S.n1568 0.002
R8304 S.n1056 S.n1043 0.002
R8305 S.n1209 S.n1196 0.002
R8306 S.n1767 S.n1766 0.002
R8307 S.n1410 S.n1409 0.002
R8308 S.n2328 S.n2327 0.002
R8309 S.n2003 S.n2002 0.002
R8310 S.n2883 S.n2882 0.002
R8311 S.n2530 S.n2529 0.002
R8312 S.n3411 S.n3410 0.002
R8313 S.n3047 S.n3046 0.002
R8314 S.n1268 S.n1255 0.002
R8315 S.n830 S.n829 0.002
R8316 S.n1832 S.n1831 0.002
R8317 S.n1373 S.n1372 0.002
R8318 S.n2392 S.n2391 0.002
R8319 S.n1967 S.n1966 0.002
R8320 S.n1301 S.n1300 0.002
R8321 S.n794 S.n793 0.002
R8322 S.n5437 S.n5436 0.002
R8323 S.n1685 S.n1684 0.002
R8324 S.n2248 S.n2247 0.002
R8325 S.n2798 S.n2797 0.002
R8326 S.n3326 S.n3325 0.002
R8327 S.n3841 S.n3840 0.002
R8328 S.n4341 S.n4340 0.002
R8329 S.n4445 S.n4444 0.002
R8330 S.n3760 S.n3759 0.002
R8331 S.n3393 S.n3392 0.002
R8332 S.n2865 S.n2864 0.002
R8333 S.n2717 S.n2716 0.002
R8334 S.n2374 S.n2373 0.002
R8335 S.n1814 S.n1813 0.002
R8336 S.n1604 S.n1603 0.002
R8337 S.n1283 S.n1282 0.002
R8338 S.n5557 S.n5549 0.002
R8339 S.n5300 S.n5293 0.002
R8340 S.n5087 S.n5079 0.002
R8341 S.n5232 S.n5225 0.002
R8342 S.n4636 S.n4628 0.002
R8343 S.n4217 S.n4216 0.002
R8344 S.n5541 S.n5533 0.002
R8345 S.n5315 S.n5308 0.002
R8346 S.n5071 S.n5063 0.002
R8347 S.n5217 S.n5210 0.002
R8348 S.n4620 S.n4612 0.002
R8349 S.n4779 S.n4772 0.002
R8350 S.n4201 S.n4193 0.002
R8351 S.n3719 S.n3718 0.002
R8352 S.n5525 S.n5517 0.002
R8353 S.n5330 S.n5323 0.002
R8354 S.n5055 S.n5047 0.002
R8355 S.n5202 S.n5195 0.002
R8356 S.n4604 S.n4596 0.002
R8357 S.n4764 S.n4757 0.002
R8358 S.n4185 S.n4177 0.002
R8359 S.n3954 S.n3947 0.002
R8360 S.n3703 S.n3695 0.002
R8361 S.n3209 S.n3208 0.002
R8362 S.n5509 S.n5501 0.002
R8363 S.n5345 S.n5338 0.002
R8364 S.n5039 S.n5031 0.002
R8365 S.n5187 S.n5180 0.002
R8366 S.n4588 S.n4580 0.002
R8367 S.n4749 S.n4742 0.002
R8368 S.n4169 S.n4161 0.002
R8369 S.n3969 S.n3962 0.002
R8370 S.n3687 S.n3679 0.002
R8371 S.n3469 S.n3462 0.002
R8372 S.n3193 S.n3185 0.002
R8373 S.n2676 S.n2675 0.002
R8374 S.n5493 S.n5485 0.002
R8375 S.n5360 S.n5353 0.002
R8376 S.n5023 S.n5015 0.002
R8377 S.n5172 S.n5165 0.002
R8378 S.n4572 S.n4564 0.002
R8379 S.n4734 S.n4727 0.002
R8380 S.n4153 S.n4145 0.002
R8381 S.n3984 S.n3977 0.002
R8382 S.n3671 S.n3663 0.002
R8383 S.n3484 S.n3477 0.002
R8384 S.n3177 S.n3169 0.002
R8385 S.n2973 S.n2966 0.002
R8386 S.n2660 S.n2652 0.002
R8387 S.n2133 S.n2132 0.002
R8388 S.n5589 S.n5376 0.002
R8389 S.n5592 S.n5368 0.002
R8390 S.n5155 S.n5142 0.002
R8391 S.n5157 S.n5134 0.002
R8392 S.n4556 S.n4549 0.002
R8393 S.n4719 S.n4711 0.002
R8394 S.n4137 S.n4130 0.002
R8395 S.n4000 S.n3992 0.002
R8396 S.n3655 S.n3648 0.002
R8397 S.n3500 S.n3492 0.002
R8398 S.n3161 S.n3154 0.002
R8399 S.n2989 S.n2981 0.002
R8400 S.n2644 S.n2637 0.002
R8401 S.n2452 S.n2444 0.002
R8402 S.n2117 S.n2110 0.002
R8403 S.n1545 S.n1544 0.002
R8404 S.n5477 S.n5468 0.002
R8405 S.n5611 S.n5600 0.002
R8406 S.n5124 S.n4939 0.002
R8407 S.n5126 S.n4931 0.002
R8408 S.n4541 S.n4534 0.002
R8409 S.n4703 S.n4695 0.002
R8410 S.n4122 S.n4115 0.002
R8411 S.n4016 S.n4008 0.002
R8412 S.n3640 S.n3633 0.002
R8413 S.n3516 S.n3508 0.002
R8414 S.n3146 S.n3139 0.002
R8415 S.n3005 S.n2997 0.002
R8416 S.n2629 S.n2622 0.002
R8417 S.n2468 S.n2460 0.002
R8418 S.n2102 S.n2095 0.002
R8419 S.n1925 S.n1917 0.002
R8420 S.n1528 S.n1520 0.002
R8421 S.n971 S.n970 0.002
R8422 S.n4976 S.n4965 0.002
R8423 S.n4879 S.n4864 0.002
R8424 S.n4525 S.n4514 0.002
R8425 S.n4432 S.n4417 0.002
R8426 S.n4106 S.n4095 0.002
R8427 S.n4305 S.n4290 0.002
R8428 S.n3624 S.n3613 0.002
R8429 S.n3809 S.n3794 0.002
R8430 S.n3130 S.n3119 0.002
R8431 S.n3294 S.n3279 0.002
R8432 S.n2613 S.n2602 0.002
R8433 S.n2766 S.n2751 0.002
R8434 S.n2086 S.n2075 0.002
R8435 S.n2216 S.n2202 0.002
R8436 S.n1495 S.n1483 0.002
R8437 S.n1653 S.n1638 0.002
R8438 S.n954 S.n943 0.002
R8439 S.n2511 S.n2500 0.002
R8440 S.n2915 S.n2900 0.002
R8441 S.n1986 S.n1975 0.002
R8442 S.n2359 S.n2345 0.002
R8443 S.n1393 S.n1381 0.002
R8444 S.n1799 S.n1784 0.002
R8445 S.n849 S.n838 0.002
R8446 S.n1179 S.n1178 0.002
R8447 S.n230 S.n229 0.002
R8448 S.n213 S.n212 0.002
R8449 S.n1354 S.n1342 0.002
R8450 S.n1864 S.n1849 0.002
R8451 S.n813 S.n802 0.002
R8452 S.n1238 S.n1237 0.002
R8453 S.n195 S.n194 0.002
R8454 S.n178 S.n177 0.002
R8455 S.n160 S.n159 0.002
R8456 S.n144 S.n143 0.002
R8457 S.n5416 S.n5404 0.002
R8458 S.n5683 S.n5682 0.002
R8459 S.n4990 S.n4989 0.002
R8460 S.n4811 S.n4810 0.002
R8461 S.n5108 S.n5099 0.002
R8462 S.n4660 S.n4648 0.002
R8463 S.n4814 S.n4813 0.002
R8464 S.n659 S.n644 0.002
R8465 S.n351 S.n350 0.002
R8466 S.n1316 S.n1315 0.002
R8467 S.n490 S.n489 0.002
R8468 S.t240 S.n5826 0.002
R8469 S.t240 S.n5841 0.002
R8470 S.n5658 S.n5640 0.002
R8471 S.n3261 S.n3244 0.002
R8472 S.n2184 S.n2168 0.002
R8473 S.n1025 S.n1010 0.002
R8474 S.n583 S.n582 0.002
R8475 S.n5630 S.n5629 0.002
R8476 S.n5007 S.n5006 0.002
R8477 S.n4923 S.n4922 0.002
R8478 S.n4677 S.n4676 0.002
R8479 S.n4687 S.n4686 0.002
R8480 S.n4234 S.n4233 0.002
R8481 S.n4244 S.n4243 0.002
R8482 S.n3736 S.n3735 0.002
R8483 S.n3746 S.n3745 0.002
R8484 S.n3226 S.n3225 0.002
R8485 S.n3236 S.n3235 0.002
R8486 S.n2693 S.n2692 0.002
R8487 S.n2703 S.n2702 0.002
R8488 S.n2150 S.n2149 0.002
R8489 S.n2160 S.n2159 0.002
R8490 S.n1512 S.n1511 0.002
R8491 S.n1590 S.n1589 0.002
R8492 S.n988 S.n987 0.002
R8493 S.n4904 S.n4903 0.002
R8494 S.n4400 S.n4399 0.002
R8495 S.n4329 S.n4328 0.002
R8496 S.n3829 S.n3828 0.002
R8497 S.n3314 S.n3313 0.002
R8498 S.n2786 S.n2785 0.002
R8499 S.n2236 S.n2235 0.002
R8500 S.n1673 S.n1672 0.002
R8501 S.n5460 S.n5459 0.002
R8502 S.n5573 S.n5564 0.002
R8503 S.n4217 S.n4208 0.002
R8504 S.n4636 S.n4635 0.002
R8505 S.n5087 S.n5086 0.002
R8506 S.n5557 S.n5556 0.002
R8507 S.n3719 S.n3710 0.002
R8508 S.n4201 S.n4200 0.002
R8509 S.n4620 S.n4619 0.002
R8510 S.n5071 S.n5070 0.002
R8511 S.n5541 S.n5540 0.002
R8512 S.n3209 S.n3200 0.002
R8513 S.n3703 S.n3702 0.002
R8514 S.n4185 S.n4184 0.002
R8515 S.n4604 S.n4603 0.002
R8516 S.n5055 S.n5054 0.002
R8517 S.n5525 S.n5524 0.002
R8518 S.n2676 S.n2667 0.002
R8519 S.n3193 S.n3192 0.002
R8520 S.n3687 S.n3686 0.002
R8521 S.n4169 S.n4168 0.002
R8522 S.n4588 S.n4587 0.002
R8523 S.n5039 S.n5038 0.002
R8524 S.n5509 S.n5508 0.002
R8525 S.n2133 S.n2124 0.002
R8526 S.n2660 S.n2659 0.002
R8527 S.n3177 S.n3176 0.002
R8528 S.n3671 S.n3670 0.002
R8529 S.n4153 S.n4152 0.002
R8530 S.n4572 S.n4571 0.002
R8531 S.n5023 S.n5022 0.002
R8532 S.n5493 S.n5492 0.002
R8533 S.n1545 S.n1317 0.002
R8534 S.n5156 S.n5155 0.002
R8535 S.n5591 S.n5589 0.002
R8536 S.n971 S.n962 0.002
R8537 S.n1528 S.n1527 0.002
R8538 S.n5125 S.n5124 0.002
R8539 S.n5477 S.n5476 0.002
R8540 S.n5460 S.n5451 0.002
R8541 S.n5007 S.n4998 0.002
R8542 S.n4678 S.n4677 0.002
R8543 S.n4235 S.n4234 0.002
R8544 S.n3737 S.n3736 0.002
R8545 S.n3227 S.n3226 0.002
R8546 S.n2694 S.n2693 0.002
R8547 S.n2151 S.n2150 0.002
R8548 S.n1512 S.n1503 0.002
R8549 S.n989 S.n988 0.002
R8550 S.n293 S.n281 0.002
R8551 S.n4065 S.n4064 0.002
R8552 S.n3585 S.n3584 0.002
R8553 S.n3091 S.n3090 0.002
R8554 S.n2574 S.n2573 0.002
R8555 S.n2047 S.n2046 0.002
R8556 S.n1455 S.n1454 0.002
R8557 S.n914 S.n913 0.002
R8558 S.n254 S.n237 0.002
R8559 S.n5437 S.n5435 0.002
R8560 S.n5658 S.n5639 0.002
R8561 S.n4976 S.n4964 0.002
R8562 S.n4879 S.n4854 0.002
R8563 S.n4525 S.n4513 0.002
R8564 S.n4432 S.n4407 0.002
R8565 S.n4106 S.n4094 0.002
R8566 S.n4305 S.n4280 0.002
R8567 S.n3624 S.n3612 0.002
R8568 S.n3809 S.n3784 0.002
R8569 S.n3130 S.n3118 0.002
R8570 S.n3294 S.n3269 0.002
R8571 S.n2613 S.n2601 0.002
R8572 S.n2766 S.n2741 0.002
R8573 S.n2086 S.n2074 0.002
R8574 S.n2216 S.n2192 0.002
R8575 S.n1495 S.n1482 0.002
R8576 S.n1653 S.n1628 0.002
R8577 S.n954 S.n942 0.002
R8578 S.n1056 S.n1033 0.002
R8579 S.n377 S.n358 0.002
R8580 S.n401 S.n380 0.002
R8581 S.n4272 S.n4251 0.002
R8582 S.n3559 S.n3547 0.002
R8583 S.n3896 S.n3871 0.002
R8584 S.n3066 S.n3054 0.002
R8585 S.n3378 S.n3353 0.002
R8586 S.n2549 S.n2537 0.002
R8587 S.n2850 S.n2825 0.002
R8588 S.n2022 S.n2010 0.002
R8589 S.n2299 S.n2275 0.002
R8590 S.n1430 S.n1417 0.002
R8591 S.n1738 S.n1712 0.002
R8592 S.n890 S.n879 0.002
R8593 S.n1151 S.n1130 0.002
R8594 S.n325 S.n313 0.002
R8595 S.n310 S.n110 0.002
R8596 S.n3261 S.n3243 0.002
R8597 S.n2511 S.n2499 0.002
R8598 S.n2915 S.n2890 0.002
R8599 S.n1986 S.n1974 0.002
R8600 S.n2359 S.n2335 0.002
R8601 S.n1393 S.n1380 0.002
R8602 S.n1799 S.n1774 0.002
R8603 S.n849 S.n837 0.002
R8604 S.n1209 S.n1186 0.002
R8605 S.n213 S.n202 0.002
R8606 S.n103 S.n95 0.002
R8607 S.n2184 S.n2167 0.002
R8608 S.n1354 S.n1341 0.002
R8609 S.n1864 S.n1839 0.002
R8610 S.n813 S.n801 0.002
R8611 S.n1268 S.n1245 0.002
R8612 S.n178 S.n167 0.002
R8613 S.n71 S.n63 0.002
R8614 S.n1025 S.n1009 0.002
R8615 S.n144 S.n135 0.002
R8616 S.n39 S.n31 0.002
R8617 S.n5844 S.n5842 0.002
R8618 S.n730 S.n729 0.001
R8619 S.n1129 S.n1128 0.001
R8620 S.n1051 S.n1050 0.001
R8621 S.n1204 S.n1203 0.001
R8622 S.n584 S.n583 0.001
R8623 S.t191 S.n584 0.001
R8624 S.n4851 S.n4850 0.001
R8625 S.n3820 S.n3819 0.001
R8626 S.n3305 S.n3304 0.001
R8627 S.n2777 S.n2776 0.001
R8628 S.n2227 S.n2226 0.001
R8629 S.n1664 S.n1663 0.001
R8630 S.n1067 S.n1066 0.001
R8631 S.n5812 S.n5810 0.001
R8632 S.n5842 S.t240 0.001
R8633 S.n1738 S.n1723 0.001
R8634 S.n3775 S.n3774 0.001
R8635 S.n2732 S.n2731 0.001
R8636 S.n1619 S.n1618 0.001
R8637 S.n4973 S.n4972 0.001
R8638 S.n4522 S.n4521 0.001
R8639 S.n2508 S.n2507 0.001
R8640 S.n1983 S.n1982 0.001
R8641 S.n3556 S.n3555 0.001
R8642 S.n3063 S.n3062 0.001
R8643 S.n1351 S.n1350 0.001
R8644 S.n810 S.n809 0.001
R8645 S.n429 S.n428 0.001
R8646 S.n5807 S.n5806 0.001
R8647 S.n5809 S.n5808 0.001
R8648 S.n457 S.n456 0.001
R8649 S.n124 S.n123 0.001
R8650 S.n748 S.n747 0.001
R8651 S.n771 S.n770 0.001
R8652 S.n1557 S.n1556 0.001
R8653 S.n1331 S.n1330 0.001
R8654 S.n1890 S.n1889 0.001
R8655 S.n1944 S.n1943 0.001
R8656 S.n2418 S.n2417 0.001
R8657 S.n2489 S.n2488 0.001
R8658 S.n2940 S.n2939 0.001
R8659 S.n3024 S.n3023 0.001
R8660 S.n3436 S.n3435 0.001
R8661 S.n3537 S.n3536 0.001
R8662 S.n3921 S.n3920 0.001
R8663 S.n4035 S.n4034 0.001
R8664 S.n4827 S.n4826 0.001
R8665 S.n4481 S.n4480 0.001
R8666 S.n4845 S.n4844 0.001
R8667 S.n4953 S.n4952 0.001
R8668 S.n5699 S.n5698 0.001
R8669 S.n5393 S.n5391 0.001
R8670 S.n5714 S.n5713 0.001
R8671 S.n951 S.n950 0.001
R8672 S.n1650 S.n1649 0.001
R8673 S.n1492 S.n1491 0.001
R8674 S.n2213 S.n2212 0.001
R8675 S.n2083 S.n2082 0.001
R8676 S.n2763 S.n2762 0.001
R8677 S.n2610 S.n2609 0.001
R8678 S.n3291 S.n3290 0.001
R8679 S.n3127 S.n3126 0.001
R8680 S.n3806 S.n3805 0.001
R8681 S.n3621 S.n3620 0.001
R8682 S.n4302 S.n4301 0.001
R8683 S.n4103 S.n4102 0.001
R8684 S.n878 S.n877 0.001
R8685 S.n1735 S.n1734 0.001
R8686 S.n1427 S.n1426 0.001
R8687 S.n2296 S.n2295 0.001
R8688 S.n2019 S.n2018 0.001
R8689 S.n2847 S.n2846 0.001
R8690 S.n2546 S.n2545 0.001
R8691 S.n846 S.n845 0.001
R8692 S.n1796 S.n1795 0.001
R8693 S.n1390 S.n1389 0.001
R8694 S.n5668 S.n5667 0.001
R8695 S.n2310 S.n2309 0.001
R8696 S.n1749 S.n1748 0.001
R8697 S.n1163 S.n1162 0.001
R8698 S.n1221 S.n1220 0.001
R8699 S.n1546 S.n1545 0.001
R8700 S.n971 S.n963 0.001
R8701 S.n293 S.n282 0.001
R8702 S.n731 S.n730 0.001
R8703 S.t191 S.n479 0.001
R8704 S.t191 S.n631 0.001
R8705 S.t191 S.n661 0.001
R8706 S.t191 S.n520 0.001
R8707 S.t191 S.n558 0.001
R8708 S.t191 S.n691 0.001
R8709 S.t191 S.n617 0.001
R8710 S.t191 S.n605 0.001
R8711 S.t191 S.n593 0.001
R8712 S.t191 S.n570 0.001
R8713 S.n3896 S.n3881 0.001
R8714 S.n3378 S.n3363 0.001
R8715 S.n2850 S.n2835 0.001
R8716 S.n2299 S.n2285 0.001
R8717 S.n5399 S.n5398 0.001
R8718 S.n3030 S.n3029 0.001
R8719 S.n4041 S.n4040 0.001
R8720 S.n4486 S.n4485 0.001
R8721 S.n4959 S.n4958 0.001
R8722 S.n3542 S.n3541 0.001
R8723 S.n1950 S.n1949 0.001
R8724 S.n2494 S.n2493 0.001
R8725 S.n777 S.n776 0.001
R8726 S.n1336 S.n1335 0.001
R8727 S.n130 S.n129 0.001
R8728 S.n5709 S.n5692 0.001
R8729 S.n490 S.n488 0.001
R8730 S.n388 S.n387 0.001
R8731 S.n4272 S.n4253 0.001
R8732 S.n91 S.n90 0.001
R8733 S.n60 S.n59 0.001
R8734 S.n28 S.n27 0.001
R8735 S.n5433 S.n5432 0.001
R8736 S.n5445 S.n5442 0.001
R8737 S.t52 S.n5445 0.001
R8738 S.n5692 S.t34 0.001
R8739 S.t52 S.n5399 0.001
R8740 S.t27 S.n3030 0.001
R8741 S.t6 S.n3542 0.001
R8742 S.t65 S.n4041 0.001
R8743 S.t4 S.n4486 0.001
R8744 S.t45 S.n4959 0.001
R8745 S.t56 S.n1950 0.001
R8746 S.t68 S.n2494 0.001
R8747 S.t14 S.n777 0.001
R8748 S.t32 S.n1336 0.001
R8749 S.t213 S.n130 0.001
R8750 S.n490 S.n487 0.001
R8751 S.n2407 S.n2406 0.001
R8752 S.n1879 S.n1878 0.001
R8753 S.n378 S.n377 0.001
R8754 S.n311 S.n310 0.001
R8755 S.n490 S.n484 0.001
R8756 S.n490 S.n483 0.001
R8757 S.n490 S.n482 0.001
R8758 S.n490 S.n486 0.001
R8759 S.n458 S.n457 0.001
R8760 S.n123 S.n122 0.001
R8761 S.n749 S.n748 0.001
R8762 S.n770 S.n769 0.001
R8763 S.n1558 S.n1557 0.001
R8764 S.n1330 S.n1329 0.001
R8765 S.n1891 S.n1890 0.001
R8766 S.n1943 S.n1942 0.001
R8767 S.n2419 S.n2418 0.001
R8768 S.n2488 S.n2487 0.001
R8769 S.n2941 S.n2940 0.001
R8770 S.n3023 S.n3022 0.001
R8771 S.n3437 S.n3436 0.001
R8772 S.n3536 S.n3535 0.001
R8773 S.n3922 S.n3921 0.001
R8774 S.n4034 S.n4033 0.001
R8775 S.n4828 S.n4827 0.001
R8776 S.n4480 S.n4479 0.001
R8777 S.n4846 S.n4845 0.001
R8778 S.n4952 S.n4951 0.001
R8779 S.n5700 S.n5699 0.001
R8780 S.n5391 S.n5390 0.001
R8781 S.n5715 S.n5714 0.001
R8782 S.n5812 S.n5809 0.001
R8783 S.n5812 S.n5807 0.001
R8784 S.n213 S.n205 0.001
R8785 S.n178 S.n170 0.001
R8786 S.n144 S.n136 0.001
R8787 S.n4212 S.n4211 0.001
R8788 S.n4794 S.n4793 0.001
R8789 S.n5555 S.n5554 0.001
R8790 S.n5299 S.n5298 0.001
R8791 S.n5085 S.n5084 0.001
R8792 S.n5231 S.n5230 0.001
R8793 S.n4634 S.n4633 0.001
R8794 S.n5568 S.n5567 0.001
R8795 S.n5280 S.n5279 0.001
R8796 S.n5103 S.n5102 0.001
R8797 S.n5246 S.n5245 0.001
R8798 S.n4652 S.n4651 0.001
R8799 S.n3714 S.n3713 0.001
R8800 S.n3938 S.n3937 0.001
R8801 S.n5539 S.n5538 0.001
R8802 S.n5314 S.n5313 0.001
R8803 S.n5069 S.n5068 0.001
R8804 S.n5216 S.n5215 0.001
R8805 S.n4618 S.n4617 0.001
R8806 S.n4778 S.n4777 0.001
R8807 S.n4199 S.n4198 0.001
R8808 S.n3204 S.n3203 0.001
R8809 S.n3453 S.n3452 0.001
R8810 S.n5523 S.n5522 0.001
R8811 S.n5329 S.n5328 0.001
R8812 S.n5053 S.n5052 0.001
R8813 S.n5201 S.n5200 0.001
R8814 S.n4602 S.n4601 0.001
R8815 S.n4763 S.n4762 0.001
R8816 S.n4183 S.n4182 0.001
R8817 S.n3953 S.n3952 0.001
R8818 S.n3701 S.n3700 0.001
R8819 S.n2671 S.n2670 0.001
R8820 S.n2957 S.n2956 0.001
R8821 S.n5507 S.n5506 0.001
R8822 S.n5344 S.n5343 0.001
R8823 S.n5037 S.n5036 0.001
R8824 S.n5186 S.n5185 0.001
R8825 S.n4586 S.n4585 0.001
R8826 S.n4748 S.n4747 0.001
R8827 S.n4167 S.n4166 0.001
R8828 S.n3968 S.n3967 0.001
R8829 S.n3685 S.n3684 0.001
R8830 S.n3468 S.n3467 0.001
R8831 S.n3191 S.n3190 0.001
R8832 S.n2128 S.n2127 0.001
R8833 S.n2435 S.n2434 0.001
R8834 S.n5491 S.n5490 0.001
R8835 S.n5359 S.n5358 0.001
R8836 S.n5021 S.n5020 0.001
R8837 S.n5171 S.n5170 0.001
R8838 S.n4570 S.n4569 0.001
R8839 S.n4733 S.n4732 0.001
R8840 S.n4151 S.n4150 0.001
R8841 S.n3983 S.n3982 0.001
R8842 S.n3669 S.n3668 0.001
R8843 S.n3483 S.n3482 0.001
R8844 S.n3175 S.n3174 0.001
R8845 S.n2972 S.n2971 0.001
R8846 S.n2658 S.n2657 0.001
R8847 S.n1320 S.n1319 0.001
R8848 S.n1907 S.n1906 0.001
R8849 S.n5588 S.n5587 0.001
R8850 S.n5374 S.n5373 0.001
R8851 S.n5154 S.n5153 0.001
R8852 S.n5140 S.n5139 0.001
R8853 S.n4555 S.n4554 0.001
R8854 S.n4717 S.n4716 0.001
R8855 S.n4136 S.n4135 0.001
R8856 S.n3998 S.n3997 0.001
R8857 S.n3654 S.n3653 0.001
R8858 S.n3498 S.n3497 0.001
R8859 S.n3160 S.n3159 0.001
R8860 S.n2987 S.n2986 0.001
R8861 S.n2643 S.n2642 0.001
R8862 S.n2450 S.n2449 0.001
R8863 S.n2116 S.n2115 0.001
R8864 S.n966 S.n965 0.001
R8865 S.n1574 S.n1573 0.001
R8866 S.n5474 S.n5473 0.001
R8867 S.n5606 S.n5605 0.001
R8868 S.n5123 S.n5122 0.001
R8869 S.n4937 S.n4936 0.001
R8870 S.n4540 S.n4539 0.001
R8871 S.n4701 S.n4700 0.001
R8872 S.n4121 S.n4120 0.001
R8873 S.n4014 S.n4013 0.001
R8874 S.n3639 S.n3638 0.001
R8875 S.n3514 S.n3513 0.001
R8876 S.n3145 S.n3144 0.001
R8877 S.n3003 S.n3002 0.001
R8878 S.n2628 S.n2627 0.001
R8879 S.n2466 S.n2465 0.001
R8880 S.n2101 S.n2100 0.001
R8881 S.n1923 S.n1922 0.001
R8882 S.n1526 S.n1525 0.001
R8883 S.n383 S.n382 0.001
R8884 S.n1049 S.n1048 0.001
R8885 S.n5646 S.n5645 0.001
R8886 S.n4971 S.n4970 0.001
R8887 S.n4870 S.n4869 0.001
R8888 S.n4520 S.n4519 0.001
R8889 S.n4423 S.n4422 0.001
R8890 S.n4101 S.n4100 0.001
R8891 S.n4296 S.n4295 0.001
R8892 S.n3619 S.n3618 0.001
R8893 S.n3800 S.n3799 0.001
R8894 S.n3125 S.n3124 0.001
R8895 S.n3285 S.n3284 0.001
R8896 S.n2608 S.n2607 0.001
R8897 S.n2757 S.n2756 0.001
R8898 S.n2081 S.n2080 0.001
R8899 S.n2208 S.n2207 0.001
R8900 S.n1489 S.n1488 0.001
R8901 S.n1644 S.n1643 0.001
R8902 S.n949 S.n948 0.001
R8903 S.n361 S.n360 0.001
R8904 S.n285 S.n284 0.001
R8905 S.n5455 S.n5454 0.001
R8906 S.n5625 S.n5624 0.001
R8907 S.n5002 S.n5001 0.001
R8908 S.n4918 S.n4917 0.001
R8909 S.n4468 S.n4467 0.001
R8910 S.n4682 S.n4681 0.001
R8911 S.n4026 S.n4025 0.001
R8912 S.n4239 S.n4238 0.001
R8913 S.n3526 S.n3525 0.001
R8914 S.n3741 S.n3740 0.001
R8915 S.n3015 S.n3014 0.001
R8916 S.n3231 S.n3230 0.001
R8917 S.n2478 S.n2477 0.001
R8918 S.n2698 S.n2697 0.001
R8919 S.n1935 S.n1934 0.001
R8920 S.n2155 S.n2154 0.001
R8921 S.n1507 S.n1506 0.001
R8922 S.n1585 S.n1584 0.001
R8923 S.n762 S.n761 0.001
R8924 S.n993 S.n992 0.001
R8925 S.n98 S.n97 0.001
R8926 S.n1202 S.n1201 0.001
R8927 S.n3250 S.n3249 0.001
R8928 S.n2506 S.n2505 0.001
R8929 S.n2906 S.n2905 0.001
R8930 S.n1981 S.n1980 0.001
R8931 S.n2351 S.n2350 0.001
R8932 S.n1387 S.n1386 0.001
R8933 S.n1790 S.n1789 0.001
R8934 S.n844 S.n843 0.001
R8935 S.n13 S.n12 0.001
R8936 S.n3764 S.n3763 0.001
R8937 S.n3042 S.n3041 0.001
R8938 S.n3397 S.n3396 0.001
R8939 S.n2525 S.n2524 0.001
R8940 S.n2869 S.n2868 0.001
R8941 S.n1998 S.n1997 0.001
R8942 S.n2314 S.n2313 0.001
R8943 S.n1405 S.n1404 0.001
R8944 S.n1753 S.n1752 0.001
R8945 S.n861 S.n860 0.001
R8946 S.n882 S.n881 0.001
R8947 S.n1133 S.n1132 0.001
R8948 S.n113 S.n112 0.001
R8949 S.n316 S.n315 0.001
R8950 S.n1729 S.n1728 0.001
R8951 S.n2291 S.n2290 0.001
R8952 S.n2841 S.n2840 0.001
R8953 S.n3369 S.n3368 0.001
R8954 S.n3887 S.n3886 0.001
R8955 S.n4261 S.n4260 0.001
R8956 S.n3554 S.n3553 0.001
R8957 S.n3061 S.n3060 0.001
R8958 S.n2544 S.n2543 0.001
R8959 S.n2017 S.n2016 0.001
R8960 S.n1424 S.n1423 0.001
R8961 S.n1105 S.n1104 0.001
R8962 S.n241 S.n240 0.001
R8963 S.n647 S.n646 0.001
R8964 S.n4453 S.n4452 0.001
R8965 S.n4062 S.n4061 0.001
R8966 S.n4349 S.n4348 0.001
R8967 S.n3582 S.n3581 0.001
R8968 S.n3849 S.n3848 0.001
R8969 S.n3089 S.n3088 0.001
R8970 S.n3334 S.n3333 0.001
R8971 S.n2572 S.n2571 0.001
R8972 S.n2806 S.n2805 0.001
R8973 S.n2045 S.n2044 0.001
R8974 S.n2256 S.n2255 0.001
R8975 S.n1453 S.n1452 0.001
R8976 S.n1693 S.n1692 0.001
R8977 S.n912 S.n911 0.001
R8978 S.n1071 S.n1070 0.001
R8979 S.n265 S.n264 0.001
R8980 S.n932 S.n931 0.001
R8981 S.n1668 S.n1667 0.001
R8982 S.n1467 S.n1466 0.001
R8983 S.n2231 S.n2230 0.001
R8984 S.n2059 S.n2058 0.001
R8985 S.n2781 S.n2780 0.001
R8986 S.n2586 S.n2585 0.001
R8987 S.n3309 S.n3308 0.001
R8988 S.n3103 S.n3102 0.001
R8989 S.n3824 S.n3823 0.001
R8990 S.n3597 S.n3596 0.001
R8991 S.n4324 S.n4323 0.001
R8992 S.n4079 S.n4078 0.001
R8993 S.n4395 S.n4394 0.001
R8994 S.n4498 S.n4497 0.001
R8995 S.n4899 S.n4898 0.001
R8996 S.n340 S.n339 0.001
R8997 S.n1166 S.n1165 0.001
R8998 S.n225 S.n224 0.001
R8999 S.n208 S.n207 0.001
R9000 S.n66 S.n65 0.001
R9001 S.n1261 S.n1260 0.001
R9002 S.n2174 S.n2173 0.001
R9003 S.n1348 S.n1347 0.001
R9004 S.n1855 S.n1854 0.001
R9005 S.n808 S.n807 0.001
R9006 S.n507 S.n506 0.001
R9007 S.n2721 S.n2720 0.001
R9008 S.n1962 S.n1961 0.001
R9009 S.n2378 S.n2377 0.001
R9010 S.n1368 S.n1367 0.001
R9011 S.n1818 S.n1817 0.001
R9012 S.n825 S.n824 0.001
R9013 S.n1224 S.n1223 0.001
R9014 S.n190 S.n189 0.001
R9015 S.n173 S.n172 0.001
R9016 S.n34 S.n33 0.001
R9017 S.n1016 S.n1015 0.001
R9018 S.n545 S.n544 0.001
R9019 S.n1608 S.n1607 0.001
R9020 S.n789 S.n788 0.001
R9021 S.n1287 S.n1286 0.001
R9022 S.n155 S.n154 0.001
R9023 S.n139 S.n138 0.001
R9024 S.n422 S.n421 0.001
R9025 S.n5678 S.n5677 0.001
R9026 S.n4985 S.n4984 0.001
R9027 S.n491 S.n490 0.001
R9028 S.n490 S.n485 0.001
R9029 S.n5396 S.n5395 0.001
R9030 S.n4955 S.n4954 0.001
R9031 S.n4483 S.n4482 0.001
R9032 S.n4037 S.n4036 0.001
R9033 S.n3539 S.n3538 0.001
R9034 S.n3026 S.n3025 0.001
R9035 S.n2491 S.n2490 0.001
R9036 S.n1946 S.n1945 0.001
R9037 S.n1333 S.n1332 0.001
R9038 S.n773 S.n772 0.001
R9039 S.n126 S.n125 0.001
R9040 S.n4373 S.t77 0.001
R9041 S.t65 S.n4220 0.001
R9042 S.t65 S.n4223 0.001
R9043 S.t20 S.n4798 0.001
R9044 S.t20 S.n4801 0.001
R9045 S.t52 S.n5560 0.001
R9046 S.t52 S.n5563 0.001
R9047 S.t34 S.n5306 0.001
R9048 S.t34 S.n5303 0.001
R9049 S.n5303 S.n5300 0.001
R9050 S.t45 S.n5090 0.001
R9051 S.t45 S.n5093 0.001
R9052 S.t36 S.n5235 0.001
R9053 S.t36 S.n5238 0.001
R9054 S.t4 S.n4639 0.001
R9055 S.t4 S.n4642 0.001
R9056 S.n4804 S.t20 0.001
R9057 S.n4834 S.n4806 0.001
R9058 S.t52 S.n5576 0.001
R9059 S.t52 S.n5579 0.001
R9060 S.t34 S.n5291 0.001
R9061 S.t34 S.n5288 0.001
R9062 S.n5288 S.n5285 0.001
R9063 S.t45 S.n5111 0.001
R9064 S.t45 S.n5114 0.001
R9065 S.t36 S.n5255 0.001
R9066 S.t36 S.n5258 0.001
R9067 S.t4 S.n4663 0.001
R9068 S.t4 S.n4666 0.001
R9069 S.n4378 S.n4373 0.001
R9070 S.n3905 S.t200 0.001
R9071 S.t6 S.n3722 0.001
R9072 S.t6 S.n3725 0.001
R9073 S.t77 S.n3945 0.001
R9074 S.t77 S.n3942 0.001
R9075 S.n3942 S.n3939 0.001
R9076 S.t52 S.n5544 0.001
R9077 S.t52 S.n5547 0.001
R9078 S.t34 S.n5321 0.001
R9079 S.t34 S.n5318 0.001
R9080 S.n5318 S.n5315 0.001
R9081 S.t45 S.n5074 0.001
R9082 S.t45 S.n5077 0.001
R9083 S.t36 S.n5220 0.001
R9084 S.t36 S.n5223 0.001
R9085 S.t4 S.n4623 0.001
R9086 S.t4 S.n4626 0.001
R9087 S.t20 S.n4782 0.001
R9088 S.t20 S.n4785 0.001
R9089 S.t65 S.n4204 0.001
R9090 S.t65 S.n4207 0.001
R9091 S.n3910 S.n3905 0.001
R9092 S.n3420 S.t30 0.001
R9093 S.t27 S.n3212 0.001
R9094 S.t27 S.n3215 0.001
R9095 S.t200 S.n3460 0.001
R9096 S.t200 S.n3457 0.001
R9097 S.n3457 S.n3454 0.001
R9098 S.t52 S.n5528 0.001
R9099 S.t52 S.n5531 0.001
R9100 S.t34 S.n5336 0.001
R9101 S.t34 S.n5333 0.001
R9102 S.n5333 S.n5330 0.001
R9103 S.t45 S.n5058 0.001
R9104 S.t45 S.n5061 0.001
R9105 S.t36 S.n5205 0.001
R9106 S.t36 S.n5208 0.001
R9107 S.t4 S.n4607 0.001
R9108 S.t4 S.n4610 0.001
R9109 S.t20 S.n4767 0.001
R9110 S.t20 S.n4770 0.001
R9111 S.t65 S.n4188 0.001
R9112 S.t65 S.n4191 0.001
R9113 S.t77 S.n3960 0.001
R9114 S.t77 S.n3957 0.001
R9115 S.n3957 S.n3954 0.001
R9116 S.t6 S.n3706 0.001
R9117 S.t6 S.n3709 0.001
R9118 S.n3425 S.n3420 0.001
R9119 S.n2924 S.t256 0.001
R9120 S.t68 S.n2679 0.001
R9121 S.t68 S.n2682 0.001
R9122 S.t30 S.n2964 0.001
R9123 S.t30 S.n2961 0.001
R9124 S.n2961 S.n2958 0.001
R9125 S.t52 S.n5512 0.001
R9126 S.t52 S.n5515 0.001
R9127 S.t34 S.n5351 0.001
R9128 S.t34 S.n5348 0.001
R9129 S.n5348 S.n5345 0.001
R9130 S.t45 S.n5042 0.001
R9131 S.t45 S.n5045 0.001
R9132 S.t36 S.n5190 0.001
R9133 S.t36 S.n5193 0.001
R9134 S.t4 S.n4591 0.001
R9135 S.t4 S.n4594 0.001
R9136 S.t20 S.n4752 0.001
R9137 S.t20 S.n4755 0.001
R9138 S.t65 S.n4172 0.001
R9139 S.t65 S.n4175 0.001
R9140 S.t77 S.n3975 0.001
R9141 S.t77 S.n3972 0.001
R9142 S.n3972 S.n3969 0.001
R9143 S.t6 S.n3690 0.001
R9144 S.t6 S.n3693 0.001
R9145 S.t200 S.n3475 0.001
R9146 S.t200 S.n3472 0.001
R9147 S.n3472 S.n3469 0.001
R9148 S.t27 S.n3196 0.001
R9149 S.t27 S.n3199 0.001
R9150 S.n2929 S.n2924 0.001
R9151 S.n2401 S.t290 0.001
R9152 S.t56 S.n2136 0.001
R9153 S.t56 S.n2139 0.001
R9154 S.t256 S.n2442 0.001
R9155 S.t256 S.n2439 0.001
R9156 S.n2439 S.n2436 0.001
R9157 S.t52 S.n5496 0.001
R9158 S.t52 S.n5499 0.001
R9159 S.t34 S.n5366 0.001
R9160 S.t34 S.n5363 0.001
R9161 S.n5363 S.n5360 0.001
R9162 S.t45 S.n5026 0.001
R9163 S.t45 S.n5029 0.001
R9164 S.t36 S.n5175 0.001
R9165 S.t36 S.n5178 0.001
R9166 S.t4 S.n4575 0.001
R9167 S.t4 S.n4578 0.001
R9168 S.t20 S.n4737 0.001
R9169 S.t20 S.n4740 0.001
R9170 S.t65 S.n4156 0.001
R9171 S.t65 S.n4159 0.001
R9172 S.t77 S.n3990 0.001
R9173 S.t77 S.n3987 0.001
R9174 S.n3987 S.n3984 0.001
R9175 S.t6 S.n3674 0.001
R9176 S.t6 S.n3677 0.001
R9177 S.t200 S.n3490 0.001
R9178 S.t200 S.n3487 0.001
R9179 S.n3487 S.n3484 0.001
R9180 S.t27 S.n3180 0.001
R9181 S.t27 S.n3183 0.001
R9182 S.t30 S.n2979 0.001
R9183 S.t30 S.n2976 0.001
R9184 S.n2976 S.n2973 0.001
R9185 S.t68 S.n2663 0.001
R9186 S.t68 S.n2666 0.001
R9187 S.n2406 S.n2401 0.001
R9188 S.n1873 S.t18 0.001
R9189 S.n1537 S.t32 0.001
R9190 S.n1545 S.n1540 0.001
R9191 S.t290 S.n1915 0.001
R9192 S.t290 S.n1912 0.001
R9193 S.n1912 S.n1909 0.001
R9194 S.n5582 S.t52 0.001
R9195 S.n5589 S.n5582 0.001
R9196 S.t34 S.n5598 0.001
R9197 S.t34 S.n5595 0.001
R9198 S.n5595 S.n5592 0.001
R9199 S.n5155 S.n5148 0.001
R9200 S.t36 S.n5160 0.001
R9201 S.t36 S.n5163 0.001
R9202 S.t4 S.n4559 0.001
R9203 S.t4 S.n4562 0.001
R9204 S.t20 S.n4722 0.001
R9205 S.t20 S.n4725 0.001
R9206 S.t65 S.n4140 0.001
R9207 S.t65 S.n4143 0.001
R9208 S.t77 S.n4006 0.001
R9209 S.t77 S.n4003 0.001
R9210 S.n4003 S.n4000 0.001
R9211 S.t6 S.n3658 0.001
R9212 S.t6 S.n3661 0.001
R9213 S.t200 S.n3506 0.001
R9214 S.t200 S.n3503 0.001
R9215 S.n3503 S.n3500 0.001
R9216 S.t27 S.n3164 0.001
R9217 S.t27 S.n3167 0.001
R9218 S.t30 S.n2995 0.001
R9219 S.t30 S.n2992 0.001
R9220 S.n2992 S.n2989 0.001
R9221 S.t68 S.n2647 0.001
R9222 S.t68 S.n2650 0.001
R9223 S.t256 S.n2458 0.001
R9224 S.t256 S.n2455 0.001
R9225 S.n2455 S.n2452 0.001
R9226 S.t56 S.n2120 0.001
R9227 S.t56 S.n2123 0.001
R9228 S.n1878 S.n1873 0.001
R9229 S.n1310 S.t58 0.001
R9230 S.t14 S.n974 0.001
R9231 S.t14 S.n977 0.001
R9232 S.t18 S.n1581 0.001
R9233 S.t18 S.n1578 0.001
R9234 S.n1578 S.n1575 0.001
R9235 S.t52 S.n5480 0.001
R9236 S.t52 S.n5483 0.001
R9237 S.t34 S.n5617 0.001
R9238 S.t34 S.n5614 0.001
R9239 S.n5614 S.n5611 0.001
R9240 S.n5117 S.t45 0.001
R9241 S.n5124 S.n5117 0.001
R9242 S.t36 S.n5129 0.001
R9243 S.t36 S.n5132 0.001
R9244 S.t4 S.n4544 0.001
R9245 S.t4 S.n4547 0.001
R9246 S.t20 S.n4706 0.001
R9247 S.t20 S.n4709 0.001
R9248 S.t65 S.n4125 0.001
R9249 S.t65 S.n4128 0.001
R9250 S.t77 S.n4022 0.001
R9251 S.t77 S.n4019 0.001
R9252 S.n4019 S.n4016 0.001
R9253 S.t6 S.n3643 0.001
R9254 S.t6 S.n3646 0.001
R9255 S.t200 S.n3522 0.001
R9256 S.t200 S.n3519 0.001
R9257 S.n3519 S.n3516 0.001
R9258 S.t27 S.n3149 0.001
R9259 S.t27 S.n3152 0.001
R9260 S.t30 S.n3011 0.001
R9261 S.t30 S.n3008 0.001
R9262 S.n3008 S.n3005 0.001
R9263 S.t68 S.n2632 0.001
R9264 S.t68 S.n2635 0.001
R9265 S.t256 S.n2474 0.001
R9266 S.t256 S.n2471 0.001
R9267 S.n2471 S.n2468 0.001
R9268 S.t56 S.n2105 0.001
R9269 S.t56 S.n2108 0.001
R9270 S.t290 S.n1931 0.001
R9271 S.t290 S.n1928 0.001
R9272 S.n1928 S.n1925 0.001
R9273 S.t32 S.n1531 0.001
R9274 S.t32 S.n1534 0.001
R9275 S.n1315 S.n1310 0.001
R9276 S.n730 S.n720 0.001
R9277 S.t151 S.n407 0.001
R9278 S.t151 S.n404 0.001
R9279 S.n404 S.n401 0.001
R9280 S.t58 S.n1059 0.001
R9281 S.t58 S.n1062 0.001
R9282 S.t34 S.n5664 0.001
R9283 S.t34 S.n5661 0.001
R9284 S.n5661 S.n5658 0.001
R9285 S.t45 S.n4982 0.001
R9286 S.t45 S.n4979 0.001
R9287 S.n4979 S.n4976 0.001
R9288 S.t36 S.n4885 0.001
R9289 S.t36 S.n4882 0.001
R9290 S.n4882 S.n4879 0.001
R9291 S.t4 S.n4531 0.001
R9292 S.t4 S.n4528 0.001
R9293 S.n4528 S.n4525 0.001
R9294 S.t20 S.n4438 0.001
R9295 S.t20 S.n4435 0.001
R9296 S.n4435 S.n4432 0.001
R9297 S.t65 S.n4112 0.001
R9298 S.t65 S.n4109 0.001
R9299 S.n4109 S.n4106 0.001
R9300 S.t77 S.n4308 0.001
R9301 S.t77 S.n4311 0.001
R9302 S.t6 S.n3630 0.001
R9303 S.t6 S.n3627 0.001
R9304 S.n3627 S.n3624 0.001
R9305 S.t200 S.n3812 0.001
R9306 S.t200 S.n3815 0.001
R9307 S.t27 S.n3136 0.001
R9308 S.t27 S.n3133 0.001
R9309 S.n3133 S.n3130 0.001
R9310 S.t30 S.n3297 0.001
R9311 S.t30 S.n3300 0.001
R9312 S.t68 S.n2619 0.001
R9313 S.t68 S.n2616 0.001
R9314 S.n2616 S.n2613 0.001
R9315 S.t256 S.n2769 0.001
R9316 S.t256 S.n2772 0.001
R9317 S.t56 S.n2092 0.001
R9318 S.t56 S.n2089 0.001
R9319 S.n2089 S.n2086 0.001
R9320 S.t290 S.n2219 0.001
R9321 S.t290 S.n2222 0.001
R9322 S.t32 S.n1501 0.001
R9323 S.t32 S.n1498 0.001
R9324 S.n1498 S.n1495 0.001
R9325 S.t18 S.n1656 0.001
R9326 S.t18 S.n1659 0.001
R9327 S.t14 S.n960 0.001
R9328 S.t14 S.n957 0.001
R9329 S.n957 S.n954 0.001
R9330 S.n377 S.n367 0.001
R9331 S.t213 S.n296 0.001
R9332 S.t213 S.n299 0.001
R9333 S.t151 S.n466 0.001
R9334 S.n463 S.n441 0.001
R9335 S.t52 S.n5463 0.001
R9336 S.t52 S.n5466 0.001
R9337 S.t34 S.n5636 0.001
R9338 S.t34 S.n5633 0.001
R9339 S.n5633 S.n5630 0.001
R9340 S.t45 S.n5010 0.001
R9341 S.t45 S.n5013 0.001
R9342 S.t36 S.n4926 0.001
R9343 S.t36 S.n4929 0.001
R9344 S.n4669 S.t4 0.001
R9345 S.n4677 S.n4672 0.001
R9346 S.t20 S.n4690 0.001
R9347 S.t20 S.n4693 0.001
R9348 S.n4226 S.t65 0.001
R9349 S.n4234 S.n4229 0.001
R9350 S.t77 S.n4250 0.001
R9351 S.t77 S.n4247 0.001
R9352 S.n4247 S.n4244 0.001
R9353 S.n3728 S.t6 0.001
R9354 S.n3736 S.n3731 0.001
R9355 S.t200 S.n3752 0.001
R9356 S.t200 S.n3749 0.001
R9357 S.n3749 S.n3746 0.001
R9358 S.n3218 S.t27 0.001
R9359 S.n3226 S.n3221 0.001
R9360 S.t30 S.n3242 0.001
R9361 S.t30 S.n3239 0.001
R9362 S.n3239 S.n3236 0.001
R9363 S.n2685 S.t68 0.001
R9364 S.n2693 S.n2688 0.001
R9365 S.t256 S.n2709 0.001
R9366 S.t256 S.n2706 0.001
R9367 S.n2706 S.n2703 0.001
R9368 S.n2142 S.t56 0.001
R9369 S.n2150 S.n2145 0.001
R9370 S.t290 S.n2166 0.001
R9371 S.t290 S.n2163 0.001
R9372 S.n2163 S.n2160 0.001
R9373 S.t32 S.n1515 0.001
R9374 S.t32 S.n1518 0.001
R9375 S.t18 S.n1596 0.001
R9376 S.t18 S.n1593 0.001
R9377 S.n1593 S.n1590 0.001
R9378 S.n980 S.t14 0.001
R9379 S.n988 S.n983 0.001
R9380 S.t58 S.n1008 0.001
R9381 S.t58 S.n1005 0.001
R9382 S.n1005 S.n1002 0.001
R9383 S.t151 S.n109 0.001
R9384 S.t151 S.n106 0.001
R9385 S.n106 S.n103 0.001
R9386 S.t58 S.n1212 0.001
R9387 S.t58 S.n1215 0.001
R9388 S.t30 S.n3267 0.001
R9389 S.t30 S.n3264 0.001
R9390 S.n3264 S.n3261 0.001
R9391 S.t68 S.n2517 0.001
R9392 S.t68 S.n2514 0.001
R9393 S.n2514 S.n2511 0.001
R9394 S.t256 S.n2918 0.001
R9395 S.t256 S.n2921 0.001
R9396 S.t56 S.n1992 0.001
R9397 S.t56 S.n1989 0.001
R9398 S.n1989 S.n1986 0.001
R9399 S.t290 S.n2362 0.001
R9400 S.t290 S.n2365 0.001
R9401 S.t32 S.n1399 0.001
R9402 S.t32 S.n1396 0.001
R9403 S.n1396 S.n1393 0.001
R9404 S.t18 S.n1802 0.001
R9405 S.t18 S.n1805 0.001
R9406 S.t14 S.n855 0.001
R9407 S.t14 S.n852 0.001
R9408 S.n852 S.n849 0.001
R9409 S.n469 S.t151 0.001
R9410 S.n477 S.n472 0.001
R9411 S.t200 S.n3782 0.001
R9412 S.t200 S.n3779 0.001
R9413 S.n3779 S.n3776 0.001
R9414 S.t27 S.n3053 0.001
R9415 S.t27 S.n3050 0.001
R9416 S.n3050 S.n3047 0.001
R9417 S.t30 S.n3414 0.001
R9418 S.t30 S.n3417 0.001
R9419 S.t68 S.n2536 0.001
R9420 S.t68 S.n2533 0.001
R9421 S.n2533 S.n2530 0.001
R9422 S.t256 S.n2886 0.001
R9423 S.t256 S.n2889 0.001
R9424 S.t56 S.n2009 0.001
R9425 S.t56 S.n2006 0.001
R9426 S.n2006 S.n2003 0.001
R9427 S.t290 S.n2331 0.001
R9428 S.t290 S.n2334 0.001
R9429 S.t32 S.n1416 0.001
R9430 S.t32 S.n1413 0.001
R9431 S.n1413 S.n1410 0.001
R9432 S.t18 S.n1770 0.001
R9433 S.t18 S.n1773 0.001
R9434 S.t14 S.n874 0.001
R9435 S.t14 S.n871 0.001
R9436 S.n871 S.n868 0.001
R9437 S.t14 S.n896 0.001
R9438 S.t14 S.n893 0.001
R9439 S.n893 S.n890 0.001
R9440 S.t58 S.n1154 0.001
R9441 S.t58 S.n1157 0.001
R9442 S.n302 S.t213 0.001
R9443 S.n310 S.n305 0.001
R9444 S.t151 S.n331 0.001
R9445 S.t151 S.n328 0.001
R9446 S.n328 S.n325 0.001
R9447 S.t18 S.n1741 0.001
R9448 S.t18 S.n1744 0.001
R9449 S.t290 S.n2302 0.001
R9450 S.t290 S.n2305 0.001
R9451 S.t256 S.n2853 0.001
R9452 S.t256 S.n2856 0.001
R9453 S.t30 S.n3381 0.001
R9454 S.t30 S.n3384 0.001
R9455 S.t200 S.n3899 0.001
R9456 S.t200 S.n3902 0.001
R9457 S.t77 S.n4278 0.001
R9458 S.t77 S.n4275 0.001
R9459 S.n4275 S.n4272 0.001
R9460 S.t6 S.n3565 0.001
R9461 S.t6 S.n3562 0.001
R9462 S.n3562 S.n3559 0.001
R9463 S.t27 S.n3072 0.001
R9464 S.t27 S.n3069 0.001
R9465 S.n3069 S.n3066 0.001
R9466 S.t68 S.n2555 0.001
R9467 S.t68 S.n2552 0.001
R9468 S.n2552 S.n2549 0.001
R9469 S.t56 S.n2028 0.001
R9470 S.t56 S.n2025 0.001
R9471 S.n2025 S.n2022 0.001
R9472 S.t32 S.n1436 0.001
R9473 S.t32 S.n1433 0.001
R9474 S.n1433 S.n1430 0.001
R9475 S.t58 S.n1120 0.001
R9476 S.t58 S.n1123 0.001
R9477 S.t213 S.n260 0.001
R9478 S.t213 S.n257 0.001
R9479 S.n257 S.n254 0.001
R9480 S.n659 S.n653 0.001
R9481 S.t20 S.n4461 0.001
R9482 S.t20 S.n4464 0.001
R9483 S.t65 S.n4071 0.001
R9484 S.t65 S.n4068 0.001
R9485 S.n4068 S.n4065 0.001
R9486 S.t77 S.n4367 0.001
R9487 S.t77 S.n4370 0.001
R9488 S.t6 S.n3591 0.001
R9489 S.t6 S.n3588 0.001
R9490 S.n3588 S.n3585 0.001
R9491 S.t200 S.n3867 0.001
R9492 S.t200 S.n3870 0.001
R9493 S.t27 S.n3097 0.001
R9494 S.t27 S.n3094 0.001
R9495 S.n3094 S.n3091 0.001
R9496 S.t30 S.n3349 0.001
R9497 S.t30 S.n3352 0.001
R9498 S.t68 S.n2580 0.001
R9499 S.t68 S.n2577 0.001
R9500 S.n2577 S.n2574 0.001
R9501 S.t256 S.n2821 0.001
R9502 S.t256 S.n2824 0.001
R9503 S.t56 S.n2053 0.001
R9504 S.t56 S.n2050 0.001
R9505 S.n2050 S.n2047 0.001
R9506 S.t290 S.n2271 0.001
R9507 S.t290 S.n2274 0.001
R9508 S.t32 S.n1461 0.001
R9509 S.t32 S.n1458 0.001
R9510 S.n1458 S.n1455 0.001
R9511 S.t18 S.n1708 0.001
R9512 S.t18 S.n1711 0.001
R9513 S.t14 S.n920 0.001
R9514 S.t14 S.n917 0.001
R9515 S.n917 S.n914 0.001
R9516 S.t58 S.n1087 0.001
R9517 S.t58 S.n1090 0.001
R9518 S.t213 S.n279 0.001
R9519 S.t213 S.n276 0.001
R9520 S.n276 S.n273 0.001
R9521 S.t14 S.n941 0.001
R9522 S.t14 S.n938 0.001
R9523 S.n938 S.n935 0.001
R9524 S.t18 S.n1676 0.001
R9525 S.t18 S.n1679 0.001
R9526 S.t32 S.n1481 0.001
R9527 S.t32 S.n1478 0.001
R9528 S.n1478 S.n1475 0.001
R9529 S.t290 S.n2239 0.001
R9530 S.t290 S.n2242 0.001
R9531 S.t56 S.n2073 0.001
R9532 S.t56 S.n2070 0.001
R9533 S.n2070 S.n2067 0.001
R9534 S.t256 S.n2789 0.001
R9535 S.t256 S.n2792 0.001
R9536 S.t68 S.n2600 0.001
R9537 S.t68 S.n2597 0.001
R9538 S.n2597 S.n2594 0.001
R9539 S.t30 S.n3317 0.001
R9540 S.t30 S.n3320 0.001
R9541 S.t27 S.n3117 0.001
R9542 S.t27 S.n3114 0.001
R9543 S.n3114 S.n3111 0.001
R9544 S.t200 S.n3832 0.001
R9545 S.t200 S.n3835 0.001
R9546 S.t6 S.n3611 0.001
R9547 S.t6 S.n3608 0.001
R9548 S.n3608 S.n3605 0.001
R9549 S.t77 S.n4332 0.001
R9550 S.t77 S.n4335 0.001
R9551 S.t65 S.n4093 0.001
R9552 S.t65 S.n4090 0.001
R9553 S.n4090 S.n4087 0.001
R9554 S.t20 S.n4406 0.001
R9555 S.t20 S.n4403 0.001
R9556 S.n4403 S.n4400 0.001
R9557 S.t4 S.n4512 0.001
R9558 S.t4 S.n4509 0.001
R9559 S.n4509 S.n4506 0.001
R9560 S.t36 S.n4907 0.001
R9561 S.t36 S.n4910 0.001
R9562 S.t151 S.n357 0.001
R9563 S.t151 S.n354 0.001
R9564 S.n354 S.n351 0.001
R9565 S.t58 S.n1182 0.001
R9566 S.t58 S.n1185 0.001
R9567 S.t213 S.n236 0.001
R9568 S.t213 S.n233 0.001
R9569 S.n233 S.n230 0.001
R9570 S.t213 S.n219 0.001
R9571 S.t213 S.n216 0.001
R9572 S.n216 S.n213 0.001
R9573 S.t151 S.n77 0.001
R9574 S.t151 S.n74 0.001
R9575 S.n74 S.n71 0.001
R9576 S.t58 S.n1271 0.001
R9577 S.t58 S.n1274 0.001
R9578 S.t290 S.n2190 0.001
R9579 S.t290 S.n2187 0.001
R9580 S.n2187 S.n2184 0.001
R9581 S.t32 S.n1360 0.001
R9582 S.t32 S.n1357 0.001
R9583 S.n1357 S.n1354 0.001
R9584 S.t18 S.n1867 0.001
R9585 S.t18 S.n1870 0.001
R9586 S.t14 S.n819 0.001
R9587 S.t14 S.n816 0.001
R9588 S.n816 S.n813 0.001
R9589 S.n518 S.n513 0.001
R9590 S.t256 S.n2739 0.001
R9591 S.t256 S.n2736 0.001
R9592 S.n2736 S.n2733 0.001
R9593 S.t56 S.n1973 0.001
R9594 S.t56 S.n1970 0.001
R9595 S.n1970 S.n1967 0.001
R9596 S.t290 S.n2395 0.001
R9597 S.t290 S.n2398 0.001
R9598 S.t32 S.n1379 0.001
R9599 S.t32 S.n1376 0.001
R9600 S.n1376 S.n1373 0.001
R9601 S.t18 S.n1835 0.001
R9602 S.t18 S.n1838 0.001
R9603 S.t14 S.n836 0.001
R9604 S.t14 S.n833 0.001
R9605 S.n833 S.n830 0.001
R9606 S.t58 S.n1241 0.001
R9607 S.t58 S.n1244 0.001
R9608 S.t213 S.n201 0.001
R9609 S.t213 S.n198 0.001
R9610 S.n198 S.n195 0.001
R9611 S.t213 S.n184 0.001
R9612 S.t213 S.n181 0.001
R9613 S.n181 S.n178 0.001
R9614 S.t151 S.n45 0.001
R9615 S.t151 S.n42 0.001
R9616 S.n42 S.n39 0.001
R9617 S.t58 S.n1031 0.001
R9618 S.t58 S.n1028 0.001
R9619 S.n1028 S.n1025 0.001
R9620 S.n556 S.n551 0.001
R9621 S.t18 S.n1626 0.001
R9622 S.t18 S.n1623 0.001
R9623 S.n1623 S.n1620 0.001
R9624 S.t14 S.n800 0.001
R9625 S.t14 S.n797 0.001
R9626 S.n797 S.n794 0.001
R9627 S.t58 S.n1304 0.001
R9628 S.t58 S.n1307 0.001
R9629 S.t213 S.n166 0.001
R9630 S.t213 S.n163 0.001
R9631 S.n163 S.n160 0.001
R9632 S.t213 S.n150 0.001
R9633 S.t213 S.n147 0.001
R9634 S.n147 S.n144 0.001
R9635 S.t151 S.n411 0.001
R9636 S.t151 S.n435 0.001
R9637 S.n435 S.n432 0.001
R9638 S.n5419 S.n5416 0.001
R9639 S.t52 S.n5422 0.001
R9640 S.n5261 S.t36 0.001
R9641 S.n5270 S.n5263 0.001
R9642 S.t34 S.n5686 0.001
R9643 S.t34 S.n5689 0.001
R9644 S.t45 S.n4996 0.001
R9645 S.t45 S.n4993 0.001
R9646 S.n4993 S.n4990 0.001
R9647 S.t52 S.n5448 0.001
R9648 S.n5442 S.n5441 0.001
R9649 S.t52 S.n5419 0.001
R9650 S.n5686 S.n5683 0.001
R9651 S.n5270 S.n5261 0.001
R9652 S.n720 S.t191 0.001
R9653 S.n377 S.n364 0.001
R9654 S.n1059 S.n1056 0.001
R9655 S.n1656 S.n1653 0.001
R9656 S.n2219 S.n2216 0.001
R9657 S.n2769 S.n2766 0.001
R9658 S.n3297 S.n3294 0.001
R9659 S.n3812 S.n3809 0.001
R9660 S.n4308 S.n4305 0.001
R9661 S.n4907 S.n4904 0.001
R9662 S.n4332 S.n4329 0.001
R9663 S.n3832 S.n3829 0.001
R9664 S.n3317 S.n3314 0.001
R9665 S.n2789 S.n2786 0.001
R9666 S.n2239 S.n2236 0.001
R9667 S.n1676 S.n1673 0.001
R9668 S.n1087 S.n1084 0.001
R9669 S.n4461 S.n4458 0.001
R9670 S.n4367 S.n4364 0.001
R9671 S.n3867 S.n3864 0.001
R9672 S.n3349 S.n3346 0.001
R9673 S.n2821 S.n2818 0.001
R9674 S.n2271 S.n2268 0.001
R9675 S.n1708 S.n1705 0.001
R9676 S.n1120 S.n1117 0.001
R9677 S.n659 S.n650 0.001
R9678 S.n310 S.n302 0.001
R9679 S.n1154 S.n1151 0.001
R9680 S.n1741 S.n1738 0.001
R9681 S.n2302 S.n2299 0.001
R9682 S.n2853 S.n2850 0.001
R9683 S.n3381 S.n3378 0.001
R9684 S.n3899 S.n3896 0.001
R9685 S.n3414 S.n3411 0.001
R9686 S.n2886 S.n2883 0.001
R9687 S.n2331 S.n2328 0.001
R9688 S.n1770 S.n1767 0.001
R9689 S.n1182 S.n1179 0.001
R9690 S.n477 S.n469 0.001
R9691 S.n1212 S.n1209 0.001
R9692 S.n1802 S.n1799 0.001
R9693 S.n2362 S.n2359 0.001
R9694 S.n2918 S.n2915 0.001
R9695 S.n2395 S.n2392 0.001
R9696 S.n1835 S.n1832 0.001
R9697 S.n1241 S.n1238 0.001
R9698 S.n518 S.n510 0.001
R9699 S.n1271 S.n1268 0.001
R9700 S.n1867 S.n1864 0.001
R9701 S.n1304 S.n1301 0.001
R9702 S.n556 S.n548 0.001
R9703 S.n466 S.n463 0.001
R9704 S.n5463 S.n5460 0.001
R9705 S.n5010 S.n5007 0.001
R9706 S.n4926 S.n4923 0.001
R9707 S.n4677 S.n4669 0.001
R9708 S.n4690 S.n4687 0.001
R9709 S.n4234 S.n4226 0.001
R9710 S.n3736 S.n3728 0.001
R9711 S.n3226 S.n3218 0.001
R9712 S.n2693 S.n2685 0.001
R9713 S.n2150 S.n2142 0.001
R9714 S.n1515 S.n1512 0.001
R9715 S.n988 S.n980 0.001
R9716 S.n296 S.n293 0.001
R9717 S.n1315 S.n1314 0.001
R9718 S.n5480 S.n5477 0.001
R9719 S.n5124 S.n5120 0.001
R9720 S.n5129 S.n5126 0.001
R9721 S.n4544 S.n4541 0.001
R9722 S.n4706 S.n4703 0.001
R9723 S.n4125 S.n4122 0.001
R9724 S.n3643 S.n3640 0.001
R9725 S.n3149 S.n3146 0.001
R9726 S.n2632 S.n2629 0.001
R9727 S.n2105 S.n2102 0.001
R9728 S.n1531 S.n1528 0.001
R9729 S.n974 S.n971 0.001
R9730 S.n1878 S.n1877 0.001
R9731 S.n5589 S.n5585 0.001
R9732 S.n5155 S.n5151 0.001
R9733 S.n5160 S.n5157 0.001
R9734 S.n4559 S.n4556 0.001
R9735 S.n4722 S.n4719 0.001
R9736 S.n4140 S.n4137 0.001
R9737 S.n3658 S.n3655 0.001
R9738 S.n3164 S.n3161 0.001
R9739 S.n2647 S.n2644 0.001
R9740 S.n2120 S.n2117 0.001
R9741 S.n1545 S.n1537 0.001
R9742 S.n2406 S.n2405 0.001
R9743 S.n2136 S.n2133 0.001
R9744 S.n2663 S.n2660 0.001
R9745 S.n3180 S.n3177 0.001
R9746 S.n3674 S.n3671 0.001
R9747 S.n4156 S.n4153 0.001
R9748 S.n4737 S.n4734 0.001
R9749 S.n4575 S.n4572 0.001
R9750 S.n5175 S.n5172 0.001
R9751 S.n5026 S.n5023 0.001
R9752 S.n5496 S.n5493 0.001
R9753 S.n2929 S.n2928 0.001
R9754 S.n2679 S.n2676 0.001
R9755 S.n3196 S.n3193 0.001
R9756 S.n3690 S.n3687 0.001
R9757 S.n4172 S.n4169 0.001
R9758 S.n4752 S.n4749 0.001
R9759 S.n4591 S.n4588 0.001
R9760 S.n5190 S.n5187 0.001
R9761 S.n5042 S.n5039 0.001
R9762 S.n5512 S.n5509 0.001
R9763 S.n3425 S.n3424 0.001
R9764 S.n3212 S.n3209 0.001
R9765 S.n3706 S.n3703 0.001
R9766 S.n4188 S.n4185 0.001
R9767 S.n4767 S.n4764 0.001
R9768 S.n4607 S.n4604 0.001
R9769 S.n5205 S.n5202 0.001
R9770 S.n5058 S.n5055 0.001
R9771 S.n5528 S.n5525 0.001
R9772 S.n3910 S.n3909 0.001
R9773 S.n3722 S.n3719 0.001
R9774 S.n4204 S.n4201 0.001
R9775 S.n4782 S.n4779 0.001
R9776 S.n4623 S.n4620 0.001
R9777 S.n5220 S.n5217 0.001
R9778 S.n5074 S.n5071 0.001
R9779 S.n5544 S.n5541 0.001
R9780 S.n4378 S.n4377 0.001
R9781 S.n4220 S.n4217 0.001
R9782 S.n4798 S.n4795 0.001
R9783 S.n4639 S.n4636 0.001
R9784 S.n5235 S.n5232 0.001
R9785 S.n5090 S.n5087 0.001
R9786 S.n5560 S.n5557 0.001
R9787 S.n4834 S.n4804 0.001
R9788 S.n4663 S.n4660 0.001
R9789 S.n5255 S.n5252 0.001
R9790 S.n5111 S.n5108 0.001
R9791 S.n5576 S.n5573 0.001
R9792 S.n5813 S.n5812 0.001
R9793 S.n5812 S.n5805 0.001
R9794 S.n460 S.n459 0.001
R9795 S.n751 S.n750 0.001
R9796 S.n1560 S.n1559 0.001
R9797 S.n1893 S.n1892 0.001
R9798 S.n2421 S.n2420 0.001
R9799 S.n2943 S.n2942 0.001
R9800 S.n3439 S.n3438 0.001
R9801 S.n3924 S.n3923 0.001
R9802 S.n4830 S.n4829 0.001
R9803 S.n4848 S.n4847 0.001
R9804 S.n5702 S.n5701 0.001
R9805 S.n5390 S.n5389 0.001
R9806 S.n5717 S.n5716 0.001
R9807 S.n577 S.n576 0.001
R9808 S.n580 S.n579 0.001
R9809 S.n5716 S.n5715 0.001
R9810 S.n459 S.n458 0.001
R9811 S.n750 S.n749 0.001
R9812 S.n1559 S.n1558 0.001
R9813 S.n1892 S.n1891 0.001
R9814 S.n2420 S.n2419 0.001
R9815 S.n2942 S.n2941 0.001
R9816 S.n3438 S.n3437 0.001
R9817 S.n3923 S.n3922 0.001
R9818 S.n4829 S.n4828 0.001
R9819 S.n4847 S.n4846 0.001
R9820 S.n5707 S.n5705 0.001
R9821 S.n4849 S.n4839 0.001
R9822 S.n461 S.n451 0.001
R9823 S.n752 S.n742 0.001
R9824 S.n1561 S.n1551 0.001
R9825 S.n1894 S.n1884 0.001
R9826 S.n2422 S.n2412 0.001
R9827 S.n2944 S.n2934 0.001
R9828 S.n3440 S.n3430 0.001
R9829 S.n3925 S.n3915 0.001
R9830 S.n4831 S.n4821 0.001
R9831 S.n5720 S.n5719 0.001
R9832 S.n5701 S.n5700 0.001
R9833 S.n5814 S.n5813 0.001
R9834 S.n5805 S.n5804 0.001
R9835 S.n5441 S.n5437 0.001
R9836 D.n1907 D.t902 7.599
R9837 D.n1897 D.t126 7.599
R9838 D.n231 D.t453 7.599
R9839 D.n222 D.t183 7.599
R9840 D.n28 D.t344 7.599
R9841 D.n1990 D.t500 7.599
R9842 D.n2015 D.t1001 7.599
R9843 D.n2000 D.t48 7.599
R9844 D.n3555 D.t1060 7.599
R9845 D.n3537 D.t1073 7.599
R9846 D.n3519 D.t1090 7.599
R9847 D.n3501 D.t1100 7.599
R9848 D.n3483 D.t9 7.599
R9849 D.n3465 D.t23 7.599
R9850 D.n3447 D.t31 7.599
R9851 D.n3429 D.t39 7.599
R9852 D.n3411 D.t51 7.599
R9853 D.n3392 D.t21 7.599
R9854 D.n3401 D.t694 7.599
R9855 D.n3419 D.t1005 7.599
R9856 D.n3437 D.t996 7.599
R9857 D.n3455 D.t979 7.599
R9858 D.n3473 D.t593 7.599
R9859 D.n3491 D.t637 7.599
R9860 D.n3509 D.t622 7.599
R9861 D.n3527 D.t612 7.599
R9862 D.n3545 D.t600 7.599
R9863 D.n3567 D.t947 7.599
R9864 D.n3584 D.t627 7.599
R9865 D.n3157 D.t687 7.599
R9866 D.n3177 D.t700 7.599
R9867 D.n3197 D.t717 7.599
R9868 D.n3217 D.t727 7.599
R9869 D.n3237 D.t739 7.599
R9870 D.n3257 D.t751 7.599
R9871 D.n3277 D.t763 7.599
R9872 D.n3297 D.t771 7.599
R9873 D.n3317 D.t753 7.599
R9874 D.n3305 D.t228 7.599
R9875 D.n3285 D.t620 7.599
R9876 D.n3265 D.t610 7.599
R9877 D.n3245 D.t597 7.599
R9878 D.n3225 D.t272 7.599
R9879 D.n3205 D.t256 7.599
R9880 D.n3185 D.t242 7.599
R9881 D.n3165 D.t234 7.599
R9882 D.n3142 D.t323 7.599
R9883 D.n3132 D.t864 7.599
R9884 D.n3072 D.t321 7.599
R9885 D.n3054 D.t336 7.599
R9886 D.n3036 D.t351 7.599
R9887 D.n3018 D.t363 7.599
R9888 D.n3000 D.t375 7.599
R9889 D.n2982 D.t387 7.599
R9890 D.n2964 D.t396 7.599
R9891 D.n2945 D.t378 7.599
R9892 D.n2954 D.t959 7.599
R9893 D.n2972 D.t241 7.599
R9894 D.n2990 D.t230 7.599
R9895 D.n3008 D.t276 7.599
R9896 D.n3026 D.t997 7.599
R9897 D.n3044 D.t981 7.599
R9898 D.n3062 D.t970 7.599
R9899 D.n3084 D.t830 7.599
R9900 D.n3101 D.t229 7.599
R9901 D.n2754 D.t1055 7.599
R9902 D.n2774 D.t1068 7.599
R9903 D.n2794 D.t1087 7.599
R9904 D.n2814 D.t1098 7.599
R9905 D.n2834 D.t8 7.599
R9906 D.n2854 D.t19 7.599
R9907 D.n2874 D.t1102 7.599
R9908 D.n2862 D.t582 7.599
R9909 D.n2842 D.t967 7.599
R9910 D.n2822 D.t1015 7.599
R9911 D.n2802 D.t1000 7.599
R9912 D.n2782 D.t611 7.599
R9913 D.n2762 D.t598 7.599
R9914 D.n2737 D.t219 7.599
R9915 D.n2724 D.t761 7.599
R9916 D.n2673 D.t681 7.599
R9917 D.n2655 D.t697 7.599
R9918 D.n2637 D.t712 7.599
R9919 D.n2619 D.t725 7.599
R9920 D.n2601 D.t736 7.599
R9921 D.n2582 D.t714 7.599
R9922 D.n2591 D.t211 7.599
R9923 D.n2609 D.t641 7.599
R9924 D.n2627 D.t626 7.599
R9925 D.n2645 D.t614 7.599
R9926 D.n2663 D.t231 7.599
R9927 D.n2684 D.t738 7.599
R9928 D.n2695 D.t185 7.599
R9929 D.n2431 D.t316 7.599
R9930 D.n2451 D.t332 7.599
R9931 D.n2471 D.t349 7.599
R9932 D.n2491 D.t362 7.599
R9933 D.n2511 D.t334 7.599
R9934 D.n2499 D.t972 7.599
R9935 D.n2479 D.t259 7.599
R9936 D.n2459 D.t244 7.599
R9937 D.n2439 D.t237 7.599
R9938 D.n2414 D.t156 7.599
R9939 D.n2401 D.t645 7.599
R9940 D.n2348 D.t1050 7.599
R9941 D.n2330 D.t1066 7.599
R9942 D.n2312 D.t1084 7.599
R9943 D.n2293 D.t1051 7.599
R9944 D.n2302 D.t592 7.599
R9945 D.n2320 D.t987 7.599
R9946 D.n2338 D.t974 7.599
R9947 D.n2360 D.t373 7.599
R9948 D.n2377 D.t68 7.599
R9949 D.n2182 D.t678 7.599
R9950 D.n2202 D.t695 7.599
R9951 D.n2222 D.t662 7.599
R9952 D.n2210 D.t222 7.599
R9953 D.n2190 D.t605 7.599
R9954 D.n2167 D.t887 7.599
R9955 D.n2157 D.t571 7.599
R9956 D.n2109 D.t312 7.599
R9957 D.n2090 D.t280 7.599
R9958 D.n2099 D.t952 7.599
R9959 D.n2121 D.t245 7.599
R9960 D.n2138 D.t1079 7.599
R9961 D.n1969 D.t949 7.599
R9962 D.n50 D.t1082 7.599
R9963 D.n59 D.t603 7.599
R9964 D.n68 D.t924 7.599
R9965 D.n77 D.t421 7.599
R9966 D.n86 D.t269 7.599
R9967 D.n95 D.t408 7.599
R9968 D.n104 D.t255 7.599
R9969 D.n113 D.t398 7.599
R9970 D.n122 D.t973 7.599
R9971 D.n131 D.t389 7.599
R9972 D.n140 D.t963 7.599
R9973 D.n149 D.t376 7.599
R9974 D.n158 D.t1011 7.599
R9975 D.n167 D.t366 7.599
R9976 D.n176 D.t999 7.599
R9977 D.n185 D.t355 7.599
R9978 D.n194 D.t982 7.599
R9979 D.n203 D.t340 7.599
R9980 D.n212 D.t108 7.599
R9981 D.n283 D.t481 7.599
R9982 D.n299 D.t557 7.599
R9983 D.n551 D.t948 7.599
R9984 D.n537 D.t196 7.599
R9985 D.n523 D.t755 7.599
R9986 D.n509 D.t1017 7.599
R9987 D.n495 D.t786 7.599
R9988 D.n481 D.t635 7.599
R9989 D.n467 D.t773 7.599
R9990 D.n453 D.t246 7.599
R9991 D.n439 D.t765 7.599
R9992 D.n425 D.t236 7.599
R9993 D.n411 D.t754 7.599
R9994 D.n397 D.t225 7.599
R9995 D.n383 D.t741 7.599
R9996 D.n369 D.t273 7.599
R9997 D.n355 D.t729 7.599
R9998 D.n341 D.t257 7.599
R9999 D.n327 D.t719 7.599
R10000 D.n313 D.t498 7.599
R10001 D.n574 D.t859 7.599
R10002 D.n590 D.t931 7.599
R10003 D.n814 D.t1083 7.599
R10004 D.n800 D.t296 7.599
R10005 D.n786 D.t893 7.599
R10006 D.n772 D.t58 7.599
R10007 D.n758 D.t54 7.599
R10008 D.n744 D.t628 7.599
R10009 D.n730 D.t43 7.599
R10010 D.n716 D.t615 7.599
R10011 D.n702 D.t33 7.599
R10012 D.n688 D.t607 7.599
R10013 D.n674 D.t24 7.599
R10014 D.n660 D.t594 7.599
R10015 D.n646 D.t11 7.599
R10016 D.n632 D.t640 7.599
R10017 D.n618 D.t1 7.599
R10018 D.n604 D.t876 7.599
R10019 D.n837 D.t140 7.599
R10020 D.n853 D.t203 7.599
R10021 D.n1049 D.t107 7.599
R10022 D.n1035 D.t437 7.599
R10023 D.n1021 D.t980 7.599
R10024 D.n1007 D.t289 7.599
R10025 D.n993 D.t423 7.599
R10026 D.n979 D.t1002 7.599
R10027 D.n965 D.t410 7.599
R10028 D.n951 D.t992 7.599
R10029 D.n937 D.t399 7.599
R10030 D.n923 D.t976 7.599
R10031 D.n909 D.t390 7.599
R10032 D.n895 D.t964 7.599
R10033 D.n881 D.t381 7.599
R10034 D.n867 D.t151 7.599
R10035 D.n1072 D.t524 7.599
R10036 D.n1088 D.t573 7.599
R10037 D.n1256 D.t217 7.599
R10038 D.n1242 D.t673 7.599
R10039 D.n1228 D.t30 7.599
R10040 D.n1214 D.t434 7.599
R10041 D.n1200 D.t787 7.599
R10042 D.n1186 D.t264 7.599
R10043 D.n1172 D.t775 7.599
R10044 D.n1158 D.t250 7.599
R10045 D.n1144 D.t767 7.599
R10046 D.n1130 D.t238 7.599
R10047 D.n1116 D.t758 7.599
R10048 D.n1102 D.t470 7.599
R10049 D.n1279 D.t832 7.599
R10050 D.n1295 D.t950 7.599
R10051 D.n1435 D.t360 7.599
R10052 D.n1421 D.t807 7.599
R10053 D.n1407 D.t170 7.599
R10054 D.n1393 D.t564 7.599
R10055 D.n1379 D.t55 7.599
R10056 D.n1365 D.t630 7.599
R10057 D.n1351 D.t45 7.599
R10058 D.n1337 D.t619 7.599
R10059 D.n1323 D.t35 7.599
R10060 D.n1309 D.t851 7.599
R10061 D.n1459 D.t114 7.599
R10062 D.n1475 D.t220 7.599
R10063 D.n1587 D.t490 7.599
R10064 D.n1573 D.t939 7.599
R10065 D.n1559 D.t247 7.599
R10066 D.n1545 D.t666 7.599
R10067 D.n1531 D.t426 7.599
R10068 D.n1517 D.t1004 7.599
R10069 D.n1503 D.t413 7.599
R10070 D.n1489 D.t129 7.599
R10071 D.n1611 D.t506 7.599
R10072 D.n1627 D.t591 7.599
R10073 D.n1711 D.t585 7.599
R10074 D.n1697 D.t1054 7.599
R10075 D.n1683 D.t401 7.599
R10076 D.n1669 D.t803 7.599
R10077 D.n1655 D.t790 7.599
R10078 D.n1641 D.t516 7.599
R10079 D.n1735 D.t883 7.599
R10080 D.n1751 D.t968 7.599
R10081 D.n1807 D.t726 7.599
R10082 D.n1793 D.t83 7.599
R10083 D.n1779 D.t546 7.599
R10084 D.n1765 D.t715 7.599
R10085 D.n1830 D.t847 7.599
R10086 D.n1846 D.t566 7.599
R10087 D.n1874 D.t863 7.599
R10088 D.n1860 D.t1099 7.599
R10089 D.n1911 D.t353 7.493
R10090 D.n1901 D.t756 7.493
R10091 D.n234 D.t135 7.493
R10092 D.n225 D.t984 7.493
R10093 D.n32 D.t207 7.493
R10094 D.n1952 D.t275 7.493
R10095 D.n2036 D.t281 7.493
R10096 D.n2019 D.t587 7.493
R10097 D.n2004 D.t975 7.493
R10098 D.n3558 D.t409 7.493
R10099 D.n3540 D.t881 7.493
R10100 D.n3522 D.t891 7.493
R10101 D.n3504 D.t903 7.493
R10102 D.n3486 D.t915 7.493
R10103 D.n3468 D.t141 7.493
R10104 D.n3450 D.t153 7.493
R10105 D.n3432 D.t167 7.493
R10106 D.n3414 D.t180 7.493
R10107 D.n3395 D.t937 7.493
R10108 D.n3369 D.t460 7.493
R10109 D.n3405 D.t828 7.493
R10110 D.n3423 D.t813 7.493
R10111 D.n3441 D.t802 7.493
R10112 D.n3459 D.t795 7.493
R10113 D.n3477 D.t783 7.493
R10114 D.n3495 D.t770 7.493
R10115 D.n3513 D.t760 7.493
R10116 D.n3531 D.t748 7.493
R10117 D.n3549 D.t737 7.493
R10118 D.n3571 D.t590 7.493
R10119 D.n3160 D.t900 7.493
R10120 D.n3180 D.t514 7.493
R10121 D.n3200 D.t527 7.493
R10122 D.n3220 D.t538 7.493
R10123 D.n3240 D.t921 7.493
R10124 D.n3260 D.t877 7.493
R10125 D.n3280 D.t889 7.493
R10126 D.n3300 D.t899 7.493
R10127 D.n3320 D.t511 7.493
R10128 D.n3334 D.t32 7.493
R10129 D.n3309 D.t451 7.493
R10130 D.n3289 D.t440 7.493
R10131 D.n3269 D.t430 7.493
R10132 D.n3249 D.t419 7.493
R10133 D.n3229 D.t406 7.493
R10134 D.n3209 D.t394 7.493
R10135 D.n3189 D.t385 7.493
R10136 D.n3169 D.t374 7.493
R10137 D.n3146 D.t386 7.493
R10138 D.n3075 D.t260 7.493
R10139 D.n3057 D.t143 7.493
R10140 D.n3039 D.t154 7.493
R10141 D.n3021 D.t544 7.493
R10142 D.n3003 D.t553 7.493
R10143 D.n2985 D.t512 7.493
R10144 D.n2967 D.t522 7.493
R10145 D.n2948 D.t119 7.493
R10146 D.n2926 D.t752 7.493
R10147 D.n2958 D.t69 7.493
R10148 D.n2976 D.t61 7.493
R10149 D.n2994 D.t49 7.493
R10150 D.n3012 D.t37 7.493
R10151 D.n3030 D.t27 7.493
R10152 D.n3048 D.t17 7.493
R10153 D.n3066 D.t7 7.493
R10154 D.n3088 D.t886 7.493
R10155 D.n2757 D.t789 7.493
R10156 D.n2777 D.t878 7.493
R10157 D.n2797 D.t163 7.493
R10158 D.n2817 D.t175 7.493
R10159 D.n2837 D.t188 7.493
R10160 D.n2857 D.t138 7.493
R10161 D.n2877 D.t836 7.493
R10162 D.n2891 D.t377 7.493
R10163 D.n2866 D.t792 7.493
R10164 D.n2846 D.t779 7.493
R10165 D.n2826 D.t769 7.493
R10166 D.n2806 D.t759 7.493
R10167 D.n2786 D.t747 7.493
R10168 D.n2766 D.t735 7.493
R10169 D.n2741 D.t235 7.493
R10170 D.n2676 D.t201 7.493
R10171 D.n2658 D.t884 7.493
R10172 D.n2640 D.t895 7.493
R10173 D.n2622 D.t909 7.493
R10174 D.n2604 D.t919 7.493
R10175 D.n2585 D.t459 7.493
R10176 D.n2563 D.t1101 7.493
R10177 D.n2595 D.t415 7.493
R10178 D.n2613 D.t403 7.493
R10179 D.n2631 D.t391 7.493
R10180 D.n2649 D.t384 7.493
R10181 D.n2667 D.t372 7.493
R10182 D.n2688 D.t750 7.493
R10183 D.n2434 D.t424 7.493
R10184 D.n2454 D.t518 7.493
R10185 D.n2474 D.t532 7.493
R10186 D.n2494 D.t543 7.493
R10187 D.n2514 D.t147 7.493
R10188 D.n2528 D.t713 7.493
R10189 D.n2503 D.t36 7.493
R10190 D.n2483 D.t25 7.493
R10191 D.n2463 D.t15 7.493
R10192 D.n2443 D.t5 7.493
R10193 D.n2418 D.t155 7.493
R10194 D.n2351 D.t935 7.493
R10195 D.n2333 D.t146 7.493
R10196 D.n2315 D.t161 7.493
R10197 D.n2296 D.t865 7.493
R10198 D.n2274 D.t333 7.493
R10199 D.n2306 D.t757 7.493
R10200 D.n2324 D.t744 7.493
R10201 D.n2342 D.t732 7.493
R10202 D.n2364 D.t601 7.493
R10203 D.n2185 D.t322 7.493
R10204 D.n2205 D.t880 7.493
R10205 D.n2225 D.t484 7.493
R10206 D.n2239 D.t1049 7.493
R10207 D.n2214 D.t382 7.493
R10208 D.n2194 D.t369 7.493
R10209 D.n2171 D.t22 7.493
R10210 D.n2112 D.t835 7.493
R10211 D.n2093 D.t94 7.493
R10212 D.n2071 D.t663 7.493
R10213 D.n2103 D.t2 7.493
R10214 D.n2125 D.t528 7.493
R10215 D.n54 D.t691 7.493
R10216 D.n63 D.t40 7.493
R10217 D.n72 D.t96 7.493
R10218 D.n81 D.t548 7.493
R10219 D.n90 D.t82 7.493
R10220 D.n99 D.t537 7.493
R10221 D.n108 D.t72 7.493
R10222 D.n117 D.t525 7.493
R10223 D.n126 D.t63 7.493
R10224 D.n135 D.t132 7.493
R10225 D.n144 D.t50 7.493
R10226 D.n153 D.t186 7.493
R10227 D.n162 D.t38 7.493
R10228 D.n171 D.t171 7.493
R10229 D.n180 D.t29 7.493
R10230 D.n189 D.t160 7.493
R10231 D.n198 D.t18 7.493
R10232 D.n207 D.t341 7.493
R10233 D.n216 D.t941 7.493
R10234 D.n286 D.t206 7.493
R10235 D.n302 D.t704 7.493
R10236 D.n554 D.t422 7.493
R10237 D.n540 D.t824 7.493
R10238 D.n526 D.t187 7.493
R10239 D.n512 D.t471 7.493
R10240 D.n498 D.t914 7.493
R10241 D.n484 D.t454 7.493
R10242 D.n470 D.t901 7.493
R10243 D.n456 D.t442 7.493
R10244 D.n442 D.t519 7.493
R10245 D.n428 D.t432 7.493
R10246 D.n414 D.t508 7.493
R10247 D.n400 D.t420 7.493
R10248 D.n386 D.t552 7.493
R10249 D.n372 D.t407 7.493
R10250 D.n358 D.t541 7.493
R10251 D.n344 D.t395 7.493
R10252 D.n330 D.t720 7.493
R10253 D.n316 D.t210 7.493
R10254 D.n577 D.t578 7.493
R10255 D.n593 D.t1093 7.493
R10256 D.n817 D.t558 7.493
R10257 D.n803 D.t945 7.493
R10258 D.n789 D.t265 7.493
R10259 D.n775 D.t833 7.493
R10260 D.n761 D.t181 7.493
R10261 D.n747 D.t816 7.493
R10262 D.n733 D.t898 7.493
R10263 D.n719 D.t804 7.493
R10264 D.n705 D.t885 7.493
R10265 D.n691 D.t797 7.493
R10266 D.n677 D.t874 7.493
R10267 D.n663 D.t785 7.493
R10268 D.n649 D.t917 7.493
R10269 D.n635 D.t772 7.493
R10270 D.n621 D.t0 7.493
R10271 D.n607 D.t581 7.493
R10272 D.n840 D.t955 7.493
R10273 D.n856 D.t368 7.493
R10274 D.n1052 D.t648 7.493
R10275 D.n1038 D.t1072 7.493
R10276 D.n1024 D.t416 7.493
R10277 D.n1010 D.t100 7.493
R10278 D.n996 D.t177 7.493
R10279 D.n982 D.t86 7.493
R10280 D.n968 D.t165 7.493
R10281 D.n954 D.t74 7.493
R10282 D.n940 D.t150 7.493
R10283 D.n926 D.t64 7.493
R10284 D.n912 D.t137 7.493
R10285 D.n898 D.t53 7.493
R10286 D.n884 D.t380 7.493
R10287 D.n870 D.t958 7.493
R10288 D.n1075 D.t223 7.493
R10289 D.n1091 D.t743 7.493
R10290 D.n1259 D.t793 7.493
R10291 D.n1245 D.t97 7.493
R10292 D.n1231 D.t639 7.493
R10293 D.n1217 D.t473 7.493
R10294 D.n1203 D.t545 7.493
R10295 D.n1189 D.t457 7.493
R10296 D.n1175 D.t534 7.493
R10297 D.n1161 D.t443 7.493
R10298 D.n1147 D.t520 7.493
R10299 D.n1133 D.t433 7.493
R10300 D.n1119 D.t693 7.493
R10301 D.n1105 D.t227 7.493
R10302 D.n1282 D.t596 7.493
R10303 D.n1298 D.t1064 7.493
R10304 D.n1438 D.t1030 7.493
R10305 D.n1424 D.t213 7.493
R10306 D.n1410 D.t788 7.493
R10307 D.n1396 D.t837 7.493
R10308 D.n1382 D.t912 7.493
R10309 D.n1368 D.t819 7.493
R10310 D.n1354 D.t897 7.493
R10311 D.n1340 D.t806 7.493
R10312 D.n1326 D.t1081 7.493
R10313 D.n1312 D.t609 7.493
R10314 D.n1462 D.t978 7.493
R10315 D.n1478 D.t347 7.493
R10316 D.n1590 D.t65 7.493
R10317 D.n1576 D.t348 7.493
R10318 D.n1562 D.t926 7.493
R10319 D.n1548 D.t103 7.493
R10320 D.n1534 D.t179 7.493
R10321 D.n1520 D.t88 7.493
R10322 D.n1506 D.t361 7.493
R10323 D.n1492 D.t991 7.493
R10324 D.n1614 D.t249 7.493
R10325 D.n1630 D.t722 7.493
R10326 D.n1714 D.t198 7.493
R10327 D.n1700 D.t480 7.493
R10328 D.n1686 D.t1024 7.493
R10329 D.n1672 D.t477 7.493
R10330 D.n1658 D.t734 7.493
R10331 D.n1644 D.t268 7.493
R10332 D.n1738 D.t634 7.493
R10333 D.n1754 D.t6 7.493
R10334 D.n1810 D.t303 7.493
R10335 D.n1796 D.t580 7.493
R10336 D.n1782 D.t944 7.493
R10337 D.n1768 D.t653 7.493
R10338 D.n1833 D.t1023 7.493
R10339 D.n1849 D.t1071 7.493
R10340 D.n1877 D.t215 7.493
R10341 D.n1863 D.t604 7.493
R10342 D.n1925 D.t166 7.099
R10343 D.n1889 D.t26 7.099
R10344 D.n1910 D.t872 7.099
R10345 D.n1900 D.t933 7.099
R10346 D.n233 D.t134 7.099
R10347 D.n224 D.t961 7.099
R10348 D.n31 D.t297 7.099
R10349 D.n2018 D.t194 7.099
R10350 D.n2003 D.t822 7.099
R10351 D.n3557 D.t75 7.099
R10352 D.n3539 D.t1031 7.099
R10353 D.n3521 D.t1046 7.099
R10354 D.n3503 D.t1062 7.099
R10355 D.n3485 D.t1080 7.099
R10356 D.n3467 D.t1016 7.099
R10357 D.n3449 D.t1032 7.099
R10358 D.n3431 D.t1048 7.099
R10359 D.n3413 D.t1065 7.099
R10360 D.n3394 D.t1018 7.099
R10361 D.n3404 D.t339 7.099
R10362 D.n3422 D.t731 7.099
R10363 D.n3440 D.t721 7.099
R10364 D.n3458 D.t706 7.099
R10365 D.n3476 D.t314 7.099
R10366 D.n3494 D.t298 7.099
R10367 D.n3512 D.t279 7.099
R10368 D.n3530 D.t266 7.099
R10369 D.n3548 D.t253 7.099
R10370 D.n3570 D.t599 7.099
R10371 D.n3159 D.t575 7.099
R10372 D.n3179 D.t659 7.099
R10373 D.n3199 D.t674 7.099
R10374 D.n3219 D.t690 7.099
R10375 D.n3239 D.t708 7.099
R10376 D.n3259 D.t642 7.099
R10377 D.n3279 D.t660 7.099
R10378 D.n3299 D.t677 7.099
R10379 D.n3319 D.t647 7.099
R10380 D.n3308 D.t1058 7.099
R10381 D.n3288 D.t358 7.099
R10382 D.n3268 D.t342 7.099
R10383 D.n3248 D.t327 7.099
R10384 D.n3228 D.t1034 7.099
R10385 D.n3208 D.t1019 7.099
R10386 D.n3188 D.t1003 7.099
R10387 D.n3168 D.t994 7.099
R10388 D.n3145 D.t3 7.099
R10389 D.n3074 D.t1094 7.099
R10390 D.n3056 D.t291 7.099
R10391 D.n3038 D.t307 7.099
R10392 D.n3020 D.t326 7.099
R10393 D.n3002 D.t345 7.099
R10394 D.n2984 D.t274 7.099
R10395 D.n2966 D.t292 7.099
R10396 D.n2947 D.t261 7.099
R10397 D.n2957 D.t669 7.099
R10398 D.n2975 D.t1075 7.099
R10399 D.n2993 D.t1061 7.099
R10400 D.n3011 D.t1045 7.099
R10401 D.n3029 D.t644 7.099
R10402 D.n3047 D.t629 7.099
R10403 D.n3065 D.t617 7.099
R10404 D.n3087 D.t521 7.099
R10405 D.n2756 D.t509 7.099
R10406 D.n2776 D.t1028 7.099
R10407 D.n2796 D.t1043 7.099
R10408 D.n2816 D.t1059 7.099
R10409 D.n2836 D.t1077 7.099
R10410 D.n2856 D.t1012 7.099
R10411 D.n2876 D.t988 7.099
R10412 D.n2865 D.t285 7.099
R10413 D.n2845 D.t688 7.099
R10414 D.n2825 D.t671 7.099
R10415 D.n2805 D.t657 7.099
R10416 D.n2785 D.t263 7.099
R10417 D.n2765 D.t248 7.099
R10418 D.n2740 D.t983 7.099
R10419 D.n2675 D.t971 7.099
R10420 D.n2657 D.t658 7.099
R10421 D.n2639 D.t670 7.099
R10422 D.n2621 D.t686 7.099
R10423 D.n2603 D.t705 7.099
R10424 D.n2584 D.t606 7.099
R10425 D.n2594 D.t1008 7.099
R10426 D.n2612 D.t305 7.099
R10427 D.n2630 D.t286 7.099
R10428 D.n2648 D.t270 7.099
R10429 D.n2666 D.t990 7.099
R10430 D.n2687 D.t412 7.099
R10431 D.n2433 D.t397 7.099
R10432 D.n2453 D.t287 7.099
R10433 D.n2473 D.t304 7.099
R10434 D.n2493 D.t320 7.099
R10435 D.n2513 D.t288 7.099
R10436 D.n2502 D.t618 7.099
R10437 D.n2482 D.t1025 7.099
R10438 D.n2462 D.t1006 7.099
R10439 D.n2442 D.t998 7.099
R10440 D.n2417 D.t927 7.099
R10441 D.n2350 D.t918 7.099
R10442 D.n2332 D.t1026 7.099
R10443 D.n2314 D.t1041 7.099
R10444 D.n2295 D.t1010 7.099
R10445 D.n2305 D.t240 7.099
R10446 D.n2323 D.t631 7.099
R10447 D.n2341 D.t621 7.099
R10448 D.n2363 D.t41 7.099
R10449 D.n2184 D.t284 7.099
R10450 D.n2204 D.t656 7.099
R10451 D.n2224 D.t623 7.099
R10452 D.n2213 D.t965 7.099
R10453 D.n2193 D.t252 7.099
R10454 D.n2170 D.t559 7.099
R10455 D.n2111 D.t805 7.099
R10456 D.n2092 D.t243 7.099
R10457 D.n2102 D.t589 7.099
R10458 D.n2124 D.t1042 7.099
R10459 D.n53 D.t784 7.099
R10460 D.n62 D.t561 7.099
R10461 D.n71 D.t14 7.099
R10462 D.n80 D.t329 7.099
R10463 D.n89 D.t4 7.099
R10464 D.n98 D.t315 7.099
R10465 D.n107 D.t1095 7.099
R10466 D.n116 D.t295 7.099
R10467 D.n125 D.t698 7.099
R10468 D.n134 D.t277 7.099
R10469 D.n143 D.t679 7.099
R10470 D.n152 D.t346 7.099
R10471 D.n161 D.t664 7.099
R10472 D.n170 D.t328 7.099
R10473 D.n179 D.t649 7.099
R10474 D.n188 D.t310 7.099
R10475 D.n197 D.t632 7.099
R10476 D.n206 D.t294 7.099
R10477 D.n215 D.t868 7.099
R10478 D.n285 D.t130 7.099
R10479 D.n301 D.t533 7.099
R10480 D.n273 D.t13 7.099
R10481 D.n553 D.t934 7.099
R10482 D.n539 D.t969 7.099
R10483 D.n525 D.t654 7.099
R10484 D.n511 D.t383 7.099
R10485 D.n497 D.t696 7.099
R10486 D.n483 D.t371 7.099
R10487 D.n469 D.t680 7.099
R10488 D.n455 D.t1088 7.099
R10489 D.n441 D.t661 7.099
R10490 D.n427 D.t1069 7.099
R10491 D.n413 D.t646 7.099
R10492 D.n399 D.t1052 7.099
R10493 D.n385 D.t709 7.099
R10494 D.n371 D.t1036 7.099
R10495 D.n357 D.t692 7.099
R10496 D.n343 D.t1021 7.099
R10497 D.n329 D.t676 7.099
R10498 D.n315 D.t145 7.099
R10499 D.n576 D.t517 7.099
R10500 D.n592 D.t906 7.099
R10501 D.n567 D.t209 7.099
R10502 D.n816 D.t1039 7.099
R10503 D.n802 D.t20 7.099
R10504 D.n788 D.t796 7.099
R10505 D.n774 D.t746 7.099
R10506 D.n760 D.t1067 7.099
R10507 D.n746 D.t364 7.099
R10508 D.n732 D.t1053 7.099
R10509 D.n718 D.t352 7.099
R10510 D.n704 D.t1035 7.099
R10511 D.n690 D.t337 7.099
R10512 D.n676 D.t1020 7.099
R10513 D.n662 D.t317 7.099
R10514 D.n648 D.t1086 7.099
R10515 D.n634 D.t300 7.099
R10516 D.n620 D.t1063 7.099
R10517 D.n606 D.t531 7.099
R10518 D.n839 D.t894 7.099
R10519 D.n855 D.t190 7.099
R10520 D.n830 D.t343 7.099
R10521 D.n1051 D.t73 7.099
R10522 D.n1037 D.t158 7.099
R10523 D.n1023 D.t930 7.099
R10524 D.n1009 D.t740 7.099
R10525 D.n995 D.t335 7.099
R10526 D.n981 D.t728 7.099
R10527 D.n967 D.t319 7.099
R10528 D.n953 D.t718 7.099
R10529 D.n939 D.t299 7.099
R10530 D.n925 D.t701 7.099
R10531 D.n911 D.t282 7.099
R10532 D.n897 D.t682 7.099
R10533 D.n883 D.t350 7.099
R10534 D.n869 D.t910 7.099
R10535 D.n1074 D.t176 7.099
R10536 D.n1090 D.t563 7.099
R10537 D.n1065 D.t474 7.099
R10538 D.n1258 D.t202 7.099
R10539 D.n1244 D.t393 7.099
R10540 D.n1230 D.t1033 7.099
R10541 D.n1216 D.t10 7.099
R10542 D.n1202 D.t699 7.099
R10543 D.n1188 D.t1103 7.099
R10544 D.n1174 D.t684 7.099
R10545 D.n1160 D.t1091 7.099
R10546 D.n1146 D.t665 7.099
R10547 D.n1132 D.t1074 7.099
R10548 D.n1118 D.t652 7.099
R10549 D.n1104 D.t189 7.099
R10550 D.n1281 D.t554 7.099
R10551 D.n1297 D.t888 7.099
R10552 D.n1272 D.t716 7.099
R10553 D.n1437 D.t311 7.099
R10554 D.n1423 D.t536 7.099
R10555 D.n1409 D.t66 7.099
R10556 D.n1395 D.t379 7.099
R10557 D.n1381 D.t1070 7.099
R10558 D.n1367 D.t367 7.099
R10559 D.n1353 D.t1057 7.099
R10560 D.n1339 D.t357 7.099
R10561 D.n1325 D.t1038 7.099
R10562 D.n1311 D.t562 7.099
R10563 D.n1461 D.t928 7.099
R10564 D.n1477 D.t169 7.099
R10565 D.n1452 D.t848 7.099
R10566 D.n1589 D.t448 7.099
R10567 D.n1575 D.t613 7.099
R10568 D.n1561 D.t200 7.099
R10569 D.n1547 D.t742 7.099
R10570 D.n1533 D.t338 7.099
R10571 D.n1519 D.t730 7.099
R10572 D.n1505 D.t325 7.099
R10573 D.n1491 D.t936 7.099
R10574 D.n1613 D.t199 7.099
R10575 D.n1629 D.t550 7.099
R10576 D.n1604 D.t954 7.099
R10577 D.n1713 D.t569 7.099
R10578 D.n1699 D.t766 7.099
R10579 D.n1685 D.t306 7.099
R10580 D.n1671 D.t12 7.099
R10581 D.n1657 D.t703 7.099
R10582 D.n1643 D.t205 7.099
R10583 D.n1737 D.t570 7.099
R10584 D.n1753 D.t923 7.099
R10585 D.n1728 D.t1097 7.099
R10586 D.n1809 D.t689 7.099
R10587 D.n1795 D.t905 7.099
R10588 D.n1781 D.t444 7.099
R10589 D.n1767 D.t576 7.099
R10590 D.n1832 D.t946 7.099
R10591 D.n1848 D.t489 7.099
R10592 D.n1823 D.t121 7.099
R10593 D.n1876 D.t820 7.099
R10594 D.n1862 D.t798 7.099
R10595 D.n238 D.t168 7.065
R10596 D.n1893 D.t672 7.065
R10597 D.n1953 D.t966 7.065
R10598 D.n2037 D.t195 7.065
R10599 D.n3370 D.t685 7.065
R10600 D.n3335 D.t302 7.065
R10601 D.n2927 D.t574 7.065
R10602 D.n2892 D.t204 7.065
R10603 D.n2564 D.t932 7.065
R10604 D.n2529 D.t560 7.065
R10605 D.n2275 D.t212 7.065
R10606 D.n2240 D.t942 7.065
R10607 D.n2072 D.t567 7.065
R10608 D.n263 D.t840 7.038
R10609 D.n1926 D.t34 7.037
R10610 D.n1890 D.t986 7.037
R10611 D.n1991 D.t911 7.037
R10612 D.n3585 D.t733 7.037
R10613 D.n3133 D.t370 7.037
R10614 D.n3102 D.t907 7.037
R10615 D.n2725 D.t542 7.037
R10616 D.n2696 D.t173 7.037
R10617 D.n2402 D.t904 7.037
R10618 D.n2378 D.t913 7.037
R10619 D.n2158 D.t547 7.037
R10620 D.n2139 D.t178 7.037
R10621 D.n1970 D.t133 7.037
R10622 D.n274 D.t1078 7.037
R10623 D.n568 D.t104 7.037
R10624 D.n831 D.t216 7.037
R10625 D.n1066 D.t354 7.037
R10626 D.n1273 D.t486 7.037
R10627 D.n1453 D.t583 7.037
R10628 D.n1605 D.t724 7.037
R10629 D.n1729 D.t858 7.037
R10630 D.n1824 D.t957 7.037
R10631 D.n292 D.t551 7.031
R10632 D.n583 D.t925 7.031
R10633 D.n846 D.t197 7.031
R10634 D.n1081 D.t568 7.031
R10635 D.n1288 D.t943 7.031
R10636 D.n1468 D.t214 7.031
R10637 D.n1620 D.t586 7.031
R10638 D.n1744 D.t962 7.031
R10639 D.n1839 D.t233 7.031
R10640 D.n1931 D.t989 7.031
R10641 D.n1908 D.t710 7.007
R10642 D.n1898 D.t239 7.007
R10643 D.n230 D.t1027 7.007
R10644 D.n221 D.t172 7.007
R10645 D.n29 D.t556 7.007
R10646 D.n2016 D.t164 7.007
R10647 D.n2001 D.t418 7.007
R10648 D.n3554 D.t356 7.007
R10649 D.n3536 D.t458 7.007
R10650 D.n3518 D.t475 7.007
R10651 D.n3500 D.t493 7.007
R10652 D.n3482 D.t507 7.007
R10653 D.n3464 D.t447 7.007
R10654 D.n3446 D.t461 7.007
R10655 D.n3428 D.t476 7.007
R10656 D.n3410 D.t494 7.007
R10657 D.n3391 D.t182 7.007
R10658 D.n3402 D.t846 7.007
R10659 D.n3420 D.t149 7.007
R10660 D.n3438 D.t128 7.007
R10661 D.n3456 D.t113 7.007
R10662 D.n3474 D.t99 7.007
R10663 D.n3492 D.t809 7.007
R10664 D.n3510 D.t799 7.007
R10665 D.n3528 D.t791 7.007
R10666 D.n3546 D.t777 7.007
R10667 D.n3568 D.t431 7.007
R10668 D.n3156 D.t869 7.007
R10669 D.n3176 D.t87 7.007
R10670 D.n3196 D.t101 7.007
R10671 D.n3216 D.t116 7.007
R10672 D.n3236 D.t131 7.007
R10673 D.n3256 D.t76 7.007
R10674 D.n3276 D.t89 7.007
R10675 D.n3296 D.t102 7.007
R10676 D.n3316 D.t780 7.007
R10677 D.n3306 D.t467 7.007
R10678 D.n3286 D.t867 7.007
R10679 D.n3266 D.t850 7.007
R10680 D.n3246 D.t831 7.007
R10681 D.n3226 D.t818 7.007
R10682 D.n3206 D.t436 7.007
R10683 D.n3186 D.t427 7.007
R10684 D.n3166 D.t411 7.007
R10685 D.n3143 D.t995 7.007
R10686 D.n3071 D.t232 7.007
R10687 D.n3053 D.t817 7.007
R10688 D.n3035 D.t834 7.007
R10689 D.n3017 D.t852 7.007
R10690 D.n2999 D.t870 7.007
R10691 D.n2981 D.t808 7.007
R10692 D.n2963 D.t823 7.007
R10693 D.n2944 D.t404 7.007
R10694 D.n2955 D.t81 7.007
R10695 D.n2973 D.t485 7.007
R10696 D.n2991 D.t469 7.007
R10697 D.n3009 D.t456 7.007
R10698 D.n3027 D.t441 7.007
R10699 D.n3045 D.t57 7.007
R10700 D.n3063 D.t44 7.007
R10701 D.n3085 D.t402 7.007
R10702 D.n2753 D.t762 7.007
R10703 D.n2773 D.t455 7.007
R10704 D.n2793 D.t472 7.007
R10705 D.n2813 D.t487 7.007
R10706 D.n2833 D.t504 7.007
R10707 D.n2853 D.t445 7.007
R10708 D.n2873 D.t28 7.007
R10709 D.n2863 D.t801 7.007
R10710 D.n2843 D.t95 7.007
R10711 D.n2823 D.t85 7.007
R10712 D.n2803 D.t70 7.007
R10713 D.n2783 D.t62 7.007
R10714 D.n2763 D.t774 7.007
R10715 D.n2738 D.t908 7.007
R10716 D.n2672 D.t184 7.007
R10717 D.n2654 D.t84 7.007
R10718 D.n2636 D.t98 7.007
R10719 D.n2618 D.t112 7.007
R10720 D.n2600 D.t127 7.007
R10721 D.n2581 D.t745 7.007
R10722 D.n2592 D.t428 7.007
R10723 D.n2610 D.t815 7.007
R10724 D.n2628 D.t800 7.007
R10725 D.n2646 D.t794 7.007
R10726 D.n2664 D.t782 7.007
R10727 D.n2685 D.t254 7.007
R10728 D.n2430 D.t650 7.007
R10729 D.n2450 D.t814 7.007
R10730 D.n2470 D.t829 7.007
R10731 D.n2490 D.t849 7.007
R10732 D.n2510 D.t425 7.007
R10733 D.n2500 D.t46 7.007
R10734 D.n2480 D.t438 7.007
R10735 D.n2460 D.t429 7.007
R10736 D.n2440 D.t417 7.007
R10737 D.n2415 D.t1047 7.007
R10738 D.n2347 D.t71 7.007
R10739 D.n2329 D.t452 7.007
R10740 D.n2311 D.t468 7.007
R10741 D.n2292 D.t42 7.007
R10742 D.n2303 D.t768 7.007
R10743 D.n2321 D.t59 7.007
R10744 D.n2339 D.t47 7.007
R10745 D.n2361 D.t446 7.007
R10746 D.n2181 D.t572 7.007
R10747 D.n2201 D.t79 7.007
R10748 D.n2221 D.t764 7.007
R10749 D.n2211 D.t392 7.007
R10750 D.n2191 D.t778 7.007
R10751 D.n2168 D.t938 7.007
R10752 D.n2108 D.t1085 7.007
R10753 D.n2089 D.t388 7.007
R10754 D.n2100 D.t16 7.007
R10755 D.n2122 D.t313 7.007
R10756 D.n51 D.t139 7.007
R10757 D.n60 D.t405 7.007
R10758 D.n69 D.t530 7.007
R10759 D.n78 D.t855 7.007
R10760 D.n87 D.t515 7.007
R10761 D.n96 D.t839 7.007
R10762 D.n105 D.t505 7.007
R10763 D.n114 D.t825 7.007
R10764 D.n123 D.t488 7.007
R10765 D.n132 D.t810 7.007
R10766 D.n141 D.t90 7.007
R10767 D.n150 D.t873 7.007
R10768 D.n159 D.t77 7.007
R10769 D.n168 D.t854 7.007
R10770 D.n177 D.t67 7.007
R10771 D.n186 D.t838 7.007
R10772 D.n195 D.t60 7.007
R10773 D.n204 D.t821 7.007
R10774 D.n213 D.t226 7.007
R10775 D.n290 D.t749 7.007
R10776 D.n282 D.t595 7.007
R10777 D.n298 D.t1007 7.007
R10778 D.n550 D.t781 7.007
R10779 D.n536 D.t331 7.007
R10780 D.n522 D.t549 7.007
R10781 D.n508 D.t892 7.007
R10782 D.n494 D.t120 7.007
R10783 D.n480 D.t882 7.007
R10784 D.n466 D.t106 7.007
R10785 D.n452 D.t871 7.007
R10786 D.n438 D.t91 7.007
R10787 D.n424 D.t478 7.007
R10788 D.n410 D.t78 7.007
R10789 D.n396 D.t462 7.007
R10790 D.n382 D.t136 7.007
R10791 D.n368 D.t449 7.007
R10792 D.n354 D.t117 7.007
R10793 D.n340 D.t439 7.007
R10794 D.n326 D.t105 7.007
R10795 D.n312 D.t608 7.007
R10796 D.n581 D.t271 7.007
R10797 D.n573 D.t977 7.007
R10798 D.n589 D.t283 7.007
R10799 D.n813 D.t922 7.007
R10800 D.n799 D.t465 7.007
R10801 D.n785 D.t625 7.007
R10802 D.n771 D.t162 7.007
R10803 D.n757 D.t497 7.007
R10804 D.n743 D.t148 7.007
R10805 D.n729 D.t479 7.007
R10806 D.n715 D.t861 7.007
R10807 D.n701 D.t463 7.007
R10808 D.n687 D.t841 7.007
R10809 D.n673 D.t450 7.007
R10810 D.n659 D.t826 7.007
R10811 D.n645 D.t510 7.007
R10812 D.n631 D.t811 7.007
R10813 D.n617 D.t495 7.007
R10814 D.n603 D.t993 7.007
R10815 D.n844 D.t655 7.007
R10816 D.n836 D.t251 7.007
R10817 D.n852 D.t668 7.007
R10818 D.n1048 D.t1014 7.007
R10819 D.n1034 D.t577 7.007
R10820 D.n1020 D.t776 7.007
R10821 D.n1006 D.t535 7.007
R10822 D.n992 D.t857 7.007
R10823 D.n978 D.t142 7.007
R10824 D.n964 D.t842 7.007
R10825 D.n950 D.t124 7.007
R10826 D.n936 D.t827 7.007
R10827 D.n922 D.t109 7.007
R10828 D.n908 D.t812 7.007
R10829 D.n894 D.t92 7.007
R10830 D.n880 D.t875 7.007
R10831 D.n866 D.t267 7.007
R10832 D.n1079 D.t1040 7.007
R10833 D.n1071 D.t633 7.007
R10834 D.n1087 D.t1056 7.007
R10835 D.n1255 D.t56 7.007
R10836 D.n1241 D.t707 7.007
R10837 D.n1227 D.t920 7.007
R10838 D.n1213 D.t526 7.007
R10839 D.n1199 D.t123 7.007
R10840 D.n1185 D.t513 7.007
R10841 D.n1171 D.t110 7.007
R10842 D.n1157 D.t502 7.007
R10843 D.n1143 D.t93 7.007
R10844 D.n1129 D.t482 7.007
R10845 D.n1115 D.t80 7.007
R10846 D.n1101 D.t651 7.007
R10847 D.n1286 D.t324 7.007
R10848 D.n1278 D.t1022 7.007
R10849 D.n1294 D.t258 7.007
R10850 D.n1434 D.t193 7.007
R10851 D.n1420 D.t951 7.007
R10852 D.n1406 D.t1009 7.007
R10853 D.n1392 D.t890 7.007
R10854 D.n1378 D.t501 7.007
R10855 D.n1364 D.t879 7.007
R10856 D.n1350 D.t483 7.007
R10857 D.n1336 D.t866 7.007
R10858 D.n1322 D.t466 7.007
R10859 D.n1308 D.t1037 7.007
R10860 D.n1466 D.t624 7.007
R10861 D.n1458 D.t301 7.007
R10862 D.n1474 D.t638 7.007
R10863 D.n1586 D.t290 7.007
R10864 D.n1572 D.t1089 7.007
R10865 D.n1558 D.t52 7.007
R10866 D.n1544 D.t157 7.007
R10867 D.n1530 D.t862 7.007
R10868 D.n1516 D.t144 7.007
R10869 D.n1502 D.t845 7.007
R10870 D.n1488 D.t318 7.007
R10871 D.n1618 D.t1013 7.007
R10872 D.n1610 D.t683 7.007
R10873 D.n1626 D.t1029 7.007
R10874 D.n1710 D.t435 7.007
R10875 D.n1696 D.t111 7.007
R10876 D.n1682 D.t192 7.007
R10877 D.n1668 D.t529 7.007
R10878 D.n1654 D.t125 7.007
R10879 D.n1640 D.t702 7.007
R10880 D.n1742 D.t293 7.007
R10881 D.n1734 D.t1076 7.007
R10882 D.n1750 D.t309 7.007
R10883 D.n1806 D.t565 7.007
R10884 D.n1792 D.t218 7.007
R10885 D.n1778 D.t278 7.007
R10886 D.n1764 D.t1092 7.007
R10887 D.n1837 D.t675 7.007
R10888 D.n1829 D.t359 7.007
R10889 D.n1845 D.t330 7.007
R10890 D.n1873 D.t667 7.007
R10891 D.n1859 D.t159 7.007
R10892 D.n1892 D.t464 7.007
R10893 D.n1929 D.t843 7.007
R10894 D.n291 D.t492 6.598
R10895 D.n582 D.t896 6.598
R10896 D.n845 D.t174 6.598
R10897 D.n1080 D.t555 6.598
R10898 D.n1287 D.t929 6.598
R10899 D.n1467 D.t152 6.598
R10900 D.n1619 D.t539 6.598
R10901 D.n1743 D.t916 6.598
R10902 D.n1838 D.t191 6.598
R10903 D.n1930 D.t960 6.598
R10904 D.n263 D.t723 6.568
R10905 D.n1954 D.t636 6.564
R10906 D.n2038 D.t940 6.564
R10907 D.n3371 D.t400 6.564
R10908 D.n3336 D.t643 6.564
R10909 D.n2928 D.t262 6.564
R10910 D.n2893 D.t985 6.564
R10911 D.n2565 D.t602 6.564
R10912 D.n2530 D.t224 6.564
R10913 D.n2276 D.t956 6.564
R10914 D.n2241 D.t579 6.564
R10915 D.n2073 D.t208 6.564
R10916 D.n1894 D.t584 6.564
R10917 D.n238 D.t308 6.528
R10918 D.n1924 D.t616 6.524
R10919 D.n1891 D.t540 6.524
R10920 D.n1989 D.t115 6.524
R10921 D.n3583 D.t1044 6.524
R10922 D.n3134 D.t860 6.524
R10923 D.n3100 D.t499 6.524
R10924 D.n2726 D.t122 6.524
R10925 D.n2697 D.t856 6.524
R10926 D.n2403 D.t496 6.524
R10927 D.n2376 D.t118 6.524
R10928 D.n2159 D.t853 6.524
R10929 D.n2137 D.t491 6.524
R10930 D.n1971 D.t414 6.524
R10931 D.n275 D.t523 6.524
R10932 D.n569 D.t711 6.524
R10933 D.n832 D.t844 6.524
R10934 D.n1067 D.t953 6.524
R10935 D.n1274 D.t1096 6.524
R10936 D.n1454 D.t221 6.524
R10937 D.n1606 D.t365 6.524
R10938 D.n1730 D.t503 6.524
R10939 D.n1825 D.t588 6.524
R10940 D.n1918 D.n1915 0.344
R10941 D.n1451 D.n1450 0.327
R10942 D.n1603 D.n1602 0.327
R10943 D.n1727 D.n1726 0.327
R10944 D.n268 D.n267 0.31
R10945 D.n1918 D.n1917 0.225
R10946 D.n280 D.n279 0.225
R10947 D.n571 D.n570 0.225
R10948 D.n834 D.n833 0.225
R10949 D.n1069 D.n1068 0.225
R10950 D.n1276 D.n1275 0.225
R10951 D.n1456 D.n1455 0.225
R10952 D.n1608 D.n1607 0.225
R10953 D.n1732 D.n1731 0.225
R10954 D.n1827 D.n1826 0.225
R10955 D.n1920 D.n1919 0.225
R10956 D.n3574 D.n3573 0.21
R10957 D.n3151 D.n3150 0.21
R10958 D.n2748 D.n2747 0.21
R10959 D.n2691 D.n2690 0.21
R10960 D.n2425 D.n2424 0.21
R10961 D.n2176 D.n2175 0.21
R10962 D.n2011 D.n2010 0.21
R10963 D.n1980 D.n1979 0.205
R10964 D.n1951 D.n1950 0.192
R10965 D.n1958 D.n1957 0.174
R10966 D.n1982 D.n1981 0.163
R10967 D.n1934 D.n1933 0.144
R10968 D.n2048 D.n2047 0.143
R10969 D.n3389 D.n3355 0.143
R10970 D.n3389 D.n3388 0.143
R10971 D.n3346 D.n3129 0.143
R10972 D.n3346 D.n3345 0.143
R10973 D.n2942 D.n2912 0.143
R10974 D.n2942 D.n2941 0.143
R10975 D.n2903 D.n2720 0.143
R10976 D.n2903 D.n2902 0.143
R10977 D.n2579 D.n2549 0.143
R10978 D.n2579 D.n2578 0.143
R10979 D.n2540 D.n2397 0.143
R10980 D.n2540 D.n2539 0.143
R10981 D.n2290 D.n2260 0.143
R10982 D.n2290 D.n2289 0.143
R10983 D.n2251 D.n2154 0.143
R10984 D.n2251 D.n2250 0.143
R10985 D.n2087 D.n2057 0.143
R10986 D.n2087 D.n2086 0.143
R10987 D.n2048 D.n1983 0.143
R10988 D.n1962 D.n1961 0.143
R10989 D.n3140 D.n3130 0.14
R10990 D.n2165 D.n2155 0.14
R10991 D.n1960 D.n1958 0.133
R10992 D.n3612 D.n3611 0.133
R10993 D.n3125 D.n3124 0.133
R10994 D.n2716 D.n2715 0.133
R10995 D.n2393 D.n2392 0.133
R10996 D.n2150 D.n2149 0.133
R10997 D.n3580 D.n3577 0.131
R10998 D.n3589 D.n3588 0.131
R10999 D.n3097 D.n3093 0.131
R11000 D.n3106 D.n3105 0.131
R11001 D.n2373 D.n2369 0.131
R11002 D.n2382 D.n2381 0.131
R11003 D.n2134 D.n2130 0.131
R11004 D.n2143 D.n2142 0.131
R11005 D.n1997 D.n1996 0.123
R11006 D.n2734 D.n2733 0.123
R11007 D.n2411 D.n2410 0.123
R11008 D.n3138 D.n3137 0.115
R11009 D.n2702 D.n2701 0.115
R11010 D.n2163 D.n2162 0.115
R11011 D.n1934 D.n1922 0.115
R11012 D.n3333 D.n3324 0.113
R11013 D.n2890 D.n2881 0.113
R11014 D.n2527 D.n2518 0.113
R11015 D.n2238 D.n2229 0.113
R11016 D.n2033 D.n2024 0.113
R11017 D.n1943 D.n565 0.111
R11018 D.n1942 D.n828 0.111
R11019 D.n1941 D.n1063 0.111
R11020 D.n1940 D.n1270 0.111
R11021 D.n1939 D.n1449 0.111
R11022 D.n1938 D.n1601 0.111
R11023 D.n1937 D.n1725 0.111
R11024 D.n1936 D.n1821 0.111
R11025 D.n1935 D.n1888 0.11
R11026 D.n1998 D.n1985 0.109
R11027 D.n3565 D.n3562 0.109
R11028 D.n3082 D.n3079 0.109
R11029 D.n2735 D.n2722 0.109
R11030 D.n2412 D.n2399 0.109
R11031 D.n2358 D.n2355 0.109
R11032 D.n2119 D.n2116 0.109
R11033 D.n1947 D.n1945 0.109
R11034 D.n2010 D.n2007 0.109
R11035 D.n2747 D.n2744 0.109
R11036 D.n2424 D.n2421 0.109
R11037 D.n3352 D.n3351 0.105
R11038 D.n2909 D.n2908 0.105
R11039 D.n2546 D.n2545 0.105
R11040 D.n2257 D.n2256 0.105
R11041 D.n2054 D.n2053 0.105
R11042 D.n3354 D.n3353 0.105
R11043 D.n2911 D.n2910 0.105
R11044 D.n2548 D.n2547 0.105
R11045 D.n2259 D.n2258 0.105
R11046 D.n2056 D.n2055 0.105
R11047 D.n1988 D.n1987 0.102
R11048 D.n3587 D.n3586 0.102
R11049 D.n3582 D.n3581 0.102
R11050 D.n3104 D.n3103 0.102
R11051 D.n3099 D.n3098 0.102
R11052 D.n2728 D.n2727 0.102
R11053 D.n2405 D.n2404 0.102
R11054 D.n2380 D.n2379 0.102
R11055 D.n2375 D.n2374 0.102
R11056 D.n2141 D.n2140 0.102
R11057 D.n2136 D.n2135 0.102
R11058 D.n1973 D.n1972 0.102
R11059 D.n1979 D.n1964 0.101
R11060 D.n3376 D.n3375 0.096
R11061 D.n278 D.n277 0.092
R11062 D.n10 D.n9 0.092
R11063 D.n268 D.n265 0.091
R11064 D.n1944 D.n271 0.085
R11065 D.n3580 D.n3579 0.084
R11066 D.n3097 D.n3096 0.084
R11067 D.n2732 D.n2731 0.084
R11068 D.n2409 D.n2408 0.084
R11069 D.n2373 D.n2372 0.084
R11070 D.n2134 D.n2133 0.084
R11071 D.n1995 D.n1994 0.084
R11072 D.n240 D.n239 0.079
R11073 D.n3566 D.n3565 0.078
R11074 D.n3153 D.n3140 0.078
R11075 D.n3083 D.n3082 0.078
R11076 D.n2750 D.n2735 0.078
R11077 D.n2683 D.n2682 0.078
R11078 D.n2427 D.n2412 0.078
R11079 D.n2359 D.n2358 0.078
R11080 D.n2178 D.n2165 0.078
R11081 D.n2120 D.n2119 0.078
R11082 D.n2013 D.n1998 0.078
R11083 D.n1933 D.n1932 0.077
R11084 D.n1905 D.n1895 0.077
R11085 D.n3136 D.n3135 0.077
R11086 D.n2699 D.n2698 0.077
R11087 D.n2694 D.n2693 0.077
R11088 D.n2161 D.n2160 0.077
R11089 D.n3 D.n2 0.075
R11090 D.n24 D.n16 0.075
R11091 D.n3323 D.n3313 0.074
R11092 D.n3303 D.n3293 0.074
R11093 D.n3283 D.n3273 0.074
R11094 D.n3263 D.n3253 0.074
R11095 D.n3243 D.n3233 0.074
R11096 D.n3223 D.n3213 0.074
R11097 D.n3203 D.n3193 0.074
R11098 D.n3183 D.n3173 0.074
R11099 D.n2880 D.n2870 0.074
R11100 D.n2860 D.n2850 0.074
R11101 D.n2840 D.n2830 0.074
R11102 D.n2820 D.n2810 0.074
R11103 D.n2800 D.n2790 0.074
R11104 D.n2780 D.n2770 0.074
R11105 D.n2517 D.n2507 0.074
R11106 D.n2497 D.n2487 0.074
R11107 D.n2477 D.n2467 0.074
R11108 D.n2457 D.n2447 0.074
R11109 D.n2228 D.n2218 0.074
R11110 D.n2208 D.n2198 0.074
R11111 D.n2043 D.n2042 0.073
R11112 D.n3364 D.n3363 0.073
R11113 D.n3363 D.n3362 0.073
R11114 D.n3384 D.n3383 0.073
R11115 D.n3383 D.n3382 0.073
R11116 D.n3329 D.n3328 0.073
R11117 D.n3341 D.n3340 0.073
R11118 D.n2921 D.n2920 0.073
R11119 D.n2920 D.n2919 0.073
R11120 D.n2937 D.n2936 0.073
R11121 D.n2936 D.n2935 0.073
R11122 D.n2886 D.n2885 0.073
R11123 D.n2898 D.n2897 0.073
R11124 D.n2558 D.n2557 0.073
R11125 D.n2557 D.n2556 0.073
R11126 D.n2574 D.n2573 0.073
R11127 D.n2573 D.n2572 0.073
R11128 D.n2523 D.n2522 0.073
R11129 D.n2535 D.n2534 0.073
R11130 D.n2269 D.n2268 0.073
R11131 D.n2268 D.n2267 0.073
R11132 D.n2285 D.n2284 0.073
R11133 D.n2284 D.n2283 0.073
R11134 D.n2234 D.n2233 0.073
R11135 D.n2246 D.n2245 0.073
R11136 D.n2066 D.n2065 0.073
R11137 D.n2065 D.n2064 0.073
R11138 D.n2082 D.n2081 0.073
R11139 D.n2081 D.n2080 0.073
R11140 D.n2029 D.n2028 0.073
R11141 D.n3163 D.n3153 0.073
R11142 D.n2760 D.n2750 0.073
R11143 D.n2437 D.n2427 0.073
R11144 D.n2188 D.n2178 0.073
R11145 D.n2703 D.n2702 0.072
R11146 D.n42 D.n34 0.072
R11147 D.n2023 D.n2013 0.072
R11148 D.n1915 D.n1905 0.072
R11149 D.n3173 D.n3163 0.072
R11150 D.n3193 D.n3183 0.072
R11151 D.n3213 D.n3203 0.072
R11152 D.n3233 D.n3223 0.072
R11153 D.n3253 D.n3243 0.072
R11154 D.n3273 D.n3263 0.072
R11155 D.n3293 D.n3283 0.072
R11156 D.n3313 D.n3303 0.072
R11157 D.n2770 D.n2760 0.072
R11158 D.n2790 D.n2780 0.072
R11159 D.n2810 D.n2800 0.072
R11160 D.n2830 D.n2820 0.072
R11161 D.n2850 D.n2840 0.072
R11162 D.n2870 D.n2860 0.072
R11163 D.n2447 D.n2437 0.072
R11164 D.n2467 D.n2457 0.072
R11165 D.n2487 D.n2477 0.072
R11166 D.n2507 D.n2497 0.072
R11167 D.n2198 D.n2188 0.072
R11168 D.n2218 D.n2208 0.072
R11169 D.n3591 D.n3590 0.071
R11170 D.n46 D.n45 0.068
R11171 D.n10 D.n3 0.064
R11172 D.n268 D.n12 0.06
R11173 D.n3108 D.n3107 0.059
R11174 D.n2384 D.n2383 0.059
R11175 D.n2145 D.n2144 0.059
R11176 D.n3614 D.n3613 0.057
R11177 D.n294 D.n293 0.056
R11178 D.n585 D.n584 0.056
R11179 D.n848 D.n847 0.056
R11180 D.n1083 D.n1082 0.056
R11181 D.n1290 D.n1289 0.056
R11182 D.n1470 D.n1469 0.056
R11183 D.n1622 D.n1621 0.056
R11184 D.n1746 D.n1745 0.056
R11185 D.n1841 D.n1840 0.056
R11186 D.n12 D.n10 0.055
R11187 D.n277 D.n276 0.055
R11188 D.n1880 D.n1879 0.055
R11189 D.n1960 D.n1959 0.053
R11190 D.n1882 D.n1881 0.053
R11191 D.n49 D.n48 0.053
R11192 D.n2024 D.n2023 0.053
R11193 D.n3398 D.n3397 0.053
R11194 D.n3324 D.n3323 0.053
R11195 D.n2951 D.n2950 0.053
R11196 D.n2881 D.n2880 0.053
R11197 D.n2588 D.n2587 0.053
R11198 D.n2518 D.n2517 0.053
R11199 D.n2299 D.n2298 0.053
R11200 D.n2229 D.n2228 0.053
R11201 D.n2096 D.n2095 0.053
R11202 D.n1912 D.n1911 0.052
R11203 D.n1902 D.n1901 0.052
R11204 D.n235 D.n234 0.052
R11205 D.n226 D.n225 0.052
R11206 D.n33 D.n32 0.052
R11207 D.n2020 D.n2019 0.052
R11208 D.n2005 D.n2004 0.052
R11209 D.n3559 D.n3558 0.052
R11210 D.n3541 D.n3540 0.052
R11211 D.n3523 D.n3522 0.052
R11212 D.n3505 D.n3504 0.052
R11213 D.n3487 D.n3486 0.052
R11214 D.n3469 D.n3468 0.052
R11215 D.n3451 D.n3450 0.052
R11216 D.n3433 D.n3432 0.052
R11217 D.n3415 D.n3414 0.052
R11218 D.n3396 D.n3395 0.052
R11219 D.n3406 D.n3405 0.052
R11220 D.n3424 D.n3423 0.052
R11221 D.n3442 D.n3441 0.052
R11222 D.n3460 D.n3459 0.052
R11223 D.n3478 D.n3477 0.052
R11224 D.n3496 D.n3495 0.052
R11225 D.n3514 D.n3513 0.052
R11226 D.n3532 D.n3531 0.052
R11227 D.n3550 D.n3549 0.052
R11228 D.n3572 D.n3571 0.052
R11229 D.n3161 D.n3160 0.052
R11230 D.n3181 D.n3180 0.052
R11231 D.n3201 D.n3200 0.052
R11232 D.n3221 D.n3220 0.052
R11233 D.n3241 D.n3240 0.052
R11234 D.n3261 D.n3260 0.052
R11235 D.n3281 D.n3280 0.052
R11236 D.n3301 D.n3300 0.052
R11237 D.n3321 D.n3320 0.052
R11238 D.n3310 D.n3309 0.052
R11239 D.n3290 D.n3289 0.052
R11240 D.n3270 D.n3269 0.052
R11241 D.n3250 D.n3249 0.052
R11242 D.n3230 D.n3229 0.052
R11243 D.n3210 D.n3209 0.052
R11244 D.n3190 D.n3189 0.052
R11245 D.n3170 D.n3169 0.052
R11246 D.n3147 D.n3146 0.052
R11247 D.n3076 D.n3075 0.052
R11248 D.n3058 D.n3057 0.052
R11249 D.n3040 D.n3039 0.052
R11250 D.n3022 D.n3021 0.052
R11251 D.n3004 D.n3003 0.052
R11252 D.n2986 D.n2985 0.052
R11253 D.n2968 D.n2967 0.052
R11254 D.n2949 D.n2948 0.052
R11255 D.n2959 D.n2958 0.052
R11256 D.n2977 D.n2976 0.052
R11257 D.n2995 D.n2994 0.052
R11258 D.n3013 D.n3012 0.052
R11259 D.n3031 D.n3030 0.052
R11260 D.n3049 D.n3048 0.052
R11261 D.n3067 D.n3066 0.052
R11262 D.n3089 D.n3088 0.052
R11263 D.n2758 D.n2757 0.052
R11264 D.n2778 D.n2777 0.052
R11265 D.n2798 D.n2797 0.052
R11266 D.n2818 D.n2817 0.052
R11267 D.n2838 D.n2837 0.052
R11268 D.n2858 D.n2857 0.052
R11269 D.n2878 D.n2877 0.052
R11270 D.n2867 D.n2866 0.052
R11271 D.n2847 D.n2846 0.052
R11272 D.n2827 D.n2826 0.052
R11273 D.n2807 D.n2806 0.052
R11274 D.n2787 D.n2786 0.052
R11275 D.n2767 D.n2766 0.052
R11276 D.n2742 D.n2741 0.052
R11277 D.n2677 D.n2676 0.052
R11278 D.n2659 D.n2658 0.052
R11279 D.n2641 D.n2640 0.052
R11280 D.n2623 D.n2622 0.052
R11281 D.n2605 D.n2604 0.052
R11282 D.n2586 D.n2585 0.052
R11283 D.n2596 D.n2595 0.052
R11284 D.n2614 D.n2613 0.052
R11285 D.n2632 D.n2631 0.052
R11286 D.n2650 D.n2649 0.052
R11287 D.n2668 D.n2667 0.052
R11288 D.n2689 D.n2688 0.052
R11289 D.n2435 D.n2434 0.052
R11290 D.n2455 D.n2454 0.052
R11291 D.n2475 D.n2474 0.052
R11292 D.n2495 D.n2494 0.052
R11293 D.n2515 D.n2514 0.052
R11294 D.n2504 D.n2503 0.052
R11295 D.n2484 D.n2483 0.052
R11296 D.n2464 D.n2463 0.052
R11297 D.n2444 D.n2443 0.052
R11298 D.n2419 D.n2418 0.052
R11299 D.n2352 D.n2351 0.052
R11300 D.n2334 D.n2333 0.052
R11301 D.n2316 D.n2315 0.052
R11302 D.n2297 D.n2296 0.052
R11303 D.n2307 D.n2306 0.052
R11304 D.n2325 D.n2324 0.052
R11305 D.n2343 D.n2342 0.052
R11306 D.n2365 D.n2364 0.052
R11307 D.n2186 D.n2185 0.052
R11308 D.n2206 D.n2205 0.052
R11309 D.n2226 D.n2225 0.052
R11310 D.n2215 D.n2214 0.052
R11311 D.n2195 D.n2194 0.052
R11312 D.n2172 D.n2171 0.052
R11313 D.n2113 D.n2112 0.052
R11314 D.n2094 D.n2093 0.052
R11315 D.n2104 D.n2103 0.052
R11316 D.n2126 D.n2125 0.052
R11317 D.n55 D.n54 0.052
R11318 D.n64 D.n63 0.052
R11319 D.n73 D.n72 0.052
R11320 D.n82 D.n81 0.052
R11321 D.n91 D.n90 0.052
R11322 D.n100 D.n99 0.052
R11323 D.n109 D.n108 0.052
R11324 D.n118 D.n117 0.052
R11325 D.n127 D.n126 0.052
R11326 D.n136 D.n135 0.052
R11327 D.n145 D.n144 0.052
R11328 D.n154 D.n153 0.052
R11329 D.n163 D.n162 0.052
R11330 D.n172 D.n171 0.052
R11331 D.n181 D.n180 0.052
R11332 D.n190 D.n189 0.052
R11333 D.n199 D.n198 0.052
R11334 D.n208 D.n207 0.052
R11335 D.n217 D.n216 0.052
R11336 D.n287 D.n286 0.052
R11337 D.n303 D.n302 0.052
R11338 D.n555 D.n554 0.052
R11339 D.n541 D.n540 0.052
R11340 D.n527 D.n526 0.052
R11341 D.n513 D.n512 0.052
R11342 D.n499 D.n498 0.052
R11343 D.n485 D.n484 0.052
R11344 D.n471 D.n470 0.052
R11345 D.n457 D.n456 0.052
R11346 D.n443 D.n442 0.052
R11347 D.n429 D.n428 0.052
R11348 D.n415 D.n414 0.052
R11349 D.n401 D.n400 0.052
R11350 D.n387 D.n386 0.052
R11351 D.n373 D.n372 0.052
R11352 D.n359 D.n358 0.052
R11353 D.n345 D.n344 0.052
R11354 D.n331 D.n330 0.052
R11355 D.n317 D.n316 0.052
R11356 D.n578 D.n577 0.052
R11357 D.n594 D.n593 0.052
R11358 D.n818 D.n817 0.052
R11359 D.n804 D.n803 0.052
R11360 D.n790 D.n789 0.052
R11361 D.n776 D.n775 0.052
R11362 D.n762 D.n761 0.052
R11363 D.n748 D.n747 0.052
R11364 D.n734 D.n733 0.052
R11365 D.n720 D.n719 0.052
R11366 D.n706 D.n705 0.052
R11367 D.n692 D.n691 0.052
R11368 D.n678 D.n677 0.052
R11369 D.n664 D.n663 0.052
R11370 D.n650 D.n649 0.052
R11371 D.n636 D.n635 0.052
R11372 D.n622 D.n621 0.052
R11373 D.n608 D.n607 0.052
R11374 D.n841 D.n840 0.052
R11375 D.n857 D.n856 0.052
R11376 D.n1053 D.n1052 0.052
R11377 D.n1039 D.n1038 0.052
R11378 D.n1025 D.n1024 0.052
R11379 D.n1011 D.n1010 0.052
R11380 D.n997 D.n996 0.052
R11381 D.n983 D.n982 0.052
R11382 D.n969 D.n968 0.052
R11383 D.n955 D.n954 0.052
R11384 D.n941 D.n940 0.052
R11385 D.n927 D.n926 0.052
R11386 D.n913 D.n912 0.052
R11387 D.n899 D.n898 0.052
R11388 D.n885 D.n884 0.052
R11389 D.n871 D.n870 0.052
R11390 D.n1076 D.n1075 0.052
R11391 D.n1092 D.n1091 0.052
R11392 D.n1260 D.n1259 0.052
R11393 D.n1246 D.n1245 0.052
R11394 D.n1232 D.n1231 0.052
R11395 D.n1218 D.n1217 0.052
R11396 D.n1204 D.n1203 0.052
R11397 D.n1190 D.n1189 0.052
R11398 D.n1176 D.n1175 0.052
R11399 D.n1162 D.n1161 0.052
R11400 D.n1148 D.n1147 0.052
R11401 D.n1134 D.n1133 0.052
R11402 D.n1120 D.n1119 0.052
R11403 D.n1106 D.n1105 0.052
R11404 D.n1283 D.n1282 0.052
R11405 D.n1299 D.n1298 0.052
R11406 D.n1439 D.n1438 0.052
R11407 D.n1425 D.n1424 0.052
R11408 D.n1411 D.n1410 0.052
R11409 D.n1397 D.n1396 0.052
R11410 D.n1383 D.n1382 0.052
R11411 D.n1369 D.n1368 0.052
R11412 D.n1355 D.n1354 0.052
R11413 D.n1341 D.n1340 0.052
R11414 D.n1327 D.n1326 0.052
R11415 D.n1313 D.n1312 0.052
R11416 D.n1463 D.n1462 0.052
R11417 D.n1479 D.n1478 0.052
R11418 D.n1591 D.n1590 0.052
R11419 D.n1577 D.n1576 0.052
R11420 D.n1563 D.n1562 0.052
R11421 D.n1549 D.n1548 0.052
R11422 D.n1535 D.n1534 0.052
R11423 D.n1521 D.n1520 0.052
R11424 D.n1507 D.n1506 0.052
R11425 D.n1493 D.n1492 0.052
R11426 D.n1615 D.n1614 0.052
R11427 D.n1631 D.n1630 0.052
R11428 D.n1715 D.n1714 0.052
R11429 D.n1701 D.n1700 0.052
R11430 D.n1687 D.n1686 0.052
R11431 D.n1673 D.n1672 0.052
R11432 D.n1659 D.n1658 0.052
R11433 D.n1645 D.n1644 0.052
R11434 D.n1739 D.n1738 0.052
R11435 D.n1755 D.n1754 0.052
R11436 D.n1811 D.n1810 0.052
R11437 D.n1797 D.n1796 0.052
R11438 D.n1783 D.n1782 0.052
R11439 D.n1769 D.n1768 0.052
R11440 D.n1834 D.n1833 0.052
R11441 D.n1850 D.n1849 0.052
R11442 D.n1878 D.n1877 0.052
R11443 D.n1864 D.n1863 0.052
R11444 D.n1917 D.n1916 0.051
R11445 D.n5 D.n4 0.051
R11446 D.n6 D.n5 0.051
R11447 D.n7 D.n6 0.051
R11448 D.n8 D.n7 0.051
R11449 D.n9 D.n8 0.051
R11450 D.n279 D.n278 0.051
R11451 D.n1909 D.n1908 0.051
R11452 D.n1899 D.n1898 0.051
R11453 D.n232 D.n230 0.051
R11454 D.n223 D.n221 0.051
R11455 D.n30 D.n29 0.051
R11456 D.n2017 D.n2016 0.051
R11457 D.n2002 D.n2001 0.051
R11458 D.n3556 D.n3554 0.051
R11459 D.n3538 D.n3536 0.051
R11460 D.n3520 D.n3518 0.051
R11461 D.n3502 D.n3500 0.051
R11462 D.n3484 D.n3482 0.051
R11463 D.n3466 D.n3464 0.051
R11464 D.n3448 D.n3446 0.051
R11465 D.n3430 D.n3428 0.051
R11466 D.n3412 D.n3410 0.051
R11467 D.n3393 D.n3391 0.051
R11468 D.n3403 D.n3402 0.051
R11469 D.n3421 D.n3420 0.051
R11470 D.n3439 D.n3438 0.051
R11471 D.n3457 D.n3456 0.051
R11472 D.n3475 D.n3474 0.051
R11473 D.n3493 D.n3492 0.051
R11474 D.n3511 D.n3510 0.051
R11475 D.n3529 D.n3528 0.051
R11476 D.n3547 D.n3546 0.051
R11477 D.n3569 D.n3568 0.051
R11478 D.n3158 D.n3156 0.051
R11479 D.n3178 D.n3176 0.051
R11480 D.n3198 D.n3196 0.051
R11481 D.n3218 D.n3216 0.051
R11482 D.n3238 D.n3236 0.051
R11483 D.n3258 D.n3256 0.051
R11484 D.n3278 D.n3276 0.051
R11485 D.n3298 D.n3296 0.051
R11486 D.n3318 D.n3316 0.051
R11487 D.n3307 D.n3306 0.051
R11488 D.n3287 D.n3286 0.051
R11489 D.n3267 D.n3266 0.051
R11490 D.n3247 D.n3246 0.051
R11491 D.n3227 D.n3226 0.051
R11492 D.n3207 D.n3206 0.051
R11493 D.n3187 D.n3186 0.051
R11494 D.n3167 D.n3166 0.051
R11495 D.n3144 D.n3143 0.051
R11496 D.n3073 D.n3071 0.051
R11497 D.n3055 D.n3053 0.051
R11498 D.n3037 D.n3035 0.051
R11499 D.n3019 D.n3017 0.051
R11500 D.n3001 D.n2999 0.051
R11501 D.n2983 D.n2981 0.051
R11502 D.n2965 D.n2963 0.051
R11503 D.n2946 D.n2944 0.051
R11504 D.n2956 D.n2955 0.051
R11505 D.n2974 D.n2973 0.051
R11506 D.n2992 D.n2991 0.051
R11507 D.n3010 D.n3009 0.051
R11508 D.n3028 D.n3027 0.051
R11509 D.n3046 D.n3045 0.051
R11510 D.n3064 D.n3063 0.051
R11511 D.n3086 D.n3085 0.051
R11512 D.n2755 D.n2753 0.051
R11513 D.n2775 D.n2773 0.051
R11514 D.n2795 D.n2793 0.051
R11515 D.n2815 D.n2813 0.051
R11516 D.n2835 D.n2833 0.051
R11517 D.n2855 D.n2853 0.051
R11518 D.n2875 D.n2873 0.051
R11519 D.n2864 D.n2863 0.051
R11520 D.n2844 D.n2843 0.051
R11521 D.n2824 D.n2823 0.051
R11522 D.n2804 D.n2803 0.051
R11523 D.n2784 D.n2783 0.051
R11524 D.n2764 D.n2763 0.051
R11525 D.n2739 D.n2738 0.051
R11526 D.n2674 D.n2672 0.051
R11527 D.n2656 D.n2654 0.051
R11528 D.n2638 D.n2636 0.051
R11529 D.n2620 D.n2618 0.051
R11530 D.n2602 D.n2600 0.051
R11531 D.n2583 D.n2581 0.051
R11532 D.n2593 D.n2592 0.051
R11533 D.n2611 D.n2610 0.051
R11534 D.n2629 D.n2628 0.051
R11535 D.n2647 D.n2646 0.051
R11536 D.n2665 D.n2664 0.051
R11537 D.n2686 D.n2685 0.051
R11538 D.n2432 D.n2430 0.051
R11539 D.n2452 D.n2450 0.051
R11540 D.n2472 D.n2470 0.051
R11541 D.n2492 D.n2490 0.051
R11542 D.n2512 D.n2510 0.051
R11543 D.n2501 D.n2500 0.051
R11544 D.n2481 D.n2480 0.051
R11545 D.n2461 D.n2460 0.051
R11546 D.n2441 D.n2440 0.051
R11547 D.n2416 D.n2415 0.051
R11548 D.n2349 D.n2347 0.051
R11549 D.n2331 D.n2329 0.051
R11550 D.n2313 D.n2311 0.051
R11551 D.n2294 D.n2292 0.051
R11552 D.n2304 D.n2303 0.051
R11553 D.n2322 D.n2321 0.051
R11554 D.n2340 D.n2339 0.051
R11555 D.n2362 D.n2361 0.051
R11556 D.n2183 D.n2181 0.051
R11557 D.n2203 D.n2201 0.051
R11558 D.n2223 D.n2221 0.051
R11559 D.n2212 D.n2211 0.051
R11560 D.n2192 D.n2191 0.051
R11561 D.n2169 D.n2168 0.051
R11562 D.n2110 D.n2108 0.051
R11563 D.n2091 D.n2089 0.051
R11564 D.n2101 D.n2100 0.051
R11565 D.n2123 D.n2122 0.051
R11566 D.n52 D.n51 0.051
R11567 D.n61 D.n60 0.051
R11568 D.n70 D.n69 0.051
R11569 D.n79 D.n78 0.051
R11570 D.n88 D.n87 0.051
R11571 D.n97 D.n96 0.051
R11572 D.n106 D.n105 0.051
R11573 D.n115 D.n114 0.051
R11574 D.n124 D.n123 0.051
R11575 D.n133 D.n132 0.051
R11576 D.n142 D.n141 0.051
R11577 D.n151 D.n150 0.051
R11578 D.n160 D.n159 0.051
R11579 D.n169 D.n168 0.051
R11580 D.n178 D.n177 0.051
R11581 D.n187 D.n186 0.051
R11582 D.n196 D.n195 0.051
R11583 D.n205 D.n204 0.051
R11584 D.n214 D.n213 0.051
R11585 D.n284 D.n282 0.051
R11586 D.n300 D.n298 0.051
R11587 D.n552 D.n550 0.051
R11588 D.n538 D.n536 0.051
R11589 D.n524 D.n522 0.051
R11590 D.n510 D.n508 0.051
R11591 D.n496 D.n494 0.051
R11592 D.n482 D.n480 0.051
R11593 D.n468 D.n466 0.051
R11594 D.n454 D.n452 0.051
R11595 D.n440 D.n438 0.051
R11596 D.n426 D.n424 0.051
R11597 D.n412 D.n410 0.051
R11598 D.n398 D.n396 0.051
R11599 D.n384 D.n382 0.051
R11600 D.n370 D.n368 0.051
R11601 D.n356 D.n354 0.051
R11602 D.n342 D.n340 0.051
R11603 D.n328 D.n326 0.051
R11604 D.n314 D.n312 0.051
R11605 D.n575 D.n573 0.051
R11606 D.n591 D.n589 0.051
R11607 D.n815 D.n813 0.051
R11608 D.n801 D.n799 0.051
R11609 D.n787 D.n785 0.051
R11610 D.n773 D.n771 0.051
R11611 D.n759 D.n757 0.051
R11612 D.n745 D.n743 0.051
R11613 D.n731 D.n729 0.051
R11614 D.n717 D.n715 0.051
R11615 D.n703 D.n701 0.051
R11616 D.n689 D.n687 0.051
R11617 D.n675 D.n673 0.051
R11618 D.n661 D.n659 0.051
R11619 D.n647 D.n645 0.051
R11620 D.n633 D.n631 0.051
R11621 D.n619 D.n617 0.051
R11622 D.n605 D.n603 0.051
R11623 D.n838 D.n836 0.051
R11624 D.n854 D.n852 0.051
R11625 D.n1050 D.n1048 0.051
R11626 D.n1036 D.n1034 0.051
R11627 D.n1022 D.n1020 0.051
R11628 D.n1008 D.n1006 0.051
R11629 D.n994 D.n992 0.051
R11630 D.n980 D.n978 0.051
R11631 D.n966 D.n964 0.051
R11632 D.n952 D.n950 0.051
R11633 D.n938 D.n936 0.051
R11634 D.n924 D.n922 0.051
R11635 D.n910 D.n908 0.051
R11636 D.n896 D.n894 0.051
R11637 D.n882 D.n880 0.051
R11638 D.n868 D.n866 0.051
R11639 D.n1073 D.n1071 0.051
R11640 D.n1089 D.n1087 0.051
R11641 D.n1257 D.n1255 0.051
R11642 D.n1243 D.n1241 0.051
R11643 D.n1229 D.n1227 0.051
R11644 D.n1215 D.n1213 0.051
R11645 D.n1201 D.n1199 0.051
R11646 D.n1187 D.n1185 0.051
R11647 D.n1173 D.n1171 0.051
R11648 D.n1159 D.n1157 0.051
R11649 D.n1145 D.n1143 0.051
R11650 D.n1131 D.n1129 0.051
R11651 D.n1117 D.n1115 0.051
R11652 D.n1103 D.n1101 0.051
R11653 D.n1280 D.n1278 0.051
R11654 D.n1296 D.n1294 0.051
R11655 D.n1436 D.n1434 0.051
R11656 D.n1422 D.n1420 0.051
R11657 D.n1408 D.n1406 0.051
R11658 D.n1394 D.n1392 0.051
R11659 D.n1380 D.n1378 0.051
R11660 D.n1366 D.n1364 0.051
R11661 D.n1352 D.n1350 0.051
R11662 D.n1338 D.n1336 0.051
R11663 D.n1324 D.n1322 0.051
R11664 D.n1310 D.n1308 0.051
R11665 D.n1460 D.n1458 0.051
R11666 D.n1476 D.n1474 0.051
R11667 D.n1588 D.n1586 0.051
R11668 D.n1574 D.n1572 0.051
R11669 D.n1560 D.n1558 0.051
R11670 D.n1546 D.n1544 0.051
R11671 D.n1532 D.n1530 0.051
R11672 D.n1518 D.n1516 0.051
R11673 D.n1504 D.n1502 0.051
R11674 D.n1490 D.n1488 0.051
R11675 D.n1612 D.n1610 0.051
R11676 D.n1628 D.n1626 0.051
R11677 D.n1712 D.n1710 0.051
R11678 D.n1698 D.n1696 0.051
R11679 D.n1684 D.n1682 0.051
R11680 D.n1670 D.n1668 0.051
R11681 D.n1656 D.n1654 0.051
R11682 D.n1642 D.n1640 0.051
R11683 D.n1736 D.n1734 0.051
R11684 D.n1752 D.n1750 0.051
R11685 D.n1808 D.n1806 0.051
R11686 D.n1794 D.n1792 0.051
R11687 D.n1780 D.n1778 0.051
R11688 D.n1766 D.n1764 0.051
R11689 D.n1831 D.n1829 0.051
R11690 D.n1847 D.n1845 0.051
R11691 D.n1875 D.n1873 0.051
R11692 D.n1861 D.n1859 0.051
R11693 D.n1950 D.n1949 0.051
R11694 D.n1928 D.n1924 0.05
R11695 D.n1921 D.n1891 0.05
R11696 D.n1993 D.n1989 0.05
R11697 D.n3590 D.n3583 0.05
R11698 D.n3137 D.n3134 0.05
R11699 D.n3107 D.n3100 0.05
R11700 D.n2730 D.n2726 0.05
R11701 D.n2702 D.n2697 0.05
R11702 D.n2407 D.n2403 0.05
R11703 D.n2383 D.n2376 0.05
R11704 D.n2162 D.n2159 0.05
R11705 D.n2144 D.n2137 0.05
R11706 D.n1977 D.n1971 0.05
R11707 D.n565 D.n275 0.05
R11708 D.n828 D.n569 0.05
R11709 D.n1063 D.n832 0.05
R11710 D.n1270 D.n1067 0.05
R11711 D.n1449 D.n1274 0.05
R11712 D.n1601 D.n1454 0.05
R11713 D.n1725 D.n1606 0.05
R11714 D.n1821 D.n1730 0.05
R11715 D.n1888 D.n1825 0.05
R11716 D.n562 D.n548 0.049
R11717 D.n548 D.n534 0.049
R11718 D.n534 D.n520 0.049
R11719 D.n520 D.n506 0.049
R11720 D.n506 D.n492 0.049
R11721 D.n492 D.n478 0.049
R11722 D.n478 D.n464 0.049
R11723 D.n464 D.n450 0.049
R11724 D.n450 D.n436 0.049
R11725 D.n436 D.n422 0.049
R11726 D.n422 D.n408 0.049
R11727 D.n408 D.n394 0.049
R11728 D.n394 D.n380 0.049
R11729 D.n380 D.n366 0.049
R11730 D.n366 D.n352 0.049
R11731 D.n352 D.n338 0.049
R11732 D.n338 D.n324 0.049
R11733 D.n324 D.n310 0.049
R11734 D.n310 D.n296 0.049
R11735 D.n825 D.n811 0.049
R11736 D.n811 D.n797 0.049
R11737 D.n797 D.n783 0.049
R11738 D.n783 D.n769 0.049
R11739 D.n769 D.n755 0.049
R11740 D.n755 D.n741 0.049
R11741 D.n741 D.n727 0.049
R11742 D.n727 D.n713 0.049
R11743 D.n713 D.n699 0.049
R11744 D.n699 D.n685 0.049
R11745 D.n685 D.n671 0.049
R11746 D.n671 D.n657 0.049
R11747 D.n657 D.n643 0.049
R11748 D.n643 D.n629 0.049
R11749 D.n629 D.n615 0.049
R11750 D.n615 D.n601 0.049
R11751 D.n601 D.n587 0.049
R11752 D.n1060 D.n1046 0.049
R11753 D.n1046 D.n1032 0.049
R11754 D.n1032 D.n1018 0.049
R11755 D.n1018 D.n1004 0.049
R11756 D.n1004 D.n990 0.049
R11757 D.n990 D.n976 0.049
R11758 D.n976 D.n962 0.049
R11759 D.n962 D.n948 0.049
R11760 D.n948 D.n934 0.049
R11761 D.n934 D.n920 0.049
R11762 D.n920 D.n906 0.049
R11763 D.n906 D.n892 0.049
R11764 D.n892 D.n878 0.049
R11765 D.n878 D.n864 0.049
R11766 D.n864 D.n850 0.049
R11767 D.n1267 D.n1253 0.049
R11768 D.n1253 D.n1239 0.049
R11769 D.n1239 D.n1225 0.049
R11770 D.n1225 D.n1211 0.049
R11771 D.n1211 D.n1197 0.049
R11772 D.n1197 D.n1183 0.049
R11773 D.n1183 D.n1169 0.049
R11774 D.n1169 D.n1155 0.049
R11775 D.n1155 D.n1141 0.049
R11776 D.n1141 D.n1127 0.049
R11777 D.n1127 D.n1113 0.049
R11778 D.n1113 D.n1099 0.049
R11779 D.n1099 D.n1085 0.049
R11780 D.n1446 D.n1432 0.049
R11781 D.n1432 D.n1418 0.049
R11782 D.n1418 D.n1404 0.049
R11783 D.n1404 D.n1390 0.049
R11784 D.n1390 D.n1376 0.049
R11785 D.n1376 D.n1362 0.049
R11786 D.n1362 D.n1348 0.049
R11787 D.n1348 D.n1334 0.049
R11788 D.n1334 D.n1320 0.049
R11789 D.n1320 D.n1306 0.049
R11790 D.n1306 D.n1292 0.049
R11791 D.n1598 D.n1584 0.049
R11792 D.n1584 D.n1570 0.049
R11793 D.n1570 D.n1556 0.049
R11794 D.n1556 D.n1542 0.049
R11795 D.n1542 D.n1528 0.049
R11796 D.n1528 D.n1514 0.049
R11797 D.n1514 D.n1500 0.049
R11798 D.n1500 D.n1486 0.049
R11799 D.n1486 D.n1472 0.049
R11800 D.n1722 D.n1708 0.049
R11801 D.n1708 D.n1694 0.049
R11802 D.n1694 D.n1680 0.049
R11803 D.n1680 D.n1666 0.049
R11804 D.n1666 D.n1652 0.049
R11805 D.n1652 D.n1638 0.049
R11806 D.n1638 D.n1624 0.049
R11807 D.n1818 D.n1804 0.049
R11808 D.n1804 D.n1790 0.049
R11809 D.n1790 D.n1776 0.049
R11810 D.n1776 D.n1762 0.049
R11811 D.n1762 D.n1748 0.049
R11812 D.n1887 D.n1871 0.049
R11813 D.n1871 D.n1857 0.049
R11814 D.n1857 D.n1843 0.049
R11815 D.n12 D.n11 0.049
R11816 D.n241 D.n240 0.049
R11817 D.n242 D.n241 0.049
R11818 D.n243 D.n242 0.049
R11819 D.n244 D.n243 0.049
R11820 D.n245 D.n244 0.049
R11821 D.n246 D.n245 0.049
R11822 D.n247 D.n246 0.049
R11823 D.n248 D.n247 0.049
R11824 D.n249 D.n248 0.049
R11825 D.n250 D.n249 0.049
R11826 D.n251 D.n250 0.049
R11827 D.n252 D.n251 0.049
R11828 D.n253 D.n252 0.049
R11829 D.n254 D.n253 0.049
R11830 D.n255 D.n254 0.049
R11831 D.n256 D.n255 0.049
R11832 D.n257 D.n256 0.049
R11833 D.n258 D.n257 0.049
R11834 D.n259 D.n258 0.049
R11835 D.n260 D.n259 0.049
R11836 D.n261 D.n260 0.049
R11837 D.n3592 D.n3591 0.049
R11838 D.n3593 D.n3592 0.049
R11839 D.n3594 D.n3593 0.049
R11840 D.n3595 D.n3594 0.049
R11841 D.n3596 D.n3595 0.049
R11842 D.n3597 D.n3596 0.049
R11843 D.n3598 D.n3597 0.049
R11844 D.n3599 D.n3598 0.049
R11845 D.n3600 D.n3599 0.049
R11846 D.n3601 D.n3600 0.049
R11847 D.n3602 D.n3601 0.049
R11848 D.n3603 D.n3602 0.049
R11849 D.n3604 D.n3603 0.049
R11850 D.n3605 D.n3604 0.049
R11851 D.n3606 D.n3605 0.049
R11852 D.n3607 D.n3606 0.049
R11853 D.n3608 D.n3607 0.049
R11854 D.n3609 D.n3608 0.049
R11855 D.n3610 D.n3609 0.049
R11856 D.n3109 D.n3108 0.049
R11857 D.n3110 D.n3109 0.049
R11858 D.n3111 D.n3110 0.049
R11859 D.n3112 D.n3111 0.049
R11860 D.n3113 D.n3112 0.049
R11861 D.n3114 D.n3113 0.049
R11862 D.n3115 D.n3114 0.049
R11863 D.n3116 D.n3115 0.049
R11864 D.n3117 D.n3116 0.049
R11865 D.n3118 D.n3117 0.049
R11866 D.n3119 D.n3118 0.049
R11867 D.n3120 D.n3119 0.049
R11868 D.n3121 D.n3120 0.049
R11869 D.n3122 D.n3121 0.049
R11870 D.n3123 D.n3122 0.049
R11871 D.n2704 D.n2703 0.049
R11872 D.n2705 D.n2704 0.049
R11873 D.n2706 D.n2705 0.049
R11874 D.n2707 D.n2706 0.049
R11875 D.n2708 D.n2707 0.049
R11876 D.n2709 D.n2708 0.049
R11877 D.n2710 D.n2709 0.049
R11878 D.n2711 D.n2710 0.049
R11879 D.n2712 D.n2711 0.049
R11880 D.n2713 D.n2712 0.049
R11881 D.n2714 D.n2713 0.049
R11882 D.n2385 D.n2384 0.049
R11883 D.n2386 D.n2385 0.049
R11884 D.n2387 D.n2386 0.049
R11885 D.n2388 D.n2387 0.049
R11886 D.n2389 D.n2388 0.049
R11887 D.n2390 D.n2389 0.049
R11888 D.n2391 D.n2390 0.049
R11889 D.n2146 D.n2145 0.049
R11890 D.n2147 D.n2146 0.049
R11891 D.n2148 D.n2147 0.049
R11892 D.n3611 D.n3610 0.049
R11893 D.n3124 D.n3123 0.049
R11894 D.n2715 D.n2714 0.049
R11895 D.n2392 D.n2391 0.049
R11896 D.n2149 D.n2148 0.049
R11897 D.n565 D.n562 0.047
R11898 D.n828 D.n825 0.047
R11899 D.n1063 D.n1060 0.047
R11900 D.n1270 D.n1267 0.047
R11901 D.n1449 D.n1446 0.047
R11902 D.n1601 D.n1598 0.047
R11903 D.n1725 D.n1722 0.047
R11904 D.n1821 D.n1818 0.047
R11905 D.n1888 D.n1887 0.047
R11906 D.n1957 D.n1956 0.045
R11907 D.n2040 D.n2039 0.045
R11908 D.n3357 D.n3356 0.045
R11909 D.n3373 D.n3372 0.045
R11910 D.n3326 D.n3325 0.045
R11911 D.n3338 D.n3337 0.045
R11912 D.n2914 D.n2913 0.045
R11913 D.n2930 D.n2929 0.045
R11914 D.n2883 D.n2882 0.045
R11915 D.n2895 D.n2894 0.045
R11916 D.n2551 D.n2550 0.045
R11917 D.n2567 D.n2566 0.045
R11918 D.n2520 D.n2519 0.045
R11919 D.n2532 D.n2531 0.045
R11920 D.n2262 D.n2261 0.045
R11921 D.n2278 D.n2277 0.045
R11922 D.n2231 D.n2230 0.045
R11923 D.n2243 D.n2242 0.045
R11924 D.n2059 D.n2058 0.045
R11925 D.n2075 D.n2074 0.045
R11926 D.n2026 D.n2025 0.045
R11927 D.n1950 D.n1947 0.044
R11928 D.n262 D.n261 0.044
R11929 D.n2010 D.n2009 0.043
R11930 D.n3150 D.n3149 0.043
R11931 D.n3095 D.n3094 0.043
R11932 D.n2747 D.n2746 0.043
R11933 D.n2424 D.n2423 0.043
R11934 D.n2371 D.n2370 0.043
R11935 D.n2175 D.n2174 0.043
R11936 D.n2132 D.n2131 0.043
R11937 D.n3565 D.n3564 0.043
R11938 D.n3140 D.n3139 0.043
R11939 D.n3082 D.n3081 0.043
R11940 D.n2735 D.n2734 0.043
R11941 D.n2682 D.n2681 0.043
R11942 D.n2412 D.n2411 0.043
R11943 D.n2358 D.n2357 0.043
R11944 D.n2165 D.n2164 0.043
R11945 D.n2119 D.n2118 0.043
R11946 D.n1998 D.n1997 0.043
R11947 D.n309 D.n308 0.042
R11948 D.n323 D.n322 0.042
R11949 D.n337 D.n336 0.042
R11950 D.n351 D.n350 0.042
R11951 D.n365 D.n364 0.042
R11952 D.n379 D.n378 0.042
R11953 D.n393 D.n392 0.042
R11954 D.n407 D.n406 0.042
R11955 D.n421 D.n420 0.042
R11956 D.n435 D.n434 0.042
R11957 D.n449 D.n448 0.042
R11958 D.n463 D.n462 0.042
R11959 D.n477 D.n476 0.042
R11960 D.n491 D.n490 0.042
R11961 D.n505 D.n504 0.042
R11962 D.n519 D.n518 0.042
R11963 D.n533 D.n532 0.042
R11964 D.n547 D.n546 0.042
R11965 D.n561 D.n560 0.042
R11966 D.n600 D.n599 0.042
R11967 D.n614 D.n613 0.042
R11968 D.n628 D.n627 0.042
R11969 D.n642 D.n641 0.042
R11970 D.n656 D.n655 0.042
R11971 D.n670 D.n669 0.042
R11972 D.n684 D.n683 0.042
R11973 D.n698 D.n697 0.042
R11974 D.n712 D.n711 0.042
R11975 D.n726 D.n725 0.042
R11976 D.n740 D.n739 0.042
R11977 D.n754 D.n753 0.042
R11978 D.n768 D.n767 0.042
R11979 D.n782 D.n781 0.042
R11980 D.n796 D.n795 0.042
R11981 D.n810 D.n809 0.042
R11982 D.n824 D.n823 0.042
R11983 D.n863 D.n862 0.042
R11984 D.n877 D.n876 0.042
R11985 D.n891 D.n890 0.042
R11986 D.n905 D.n904 0.042
R11987 D.n919 D.n918 0.042
R11988 D.n933 D.n932 0.042
R11989 D.n947 D.n946 0.042
R11990 D.n961 D.n960 0.042
R11991 D.n975 D.n974 0.042
R11992 D.n989 D.n988 0.042
R11993 D.n1003 D.n1002 0.042
R11994 D.n1017 D.n1016 0.042
R11995 D.n1031 D.n1030 0.042
R11996 D.n1045 D.n1044 0.042
R11997 D.n1059 D.n1058 0.042
R11998 D.n1098 D.n1097 0.042
R11999 D.n1112 D.n1111 0.042
R12000 D.n1126 D.n1125 0.042
R12001 D.n1140 D.n1139 0.042
R12002 D.n1154 D.n1153 0.042
R12003 D.n1168 D.n1167 0.042
R12004 D.n1182 D.n1181 0.042
R12005 D.n1196 D.n1195 0.042
R12006 D.n1210 D.n1209 0.042
R12007 D.n1224 D.n1223 0.042
R12008 D.n1238 D.n1237 0.042
R12009 D.n1252 D.n1251 0.042
R12010 D.n1266 D.n1265 0.042
R12011 D.n1305 D.n1304 0.042
R12012 D.n1319 D.n1318 0.042
R12013 D.n1333 D.n1332 0.042
R12014 D.n1347 D.n1346 0.042
R12015 D.n1361 D.n1360 0.042
R12016 D.n1375 D.n1374 0.042
R12017 D.n1389 D.n1388 0.042
R12018 D.n1403 D.n1402 0.042
R12019 D.n1417 D.n1416 0.042
R12020 D.n1431 D.n1430 0.042
R12021 D.n1445 D.n1444 0.042
R12022 D.n1485 D.n1484 0.042
R12023 D.n1499 D.n1498 0.042
R12024 D.n1513 D.n1512 0.042
R12025 D.n1527 D.n1526 0.042
R12026 D.n1541 D.n1540 0.042
R12027 D.n1555 D.n1554 0.042
R12028 D.n1569 D.n1568 0.042
R12029 D.n1583 D.n1582 0.042
R12030 D.n1597 D.n1596 0.042
R12031 D.n1637 D.n1636 0.042
R12032 D.n1651 D.n1650 0.042
R12033 D.n1665 D.n1664 0.042
R12034 D.n1679 D.n1678 0.042
R12035 D.n1693 D.n1692 0.042
R12036 D.n1707 D.n1706 0.042
R12037 D.n1721 D.n1720 0.042
R12038 D.n1761 D.n1760 0.042
R12039 D.n1775 D.n1774 0.042
R12040 D.n1789 D.n1788 0.042
R12041 D.n1803 D.n1802 0.042
R12042 D.n1817 D.n1816 0.042
R12043 D.n1856 D.n1855 0.042
R12044 D.n1870 D.n1869 0.042
R12045 D.n1886 D.n1885 0.042
R12046 D.n3362 D.n3361 0.041
R12047 D.n2919 D.n2918 0.041
R12048 D.n2556 D.n2555 0.041
R12049 D.n2267 D.n2266 0.041
R12050 D.n2064 D.n2063 0.041
R12051 D.n3382 D.n3381 0.041
R12052 D.n2935 D.n2934 0.041
R12053 D.n2572 D.n2571 0.041
R12054 D.n2283 D.n2282 0.041
R12055 D.n2080 D.n2079 0.041
R12056 D.n2046 D.n2045 0.039
R12057 D.n2048 D.n2046 0.039
R12058 D.n2007 D.n2006 0.039
R12059 D.n3367 D.n3366 0.039
R12060 D.n3387 D.n3386 0.039
R12061 D.n3389 D.n3387 0.039
R12062 D.n3577 D.n3576 0.039
R12063 D.n3332 D.n3331 0.039
R12064 D.n3344 D.n3343 0.039
R12065 D.n3346 D.n3344 0.039
R12066 D.n2924 D.n2923 0.039
R12067 D.n2940 D.n2939 0.039
R12068 D.n2942 D.n2940 0.039
R12069 D.n3093 D.n3092 0.039
R12070 D.n2889 D.n2888 0.039
R12071 D.n2901 D.n2900 0.039
R12072 D.n2903 D.n2901 0.039
R12073 D.n2744 D.n2743 0.039
R12074 D.n2722 D.n2721 0.039
R12075 D.n2561 D.n2560 0.039
R12076 D.n2577 D.n2576 0.039
R12077 D.n2579 D.n2577 0.039
R12078 D.n2526 D.n2525 0.039
R12079 D.n2538 D.n2537 0.039
R12080 D.n2540 D.n2538 0.039
R12081 D.n2421 D.n2420 0.039
R12082 D.n2399 D.n2398 0.039
R12083 D.n2272 D.n2271 0.039
R12084 D.n2288 D.n2287 0.039
R12085 D.n2290 D.n2288 0.039
R12086 D.n2369 D.n2368 0.039
R12087 D.n2237 D.n2236 0.039
R12088 D.n2249 D.n2248 0.039
R12089 D.n2251 D.n2249 0.039
R12090 D.n2069 D.n2068 0.039
R12091 D.n2085 D.n2084 0.039
R12092 D.n2087 D.n2085 0.039
R12093 D.n2130 D.n2129 0.039
R12094 D.n1985 D.n1984 0.039
R12095 D.n2032 D.n2031 0.039
R12096 D.n1949 D.n1948 0.039
R12097 D.n1956 D.n1955 0.039
R12098 D.n1976 D.n1975 0.039
R12099 D.n47 D.n26 0.039
R12100 D D.n3614 0.038
R12101 D D.n1944 0.037
R12102 D.n1962 D.n1951 0.035
R12103 D.n1981 D.n1980 0.034
R12104 D.n293 D.n292 0.034
R12105 D.n584 D.n583 0.034
R12106 D.n847 D.n846 0.034
R12107 D.n1082 D.n1081 0.034
R12108 D.n1289 D.n1288 0.034
R12109 D.n1469 D.n1468 0.034
R12110 D.n1621 D.n1620 0.034
R12111 D.n1745 D.n1744 0.034
R12112 D.n1840 D.n1839 0.034
R12113 D.n1932 D.n1931 0.034
R12114 D.n3379 D.n3378 0.034
R12115 D.n1962 D.n1954 0.033
R12116 D.n2048 D.n2038 0.033
R12117 D.n3389 D.n3371 0.033
R12118 D.n3346 D.n3336 0.033
R12119 D.n2942 D.n2928 0.033
R12120 D.n2903 D.n2893 0.033
R12121 D.n2579 D.n2565 0.033
R12122 D.n2540 D.n2530 0.033
R12123 D.n2290 D.n2276 0.033
R12124 D.n2251 D.n2241 0.033
R12125 D.n2087 D.n2073 0.033
R12126 D.n1895 D.n1894 0.033
R12127 D.n3614 D.n3612 0.032
R12128 D.n271 D.n270 0.031
R12129 D.n1935 D.n1934 0.031
R12130 D.n1936 D.n1935 0.031
R12131 D.n1937 D.n1936 0.031
R12132 D.n1938 D.n1937 0.031
R12133 D.n1939 D.n1938 0.031
R12134 D.n1940 D.n1939 0.031
R12135 D.n1941 D.n1940 0.031
R12136 D.n1942 D.n1941 0.031
R12137 D.n1943 D.n1942 0.031
R12138 D.n1944 D.n1943 0.031
R12139 D.n1993 D.n1988 0.03
R12140 D.n3590 D.n3582 0.03
R12141 D.n3590 D.n3587 0.03
R12142 D.n3107 D.n3099 0.03
R12143 D.n3107 D.n3104 0.03
R12144 D.n2730 D.n2728 0.03
R12145 D.n2730 D.n2723 0.03
R12146 D.n2407 D.n2405 0.03
R12147 D.n2407 D.n2400 0.03
R12148 D.n2383 D.n2375 0.03
R12149 D.n2383 D.n2380 0.03
R12150 D.n2144 D.n2136 0.03
R12151 D.n2144 D.n2141 0.03
R12152 D.n1993 D.n1992 0.03
R12153 D.n1977 D.n1968 0.03
R12154 D.n1977 D.n1973 0.03
R12155 D.n3126 D.n3125 0.029
R12156 D.n2717 D.n2716 0.029
R12157 D.n2394 D.n2393 0.029
R12158 D.n2151 D.n2150 0.029
R12159 D.n3612 D.n3354 0.029
R12160 D.n3125 D.n2911 0.029
R12161 D.n2716 D.n2548 0.029
R12162 D.n2393 D.n2259 0.029
R12163 D.n2150 D.n2056 0.029
R12164 D.n25 D.n15 0.029
R12165 D.n23 D.n22 0.028
R12166 D.n41 D.n40 0.028
R12167 D.n23 D.n17 0.027
R12168 D.n3389 D.n3368 0.027
R12169 D.n3346 D.n3333 0.027
R12170 D.n2942 D.n2925 0.027
R12171 D.n2903 D.n2890 0.027
R12172 D.n2579 D.n2562 0.027
R12173 D.n2540 D.n2527 0.027
R12174 D.n2290 D.n2273 0.027
R12175 D.n2251 D.n2238 0.027
R12176 D.n2087 D.n2070 0.027
R12177 D.n2048 D.n2033 0.027
R12178 D.n1962 D.n1960 0.027
R12179 D.n47 D.n27 0.027
R12180 D.n3 D.n0 0.026
R12181 D.n41 D.n35 0.026
R12182 D.n561 D.n557 0.025
R12183 D.n547 D.n543 0.025
R12184 D.n533 D.n529 0.025
R12185 D.n519 D.n515 0.025
R12186 D.n505 D.n501 0.025
R12187 D.n491 D.n487 0.025
R12188 D.n477 D.n473 0.025
R12189 D.n463 D.n459 0.025
R12190 D.n449 D.n445 0.025
R12191 D.n435 D.n431 0.025
R12192 D.n421 D.n417 0.025
R12193 D.n407 D.n403 0.025
R12194 D.n393 D.n389 0.025
R12195 D.n379 D.n375 0.025
R12196 D.n365 D.n361 0.025
R12197 D.n351 D.n347 0.025
R12198 D.n337 D.n333 0.025
R12199 D.n323 D.n319 0.025
R12200 D.n309 D.n305 0.025
R12201 D.n295 D.n289 0.025
R12202 D.n824 D.n820 0.025
R12203 D.n810 D.n806 0.025
R12204 D.n796 D.n792 0.025
R12205 D.n782 D.n778 0.025
R12206 D.n768 D.n764 0.025
R12207 D.n754 D.n750 0.025
R12208 D.n740 D.n736 0.025
R12209 D.n726 D.n722 0.025
R12210 D.n712 D.n708 0.025
R12211 D.n698 D.n694 0.025
R12212 D.n684 D.n680 0.025
R12213 D.n670 D.n666 0.025
R12214 D.n656 D.n652 0.025
R12215 D.n642 D.n638 0.025
R12216 D.n628 D.n624 0.025
R12217 D.n614 D.n610 0.025
R12218 D.n600 D.n596 0.025
R12219 D.n586 D.n580 0.025
R12220 D.n1059 D.n1055 0.025
R12221 D.n1045 D.n1041 0.025
R12222 D.n1031 D.n1027 0.025
R12223 D.n1017 D.n1013 0.025
R12224 D.n1003 D.n999 0.025
R12225 D.n989 D.n985 0.025
R12226 D.n975 D.n971 0.025
R12227 D.n961 D.n957 0.025
R12228 D.n947 D.n943 0.025
R12229 D.n933 D.n929 0.025
R12230 D.n919 D.n915 0.025
R12231 D.n905 D.n901 0.025
R12232 D.n891 D.n887 0.025
R12233 D.n877 D.n873 0.025
R12234 D.n863 D.n859 0.025
R12235 D.n849 D.n843 0.025
R12236 D.n1266 D.n1262 0.025
R12237 D.n1252 D.n1248 0.025
R12238 D.n1238 D.n1234 0.025
R12239 D.n1224 D.n1220 0.025
R12240 D.n1210 D.n1206 0.025
R12241 D.n1196 D.n1192 0.025
R12242 D.n1182 D.n1178 0.025
R12243 D.n1168 D.n1164 0.025
R12244 D.n1154 D.n1150 0.025
R12245 D.n1140 D.n1136 0.025
R12246 D.n1126 D.n1122 0.025
R12247 D.n1112 D.n1108 0.025
R12248 D.n1098 D.n1094 0.025
R12249 D.n1084 D.n1078 0.025
R12250 D.n1445 D.n1441 0.025
R12251 D.n1431 D.n1427 0.025
R12252 D.n1417 D.n1413 0.025
R12253 D.n1403 D.n1399 0.025
R12254 D.n1389 D.n1385 0.025
R12255 D.n1375 D.n1371 0.025
R12256 D.n1361 D.n1357 0.025
R12257 D.n1347 D.n1343 0.025
R12258 D.n1333 D.n1329 0.025
R12259 D.n1319 D.n1315 0.025
R12260 D.n1305 D.n1301 0.025
R12261 D.n1291 D.n1285 0.025
R12262 D.n1597 D.n1593 0.025
R12263 D.n1583 D.n1579 0.025
R12264 D.n1569 D.n1565 0.025
R12265 D.n1555 D.n1551 0.025
R12266 D.n1541 D.n1537 0.025
R12267 D.n1527 D.n1523 0.025
R12268 D.n1513 D.n1509 0.025
R12269 D.n1499 D.n1495 0.025
R12270 D.n1485 D.n1481 0.025
R12271 D.n1471 D.n1465 0.025
R12272 D.n1721 D.n1717 0.025
R12273 D.n1707 D.n1703 0.025
R12274 D.n1693 D.n1689 0.025
R12275 D.n1679 D.n1675 0.025
R12276 D.n1665 D.n1661 0.025
R12277 D.n1651 D.n1647 0.025
R12278 D.n1637 D.n1633 0.025
R12279 D.n1623 D.n1617 0.025
R12280 D.n1817 D.n1813 0.025
R12281 D.n1803 D.n1799 0.025
R12282 D.n1789 D.n1785 0.025
R12283 D.n1775 D.n1771 0.025
R12284 D.n1761 D.n1757 0.025
R12285 D.n1747 D.n1741 0.025
R12286 D.n1886 D.n1882 0.025
R12287 D.n1870 D.n1866 0.025
R12288 D.n1856 D.n1852 0.025
R12289 D.n1842 D.n1836 0.025
R12290 D.n265 D.n264 0.024
R12291 D.n26 D.n25 0.023
R12292 D.n2043 D.n2040 0.023
R12293 D.n2045 D.n2044 0.023
R12294 D.n3364 D.n3357 0.023
R12295 D.n3366 D.n3365 0.023
R12296 D.n3384 D.n3373 0.023
R12297 D.n3386 D.n3385 0.023
R12298 D.n3329 D.n3326 0.023
R12299 D.n3331 D.n3330 0.023
R12300 D.n3341 D.n3338 0.023
R12301 D.n3343 D.n3342 0.023
R12302 D.n2921 D.n2914 0.023
R12303 D.n2923 D.n2922 0.023
R12304 D.n2937 D.n2930 0.023
R12305 D.n2939 D.n2938 0.023
R12306 D.n2886 D.n2883 0.023
R12307 D.n2888 D.n2887 0.023
R12308 D.n2898 D.n2895 0.023
R12309 D.n2900 D.n2899 0.023
R12310 D.n2558 D.n2551 0.023
R12311 D.n2560 D.n2559 0.023
R12312 D.n2574 D.n2567 0.023
R12313 D.n2576 D.n2575 0.023
R12314 D.n2523 D.n2520 0.023
R12315 D.n2525 D.n2524 0.023
R12316 D.n2535 D.n2532 0.023
R12317 D.n2537 D.n2536 0.023
R12318 D.n2269 D.n2262 0.023
R12319 D.n2271 D.n2270 0.023
R12320 D.n2285 D.n2278 0.023
R12321 D.n2287 D.n2286 0.023
R12322 D.n2234 D.n2231 0.023
R12323 D.n2236 D.n2235 0.023
R12324 D.n2246 D.n2243 0.023
R12325 D.n2248 D.n2247 0.023
R12326 D.n2066 D.n2059 0.023
R12327 D.n2068 D.n2067 0.023
R12328 D.n2082 D.n2075 0.023
R12329 D.n2084 D.n2083 0.023
R12330 D.n2031 D.n2030 0.023
R12331 D.n2029 D.n2026 0.023
R12332 D.n44 D.n43 0.023
R12333 D.n565 D.n564 0.023
R12334 D.n309 D.n307 0.023
R12335 D.n323 D.n321 0.023
R12336 D.n337 D.n335 0.023
R12337 D.n351 D.n349 0.023
R12338 D.n365 D.n363 0.023
R12339 D.n379 D.n377 0.023
R12340 D.n393 D.n391 0.023
R12341 D.n407 D.n405 0.023
R12342 D.n421 D.n419 0.023
R12343 D.n435 D.n433 0.023
R12344 D.n449 D.n447 0.023
R12345 D.n463 D.n461 0.023
R12346 D.n477 D.n475 0.023
R12347 D.n491 D.n489 0.023
R12348 D.n505 D.n503 0.023
R12349 D.n519 D.n517 0.023
R12350 D.n533 D.n531 0.023
R12351 D.n547 D.n545 0.023
R12352 D.n561 D.n559 0.023
R12353 D.n828 D.n827 0.023
R12354 D.n600 D.n598 0.023
R12355 D.n614 D.n612 0.023
R12356 D.n628 D.n626 0.023
R12357 D.n642 D.n640 0.023
R12358 D.n656 D.n654 0.023
R12359 D.n670 D.n668 0.023
R12360 D.n684 D.n682 0.023
R12361 D.n698 D.n696 0.023
R12362 D.n712 D.n710 0.023
R12363 D.n726 D.n724 0.023
R12364 D.n740 D.n738 0.023
R12365 D.n754 D.n752 0.023
R12366 D.n768 D.n766 0.023
R12367 D.n782 D.n780 0.023
R12368 D.n796 D.n794 0.023
R12369 D.n810 D.n808 0.023
R12370 D.n824 D.n822 0.023
R12371 D.n1063 D.n1062 0.023
R12372 D.n863 D.n861 0.023
R12373 D.n877 D.n875 0.023
R12374 D.n891 D.n889 0.023
R12375 D.n905 D.n903 0.023
R12376 D.n919 D.n917 0.023
R12377 D.n933 D.n931 0.023
R12378 D.n947 D.n945 0.023
R12379 D.n961 D.n959 0.023
R12380 D.n975 D.n973 0.023
R12381 D.n989 D.n987 0.023
R12382 D.n1003 D.n1001 0.023
R12383 D.n1017 D.n1015 0.023
R12384 D.n1031 D.n1029 0.023
R12385 D.n1045 D.n1043 0.023
R12386 D.n1059 D.n1057 0.023
R12387 D.n1270 D.n1269 0.023
R12388 D.n1098 D.n1096 0.023
R12389 D.n1112 D.n1110 0.023
R12390 D.n1126 D.n1124 0.023
R12391 D.n1140 D.n1138 0.023
R12392 D.n1154 D.n1152 0.023
R12393 D.n1168 D.n1166 0.023
R12394 D.n1182 D.n1180 0.023
R12395 D.n1196 D.n1194 0.023
R12396 D.n1210 D.n1208 0.023
R12397 D.n1224 D.n1222 0.023
R12398 D.n1238 D.n1236 0.023
R12399 D.n1252 D.n1250 0.023
R12400 D.n1266 D.n1264 0.023
R12401 D.n1449 D.n1448 0.023
R12402 D.n1305 D.n1303 0.023
R12403 D.n1319 D.n1317 0.023
R12404 D.n1333 D.n1331 0.023
R12405 D.n1347 D.n1345 0.023
R12406 D.n1361 D.n1359 0.023
R12407 D.n1375 D.n1373 0.023
R12408 D.n1389 D.n1387 0.023
R12409 D.n1403 D.n1401 0.023
R12410 D.n1417 D.n1415 0.023
R12411 D.n1431 D.n1429 0.023
R12412 D.n1445 D.n1443 0.023
R12413 D.n1601 D.n1600 0.023
R12414 D.n1485 D.n1483 0.023
R12415 D.n1499 D.n1497 0.023
R12416 D.n1513 D.n1511 0.023
R12417 D.n1527 D.n1525 0.023
R12418 D.n1541 D.n1539 0.023
R12419 D.n1555 D.n1553 0.023
R12420 D.n1569 D.n1567 0.023
R12421 D.n1583 D.n1581 0.023
R12422 D.n1597 D.n1595 0.023
R12423 D.n1725 D.n1724 0.023
R12424 D.n1637 D.n1635 0.023
R12425 D.n1651 D.n1649 0.023
R12426 D.n1665 D.n1663 0.023
R12427 D.n1679 D.n1677 0.023
R12428 D.n1693 D.n1691 0.023
R12429 D.n1707 D.n1705 0.023
R12430 D.n1721 D.n1719 0.023
R12431 D.n1821 D.n1820 0.023
R12432 D.n1761 D.n1759 0.023
R12433 D.n1775 D.n1773 0.023
R12434 D.n1789 D.n1787 0.023
R12435 D.n1803 D.n1801 0.023
R12436 D.n1817 D.n1815 0.023
R12437 D.n1856 D.n1854 0.023
R12438 D.n1870 D.n1868 0.023
R12439 D.n1886 D.n1884 0.023
R12440 D.n1979 D.n1978 0.023
R12441 D.n1947 D.n1946 0.021
R12442 D.n1975 D.n1974 0.021
R12443 D.n46 D.n44 0.021
R12444 D.n3351 D.n3348 0.02
R12445 D.n2908 D.n2905 0.02
R12446 D.n2545 D.n2542 0.02
R12447 D.n2256 D.n2253 0.02
R12448 D.n2053 D.n2050 0.02
R12449 D.n565 D.n272 0.019
R12450 D.n828 D.n566 0.019
R12451 D.n1063 D.n829 0.019
R12452 D.n1270 D.n1064 0.019
R12453 D.n1449 D.n1271 0.019
R12454 D.n1601 D.n1451 0.019
R12455 D.n1725 D.n1603 0.019
R12456 D.n1821 D.n1727 0.019
R12457 D.n1978 D.n1977 0.017
R12458 D.n1914 D.n1913 0.016
R12459 D.n1921 D.n1920 0.016
R12460 D.n47 D.n46 0.016
R12461 D.n1993 D.n1986 0.016
R12462 D.n3590 D.n3580 0.016
R12463 D.n3590 D.n3589 0.016
R12464 D.n3107 D.n3097 0.016
R12465 D.n3107 D.n3106 0.016
R12466 D.n2730 D.n2729 0.016
R12467 D.n2731 D.n2730 0.016
R12468 D.n2407 D.n2406 0.016
R12469 D.n2408 D.n2407 0.016
R12470 D.n2383 D.n2373 0.016
R12471 D.n2383 D.n2382 0.016
R12472 D.n2144 D.n2134 0.016
R12473 D.n2144 D.n2143 0.016
R12474 D.n1994 D.n1993 0.016
R12475 D.n1977 D.n1967 0.016
R12476 D.n1977 D.n1976 0.016
R12477 D.n3408 D.n3407 0.016
R12478 D.n3426 D.n3425 0.016
R12479 D.n3444 D.n3443 0.016
R12480 D.n3462 D.n3461 0.016
R12481 D.n3480 D.n3479 0.016
R12482 D.n3498 D.n3497 0.016
R12483 D.n3516 D.n3515 0.016
R12484 D.n3534 D.n3533 0.016
R12485 D.n3552 D.n3551 0.016
R12486 D.n3312 D.n3311 0.016
R12487 D.n3292 D.n3291 0.016
R12488 D.n3272 D.n3271 0.016
R12489 D.n3252 D.n3251 0.016
R12490 D.n3232 D.n3231 0.016
R12491 D.n3212 D.n3211 0.016
R12492 D.n3192 D.n3191 0.016
R12493 D.n3172 D.n3171 0.016
R12494 D.n2961 D.n2960 0.016
R12495 D.n2979 D.n2978 0.016
R12496 D.n2997 D.n2996 0.016
R12497 D.n3015 D.n3014 0.016
R12498 D.n3033 D.n3032 0.016
R12499 D.n3051 D.n3050 0.016
R12500 D.n3069 D.n3068 0.016
R12501 D.n2869 D.n2868 0.016
R12502 D.n2849 D.n2848 0.016
R12503 D.n2829 D.n2828 0.016
R12504 D.n2809 D.n2808 0.016
R12505 D.n2789 D.n2788 0.016
R12506 D.n2769 D.n2768 0.016
R12507 D.n2598 D.n2597 0.016
R12508 D.n2616 D.n2615 0.016
R12509 D.n2634 D.n2633 0.016
R12510 D.n2652 D.n2651 0.016
R12511 D.n2670 D.n2669 0.016
R12512 D.n2506 D.n2505 0.016
R12513 D.n2486 D.n2485 0.016
R12514 D.n2466 D.n2465 0.016
R12515 D.n2446 D.n2445 0.016
R12516 D.n2309 D.n2308 0.016
R12517 D.n2327 D.n2326 0.016
R12518 D.n2345 D.n2344 0.016
R12519 D.n2217 D.n2216 0.016
R12520 D.n2197 D.n2196 0.016
R12521 D.n2106 D.n2105 0.016
R12522 D.n2022 D.n2021 0.016
R12523 D.n3399 D.n3390 0.016
R12524 D.n3417 D.n3409 0.016
R12525 D.n3435 D.n3427 0.016
R12526 D.n3453 D.n3445 0.016
R12527 D.n3471 D.n3463 0.016
R12528 D.n3489 D.n3481 0.016
R12529 D.n3507 D.n3499 0.016
R12530 D.n3525 D.n3517 0.016
R12531 D.n3543 D.n3535 0.016
R12532 D.n3561 D.n3553 0.016
R12533 D.n3322 D.n3315 0.016
R12534 D.n3302 D.n3295 0.016
R12535 D.n3282 D.n3275 0.016
R12536 D.n3262 D.n3255 0.016
R12537 D.n3242 D.n3235 0.016
R12538 D.n3222 D.n3215 0.016
R12539 D.n3202 D.n3195 0.016
R12540 D.n3182 D.n3175 0.016
R12541 D.n3162 D.n3155 0.016
R12542 D.n2952 D.n2943 0.016
R12543 D.n2970 D.n2962 0.016
R12544 D.n2988 D.n2980 0.016
R12545 D.n3006 D.n2998 0.016
R12546 D.n3024 D.n3016 0.016
R12547 D.n3042 D.n3034 0.016
R12548 D.n3060 D.n3052 0.016
R12549 D.n3078 D.n3070 0.016
R12550 D.n2879 D.n2872 0.016
R12551 D.n2859 D.n2852 0.016
R12552 D.n2839 D.n2832 0.016
R12553 D.n2819 D.n2812 0.016
R12554 D.n2799 D.n2792 0.016
R12555 D.n2779 D.n2772 0.016
R12556 D.n2759 D.n2752 0.016
R12557 D.n2589 D.n2580 0.016
R12558 D.n2607 D.n2599 0.016
R12559 D.n2625 D.n2617 0.016
R12560 D.n2643 D.n2635 0.016
R12561 D.n2661 D.n2653 0.016
R12562 D.n2679 D.n2671 0.016
R12563 D.n2516 D.n2509 0.016
R12564 D.n2496 D.n2489 0.016
R12565 D.n2476 D.n2469 0.016
R12566 D.n2456 D.n2449 0.016
R12567 D.n2436 D.n2429 0.016
R12568 D.n2300 D.n2291 0.016
R12569 D.n2318 D.n2310 0.016
R12570 D.n2336 D.n2328 0.016
R12571 D.n2354 D.n2346 0.016
R12572 D.n2227 D.n2220 0.016
R12573 D.n2207 D.n2200 0.016
R12574 D.n2187 D.n2180 0.016
R12575 D.n2097 D.n2088 0.016
R12576 D.n2115 D.n2107 0.016
R12577 D.n57 D.n56 0.016
R12578 D.n66 D.n65 0.016
R12579 D.n75 D.n74 0.016
R12580 D.n84 D.n83 0.016
R12581 D.n93 D.n92 0.016
R12582 D.n102 D.n101 0.016
R12583 D.n111 D.n110 0.016
R12584 D.n120 D.n119 0.016
R12585 D.n129 D.n128 0.016
R12586 D.n138 D.n137 0.016
R12587 D.n147 D.n146 0.016
R12588 D.n156 D.n155 0.016
R12589 D.n165 D.n164 0.016
R12590 D.n174 D.n173 0.016
R12591 D.n183 D.n182 0.016
R12592 D.n192 D.n191 0.016
R12593 D.n201 D.n200 0.016
R12594 D.n210 D.n209 0.016
R12595 D.n219 D.n218 0.016
R12596 D.n561 D.n549 0.016
R12597 D.n547 D.n535 0.016
R12598 D.n533 D.n521 0.016
R12599 D.n519 D.n507 0.016
R12600 D.n505 D.n493 0.016
R12601 D.n491 D.n479 0.016
R12602 D.n477 D.n465 0.016
R12603 D.n463 D.n451 0.016
R12604 D.n449 D.n437 0.016
R12605 D.n435 D.n423 0.016
R12606 D.n421 D.n409 0.016
R12607 D.n407 D.n395 0.016
R12608 D.n393 D.n381 0.016
R12609 D.n379 D.n367 0.016
R12610 D.n365 D.n353 0.016
R12611 D.n351 D.n339 0.016
R12612 D.n337 D.n325 0.016
R12613 D.n323 D.n311 0.016
R12614 D.n824 D.n812 0.016
R12615 D.n810 D.n798 0.016
R12616 D.n796 D.n784 0.016
R12617 D.n782 D.n770 0.016
R12618 D.n768 D.n756 0.016
R12619 D.n754 D.n742 0.016
R12620 D.n740 D.n728 0.016
R12621 D.n726 D.n714 0.016
R12622 D.n712 D.n700 0.016
R12623 D.n698 D.n686 0.016
R12624 D.n684 D.n672 0.016
R12625 D.n670 D.n658 0.016
R12626 D.n656 D.n644 0.016
R12627 D.n642 D.n630 0.016
R12628 D.n628 D.n616 0.016
R12629 D.n614 D.n602 0.016
R12630 D.n1059 D.n1047 0.016
R12631 D.n1045 D.n1033 0.016
R12632 D.n1031 D.n1019 0.016
R12633 D.n1017 D.n1005 0.016
R12634 D.n1003 D.n991 0.016
R12635 D.n989 D.n977 0.016
R12636 D.n975 D.n963 0.016
R12637 D.n961 D.n949 0.016
R12638 D.n947 D.n935 0.016
R12639 D.n933 D.n921 0.016
R12640 D.n919 D.n907 0.016
R12641 D.n905 D.n893 0.016
R12642 D.n891 D.n879 0.016
R12643 D.n877 D.n865 0.016
R12644 D.n1266 D.n1254 0.016
R12645 D.n1252 D.n1240 0.016
R12646 D.n1238 D.n1226 0.016
R12647 D.n1224 D.n1212 0.016
R12648 D.n1210 D.n1198 0.016
R12649 D.n1196 D.n1184 0.016
R12650 D.n1182 D.n1170 0.016
R12651 D.n1168 D.n1156 0.016
R12652 D.n1154 D.n1142 0.016
R12653 D.n1140 D.n1128 0.016
R12654 D.n1126 D.n1114 0.016
R12655 D.n1112 D.n1100 0.016
R12656 D.n1445 D.n1433 0.016
R12657 D.n1431 D.n1419 0.016
R12658 D.n1417 D.n1405 0.016
R12659 D.n1403 D.n1391 0.016
R12660 D.n1389 D.n1377 0.016
R12661 D.n1375 D.n1363 0.016
R12662 D.n1361 D.n1349 0.016
R12663 D.n1347 D.n1335 0.016
R12664 D.n1333 D.n1321 0.016
R12665 D.n1319 D.n1307 0.016
R12666 D.n1597 D.n1585 0.016
R12667 D.n1583 D.n1571 0.016
R12668 D.n1569 D.n1557 0.016
R12669 D.n1555 D.n1543 0.016
R12670 D.n1541 D.n1529 0.016
R12671 D.n1527 D.n1515 0.016
R12672 D.n1513 D.n1501 0.016
R12673 D.n1499 D.n1487 0.016
R12674 D.n1721 D.n1709 0.016
R12675 D.n1707 D.n1695 0.016
R12676 D.n1693 D.n1681 0.016
R12677 D.n1679 D.n1667 0.016
R12678 D.n1665 D.n1653 0.016
R12679 D.n1651 D.n1639 0.016
R12680 D.n1817 D.n1805 0.016
R12681 D.n1803 D.n1791 0.016
R12682 D.n1789 D.n1777 0.016
R12683 D.n1775 D.n1763 0.016
R12684 D.n1886 D.n1872 0.016
R12685 D.n1870 D.n1858 0.016
R12686 D.n565 D.n280 0.016
R12687 D.n828 D.n571 0.016
R12688 D.n1063 D.n834 0.016
R12689 D.n1270 D.n1069 0.016
R12690 D.n1449 D.n1276 0.016
R12691 D.n1601 D.n1456 0.016
R12692 D.n1725 D.n1608 0.016
R12693 D.n1821 D.n1732 0.016
R12694 D.n1888 D.n1827 0.016
R12695 D.n1921 D.n1918 0.016
R12696 D.n1928 D.n1923 0.016
R12697 D.n1928 D.n1927 0.016
R12698 D.n3128 D.n3127 0.015
R12699 D.n2719 D.n2718 0.015
R12700 D.n2396 D.n2395 0.015
R12701 D.n2153 D.n2152 0.015
R12702 D.n2035 D.n2034 0.015
R12703 D.n2009 D.n2008 0.015
R12704 D.n3579 D.n3578 0.015
R12705 D.n3564 D.n3563 0.015
R12706 D.n3149 D.n3148 0.015
R12707 D.n3139 D.n3138 0.015
R12708 D.n3096 D.n3095 0.015
R12709 D.n3081 D.n3080 0.015
R12710 D.n2746 D.n2745 0.015
R12711 D.n2734 D.n2732 0.015
R12712 D.n2701 D.n2700 0.015
R12713 D.n2681 D.n2680 0.015
R12714 D.n2423 D.n2422 0.015
R12715 D.n2411 D.n2409 0.015
R12716 D.n2372 D.n2371 0.015
R12717 D.n2357 D.n2356 0.015
R12718 D.n2174 D.n2173 0.015
R12719 D.n2164 D.n2163 0.015
R12720 D.n2133 D.n2132 0.015
R12721 D.n2118 D.n2117 0.015
R12722 D.n1997 D.n1995 0.015
R12723 D.n262 D.n13 0.014
R12724 D.n42 D.n41 0.013
R12725 D.n24 D.n23 0.013
R12726 D.n307 D.n306 0.013
R12727 D.n321 D.n320 0.013
R12728 D.n335 D.n334 0.013
R12729 D.n349 D.n348 0.013
R12730 D.n363 D.n362 0.013
R12731 D.n377 D.n376 0.013
R12732 D.n391 D.n390 0.013
R12733 D.n405 D.n404 0.013
R12734 D.n419 D.n418 0.013
R12735 D.n433 D.n432 0.013
R12736 D.n447 D.n446 0.013
R12737 D.n461 D.n460 0.013
R12738 D.n475 D.n474 0.013
R12739 D.n489 D.n488 0.013
R12740 D.n503 D.n502 0.013
R12741 D.n517 D.n516 0.013
R12742 D.n531 D.n530 0.013
R12743 D.n545 D.n544 0.013
R12744 D.n559 D.n558 0.013
R12745 D.n564 D.n563 0.013
R12746 D.n598 D.n597 0.013
R12747 D.n612 D.n611 0.013
R12748 D.n626 D.n625 0.013
R12749 D.n640 D.n639 0.013
R12750 D.n654 D.n653 0.013
R12751 D.n668 D.n667 0.013
R12752 D.n682 D.n681 0.013
R12753 D.n696 D.n695 0.013
R12754 D.n710 D.n709 0.013
R12755 D.n724 D.n723 0.013
R12756 D.n738 D.n737 0.013
R12757 D.n752 D.n751 0.013
R12758 D.n766 D.n765 0.013
R12759 D.n780 D.n779 0.013
R12760 D.n794 D.n793 0.013
R12761 D.n808 D.n807 0.013
R12762 D.n822 D.n821 0.013
R12763 D.n827 D.n826 0.013
R12764 D.n861 D.n860 0.013
R12765 D.n875 D.n874 0.013
R12766 D.n889 D.n888 0.013
R12767 D.n903 D.n902 0.013
R12768 D.n917 D.n916 0.013
R12769 D.n931 D.n930 0.013
R12770 D.n945 D.n944 0.013
R12771 D.n959 D.n958 0.013
R12772 D.n973 D.n972 0.013
R12773 D.n987 D.n986 0.013
R12774 D.n1001 D.n1000 0.013
R12775 D.n1015 D.n1014 0.013
R12776 D.n1029 D.n1028 0.013
R12777 D.n1043 D.n1042 0.013
R12778 D.n1057 D.n1056 0.013
R12779 D.n1062 D.n1061 0.013
R12780 D.n1096 D.n1095 0.013
R12781 D.n1110 D.n1109 0.013
R12782 D.n1124 D.n1123 0.013
R12783 D.n1138 D.n1137 0.013
R12784 D.n1152 D.n1151 0.013
R12785 D.n1166 D.n1165 0.013
R12786 D.n1180 D.n1179 0.013
R12787 D.n1194 D.n1193 0.013
R12788 D.n1208 D.n1207 0.013
R12789 D.n1222 D.n1221 0.013
R12790 D.n1236 D.n1235 0.013
R12791 D.n1250 D.n1249 0.013
R12792 D.n1264 D.n1263 0.013
R12793 D.n1269 D.n1268 0.013
R12794 D.n1303 D.n1302 0.013
R12795 D.n1317 D.n1316 0.013
R12796 D.n1331 D.n1330 0.013
R12797 D.n1345 D.n1344 0.013
R12798 D.n1359 D.n1358 0.013
R12799 D.n1373 D.n1372 0.013
R12800 D.n1387 D.n1386 0.013
R12801 D.n1401 D.n1400 0.013
R12802 D.n1415 D.n1414 0.013
R12803 D.n1429 D.n1428 0.013
R12804 D.n1443 D.n1442 0.013
R12805 D.n1448 D.n1447 0.013
R12806 D.n1483 D.n1482 0.013
R12807 D.n1497 D.n1496 0.013
R12808 D.n1511 D.n1510 0.013
R12809 D.n1525 D.n1524 0.013
R12810 D.n1539 D.n1538 0.013
R12811 D.n1553 D.n1552 0.013
R12812 D.n1567 D.n1566 0.013
R12813 D.n1581 D.n1580 0.013
R12814 D.n1595 D.n1594 0.013
R12815 D.n1600 D.n1599 0.013
R12816 D.n1635 D.n1634 0.013
R12817 D.n1649 D.n1648 0.013
R12818 D.n1663 D.n1662 0.013
R12819 D.n1677 D.n1676 0.013
R12820 D.n1691 D.n1690 0.013
R12821 D.n1705 D.n1704 0.013
R12822 D.n1719 D.n1718 0.013
R12823 D.n1724 D.n1723 0.013
R12824 D.n1759 D.n1758 0.013
R12825 D.n1773 D.n1772 0.013
R12826 D.n1787 D.n1786 0.013
R12827 D.n1801 D.n1800 0.013
R12828 D.n1815 D.n1814 0.013
R12829 D.n1820 D.n1819 0.013
R12830 D.n1854 D.n1853 0.013
R12831 D.n1868 D.n1867 0.013
R12832 D.n1884 D.n1883 0.013
R12833 D.n3368 D.n3367 0.012
R12834 D.n3333 D.n3332 0.012
R12835 D.n2925 D.n2924 0.012
R12836 D.n2890 D.n2889 0.012
R12837 D.n2562 D.n2561 0.012
R12838 D.n2527 D.n2526 0.012
R12839 D.n2273 D.n2272 0.012
R12840 D.n2238 D.n2237 0.012
R12841 D.n2070 D.n2069 0.012
R12842 D.n2033 D.n2032 0.012
R12843 D.n237 D.n236 0.011
R12844 D.n1915 D.n1914 0.011
R12845 D.n3399 D.n3398 0.011
R12846 D.n3417 D.n3416 0.011
R12847 D.n3435 D.n3434 0.011
R12848 D.n3453 D.n3452 0.011
R12849 D.n3471 D.n3470 0.011
R12850 D.n3489 D.n3488 0.011
R12851 D.n3507 D.n3506 0.011
R12852 D.n3525 D.n3524 0.011
R12853 D.n3543 D.n3542 0.011
R12854 D.n3561 D.n3560 0.011
R12855 D.n3323 D.n3322 0.011
R12856 D.n3303 D.n3302 0.011
R12857 D.n3283 D.n3282 0.011
R12858 D.n3263 D.n3262 0.011
R12859 D.n3243 D.n3242 0.011
R12860 D.n3223 D.n3222 0.011
R12861 D.n3203 D.n3202 0.011
R12862 D.n3183 D.n3182 0.011
R12863 D.n3163 D.n3162 0.011
R12864 D.n2952 D.n2951 0.011
R12865 D.n2970 D.n2969 0.011
R12866 D.n2988 D.n2987 0.011
R12867 D.n3006 D.n3005 0.011
R12868 D.n3024 D.n3023 0.011
R12869 D.n3042 D.n3041 0.011
R12870 D.n3060 D.n3059 0.011
R12871 D.n3078 D.n3077 0.011
R12872 D.n2880 D.n2879 0.011
R12873 D.n2860 D.n2859 0.011
R12874 D.n2840 D.n2839 0.011
R12875 D.n2820 D.n2819 0.011
R12876 D.n2800 D.n2799 0.011
R12877 D.n2780 D.n2779 0.011
R12878 D.n2760 D.n2759 0.011
R12879 D.n2589 D.n2588 0.011
R12880 D.n2607 D.n2606 0.011
R12881 D.n2625 D.n2624 0.011
R12882 D.n2643 D.n2642 0.011
R12883 D.n2661 D.n2660 0.011
R12884 D.n2679 D.n2678 0.011
R12885 D.n2517 D.n2516 0.011
R12886 D.n2497 D.n2496 0.011
R12887 D.n2477 D.n2476 0.011
R12888 D.n2457 D.n2456 0.011
R12889 D.n2437 D.n2436 0.011
R12890 D.n2300 D.n2299 0.011
R12891 D.n2318 D.n2317 0.011
R12892 D.n2336 D.n2335 0.011
R12893 D.n2354 D.n2353 0.011
R12894 D.n2228 D.n2227 0.011
R12895 D.n2208 D.n2207 0.011
R12896 D.n2188 D.n2187 0.011
R12897 D.n2097 D.n2096 0.011
R12898 D.n2115 D.n2114 0.011
R12899 D.n2023 D.n2022 0.011
R12900 D.n228 D.n227 0.011
R12901 D.n219 D.n211 0.011
R12902 D.n210 D.n202 0.011
R12903 D.n201 D.n193 0.011
R12904 D.n192 D.n184 0.011
R12905 D.n183 D.n175 0.011
R12906 D.n174 D.n166 0.011
R12907 D.n165 D.n157 0.011
R12908 D.n156 D.n148 0.011
R12909 D.n147 D.n139 0.011
R12910 D.n138 D.n130 0.011
R12911 D.n129 D.n121 0.011
R12912 D.n120 D.n112 0.011
R12913 D.n111 D.n103 0.011
R12914 D.n102 D.n94 0.011
R12915 D.n93 D.n85 0.011
R12916 D.n84 D.n76 0.011
R12917 D.n75 D.n67 0.011
R12918 D.n66 D.n58 0.011
R12919 D.n57 D.n49 0.011
R12920 D.n1905 D.n1904 0.011
R12921 D.n1888 D.n1822 0.011
R12922 D.n2 D.n1 0.01
R12923 D.n3408 D.n3400 0.01
R12924 D.n3426 D.n3418 0.01
R12925 D.n3444 D.n3436 0.01
R12926 D.n3462 D.n3454 0.01
R12927 D.n3480 D.n3472 0.01
R12928 D.n3498 D.n3490 0.01
R12929 D.n3516 D.n3508 0.01
R12930 D.n3534 D.n3526 0.01
R12931 D.n3552 D.n3544 0.01
R12932 D.n3313 D.n3312 0.01
R12933 D.n3293 D.n3292 0.01
R12934 D.n3273 D.n3272 0.01
R12935 D.n3253 D.n3252 0.01
R12936 D.n3233 D.n3232 0.01
R12937 D.n3213 D.n3212 0.01
R12938 D.n3193 D.n3192 0.01
R12939 D.n3173 D.n3172 0.01
R12940 D.n2961 D.n2953 0.01
R12941 D.n2979 D.n2971 0.01
R12942 D.n2997 D.n2989 0.01
R12943 D.n3015 D.n3007 0.01
R12944 D.n3033 D.n3025 0.01
R12945 D.n3051 D.n3043 0.01
R12946 D.n3069 D.n3061 0.01
R12947 D.n2870 D.n2869 0.01
R12948 D.n2850 D.n2849 0.01
R12949 D.n2830 D.n2829 0.01
R12950 D.n2810 D.n2809 0.01
R12951 D.n2790 D.n2789 0.01
R12952 D.n2770 D.n2769 0.01
R12953 D.n2598 D.n2590 0.01
R12954 D.n2616 D.n2608 0.01
R12955 D.n2634 D.n2626 0.01
R12956 D.n2652 D.n2644 0.01
R12957 D.n2670 D.n2662 0.01
R12958 D.n2507 D.n2506 0.01
R12959 D.n2487 D.n2486 0.01
R12960 D.n2467 D.n2466 0.01
R12961 D.n2447 D.n2446 0.01
R12962 D.n2309 D.n2301 0.01
R12963 D.n2327 D.n2319 0.01
R12964 D.n2345 D.n2337 0.01
R12965 D.n2218 D.n2217 0.01
R12966 D.n2198 D.n2197 0.01
R12967 D.n2106 D.n2098 0.01
R12968 D.n2063 D.n2062 0.01
R12969 D.n2079 D.n2078 0.01
R12970 D.n3362 D.n3359 0.01
R12971 D.n3382 D.n3379 0.01
R12972 D.n3361 D.n3360 0.01
R12973 D.n3381 D.n3380 0.01
R12974 D.n2919 D.n2916 0.01
R12975 D.n2935 D.n2932 0.01
R12976 D.n2918 D.n2917 0.01
R12977 D.n2934 D.n2933 0.01
R12978 D.n2556 D.n2553 0.01
R12979 D.n2572 D.n2569 0.01
R12980 D.n2555 D.n2554 0.01
R12981 D.n2571 D.n2570 0.01
R12982 D.n2267 D.n2264 0.01
R12983 D.n2283 D.n2280 0.01
R12984 D.n2266 D.n2265 0.01
R12985 D.n2282 D.n2281 0.01
R12986 D.n2064 D.n2061 0.01
R12987 D.n2080 D.n2077 0.01
R12988 D.n295 D.n294 0.01
R12989 D.n586 D.n585 0.01
R12990 D.n849 D.n848 0.01
R12991 D.n1084 D.n1083 0.01
R12992 D.n1291 D.n1290 0.01
R12993 D.n1471 D.n1470 0.01
R12994 D.n1623 D.n1622 0.01
R12995 D.n1747 D.n1746 0.01
R12996 D.n1842 D.n1841 0.01
R12997 D.n3575 D.n3574 0.009
R12998 D.n3152 D.n3151 0.009
R12999 D.n3091 D.n3090 0.009
R13000 D.n2749 D.n2748 0.009
R13001 D.n2692 D.n2691 0.009
R13002 D.n2426 D.n2425 0.009
R13003 D.n2367 D.n2366 0.009
R13004 D.n2177 D.n2176 0.009
R13005 D.n2128 D.n2127 0.009
R13006 D.n3377 D.n3376 0.009
R13007 D.n269 D.n268 0.009
R13008 D.n3347 D.n3346 0.009
R13009 D.n2904 D.n2903 0.009
R13010 D.n2541 D.n2540 0.009
R13011 D.n2252 D.n2251 0.009
R13012 D.n2049 D.n2048 0.009
R13013 D.n2012 D.n2011 0.009
R13014 D.n22 D.n21 0.008
R13015 D.n3575 D.n3566 0.008
R13016 D.n3153 D.n3152 0.008
R13017 D.n3091 D.n3083 0.008
R13018 D.n2750 D.n2749 0.008
R13019 D.n2692 D.n2683 0.008
R13020 D.n2427 D.n2426 0.008
R13021 D.n2367 D.n2359 0.008
R13022 D.n2178 D.n2177 0.008
R13023 D.n2128 D.n2120 0.008
R13024 D.n2013 D.n2012 0.008
R13025 D.n3137 D.n3136 0.007
R13026 D.n3137 D.n3131 0.007
R13027 D.n2702 D.n2699 0.007
R13028 D.n2702 D.n2694 0.007
R13029 D.n2162 D.n2161 0.007
R13030 D.n2162 D.n2156 0.007
R13031 D.n237 D.n229 0.006
R13032 D.n22 D.n19 0.006
R13033 D.n268 D.n262 0.006
R13034 D.n40 D.n37 0.006
R13035 D.n40 D.n39 0.006
R13036 D.n1966 D.n1965 0.006
R13037 D.n295 D.n281 0.006
R13038 D.n586 D.n572 0.006
R13039 D.n849 D.n835 0.006
R13040 D.n1084 D.n1070 0.006
R13041 D.n1291 D.n1277 0.006
R13042 D.n1471 D.n1457 0.006
R13043 D.n1623 D.n1609 0.006
R13044 D.n1747 D.n1733 0.006
R13045 D.n1842 D.n1828 0.006
R13046 D.n228 D.n220 0.006
R13047 D.n309 D.n297 0.006
R13048 D.n600 D.n588 0.006
R13049 D.n863 D.n851 0.006
R13050 D.n1098 D.n1086 0.006
R13051 D.n1305 D.n1293 0.006
R13052 D.n1485 D.n1473 0.006
R13053 D.n1637 D.n1625 0.006
R13054 D.n1761 D.n1749 0.006
R13055 D.n1856 D.n1844 0.006
R13056 D.n1904 D.n1903 0.005
R13057 D.n270 D.n269 0.005
R13058 D.n3351 D.n3350 0.005
R13059 D.n2908 D.n2907 0.005
R13060 D.n2545 D.n2544 0.005
R13061 D.n2256 D.n2255 0.005
R13062 D.n2053 D.n2052 0.005
R13063 D.n2028 D.n2027 0.004
R13064 D.n2042 D.n2041 0.004
R13065 D.n3363 D.n3358 0.004
R13066 D.n3383 D.n3374 0.004
R13067 D.n3328 D.n3327 0.004
R13068 D.n3340 D.n3339 0.004
R13069 D.n2920 D.n2915 0.004
R13070 D.n2936 D.n2931 0.004
R13071 D.n2885 D.n2884 0.004
R13072 D.n2897 D.n2896 0.004
R13073 D.n2557 D.n2552 0.004
R13074 D.n2573 D.n2568 0.004
R13075 D.n2522 D.n2521 0.004
R13076 D.n2534 D.n2533 0.004
R13077 D.n2268 D.n2263 0.004
R13078 D.n2284 D.n2279 0.004
R13079 D.n2233 D.n2232 0.004
R13080 D.n2245 D.n2244 0.004
R13081 D.n2065 D.n2060 0.004
R13082 D.n2081 D.n2076 0.004
R13083 D.n3354 D.n3126 0.004
R13084 D.n2911 D.n2717 0.004
R13085 D.n2548 D.n2394 0.004
R13086 D.n2259 D.n2151 0.004
R13087 D.n2056 D.n1982 0.004
R13088 D.n3350 D.n3349 0.004
R13089 D.n2907 D.n2906 0.004
R13090 D.n2544 D.n2543 0.004
R13091 D.n2255 D.n2254 0.004
R13092 D.n1980 D.n1963 0.004
R13093 D.n1977 D.n1966 0.004
R13094 D.n2052 D.n2051 0.004
R13095 D.n3346 D.n3128 0.004
R13096 D.n2903 D.n2719 0.004
R13097 D.n2540 D.n2396 0.004
R13098 D.n2251 D.n2153 0.004
R13099 D.n2048 D.n2035 0.004
R13100 D.n291 D.n290 0.003
R13101 D.n582 D.n581 0.003
R13102 D.n845 D.n844 0.003
R13103 D.n1080 D.n1079 0.003
R13104 D.n1287 D.n1286 0.003
R13105 D.n1467 D.n1466 0.003
R13106 D.n1619 D.n1618 0.003
R13107 D.n1743 D.n1742 0.003
R13108 D.n1838 D.n1837 0.003
R13109 D.n1930 D.n1929 0.003
R13110 D.n1893 D.n1892 0.003
R13111 D.n1953 D.n1952 0.003
R13112 D.n2037 D.n2036 0.003
R13113 D.n3370 D.n3369 0.003
R13114 D.n3335 D.n3334 0.003
R13115 D.n2927 D.n2926 0.003
R13116 D.n2892 D.n2891 0.003
R13117 D.n2564 D.n2563 0.003
R13118 D.n2529 D.n2528 0.003
R13119 D.n2275 D.n2274 0.003
R13120 D.n2240 D.n2239 0.003
R13121 D.n2072 D.n2071 0.003
R13122 D.n1909 D.n1907 0.003
R13123 D.n1899 D.n1897 0.003
R13124 D.n232 D.n231 0.003
R13125 D.n223 D.n222 0.003
R13126 D.n30 D.n28 0.003
R13127 D.n2017 D.n2015 0.003
R13128 D.n2002 D.n2000 0.003
R13129 D.n3556 D.n3555 0.003
R13130 D.n3538 D.n3537 0.003
R13131 D.n3520 D.n3519 0.003
R13132 D.n3502 D.n3501 0.003
R13133 D.n3484 D.n3483 0.003
R13134 D.n3466 D.n3465 0.003
R13135 D.n3448 D.n3447 0.003
R13136 D.n3430 D.n3429 0.003
R13137 D.n3412 D.n3411 0.003
R13138 D.n3393 D.n3392 0.003
R13139 D.n3403 D.n3401 0.003
R13140 D.n3421 D.n3419 0.003
R13141 D.n3439 D.n3437 0.003
R13142 D.n3457 D.n3455 0.003
R13143 D.n3475 D.n3473 0.003
R13144 D.n3493 D.n3491 0.003
R13145 D.n3511 D.n3509 0.003
R13146 D.n3529 D.n3527 0.003
R13147 D.n3547 D.n3545 0.003
R13148 D.n3569 D.n3567 0.003
R13149 D.n3158 D.n3157 0.003
R13150 D.n3178 D.n3177 0.003
R13151 D.n3198 D.n3197 0.003
R13152 D.n3218 D.n3217 0.003
R13153 D.n3238 D.n3237 0.003
R13154 D.n3258 D.n3257 0.003
R13155 D.n3278 D.n3277 0.003
R13156 D.n3298 D.n3297 0.003
R13157 D.n3318 D.n3317 0.003
R13158 D.n3307 D.n3305 0.003
R13159 D.n3287 D.n3285 0.003
R13160 D.n3267 D.n3265 0.003
R13161 D.n3247 D.n3245 0.003
R13162 D.n3227 D.n3225 0.003
R13163 D.n3207 D.n3205 0.003
R13164 D.n3187 D.n3185 0.003
R13165 D.n3167 D.n3165 0.003
R13166 D.n3144 D.n3142 0.003
R13167 D.n3073 D.n3072 0.003
R13168 D.n3055 D.n3054 0.003
R13169 D.n3037 D.n3036 0.003
R13170 D.n3019 D.n3018 0.003
R13171 D.n3001 D.n3000 0.003
R13172 D.n2983 D.n2982 0.003
R13173 D.n2965 D.n2964 0.003
R13174 D.n2946 D.n2945 0.003
R13175 D.n2956 D.n2954 0.003
R13176 D.n2974 D.n2972 0.003
R13177 D.n2992 D.n2990 0.003
R13178 D.n3010 D.n3008 0.003
R13179 D.n3028 D.n3026 0.003
R13180 D.n3046 D.n3044 0.003
R13181 D.n3064 D.n3062 0.003
R13182 D.n3086 D.n3084 0.003
R13183 D.n2755 D.n2754 0.003
R13184 D.n2775 D.n2774 0.003
R13185 D.n2795 D.n2794 0.003
R13186 D.n2815 D.n2814 0.003
R13187 D.n2835 D.n2834 0.003
R13188 D.n2855 D.n2854 0.003
R13189 D.n2875 D.n2874 0.003
R13190 D.n2864 D.n2862 0.003
R13191 D.n2844 D.n2842 0.003
R13192 D.n2824 D.n2822 0.003
R13193 D.n2804 D.n2802 0.003
R13194 D.n2784 D.n2782 0.003
R13195 D.n2764 D.n2762 0.003
R13196 D.n2739 D.n2737 0.003
R13197 D.n2674 D.n2673 0.003
R13198 D.n2656 D.n2655 0.003
R13199 D.n2638 D.n2637 0.003
R13200 D.n2620 D.n2619 0.003
R13201 D.n2602 D.n2601 0.003
R13202 D.n2583 D.n2582 0.003
R13203 D.n2593 D.n2591 0.003
R13204 D.n2611 D.n2609 0.003
R13205 D.n2629 D.n2627 0.003
R13206 D.n2647 D.n2645 0.003
R13207 D.n2665 D.n2663 0.003
R13208 D.n2686 D.n2684 0.003
R13209 D.n2432 D.n2431 0.003
R13210 D.n2452 D.n2451 0.003
R13211 D.n2472 D.n2471 0.003
R13212 D.n2492 D.n2491 0.003
R13213 D.n2512 D.n2511 0.003
R13214 D.n2501 D.n2499 0.003
R13215 D.n2481 D.n2479 0.003
R13216 D.n2461 D.n2459 0.003
R13217 D.n2441 D.n2439 0.003
R13218 D.n2416 D.n2414 0.003
R13219 D.n2349 D.n2348 0.003
R13220 D.n2331 D.n2330 0.003
R13221 D.n2313 D.n2312 0.003
R13222 D.n2294 D.n2293 0.003
R13223 D.n2304 D.n2302 0.003
R13224 D.n2322 D.n2320 0.003
R13225 D.n2340 D.n2338 0.003
R13226 D.n2362 D.n2360 0.003
R13227 D.n2183 D.n2182 0.003
R13228 D.n2203 D.n2202 0.003
R13229 D.n2223 D.n2222 0.003
R13230 D.n2212 D.n2210 0.003
R13231 D.n2192 D.n2190 0.003
R13232 D.n2169 D.n2167 0.003
R13233 D.n2110 D.n2109 0.003
R13234 D.n2091 D.n2090 0.003
R13235 D.n2101 D.n2099 0.003
R13236 D.n2123 D.n2121 0.003
R13237 D.n52 D.n50 0.003
R13238 D.n61 D.n59 0.003
R13239 D.n70 D.n68 0.003
R13240 D.n79 D.n77 0.003
R13241 D.n88 D.n86 0.003
R13242 D.n97 D.n95 0.003
R13243 D.n106 D.n104 0.003
R13244 D.n115 D.n113 0.003
R13245 D.n124 D.n122 0.003
R13246 D.n133 D.n131 0.003
R13247 D.n142 D.n140 0.003
R13248 D.n151 D.n149 0.003
R13249 D.n160 D.n158 0.003
R13250 D.n169 D.n167 0.003
R13251 D.n178 D.n176 0.003
R13252 D.n187 D.n185 0.003
R13253 D.n196 D.n194 0.003
R13254 D.n205 D.n203 0.003
R13255 D.n214 D.n212 0.003
R13256 D.n284 D.n283 0.003
R13257 D.n300 D.n299 0.003
R13258 D.n552 D.n551 0.003
R13259 D.n538 D.n537 0.003
R13260 D.n524 D.n523 0.003
R13261 D.n510 D.n509 0.003
R13262 D.n496 D.n495 0.003
R13263 D.n482 D.n481 0.003
R13264 D.n468 D.n467 0.003
R13265 D.n454 D.n453 0.003
R13266 D.n440 D.n439 0.003
R13267 D.n426 D.n425 0.003
R13268 D.n412 D.n411 0.003
R13269 D.n398 D.n397 0.003
R13270 D.n384 D.n383 0.003
R13271 D.n370 D.n369 0.003
R13272 D.n356 D.n355 0.003
R13273 D.n342 D.n341 0.003
R13274 D.n328 D.n327 0.003
R13275 D.n314 D.n313 0.003
R13276 D.n575 D.n574 0.003
R13277 D.n591 D.n590 0.003
R13278 D.n815 D.n814 0.003
R13279 D.n801 D.n800 0.003
R13280 D.n787 D.n786 0.003
R13281 D.n773 D.n772 0.003
R13282 D.n759 D.n758 0.003
R13283 D.n745 D.n744 0.003
R13284 D.n731 D.n730 0.003
R13285 D.n717 D.n716 0.003
R13286 D.n703 D.n702 0.003
R13287 D.n689 D.n688 0.003
R13288 D.n675 D.n674 0.003
R13289 D.n661 D.n660 0.003
R13290 D.n647 D.n646 0.003
R13291 D.n633 D.n632 0.003
R13292 D.n619 D.n618 0.003
R13293 D.n605 D.n604 0.003
R13294 D.n838 D.n837 0.003
R13295 D.n854 D.n853 0.003
R13296 D.n1050 D.n1049 0.003
R13297 D.n1036 D.n1035 0.003
R13298 D.n1022 D.n1021 0.003
R13299 D.n1008 D.n1007 0.003
R13300 D.n994 D.n993 0.003
R13301 D.n980 D.n979 0.003
R13302 D.n966 D.n965 0.003
R13303 D.n952 D.n951 0.003
R13304 D.n938 D.n937 0.003
R13305 D.n924 D.n923 0.003
R13306 D.n910 D.n909 0.003
R13307 D.n896 D.n895 0.003
R13308 D.n882 D.n881 0.003
R13309 D.n868 D.n867 0.003
R13310 D.n1073 D.n1072 0.003
R13311 D.n1089 D.n1088 0.003
R13312 D.n1257 D.n1256 0.003
R13313 D.n1243 D.n1242 0.003
R13314 D.n1229 D.n1228 0.003
R13315 D.n1215 D.n1214 0.003
R13316 D.n1201 D.n1200 0.003
R13317 D.n1187 D.n1186 0.003
R13318 D.n1173 D.n1172 0.003
R13319 D.n1159 D.n1158 0.003
R13320 D.n1145 D.n1144 0.003
R13321 D.n1131 D.n1130 0.003
R13322 D.n1117 D.n1116 0.003
R13323 D.n1103 D.n1102 0.003
R13324 D.n1280 D.n1279 0.003
R13325 D.n1296 D.n1295 0.003
R13326 D.n1436 D.n1435 0.003
R13327 D.n1422 D.n1421 0.003
R13328 D.n1408 D.n1407 0.003
R13329 D.n1394 D.n1393 0.003
R13330 D.n1380 D.n1379 0.003
R13331 D.n1366 D.n1365 0.003
R13332 D.n1352 D.n1351 0.003
R13333 D.n1338 D.n1337 0.003
R13334 D.n1324 D.n1323 0.003
R13335 D.n1310 D.n1309 0.003
R13336 D.n1460 D.n1459 0.003
R13337 D.n1476 D.n1475 0.003
R13338 D.n1588 D.n1587 0.003
R13339 D.n1574 D.n1573 0.003
R13340 D.n1560 D.n1559 0.003
R13341 D.n1546 D.n1545 0.003
R13342 D.n1532 D.n1531 0.003
R13343 D.n1518 D.n1517 0.003
R13344 D.n1504 D.n1503 0.003
R13345 D.n1490 D.n1489 0.003
R13346 D.n1612 D.n1611 0.003
R13347 D.n1628 D.n1627 0.003
R13348 D.n1712 D.n1711 0.003
R13349 D.n1698 D.n1697 0.003
R13350 D.n1684 D.n1683 0.003
R13351 D.n1670 D.n1669 0.003
R13352 D.n1656 D.n1655 0.003
R13353 D.n1642 D.n1641 0.003
R13354 D.n1736 D.n1735 0.003
R13355 D.n1752 D.n1751 0.003
R13356 D.n1808 D.n1807 0.003
R13357 D.n1794 D.n1793 0.003
R13358 D.n1780 D.n1779 0.003
R13359 D.n1766 D.n1765 0.003
R13360 D.n1831 D.n1830 0.003
R13361 D.n1847 D.n1846 0.003
R13362 D.n1875 D.n1874 0.003
R13363 D.n1861 D.n1860 0.003
R13364 D.n1926 D.n1925 0.003
R13365 D.n1890 D.n1889 0.003
R13366 D.n1912 D.n1910 0.003
R13367 D.n1902 D.n1900 0.003
R13368 D.n235 D.n233 0.003
R13369 D.n226 D.n224 0.003
R13370 D.n33 D.n31 0.003
R13371 D.n1991 D.n1990 0.003
R13372 D.n2020 D.n2018 0.003
R13373 D.n2005 D.n2003 0.003
R13374 D.n3559 D.n3557 0.003
R13375 D.n3541 D.n3539 0.003
R13376 D.n3523 D.n3521 0.003
R13377 D.n3505 D.n3503 0.003
R13378 D.n3487 D.n3485 0.003
R13379 D.n3469 D.n3467 0.003
R13380 D.n3451 D.n3449 0.003
R13381 D.n3433 D.n3431 0.003
R13382 D.n3415 D.n3413 0.003
R13383 D.n3396 D.n3394 0.003
R13384 D.n3406 D.n3404 0.003
R13385 D.n3424 D.n3422 0.003
R13386 D.n3442 D.n3440 0.003
R13387 D.n3460 D.n3458 0.003
R13388 D.n3478 D.n3476 0.003
R13389 D.n3496 D.n3494 0.003
R13390 D.n3514 D.n3512 0.003
R13391 D.n3532 D.n3530 0.003
R13392 D.n3550 D.n3548 0.003
R13393 D.n3572 D.n3570 0.003
R13394 D.n3585 D.n3584 0.003
R13395 D.n3161 D.n3159 0.003
R13396 D.n3181 D.n3179 0.003
R13397 D.n3201 D.n3199 0.003
R13398 D.n3221 D.n3219 0.003
R13399 D.n3241 D.n3239 0.003
R13400 D.n3261 D.n3259 0.003
R13401 D.n3281 D.n3279 0.003
R13402 D.n3301 D.n3299 0.003
R13403 D.n3321 D.n3319 0.003
R13404 D.n3310 D.n3308 0.003
R13405 D.n3290 D.n3288 0.003
R13406 D.n3270 D.n3268 0.003
R13407 D.n3250 D.n3248 0.003
R13408 D.n3230 D.n3228 0.003
R13409 D.n3210 D.n3208 0.003
R13410 D.n3190 D.n3188 0.003
R13411 D.n3170 D.n3168 0.003
R13412 D.n3147 D.n3145 0.003
R13413 D.n3133 D.n3132 0.003
R13414 D.n3076 D.n3074 0.003
R13415 D.n3058 D.n3056 0.003
R13416 D.n3040 D.n3038 0.003
R13417 D.n3022 D.n3020 0.003
R13418 D.n3004 D.n3002 0.003
R13419 D.n2986 D.n2984 0.003
R13420 D.n2968 D.n2966 0.003
R13421 D.n2949 D.n2947 0.003
R13422 D.n2959 D.n2957 0.003
R13423 D.n2977 D.n2975 0.003
R13424 D.n2995 D.n2993 0.003
R13425 D.n3013 D.n3011 0.003
R13426 D.n3031 D.n3029 0.003
R13427 D.n3049 D.n3047 0.003
R13428 D.n3067 D.n3065 0.003
R13429 D.n3089 D.n3087 0.003
R13430 D.n3102 D.n3101 0.003
R13431 D.n2758 D.n2756 0.003
R13432 D.n2778 D.n2776 0.003
R13433 D.n2798 D.n2796 0.003
R13434 D.n2818 D.n2816 0.003
R13435 D.n2838 D.n2836 0.003
R13436 D.n2858 D.n2856 0.003
R13437 D.n2878 D.n2876 0.003
R13438 D.n2867 D.n2865 0.003
R13439 D.n2847 D.n2845 0.003
R13440 D.n2827 D.n2825 0.003
R13441 D.n2807 D.n2805 0.003
R13442 D.n2787 D.n2785 0.003
R13443 D.n2767 D.n2765 0.003
R13444 D.n2742 D.n2740 0.003
R13445 D.n2725 D.n2724 0.003
R13446 D.n2677 D.n2675 0.003
R13447 D.n2659 D.n2657 0.003
R13448 D.n2641 D.n2639 0.003
R13449 D.n2623 D.n2621 0.003
R13450 D.n2605 D.n2603 0.003
R13451 D.n2586 D.n2584 0.003
R13452 D.n2596 D.n2594 0.003
R13453 D.n2614 D.n2612 0.003
R13454 D.n2632 D.n2630 0.003
R13455 D.n2650 D.n2648 0.003
R13456 D.n2668 D.n2666 0.003
R13457 D.n2689 D.n2687 0.003
R13458 D.n2696 D.n2695 0.003
R13459 D.n2435 D.n2433 0.003
R13460 D.n2455 D.n2453 0.003
R13461 D.n2475 D.n2473 0.003
R13462 D.n2495 D.n2493 0.003
R13463 D.n2515 D.n2513 0.003
R13464 D.n2504 D.n2502 0.003
R13465 D.n2484 D.n2482 0.003
R13466 D.n2464 D.n2462 0.003
R13467 D.n2444 D.n2442 0.003
R13468 D.n2419 D.n2417 0.003
R13469 D.n2402 D.n2401 0.003
R13470 D.n2352 D.n2350 0.003
R13471 D.n2334 D.n2332 0.003
R13472 D.n2316 D.n2314 0.003
R13473 D.n2297 D.n2295 0.003
R13474 D.n2307 D.n2305 0.003
R13475 D.n2325 D.n2323 0.003
R13476 D.n2343 D.n2341 0.003
R13477 D.n2365 D.n2363 0.003
R13478 D.n2378 D.n2377 0.003
R13479 D.n2186 D.n2184 0.003
R13480 D.n2206 D.n2204 0.003
R13481 D.n2226 D.n2224 0.003
R13482 D.n2215 D.n2213 0.003
R13483 D.n2195 D.n2193 0.003
R13484 D.n2172 D.n2170 0.003
R13485 D.n2158 D.n2157 0.003
R13486 D.n2113 D.n2111 0.003
R13487 D.n2094 D.n2092 0.003
R13488 D.n2104 D.n2102 0.003
R13489 D.n2126 D.n2124 0.003
R13490 D.n2139 D.n2138 0.003
R13491 D.n1970 D.n1969 0.003
R13492 D.n55 D.n53 0.003
R13493 D.n64 D.n62 0.003
R13494 D.n73 D.n71 0.003
R13495 D.n82 D.n80 0.003
R13496 D.n91 D.n89 0.003
R13497 D.n100 D.n98 0.003
R13498 D.n109 D.n107 0.003
R13499 D.n118 D.n116 0.003
R13500 D.n127 D.n125 0.003
R13501 D.n136 D.n134 0.003
R13502 D.n145 D.n143 0.003
R13503 D.n154 D.n152 0.003
R13504 D.n163 D.n161 0.003
R13505 D.n172 D.n170 0.003
R13506 D.n181 D.n179 0.003
R13507 D.n190 D.n188 0.003
R13508 D.n199 D.n197 0.003
R13509 D.n208 D.n206 0.003
R13510 D.n217 D.n215 0.003
R13511 D.n287 D.n285 0.003
R13512 D.n303 D.n301 0.003
R13513 D.n274 D.n273 0.003
R13514 D.n555 D.n553 0.003
R13515 D.n541 D.n539 0.003
R13516 D.n527 D.n525 0.003
R13517 D.n513 D.n511 0.003
R13518 D.n499 D.n497 0.003
R13519 D.n485 D.n483 0.003
R13520 D.n471 D.n469 0.003
R13521 D.n457 D.n455 0.003
R13522 D.n443 D.n441 0.003
R13523 D.n429 D.n427 0.003
R13524 D.n415 D.n413 0.003
R13525 D.n401 D.n399 0.003
R13526 D.n387 D.n385 0.003
R13527 D.n373 D.n371 0.003
R13528 D.n359 D.n357 0.003
R13529 D.n345 D.n343 0.003
R13530 D.n331 D.n329 0.003
R13531 D.n317 D.n315 0.003
R13532 D.n578 D.n576 0.003
R13533 D.n594 D.n592 0.003
R13534 D.n568 D.n567 0.003
R13535 D.n818 D.n816 0.003
R13536 D.n804 D.n802 0.003
R13537 D.n790 D.n788 0.003
R13538 D.n776 D.n774 0.003
R13539 D.n762 D.n760 0.003
R13540 D.n748 D.n746 0.003
R13541 D.n734 D.n732 0.003
R13542 D.n720 D.n718 0.003
R13543 D.n706 D.n704 0.003
R13544 D.n692 D.n690 0.003
R13545 D.n678 D.n676 0.003
R13546 D.n664 D.n662 0.003
R13547 D.n650 D.n648 0.003
R13548 D.n636 D.n634 0.003
R13549 D.n622 D.n620 0.003
R13550 D.n608 D.n606 0.003
R13551 D.n841 D.n839 0.003
R13552 D.n857 D.n855 0.003
R13553 D.n831 D.n830 0.003
R13554 D.n1053 D.n1051 0.003
R13555 D.n1039 D.n1037 0.003
R13556 D.n1025 D.n1023 0.003
R13557 D.n1011 D.n1009 0.003
R13558 D.n997 D.n995 0.003
R13559 D.n983 D.n981 0.003
R13560 D.n969 D.n967 0.003
R13561 D.n955 D.n953 0.003
R13562 D.n941 D.n939 0.003
R13563 D.n927 D.n925 0.003
R13564 D.n913 D.n911 0.003
R13565 D.n899 D.n897 0.003
R13566 D.n885 D.n883 0.003
R13567 D.n871 D.n869 0.003
R13568 D.n1076 D.n1074 0.003
R13569 D.n1092 D.n1090 0.003
R13570 D.n1066 D.n1065 0.003
R13571 D.n1260 D.n1258 0.003
R13572 D.n1246 D.n1244 0.003
R13573 D.n1232 D.n1230 0.003
R13574 D.n1218 D.n1216 0.003
R13575 D.n1204 D.n1202 0.003
R13576 D.n1190 D.n1188 0.003
R13577 D.n1176 D.n1174 0.003
R13578 D.n1162 D.n1160 0.003
R13579 D.n1148 D.n1146 0.003
R13580 D.n1134 D.n1132 0.003
R13581 D.n1120 D.n1118 0.003
R13582 D.n1106 D.n1104 0.003
R13583 D.n1283 D.n1281 0.003
R13584 D.n1299 D.n1297 0.003
R13585 D.n1273 D.n1272 0.003
R13586 D.n1439 D.n1437 0.003
R13587 D.n1425 D.n1423 0.003
R13588 D.n1411 D.n1409 0.003
R13589 D.n1397 D.n1395 0.003
R13590 D.n1383 D.n1381 0.003
R13591 D.n1369 D.n1367 0.003
R13592 D.n1355 D.n1353 0.003
R13593 D.n1341 D.n1339 0.003
R13594 D.n1327 D.n1325 0.003
R13595 D.n1313 D.n1311 0.003
R13596 D.n1463 D.n1461 0.003
R13597 D.n1479 D.n1477 0.003
R13598 D.n1453 D.n1452 0.003
R13599 D.n1591 D.n1589 0.003
R13600 D.n1577 D.n1575 0.003
R13601 D.n1563 D.n1561 0.003
R13602 D.n1549 D.n1547 0.003
R13603 D.n1535 D.n1533 0.003
R13604 D.n1521 D.n1519 0.003
R13605 D.n1507 D.n1505 0.003
R13606 D.n1493 D.n1491 0.003
R13607 D.n1615 D.n1613 0.003
R13608 D.n1631 D.n1629 0.003
R13609 D.n1605 D.n1604 0.003
R13610 D.n1715 D.n1713 0.003
R13611 D.n1701 D.n1699 0.003
R13612 D.n1687 D.n1685 0.003
R13613 D.n1673 D.n1671 0.003
R13614 D.n1659 D.n1657 0.003
R13615 D.n1645 D.n1643 0.003
R13616 D.n1739 D.n1737 0.003
R13617 D.n1755 D.n1753 0.003
R13618 D.n1729 D.n1728 0.003
R13619 D.n1811 D.n1809 0.003
R13620 D.n1797 D.n1795 0.003
R13621 D.n1783 D.n1781 0.003
R13622 D.n1769 D.n1767 0.003
R13623 D.n1834 D.n1832 0.003
R13624 D.n1850 D.n1848 0.003
R13625 D.n1824 D.n1823 0.003
R13626 D.n1878 D.n1876 0.003
R13627 D.n1864 D.n1862 0.003
R13628 D.n289 D.n288 0.003
R13629 D.n305 D.n304 0.003
R13630 D.n319 D.n318 0.003
R13631 D.n333 D.n332 0.003
R13632 D.n347 D.n346 0.003
R13633 D.n361 D.n360 0.003
R13634 D.n375 D.n374 0.003
R13635 D.n389 D.n388 0.003
R13636 D.n403 D.n402 0.003
R13637 D.n417 D.n416 0.003
R13638 D.n431 D.n430 0.003
R13639 D.n445 D.n444 0.003
R13640 D.n459 D.n458 0.003
R13641 D.n473 D.n472 0.003
R13642 D.n487 D.n486 0.003
R13643 D.n501 D.n500 0.003
R13644 D.n515 D.n514 0.003
R13645 D.n529 D.n528 0.003
R13646 D.n543 D.n542 0.003
R13647 D.n557 D.n556 0.003
R13648 D.n580 D.n579 0.003
R13649 D.n596 D.n595 0.003
R13650 D.n610 D.n609 0.003
R13651 D.n624 D.n623 0.003
R13652 D.n638 D.n637 0.003
R13653 D.n652 D.n651 0.003
R13654 D.n666 D.n665 0.003
R13655 D.n680 D.n679 0.003
R13656 D.n694 D.n693 0.003
R13657 D.n708 D.n707 0.003
R13658 D.n722 D.n721 0.003
R13659 D.n736 D.n735 0.003
R13660 D.n750 D.n749 0.003
R13661 D.n764 D.n763 0.003
R13662 D.n778 D.n777 0.003
R13663 D.n792 D.n791 0.003
R13664 D.n806 D.n805 0.003
R13665 D.n820 D.n819 0.003
R13666 D.n843 D.n842 0.003
R13667 D.n859 D.n858 0.003
R13668 D.n873 D.n872 0.003
R13669 D.n887 D.n886 0.003
R13670 D.n901 D.n900 0.003
R13671 D.n915 D.n914 0.003
R13672 D.n929 D.n928 0.003
R13673 D.n943 D.n942 0.003
R13674 D.n957 D.n956 0.003
R13675 D.n971 D.n970 0.003
R13676 D.n985 D.n984 0.003
R13677 D.n999 D.n998 0.003
R13678 D.n1013 D.n1012 0.003
R13679 D.n1027 D.n1026 0.003
R13680 D.n1041 D.n1040 0.003
R13681 D.n1055 D.n1054 0.003
R13682 D.n1078 D.n1077 0.003
R13683 D.n1094 D.n1093 0.003
R13684 D.n1108 D.n1107 0.003
R13685 D.n1122 D.n1121 0.003
R13686 D.n1136 D.n1135 0.003
R13687 D.n1150 D.n1149 0.003
R13688 D.n1164 D.n1163 0.003
R13689 D.n1178 D.n1177 0.003
R13690 D.n1192 D.n1191 0.003
R13691 D.n1206 D.n1205 0.003
R13692 D.n1220 D.n1219 0.003
R13693 D.n1234 D.n1233 0.003
R13694 D.n1248 D.n1247 0.003
R13695 D.n1262 D.n1261 0.003
R13696 D.n1285 D.n1284 0.003
R13697 D.n1301 D.n1300 0.003
R13698 D.n1315 D.n1314 0.003
R13699 D.n1329 D.n1328 0.003
R13700 D.n1343 D.n1342 0.003
R13701 D.n1357 D.n1356 0.003
R13702 D.n1371 D.n1370 0.003
R13703 D.n1385 D.n1384 0.003
R13704 D.n1399 D.n1398 0.003
R13705 D.n1413 D.n1412 0.003
R13706 D.n1427 D.n1426 0.003
R13707 D.n1441 D.n1440 0.003
R13708 D.n1465 D.n1464 0.003
R13709 D.n1481 D.n1480 0.003
R13710 D.n1495 D.n1494 0.003
R13711 D.n1509 D.n1508 0.003
R13712 D.n1523 D.n1522 0.003
R13713 D.n1537 D.n1536 0.003
R13714 D.n1551 D.n1550 0.003
R13715 D.n1565 D.n1564 0.003
R13716 D.n1579 D.n1578 0.003
R13717 D.n1593 D.n1592 0.003
R13718 D.n1617 D.n1616 0.003
R13719 D.n1633 D.n1632 0.003
R13720 D.n1647 D.n1646 0.003
R13721 D.n1661 D.n1660 0.003
R13722 D.n1675 D.n1674 0.003
R13723 D.n1689 D.n1688 0.003
R13724 D.n1703 D.n1702 0.003
R13725 D.n1717 D.n1716 0.003
R13726 D.n1741 D.n1740 0.003
R13727 D.n1757 D.n1756 0.003
R13728 D.n1771 D.n1770 0.003
R13729 D.n1785 D.n1784 0.003
R13730 D.n1799 D.n1798 0.003
R13731 D.n1813 D.n1812 0.003
R13732 D.n1836 D.n1835 0.003
R13733 D.n1852 D.n1851 0.003
R13734 D.n1866 D.n1865 0.003
R13735 D.n1882 D.n1880 0.003
R13736 D.n39 D.n38 0.003
R13737 D.n37 D.n36 0.003
R13738 D.n3353 D.n3352 0.003
R13739 D.n2910 D.n2909 0.003
R13740 D.n2547 D.n2546 0.003
R13741 D.n2258 D.n2257 0.003
R13742 D.n2055 D.n2054 0.003
R13743 D.n1904 D.n1896 0.003
R13744 D.n2022 D.n2014 0.003
R13745 D.n1914 D.n1906 0.003
R13746 D.n2012 D.n1999 0.003
R13747 D.n3162 D.n3154 0.003
R13748 D.n3172 D.n3164 0.003
R13749 D.n3182 D.n3174 0.003
R13750 D.n3192 D.n3184 0.003
R13751 D.n3202 D.n3194 0.003
R13752 D.n3212 D.n3204 0.003
R13753 D.n3222 D.n3214 0.003
R13754 D.n3232 D.n3224 0.003
R13755 D.n3242 D.n3234 0.003
R13756 D.n3252 D.n3244 0.003
R13757 D.n3262 D.n3254 0.003
R13758 D.n3272 D.n3264 0.003
R13759 D.n3282 D.n3274 0.003
R13760 D.n3292 D.n3284 0.003
R13761 D.n3302 D.n3294 0.003
R13762 D.n3312 D.n3304 0.003
R13763 D.n3322 D.n3314 0.003
R13764 D.n2759 D.n2751 0.003
R13765 D.n2769 D.n2761 0.003
R13766 D.n2779 D.n2771 0.003
R13767 D.n2789 D.n2781 0.003
R13768 D.n2799 D.n2791 0.003
R13769 D.n2809 D.n2801 0.003
R13770 D.n2819 D.n2811 0.003
R13771 D.n2829 D.n2821 0.003
R13772 D.n2839 D.n2831 0.003
R13773 D.n2849 D.n2841 0.003
R13774 D.n2859 D.n2851 0.003
R13775 D.n2869 D.n2861 0.003
R13776 D.n2879 D.n2871 0.003
R13777 D.n2436 D.n2428 0.003
R13778 D.n2446 D.n2438 0.003
R13779 D.n2456 D.n2448 0.003
R13780 D.n2466 D.n2458 0.003
R13781 D.n2476 D.n2468 0.003
R13782 D.n2486 D.n2478 0.003
R13783 D.n2496 D.n2488 0.003
R13784 D.n2506 D.n2498 0.003
R13785 D.n2516 D.n2508 0.003
R13786 D.n2187 D.n2179 0.003
R13787 D.n2197 D.n2189 0.003
R13788 D.n2207 D.n2199 0.003
R13789 D.n2217 D.n2209 0.003
R13790 D.n2227 D.n2219 0.003
R13791 D.n3152 D.n3141 0.003
R13792 D.n2749 D.n2736 0.003
R13793 D.n2426 D.n2413 0.003
R13794 D.n2177 D.n2166 0.003
R13795 D.n3378 D.n3377 0.002
R13796 D.n21 D.n20 0.002
R13797 D.n19 D.n18 0.002
R13798 D.n2044 D.n2043 0.001
R13799 D.n3365 D.n3364 0.001
R13800 D.n3385 D.n3384 0.001
R13801 D.n3330 D.n3329 0.001
R13802 D.n3342 D.n3341 0.001
R13803 D.n3348 D.n3347 0.001
R13804 D.n2922 D.n2921 0.001
R13805 D.n2938 D.n2937 0.001
R13806 D.n2887 D.n2886 0.001
R13807 D.n2899 D.n2898 0.001
R13808 D.n2905 D.n2904 0.001
R13809 D.n2559 D.n2558 0.001
R13810 D.n2575 D.n2574 0.001
R13811 D.n2524 D.n2523 0.001
R13812 D.n2536 D.n2535 0.001
R13813 D.n2542 D.n2541 0.001
R13814 D.n2270 D.n2269 0.001
R13815 D.n2286 D.n2285 0.001
R13816 D.n2235 D.n2234 0.001
R13817 D.n2247 D.n2246 0.001
R13818 D.n2253 D.n2252 0.001
R13819 D.n2067 D.n2066 0.001
R13820 D.n2083 D.n2082 0.001
R13821 D.n2050 D.n2049 0.001
R13822 D.n2030 D.n2029 0.001
R13823 D.n267 D.n266 0.001
R13824 D.n43 D.n42 0.001
R13825 D.n15 D.n14 0.001
R13826 D.n25 D.n24 0.001
R13827 D.n1922 D.n1921 0.001
R13828 D.n3611 D.n3389 0.001
R13829 D.n3124 D.n2942 0.001
R13830 D.n2715 D.n2579 0.001
R13831 D.n2392 D.n2290 0.001
R13832 D.n2149 D.n2087 0.001
R13833 D.n1981 D.n1962 0.001
R13834 D.n240 D.n237 0.001
R13835 D.n241 D.n228 0.001
R13836 D.n242 D.n219 0.001
R13837 D.n243 D.n210 0.001
R13838 D.n244 D.n201 0.001
R13839 D.n245 D.n192 0.001
R13840 D.n246 D.n183 0.001
R13841 D.n247 D.n174 0.001
R13842 D.n248 D.n165 0.001
R13843 D.n249 D.n156 0.001
R13844 D.n250 D.n147 0.001
R13845 D.n251 D.n138 0.001
R13846 D.n252 D.n129 0.001
R13847 D.n253 D.n120 0.001
R13848 D.n254 D.n111 0.001
R13849 D.n255 D.n102 0.001
R13850 D.n256 D.n93 0.001
R13851 D.n257 D.n84 0.001
R13852 D.n258 D.n75 0.001
R13853 D.n259 D.n66 0.001
R13854 D.n260 D.n57 0.001
R13855 D.n261 D.n47 0.001
R13856 D.n3591 D.n3575 0.001
R13857 D.n3592 D.n3561 0.001
R13858 D.n3593 D.n3552 0.001
R13859 D.n3594 D.n3543 0.001
R13860 D.n3595 D.n3534 0.001
R13861 D.n3596 D.n3525 0.001
R13862 D.n3597 D.n3516 0.001
R13863 D.n3598 D.n3507 0.001
R13864 D.n3599 D.n3498 0.001
R13865 D.n3600 D.n3489 0.001
R13866 D.n3601 D.n3480 0.001
R13867 D.n3602 D.n3471 0.001
R13868 D.n3603 D.n3462 0.001
R13869 D.n3604 D.n3453 0.001
R13870 D.n3605 D.n3444 0.001
R13871 D.n3606 D.n3435 0.001
R13872 D.n3607 D.n3426 0.001
R13873 D.n3608 D.n3417 0.001
R13874 D.n3609 D.n3408 0.001
R13875 D.n3610 D.n3399 0.001
R13876 D.n3108 D.n3091 0.001
R13877 D.n3109 D.n3078 0.001
R13878 D.n3110 D.n3069 0.001
R13879 D.n3111 D.n3060 0.001
R13880 D.n3112 D.n3051 0.001
R13881 D.n3113 D.n3042 0.001
R13882 D.n3114 D.n3033 0.001
R13883 D.n3115 D.n3024 0.001
R13884 D.n3116 D.n3015 0.001
R13885 D.n3117 D.n3006 0.001
R13886 D.n3118 D.n2997 0.001
R13887 D.n3119 D.n2988 0.001
R13888 D.n3120 D.n2979 0.001
R13889 D.n3121 D.n2970 0.001
R13890 D.n3122 D.n2961 0.001
R13891 D.n3123 D.n2952 0.001
R13892 D.n2703 D.n2692 0.001
R13893 D.n2704 D.n2679 0.001
R13894 D.n2705 D.n2670 0.001
R13895 D.n2706 D.n2661 0.001
R13896 D.n2707 D.n2652 0.001
R13897 D.n2708 D.n2643 0.001
R13898 D.n2709 D.n2634 0.001
R13899 D.n2710 D.n2625 0.001
R13900 D.n2711 D.n2616 0.001
R13901 D.n2712 D.n2607 0.001
R13902 D.n2713 D.n2598 0.001
R13903 D.n2714 D.n2589 0.001
R13904 D.n2384 D.n2367 0.001
R13905 D.n2385 D.n2354 0.001
R13906 D.n2386 D.n2345 0.001
R13907 D.n2387 D.n2336 0.001
R13908 D.n2388 D.n2327 0.001
R13909 D.n2389 D.n2318 0.001
R13910 D.n2390 D.n2309 0.001
R13911 D.n2391 D.n2300 0.001
R13912 D.n2145 D.n2128 0.001
R13913 D.n2146 D.n2115 0.001
R13914 D.n2147 D.n2106 0.001
R13915 D.n2148 D.n2097 0.001
R13916 D.n562 D.n561 0.001
R13917 D.n548 D.n547 0.001
R13918 D.n534 D.n533 0.001
R13919 D.n520 D.n519 0.001
R13920 D.n506 D.n505 0.001
R13921 D.n492 D.n491 0.001
R13922 D.n478 D.n477 0.001
R13923 D.n464 D.n463 0.001
R13924 D.n450 D.n449 0.001
R13925 D.n436 D.n435 0.001
R13926 D.n422 D.n421 0.001
R13927 D.n408 D.n407 0.001
R13928 D.n394 D.n393 0.001
R13929 D.n380 D.n379 0.001
R13930 D.n366 D.n365 0.001
R13931 D.n352 D.n351 0.001
R13932 D.n338 D.n337 0.001
R13933 D.n324 D.n323 0.001
R13934 D.n310 D.n309 0.001
R13935 D.n296 D.n295 0.001
R13936 D.n825 D.n824 0.001
R13937 D.n811 D.n810 0.001
R13938 D.n797 D.n796 0.001
R13939 D.n783 D.n782 0.001
R13940 D.n769 D.n768 0.001
R13941 D.n755 D.n754 0.001
R13942 D.n741 D.n740 0.001
R13943 D.n727 D.n726 0.001
R13944 D.n713 D.n712 0.001
R13945 D.n699 D.n698 0.001
R13946 D.n685 D.n684 0.001
R13947 D.n671 D.n670 0.001
R13948 D.n657 D.n656 0.001
R13949 D.n643 D.n642 0.001
R13950 D.n629 D.n628 0.001
R13951 D.n615 D.n614 0.001
R13952 D.n601 D.n600 0.001
R13953 D.n587 D.n586 0.001
R13954 D.n1060 D.n1059 0.001
R13955 D.n1046 D.n1045 0.001
R13956 D.n1032 D.n1031 0.001
R13957 D.n1018 D.n1017 0.001
R13958 D.n1004 D.n1003 0.001
R13959 D.n990 D.n989 0.001
R13960 D.n976 D.n975 0.001
R13961 D.n962 D.n961 0.001
R13962 D.n948 D.n947 0.001
R13963 D.n934 D.n933 0.001
R13964 D.n920 D.n919 0.001
R13965 D.n906 D.n905 0.001
R13966 D.n892 D.n891 0.001
R13967 D.n878 D.n877 0.001
R13968 D.n864 D.n863 0.001
R13969 D.n850 D.n849 0.001
R13970 D.n1267 D.n1266 0.001
R13971 D.n1253 D.n1252 0.001
R13972 D.n1239 D.n1238 0.001
R13973 D.n1225 D.n1224 0.001
R13974 D.n1211 D.n1210 0.001
R13975 D.n1197 D.n1196 0.001
R13976 D.n1183 D.n1182 0.001
R13977 D.n1169 D.n1168 0.001
R13978 D.n1155 D.n1154 0.001
R13979 D.n1141 D.n1140 0.001
R13980 D.n1127 D.n1126 0.001
R13981 D.n1113 D.n1112 0.001
R13982 D.n1099 D.n1098 0.001
R13983 D.n1085 D.n1084 0.001
R13984 D.n1446 D.n1445 0.001
R13985 D.n1432 D.n1431 0.001
R13986 D.n1418 D.n1417 0.001
R13987 D.n1404 D.n1403 0.001
R13988 D.n1390 D.n1389 0.001
R13989 D.n1376 D.n1375 0.001
R13990 D.n1362 D.n1361 0.001
R13991 D.n1348 D.n1347 0.001
R13992 D.n1334 D.n1333 0.001
R13993 D.n1320 D.n1319 0.001
R13994 D.n1306 D.n1305 0.001
R13995 D.n1292 D.n1291 0.001
R13996 D.n1598 D.n1597 0.001
R13997 D.n1584 D.n1583 0.001
R13998 D.n1570 D.n1569 0.001
R13999 D.n1556 D.n1555 0.001
R14000 D.n1542 D.n1541 0.001
R14001 D.n1528 D.n1527 0.001
R14002 D.n1514 D.n1513 0.001
R14003 D.n1500 D.n1499 0.001
R14004 D.n1486 D.n1485 0.001
R14005 D.n1472 D.n1471 0.001
R14006 D.n1722 D.n1721 0.001
R14007 D.n1708 D.n1707 0.001
R14008 D.n1694 D.n1693 0.001
R14009 D.n1680 D.n1679 0.001
R14010 D.n1666 D.n1665 0.001
R14011 D.n1652 D.n1651 0.001
R14012 D.n1638 D.n1637 0.001
R14013 D.n1624 D.n1623 0.001
R14014 D.n1818 D.n1817 0.001
R14015 D.n1804 D.n1803 0.001
R14016 D.n1790 D.n1789 0.001
R14017 D.n1776 D.n1775 0.001
R14018 D.n1762 D.n1761 0.001
R14019 D.n1748 D.n1747 0.001
R14020 D.n1887 D.n1886 0.001
R14021 D.n1871 D.n1870 0.001
R14022 D.n1857 D.n1856 0.001
R14023 D.n1843 D.n1842 0.001
R14024 D.n268 D.n263 0.001
R14025 D.n1928 D.n1926 0.001
R14026 D.n1921 D.n1890 0.001
R14027 D.n1914 D.n1912 0.001
R14028 D.n1904 D.n1902 0.001
R14029 D.n237 D.n235 0.001
R14030 D.n228 D.n226 0.001
R14031 D.n47 D.n33 0.001
R14032 D.n1993 D.n1991 0.001
R14033 D.n2022 D.n2020 0.001
R14034 D.n2012 D.n2005 0.001
R14035 D.n3561 D.n3559 0.001
R14036 D.n3543 D.n3541 0.001
R14037 D.n3525 D.n3523 0.001
R14038 D.n3507 D.n3505 0.001
R14039 D.n3489 D.n3487 0.001
R14040 D.n3471 D.n3469 0.001
R14041 D.n3453 D.n3451 0.001
R14042 D.n3435 D.n3433 0.001
R14043 D.n3417 D.n3415 0.001
R14044 D.n3399 D.n3396 0.001
R14045 D.n3408 D.n3406 0.001
R14046 D.n3426 D.n3424 0.001
R14047 D.n3444 D.n3442 0.001
R14048 D.n3462 D.n3460 0.001
R14049 D.n3480 D.n3478 0.001
R14050 D.n3498 D.n3496 0.001
R14051 D.n3516 D.n3514 0.001
R14052 D.n3534 D.n3532 0.001
R14053 D.n3552 D.n3550 0.001
R14054 D.n3575 D.n3572 0.001
R14055 D.n3590 D.n3585 0.001
R14056 D.n3162 D.n3161 0.001
R14057 D.n3182 D.n3181 0.001
R14058 D.n3202 D.n3201 0.001
R14059 D.n3222 D.n3221 0.001
R14060 D.n3242 D.n3241 0.001
R14061 D.n3262 D.n3261 0.001
R14062 D.n3282 D.n3281 0.001
R14063 D.n3302 D.n3301 0.001
R14064 D.n3322 D.n3321 0.001
R14065 D.n3312 D.n3310 0.001
R14066 D.n3292 D.n3290 0.001
R14067 D.n3272 D.n3270 0.001
R14068 D.n3252 D.n3250 0.001
R14069 D.n3232 D.n3230 0.001
R14070 D.n3212 D.n3210 0.001
R14071 D.n3192 D.n3190 0.001
R14072 D.n3172 D.n3170 0.001
R14073 D.n3152 D.n3147 0.001
R14074 D.n3137 D.n3133 0.001
R14075 D.n3078 D.n3076 0.001
R14076 D.n3060 D.n3058 0.001
R14077 D.n3042 D.n3040 0.001
R14078 D.n3024 D.n3022 0.001
R14079 D.n3006 D.n3004 0.001
R14080 D.n2988 D.n2986 0.001
R14081 D.n2970 D.n2968 0.001
R14082 D.n2952 D.n2949 0.001
R14083 D.n2961 D.n2959 0.001
R14084 D.n2979 D.n2977 0.001
R14085 D.n2997 D.n2995 0.001
R14086 D.n3015 D.n3013 0.001
R14087 D.n3033 D.n3031 0.001
R14088 D.n3051 D.n3049 0.001
R14089 D.n3069 D.n3067 0.001
R14090 D.n3091 D.n3089 0.001
R14091 D.n3107 D.n3102 0.001
R14092 D.n2759 D.n2758 0.001
R14093 D.n2779 D.n2778 0.001
R14094 D.n2799 D.n2798 0.001
R14095 D.n2819 D.n2818 0.001
R14096 D.n2839 D.n2838 0.001
R14097 D.n2859 D.n2858 0.001
R14098 D.n2879 D.n2878 0.001
R14099 D.n2869 D.n2867 0.001
R14100 D.n2849 D.n2847 0.001
R14101 D.n2829 D.n2827 0.001
R14102 D.n2809 D.n2807 0.001
R14103 D.n2789 D.n2787 0.001
R14104 D.n2769 D.n2767 0.001
R14105 D.n2749 D.n2742 0.001
R14106 D.n2730 D.n2725 0.001
R14107 D.n2679 D.n2677 0.001
R14108 D.n2661 D.n2659 0.001
R14109 D.n2643 D.n2641 0.001
R14110 D.n2625 D.n2623 0.001
R14111 D.n2607 D.n2605 0.001
R14112 D.n2589 D.n2586 0.001
R14113 D.n2598 D.n2596 0.001
R14114 D.n2616 D.n2614 0.001
R14115 D.n2634 D.n2632 0.001
R14116 D.n2652 D.n2650 0.001
R14117 D.n2670 D.n2668 0.001
R14118 D.n2692 D.n2689 0.001
R14119 D.n2702 D.n2696 0.001
R14120 D.n2436 D.n2435 0.001
R14121 D.n2456 D.n2455 0.001
R14122 D.n2476 D.n2475 0.001
R14123 D.n2496 D.n2495 0.001
R14124 D.n2516 D.n2515 0.001
R14125 D.n2506 D.n2504 0.001
R14126 D.n2486 D.n2484 0.001
R14127 D.n2466 D.n2464 0.001
R14128 D.n2446 D.n2444 0.001
R14129 D.n2426 D.n2419 0.001
R14130 D.n2407 D.n2402 0.001
R14131 D.n2354 D.n2352 0.001
R14132 D.n2336 D.n2334 0.001
R14133 D.n2318 D.n2316 0.001
R14134 D.n2300 D.n2297 0.001
R14135 D.n2309 D.n2307 0.001
R14136 D.n2327 D.n2325 0.001
R14137 D.n2345 D.n2343 0.001
R14138 D.n2367 D.n2365 0.001
R14139 D.n2383 D.n2378 0.001
R14140 D.n2187 D.n2186 0.001
R14141 D.n2207 D.n2206 0.001
R14142 D.n2227 D.n2226 0.001
R14143 D.n2217 D.n2215 0.001
R14144 D.n2197 D.n2195 0.001
R14145 D.n2177 D.n2172 0.001
R14146 D.n2162 D.n2158 0.001
R14147 D.n2115 D.n2113 0.001
R14148 D.n2097 D.n2094 0.001
R14149 D.n2106 D.n2104 0.001
R14150 D.n2128 D.n2126 0.001
R14151 D.n2144 D.n2139 0.001
R14152 D.n1977 D.n1970 0.001
R14153 D.n57 D.n55 0.001
R14154 D.n66 D.n64 0.001
R14155 D.n75 D.n73 0.001
R14156 D.n84 D.n82 0.001
R14157 D.n93 D.n91 0.001
R14158 D.n102 D.n100 0.001
R14159 D.n111 D.n109 0.001
R14160 D.n120 D.n118 0.001
R14161 D.n129 D.n127 0.001
R14162 D.n138 D.n136 0.001
R14163 D.n147 D.n145 0.001
R14164 D.n156 D.n154 0.001
R14165 D.n165 D.n163 0.001
R14166 D.n174 D.n172 0.001
R14167 D.n183 D.n181 0.001
R14168 D.n192 D.n190 0.001
R14169 D.n201 D.n199 0.001
R14170 D.n210 D.n208 0.001
R14171 D.n219 D.n217 0.001
R14172 D.n295 D.n287 0.001
R14173 D.n309 D.n303 0.001
R14174 D.n565 D.n274 0.001
R14175 D.n561 D.n555 0.001
R14176 D.n547 D.n541 0.001
R14177 D.n533 D.n527 0.001
R14178 D.n519 D.n513 0.001
R14179 D.n505 D.n499 0.001
R14180 D.n491 D.n485 0.001
R14181 D.n477 D.n471 0.001
R14182 D.n463 D.n457 0.001
R14183 D.n449 D.n443 0.001
R14184 D.n435 D.n429 0.001
R14185 D.n421 D.n415 0.001
R14186 D.n407 D.n401 0.001
R14187 D.n393 D.n387 0.001
R14188 D.n379 D.n373 0.001
R14189 D.n365 D.n359 0.001
R14190 D.n351 D.n345 0.001
R14191 D.n337 D.n331 0.001
R14192 D.n323 D.n317 0.001
R14193 D.n586 D.n578 0.001
R14194 D.n600 D.n594 0.001
R14195 D.n828 D.n568 0.001
R14196 D.n824 D.n818 0.001
R14197 D.n810 D.n804 0.001
R14198 D.n796 D.n790 0.001
R14199 D.n782 D.n776 0.001
R14200 D.n768 D.n762 0.001
R14201 D.n754 D.n748 0.001
R14202 D.n740 D.n734 0.001
R14203 D.n726 D.n720 0.001
R14204 D.n712 D.n706 0.001
R14205 D.n698 D.n692 0.001
R14206 D.n684 D.n678 0.001
R14207 D.n670 D.n664 0.001
R14208 D.n656 D.n650 0.001
R14209 D.n642 D.n636 0.001
R14210 D.n628 D.n622 0.001
R14211 D.n614 D.n608 0.001
R14212 D.n849 D.n841 0.001
R14213 D.n863 D.n857 0.001
R14214 D.n1063 D.n831 0.001
R14215 D.n1059 D.n1053 0.001
R14216 D.n1045 D.n1039 0.001
R14217 D.n1031 D.n1025 0.001
R14218 D.n1017 D.n1011 0.001
R14219 D.n1003 D.n997 0.001
R14220 D.n989 D.n983 0.001
R14221 D.n975 D.n969 0.001
R14222 D.n961 D.n955 0.001
R14223 D.n947 D.n941 0.001
R14224 D.n933 D.n927 0.001
R14225 D.n919 D.n913 0.001
R14226 D.n905 D.n899 0.001
R14227 D.n891 D.n885 0.001
R14228 D.n877 D.n871 0.001
R14229 D.n1084 D.n1076 0.001
R14230 D.n1098 D.n1092 0.001
R14231 D.n1270 D.n1066 0.001
R14232 D.n1266 D.n1260 0.001
R14233 D.n1252 D.n1246 0.001
R14234 D.n1238 D.n1232 0.001
R14235 D.n1224 D.n1218 0.001
R14236 D.n1210 D.n1204 0.001
R14237 D.n1196 D.n1190 0.001
R14238 D.n1182 D.n1176 0.001
R14239 D.n1168 D.n1162 0.001
R14240 D.n1154 D.n1148 0.001
R14241 D.n1140 D.n1134 0.001
R14242 D.n1126 D.n1120 0.001
R14243 D.n1112 D.n1106 0.001
R14244 D.n1291 D.n1283 0.001
R14245 D.n1305 D.n1299 0.001
R14246 D.n1449 D.n1273 0.001
R14247 D.n1445 D.n1439 0.001
R14248 D.n1431 D.n1425 0.001
R14249 D.n1417 D.n1411 0.001
R14250 D.n1403 D.n1397 0.001
R14251 D.n1389 D.n1383 0.001
R14252 D.n1375 D.n1369 0.001
R14253 D.n1361 D.n1355 0.001
R14254 D.n1347 D.n1341 0.001
R14255 D.n1333 D.n1327 0.001
R14256 D.n1319 D.n1313 0.001
R14257 D.n1471 D.n1463 0.001
R14258 D.n1485 D.n1479 0.001
R14259 D.n1601 D.n1453 0.001
R14260 D.n1597 D.n1591 0.001
R14261 D.n1583 D.n1577 0.001
R14262 D.n1569 D.n1563 0.001
R14263 D.n1555 D.n1549 0.001
R14264 D.n1541 D.n1535 0.001
R14265 D.n1527 D.n1521 0.001
R14266 D.n1513 D.n1507 0.001
R14267 D.n1499 D.n1493 0.001
R14268 D.n1623 D.n1615 0.001
R14269 D.n1637 D.n1631 0.001
R14270 D.n1725 D.n1605 0.001
R14271 D.n1721 D.n1715 0.001
R14272 D.n1707 D.n1701 0.001
R14273 D.n1693 D.n1687 0.001
R14274 D.n1679 D.n1673 0.001
R14275 D.n1665 D.n1659 0.001
R14276 D.n1651 D.n1645 0.001
R14277 D.n1747 D.n1739 0.001
R14278 D.n1761 D.n1755 0.001
R14279 D.n1821 D.n1729 0.001
R14280 D.n1817 D.n1811 0.001
R14281 D.n1803 D.n1797 0.001
R14282 D.n1789 D.n1783 0.001
R14283 D.n1775 D.n1769 0.001
R14284 D.n1842 D.n1834 0.001
R14285 D.n1856 D.n1850 0.001
R14286 D.n1888 D.n1824 0.001
R14287 D.n1886 D.n1878 0.001
R14288 D.n1870 D.n1864 0.001
R14289 D.n1914 D.n1909 0.001
R14290 D.n1904 D.n1899 0.001
R14291 D.n237 D.n232 0.001
R14292 D.n228 D.n223 0.001
R14293 D.n47 D.n30 0.001
R14294 D.n2022 D.n2017 0.001
R14295 D.n2012 D.n2002 0.001
R14296 D.n3561 D.n3556 0.001
R14297 D.n3543 D.n3538 0.001
R14298 D.n3525 D.n3520 0.001
R14299 D.n3507 D.n3502 0.001
R14300 D.n3489 D.n3484 0.001
R14301 D.n3471 D.n3466 0.001
R14302 D.n3453 D.n3448 0.001
R14303 D.n3435 D.n3430 0.001
R14304 D.n3417 D.n3412 0.001
R14305 D.n3399 D.n3393 0.001
R14306 D.n3408 D.n3403 0.001
R14307 D.n3426 D.n3421 0.001
R14308 D.n3444 D.n3439 0.001
R14309 D.n3462 D.n3457 0.001
R14310 D.n3480 D.n3475 0.001
R14311 D.n3498 D.n3493 0.001
R14312 D.n3516 D.n3511 0.001
R14313 D.n3534 D.n3529 0.001
R14314 D.n3552 D.n3547 0.001
R14315 D.n3575 D.n3569 0.001
R14316 D.n3162 D.n3158 0.001
R14317 D.n3182 D.n3178 0.001
R14318 D.n3202 D.n3198 0.001
R14319 D.n3222 D.n3218 0.001
R14320 D.n3242 D.n3238 0.001
R14321 D.n3262 D.n3258 0.001
R14322 D.n3282 D.n3278 0.001
R14323 D.n3302 D.n3298 0.001
R14324 D.n3322 D.n3318 0.001
R14325 D.n3312 D.n3307 0.001
R14326 D.n3292 D.n3287 0.001
R14327 D.n3272 D.n3267 0.001
R14328 D.n3252 D.n3247 0.001
R14329 D.n3232 D.n3227 0.001
R14330 D.n3212 D.n3207 0.001
R14331 D.n3192 D.n3187 0.001
R14332 D.n3172 D.n3167 0.001
R14333 D.n3152 D.n3144 0.001
R14334 D.n3078 D.n3073 0.001
R14335 D.n3060 D.n3055 0.001
R14336 D.n3042 D.n3037 0.001
R14337 D.n3024 D.n3019 0.001
R14338 D.n3006 D.n3001 0.001
R14339 D.n2988 D.n2983 0.001
R14340 D.n2970 D.n2965 0.001
R14341 D.n2952 D.n2946 0.001
R14342 D.n2961 D.n2956 0.001
R14343 D.n2979 D.n2974 0.001
R14344 D.n2997 D.n2992 0.001
R14345 D.n3015 D.n3010 0.001
R14346 D.n3033 D.n3028 0.001
R14347 D.n3051 D.n3046 0.001
R14348 D.n3069 D.n3064 0.001
R14349 D.n3091 D.n3086 0.001
R14350 D.n2759 D.n2755 0.001
R14351 D.n2779 D.n2775 0.001
R14352 D.n2799 D.n2795 0.001
R14353 D.n2819 D.n2815 0.001
R14354 D.n2839 D.n2835 0.001
R14355 D.n2859 D.n2855 0.001
R14356 D.n2879 D.n2875 0.001
R14357 D.n2869 D.n2864 0.001
R14358 D.n2849 D.n2844 0.001
R14359 D.n2829 D.n2824 0.001
R14360 D.n2809 D.n2804 0.001
R14361 D.n2789 D.n2784 0.001
R14362 D.n2769 D.n2764 0.001
R14363 D.n2749 D.n2739 0.001
R14364 D.n2679 D.n2674 0.001
R14365 D.n2661 D.n2656 0.001
R14366 D.n2643 D.n2638 0.001
R14367 D.n2625 D.n2620 0.001
R14368 D.n2607 D.n2602 0.001
R14369 D.n2589 D.n2583 0.001
R14370 D.n2598 D.n2593 0.001
R14371 D.n2616 D.n2611 0.001
R14372 D.n2634 D.n2629 0.001
R14373 D.n2652 D.n2647 0.001
R14374 D.n2670 D.n2665 0.001
R14375 D.n2692 D.n2686 0.001
R14376 D.n2436 D.n2432 0.001
R14377 D.n2456 D.n2452 0.001
R14378 D.n2476 D.n2472 0.001
R14379 D.n2496 D.n2492 0.001
R14380 D.n2516 D.n2512 0.001
R14381 D.n2506 D.n2501 0.001
R14382 D.n2486 D.n2481 0.001
R14383 D.n2466 D.n2461 0.001
R14384 D.n2446 D.n2441 0.001
R14385 D.n2426 D.n2416 0.001
R14386 D.n2354 D.n2349 0.001
R14387 D.n2336 D.n2331 0.001
R14388 D.n2318 D.n2313 0.001
R14389 D.n2300 D.n2294 0.001
R14390 D.n2309 D.n2304 0.001
R14391 D.n2327 D.n2322 0.001
R14392 D.n2345 D.n2340 0.001
R14393 D.n2367 D.n2362 0.001
R14394 D.n2187 D.n2183 0.001
R14395 D.n2207 D.n2203 0.001
R14396 D.n2227 D.n2223 0.001
R14397 D.n2217 D.n2212 0.001
R14398 D.n2197 D.n2192 0.001
R14399 D.n2177 D.n2169 0.001
R14400 D.n2115 D.n2110 0.001
R14401 D.n2097 D.n2091 0.001
R14402 D.n2106 D.n2101 0.001
R14403 D.n2128 D.n2123 0.001
R14404 D.n57 D.n52 0.001
R14405 D.n66 D.n61 0.001
R14406 D.n75 D.n70 0.001
R14407 D.n84 D.n79 0.001
R14408 D.n93 D.n88 0.001
R14409 D.n102 D.n97 0.001
R14410 D.n111 D.n106 0.001
R14411 D.n120 D.n115 0.001
R14412 D.n129 D.n124 0.001
R14413 D.n138 D.n133 0.001
R14414 D.n147 D.n142 0.001
R14415 D.n156 D.n151 0.001
R14416 D.n165 D.n160 0.001
R14417 D.n174 D.n169 0.001
R14418 D.n183 D.n178 0.001
R14419 D.n192 D.n187 0.001
R14420 D.n201 D.n196 0.001
R14421 D.n210 D.n205 0.001
R14422 D.n219 D.n214 0.001
R14423 D.n295 D.n284 0.001
R14424 D.n309 D.n300 0.001
R14425 D.n561 D.n552 0.001
R14426 D.n547 D.n538 0.001
R14427 D.n533 D.n524 0.001
R14428 D.n519 D.n510 0.001
R14429 D.n505 D.n496 0.001
R14430 D.n491 D.n482 0.001
R14431 D.n477 D.n468 0.001
R14432 D.n463 D.n454 0.001
R14433 D.n449 D.n440 0.001
R14434 D.n435 D.n426 0.001
R14435 D.n421 D.n412 0.001
R14436 D.n407 D.n398 0.001
R14437 D.n393 D.n384 0.001
R14438 D.n379 D.n370 0.001
R14439 D.n365 D.n356 0.001
R14440 D.n351 D.n342 0.001
R14441 D.n337 D.n328 0.001
R14442 D.n323 D.n314 0.001
R14443 D.n586 D.n575 0.001
R14444 D.n600 D.n591 0.001
R14445 D.n824 D.n815 0.001
R14446 D.n810 D.n801 0.001
R14447 D.n796 D.n787 0.001
R14448 D.n782 D.n773 0.001
R14449 D.n768 D.n759 0.001
R14450 D.n754 D.n745 0.001
R14451 D.n740 D.n731 0.001
R14452 D.n726 D.n717 0.001
R14453 D.n712 D.n703 0.001
R14454 D.n698 D.n689 0.001
R14455 D.n684 D.n675 0.001
R14456 D.n670 D.n661 0.001
R14457 D.n656 D.n647 0.001
R14458 D.n642 D.n633 0.001
R14459 D.n628 D.n619 0.001
R14460 D.n614 D.n605 0.001
R14461 D.n849 D.n838 0.001
R14462 D.n863 D.n854 0.001
R14463 D.n1059 D.n1050 0.001
R14464 D.n1045 D.n1036 0.001
R14465 D.n1031 D.n1022 0.001
R14466 D.n1017 D.n1008 0.001
R14467 D.n1003 D.n994 0.001
R14468 D.n989 D.n980 0.001
R14469 D.n975 D.n966 0.001
R14470 D.n961 D.n952 0.001
R14471 D.n947 D.n938 0.001
R14472 D.n933 D.n924 0.001
R14473 D.n919 D.n910 0.001
R14474 D.n905 D.n896 0.001
R14475 D.n891 D.n882 0.001
R14476 D.n877 D.n868 0.001
R14477 D.n1084 D.n1073 0.001
R14478 D.n1098 D.n1089 0.001
R14479 D.n1266 D.n1257 0.001
R14480 D.n1252 D.n1243 0.001
R14481 D.n1238 D.n1229 0.001
R14482 D.n1224 D.n1215 0.001
R14483 D.n1210 D.n1201 0.001
R14484 D.n1196 D.n1187 0.001
R14485 D.n1182 D.n1173 0.001
R14486 D.n1168 D.n1159 0.001
R14487 D.n1154 D.n1145 0.001
R14488 D.n1140 D.n1131 0.001
R14489 D.n1126 D.n1117 0.001
R14490 D.n1112 D.n1103 0.001
R14491 D.n1291 D.n1280 0.001
R14492 D.n1305 D.n1296 0.001
R14493 D.n1445 D.n1436 0.001
R14494 D.n1431 D.n1422 0.001
R14495 D.n1417 D.n1408 0.001
R14496 D.n1403 D.n1394 0.001
R14497 D.n1389 D.n1380 0.001
R14498 D.n1375 D.n1366 0.001
R14499 D.n1361 D.n1352 0.001
R14500 D.n1347 D.n1338 0.001
R14501 D.n1333 D.n1324 0.001
R14502 D.n1319 D.n1310 0.001
R14503 D.n1471 D.n1460 0.001
R14504 D.n1485 D.n1476 0.001
R14505 D.n1597 D.n1588 0.001
R14506 D.n1583 D.n1574 0.001
R14507 D.n1569 D.n1560 0.001
R14508 D.n1555 D.n1546 0.001
R14509 D.n1541 D.n1532 0.001
R14510 D.n1527 D.n1518 0.001
R14511 D.n1513 D.n1504 0.001
R14512 D.n1499 D.n1490 0.001
R14513 D.n1623 D.n1612 0.001
R14514 D.n1637 D.n1628 0.001
R14515 D.n1721 D.n1712 0.001
R14516 D.n1707 D.n1698 0.001
R14517 D.n1693 D.n1684 0.001
R14518 D.n1679 D.n1670 0.001
R14519 D.n1665 D.n1656 0.001
R14520 D.n1651 D.n1642 0.001
R14521 D.n1747 D.n1736 0.001
R14522 D.n1761 D.n1752 0.001
R14523 D.n1817 D.n1808 0.001
R14524 D.n1803 D.n1794 0.001
R14525 D.n1789 D.n1780 0.001
R14526 D.n1775 D.n1766 0.001
R14527 D.n1842 D.n1831 0.001
R14528 D.n1856 D.n1847 0.001
R14529 D.n1886 D.n1875 0.001
R14530 D.n1870 D.n1861 0.001
R14531 D.n1962 D.n1953 0.001
R14532 D.n2048 D.n2037 0.001
R14533 D.n3389 D.n3370 0.001
R14534 D.n3346 D.n3335 0.001
R14535 D.n2942 D.n2927 0.001
R14536 D.n2903 D.n2892 0.001
R14537 D.n2579 D.n2564 0.001
R14538 D.n2540 D.n2529 0.001
R14539 D.n2290 D.n2275 0.001
R14540 D.n2251 D.n2240 0.001
R14541 D.n2087 D.n2072 0.001
R14542 D.n239 D.n238 0.001
R14543 D.n1895 D.n1893 0.001
R14544 D.n293 D.n291 0.001
R14545 D.n584 D.n582 0.001
R14546 D.n847 D.n845 0.001
R14547 D.n1082 D.n1080 0.001
R14548 D.n1289 D.n1287 0.001
R14549 D.n1469 D.n1467 0.001
R14550 D.n1621 D.n1619 0.001
R14551 D.n1745 D.n1743 0.001
R14552 D.n1840 D.n1838 0.001
R14553 D.n1932 D.n1930 0.001
R14554 D.n1933 D.n1928 0.001
R14555 PW PW.n0 1.963
C0 S G 1404.81fF
C1 S D 2210.82fF
C2 G D 1015.86fF
.ends

