* NGSPICE file created from mag_files/POSTLAYOUT/pmos_flat_6x6.ext - technology: sky130A

.subckt pmos_flat_6x6 G S D PW
X0 S.t70 G D S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X1 D G S.t69 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2 S.t68 G D S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X3 D G S.t67 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4 D G S.t66 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X5 S.t65 G D S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X6 S.t64 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7 D.t6 G S.t63 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X8 S.t62 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X9 S.t61 G D S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X10 D G S.t60 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X11 S.t59 G D S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X12 S.t58 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X13 S.t57 G D.t1 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14 S.t56 G D S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X15 D G S.t55 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X16 D G S.t54 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X17 D.t1 G S.t53 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X18 S.t52 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X19 S.t51 G D.t1 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X20 S.t50 G D.t7 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X21 S.t49 G D S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.3312 ps=9.38 w=4.38 l=0.5
X22 D G S.t48 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X23 D.t1 G S.t47 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X24 D G S.t46 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X25 S.t45 G D.t5 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X26 D G S.t44 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X27 S.t43 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X28 D.t3 G S.t42 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X29 S.t41 G D S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X30 S.t40 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X31 D G S.t39 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X32 D G S.t38 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X33 D G S.t37 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X34 D G S.t36 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X35 D.t0 G S.t35 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X36 S.t34 G D.t6 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X37 D G S.t33 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X38 S.t32 G D.t1 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X39 S.t30 G D S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X40 D G S.t28 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X41 S.t27 G D S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X42 D G S.t26 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X43 S.t25 G D S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X44 D.t2 G S.t24 S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X45 S.t23 G D S.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X46 D.t4 G S.t21 S.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X47 S.t19 G D S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X48 D G S.t18 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=1.3312 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X49 S.t17 G D S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X50 D G S.t15 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X51 D G S.t13 S.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X52 S.t11 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X53 D G S.t10 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X54 S.t9 G D S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X55 D.t1 G S.t8 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X56 D G S.t7 S.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X57 S.t5 G D S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X58 D G S.t3 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X59 S.t1 G D S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
R0 D.t1 D.t5 7.599
R1 D.t1 D.t2 7.099
R2 D.n0 D.t7 7.065
R3 D.n0 D.t3 7.007
R4 D.n0 D.t4 6.564
R5 D.t6 D.t0 6.524
R6 D.t6 D.t1 0.343
R7 D.t1 D.n0 0.293
R8 D D.t6 0.182
R9 S.n81 S.n80 153.554
R10 S.n220 S.n219 153.554
R11 S.n289 S.n288 153.118
R12 S.n135 S.n134 153.118
R13 S.n188 S.n187 146.135
R14 S.n169 S.n168 146.135
R15 S.n323 S.n322 145.699
R16 S.n319 S.n318 145.699
R17 S.n73 S.n72 101.08
R18 S.n228 S.n227 101.08
R19 S.n118 S.n117 98.123
R20 S.n339 S.n338 88.439
R21 S.n304 S.n303 68.042
R22 S.n230 S.n229 65.312
R23 S.n296 S.n295 62.872
R24 S.n120 S.n119 62.872
R25 S.t20 S.t31 58.055
R26 S.n125 S.t6 50.666
R27 S.n74 S.t0 50.666
R28 S.n301 S.t2 50.666
R29 S.n231 S.t12 50.666
R30 S.t22 S.n136 48.977
R31 S.t29 S.n100 48.977
R32 S.t4 S.n258 48.977
R33 S.t14 S.n216 48.977
R34 S.t16 S.n316 48.977
R35 S.n340 S.n339 10.138
R36 S.n215 S.n214 6.541
R37 S.n199 S.t15 6.541
R38 S.n210 S.n209 6.541
R39 S.n201 S.t37 6.541
R40 S.n325 S.t60 6.541
R41 S.n323 S.t13 6.541
R42 S.n289 S.t55 6.541
R43 S.n286 S.t10 6.541
R44 S.n321 S.t46 6.541
R45 S.n308 S.t36 6.541
R46 S.n135 S.t66 6.541
R47 S.n2 S.n67 6.541
R48 S.n102 S.t54 6.541
R49 S.n104 S.t28 6.541
R50 S.n106 S.n105 6.541
R51 S.n186 S.t67 6.541
R52 S.n3 S.n36 6.541
R53 S.n138 S.t48 6.541
R54 S.n140 S.t38 6.541
R55 S.n142 S.n141 6.541
R56 S.n82 S.t7 6.541
R57 S.n4 S.n44 6.541
R58 S.n60 S.t24 6.541
R59 S.n58 S.t42 6.541
R60 S.n46 S.n45 6.541
R61 S.n167 S.t21 6.541
R62 S.n217 S.t35 6.541
R63 S.n5 S.n271 6.541
R64 S.n283 S.t63 6.541
R65 S.n285 S.t8 6.541
R66 S.n269 S.n268 6.541
R67 S.n6 S.n90 6.541
R68 S.n99 S.t47 6.541
R69 S.n97 S.t53 6.541
R70 S.n88 S.n87 6.541
R71 S.n7 S.n248 6.541
R72 S.n257 S.t44 6.541
R73 S.n194 S.t69 6.541
R74 S.n250 S.n249 6.541
R75 S.n8 S.n197 6.541
R76 S.n240 S.t26 6.541
R77 S.n242 S.t3 6.541
R78 S.n244 S.n243 6.541
R79 S.n319 S.t33 6.541
R80 S.n317 S.t18 6.541
R81 S.n133 S.t39 6.541
R82 S.t20 S.t52 6.158
R83 S.t20 S.t70 6.109
R84 S.n215 S.t59 6.105
R85 S.n199 S.n198 6.105
R86 S.n210 S.t19 6.105
R87 S.n201 S.n200 6.105
R88 S.n324 S.t61 6.105
R89 S.n192 S.t11 6.105
R90 S.n2 S.t40 6.105
R91 S.n102 S.n101 6.105
R92 S.n104 S.n103 6.105
R93 S.n106 S.t64 6.105
R94 S.n188 S.t32 6.105
R95 S.n189 S.t50 6.105
R96 S.n3 S.t45 6.105
R97 S.n138 S.n137 6.105
R98 S.n140 S.n139 6.105
R99 S.n142 S.t57 6.105
R100 S.n81 S.t51 6.105
R101 S.n68 S.t34 6.105
R102 S.n4 S.t23 6.105
R103 S.n60 S.n59 6.105
R104 S.n58 S.n57 6.105
R105 S.n46 S.t56 6.105
R106 S.n169 S.t41 6.105
R107 S.n170 S.t68 6.105
R108 S.n220 S.t27 6.105
R109 S.n221 S.t49 6.105
R110 S.n5 S.t62 6.105
R111 S.n283 S.n282 6.105
R112 S.n285 S.n284 6.105
R113 S.n269 S.t9 6.105
R114 S.n6 S.t30 6.105
R115 S.n99 S.n98 6.105
R116 S.n97 S.n96 6.105
R117 S.n88 S.t1 6.105
R118 S.n7 S.t5 6.105
R119 S.n257 S.n256 6.105
R120 S.n194 S.n193 6.105
R121 S.n250 S.t43 6.105
R122 S.n8 S.t65 6.105
R123 S.n240 S.n239 6.105
R124 S.n242 S.n241 6.105
R125 S.n244 S.t25 6.105
R126 S.n320 S.t17 6.105
R127 S.n131 S.t58 6.105
R128 S.n231 S.n230 4.263
R129 S.n121 S.n120 3.857
R130 S.n297 S.n296 3.857
R131 S.n27 S.n343 0.178
R132 S.n348 S.n347 0.143
R133 S.n26 S.n118 0.136
R134 S.n123 S.n122 0.117
R135 S.n299 S.n298 0.117
R136 S.n348 S.n307 0.114
R137 S.n1 S.n331 0.111
R138 S.n255 S.n253 0.109
R139 S.n25 S.n304 0.103
R140 S.n191 S.n190 0.099
R141 S.n312 S.n309 0.093
R142 S.n226 S.n224 0.093
R143 S S.n349 0.09
R144 S.n50 S.n48 0.087
R145 S.n311 S.n310 0.085
R146 S.n180 S.n9 0.082
R147 S.n26 S.n126 0.082
R148 S.n25 S.n302 0.082
R149 S.n346 S.n345 0.079
R150 S.n12 S.n144 0.077
R151 S.n166 S.n162 0.075
R152 S.n14 S.n112 0.074
R153 S.n236 S.n10 0.074
R154 S.n77 S.n11 0.074
R155 S.n335 S.n329 0.127
R156 S.n328 S.n327 0.071
R157 S.t16 S.n313 0.068
R158 S.n154 S.n152 0.067
R159 S.n154 S.n153 0.067
R160 S.n180 S.n178 0.067
R161 S.n180 S.n179 0.067
R162 S.n26 S.n116 0.067
R163 S.n26 S.n114 0.067
R164 S.n30 S.n29 0.066
R165 S.n181 S.n180 0.063
R166 S.n16 S.n95 0.063
R167 S.n13 S.n38 0.063
R168 S.n181 S.n174 0.062
R169 S.n148 S.n147 0.06
R170 S.n31 S.n30 0.059
R171 S.n280 S.n279 0.059
R172 S.n14 S.n133 0.055
R173 S.n290 S.n192 0.054
R174 S.n79 S.n68 0.054
R175 S.n238 S.n221 0.054
R176 S.n346 S.n27 0.054
R177 S.n22 S.n104 0.054
R178 S.n24 S.n140 0.054
R179 S.n13 S.n58 0.054
R180 S.n19 S.n285 0.054
R181 S.n16 S.n97 0.054
R182 S.t4 S.n194 0.054
R183 S.n21 S.n242 0.054
R184 S.n336 S.n308 0.053
R185 S.n305 S.n25 0.052
R186 S.n10 S.n234 0.052
R187 S.n11 S.n76 0.052
R188 S.n129 S.n128 0.052
R189 S.n116 S.n115 0.051
R190 S.n114 S.n113 0.051
R191 S.n262 S.n261 0.05
R192 S.n18 S.n281 0.05
R193 S.t22 S.n35 0.05
R194 S.n41 S.n40 0.05
R195 S.n28 S.n211 0.05
R196 S.n127 S.n26 0.049
R197 S.n155 S.n154 0.048
R198 S.n23 S.n107 0.047
R199 S.t22 S.n143 0.047
R200 S.n13 S.n47 0.047
R201 S.n18 S.n270 0.047
R202 S.n16 S.n89 0.047
R203 S.n17 S.n251 0.047
R204 S.t14 S.n245 0.047
R205 S.n14 S.n132 0.047
R206 S.n17 S.t14 0.046
R207 S.n157 S.n155 0.045
R208 S.n190 S.n146 0.044
R209 S.n281 S.n278 0.043
R210 S.n35 S.n34 0.043
R211 S.n92 S.n91 0.042
R212 S.n335 S.n326 0.041
R213 S.n76 S.n71 0.039
R214 S.n234 S.n233 0.039
R215 S.n329 S.n328 0.039
R216 S.n166 S.n165 0.038
R217 S.n226 S.n225 0.038
R218 S.n165 S.n164 0.038
R219 S.n56 S.n51 0.036
R220 S.n287 S.n286 0.035
R221 S.n83 S.n82 0.035
R222 S.n218 S.n217 0.035
R223 S.t20 S.n151 0.035
R224 S.t16 S.n325 0.035
R225 S.t20 S.n186 0.035
R226 S.t20 S.n167 0.035
R227 S.t16 S.n317 0.035
R228 S.n184 S.n183 0.035
R229 S.n315 S.n314 0.035
R230 S.n14 S.n130 0.034
R231 S.t16 S.n324 0.034
R232 S.t20 S.n189 0.034
R233 S.t20 S.n170 0.034
R234 S.t16 S.n320 0.034
R235 S.n62 S.n61 0.034
R236 S.n124 S.n121 0.033
R237 S.n75 S.n73 0.033
R238 S.n300 S.n297 0.033
R239 S.n232 S.n228 0.033
R240 S.n342 S.n340 0.033
R241 S.n185 S.n184 0.033
R242 S.n208 S.n207 0.033
R243 S.n236 S.n226 0.032
R244 S.n77 S.n69 0.032
R245 S.t4 S.n287 0.031
R246 S.t29 S.n83 0.031
R247 S.t14 S.n218 0.031
R248 S.n212 S.n203 0.031
R249 S.n349 S.n348 0.031
R250 S.n203 S.n202 0.031
R251 S.n265 S.n264 0.031
R252 S.n161 S.n160 0.029
R253 S.n54 S.n53 0.028
R254 S.n275 S.n274 0.028
R255 S.n264 S.n263 0.027
R256 S.n14 S.n63 0.027
R257 S.n255 S.n254 0.026
R258 S.n18 S.n276 0.026
R259 S.n16 S.n93 0.026
R260 S.n306 S.n292 0.026
R261 S.n27 S.n344 0.025
R262 S.n292 S.n291 0.024
R263 S.n63 S.n62 0.024
R264 S.n129 S.n127 0.023
R265 S.n51 S.n50 0.023
R266 S.n109 S.n108 0.023
R267 S.n164 S.n163 0.023
R268 S.n294 S.n293 0.023
R269 S.n65 S.n64 0.023
R270 S.n157 S.n156 0.022
R271 S.n151 S.n150 0.022
R272 S.n50 S.n49 0.022
R273 S.t14 S.n195 0.022
R274 S.n278 S.n277 0.022
R275 S.n34 S.n33 0.022
R276 S.n275 S.n273 0.021
R277 S.n40 S.n39 0.021
R278 S.n38 S.n37 0.021
R279 S.n312 S.n311 0.021
R280 S.n174 S.n173 0.021
R281 S.n281 S.n280 0.02
R282 S.n35 S.n31 0.02
R283 S.t20 S.n157 0.019
R284 S.n28 S.n208 0.019
R285 S S.n191 0.018
R286 S.n33 S.n32 0.018
R287 S.n16 S.n86 0.016
R288 S.n18 S.n267 0.016
R289 S.t20 S.n161 0.016
R290 S.n16 S.n85 0.015
R291 S.n173 S.n172 0.015
R292 S.n273 S.n272 0.015
R293 S.t16 S.n315 0.015
R294 S.n13 S.n42 0.012
R295 S.n56 S.n55 0.012
R296 S.n12 S.n145 0.011
R297 S.n13 S.n56 0.011
R298 S.n17 S.n252 0.01
R299 S.n306 S.n294 0.01
R300 S.n14 S.n65 0.01
R301 S.n14 S.n129 0.01
R302 S.n306 S.n305 0.01
R303 S.n237 S.n223 0.01
R304 S.t16 S.n312 0.009
R305 S.n17 S.n255 0.008
R306 S.n111 S.n109 0.008
R307 S.n266 S.n262 0.008
R308 S.n95 S.n94 0.008
R309 S.t20 S.n166 0.008
R310 S.n53 S.n52 0.008
R311 S.n184 S.n182 0.007
R312 S.n347 S.n337 0.007
R313 S.t20 S.n149 0.119
R314 S.n11 S.n70 0.041
R315 S.n10 S.n235 0.041
R316 S.n261 S.n260 0.005
R317 S.t20 S.n158 0.005
R318 S.n28 S.n206 0.005
R319 S.t20 S.n148 0.005
R320 S.t20 S.n185 0.005
R321 S.n211 S.n210 0.004
R322 S.n107 S.n106 0.004
R323 S.n143 S.n142 0.004
R324 S.n47 S.n46 0.004
R325 S.n270 S.n269 0.004
R326 S.n89 S.n88 0.004
R327 S.n251 S.n250 0.004
R328 S.n245 S.n244 0.004
R329 S.n132 S.n131 0.004
R330 S.n202 S.n201 0.004
R331 S.n237 S.n236 0.004
R332 S.n78 S.n77 0.004
R333 S.n18 S.n266 0.004
R334 S.n237 S.n222 0.004
R335 S.n23 S.n111 0.004
R336 S.t14 S.n8 0.004
R337 S.n17 S.n7 0.004
R338 S.n16 S.n6 0.004
R339 S.n18 S.n5 0.004
R340 S.n13 S.n4 0.004
R341 S.t22 S.n3 0.004
R342 S.n23 S.n2 0.004
R343 S.t16 S.n335 0.004
R344 S.n213 S.n199 0.004
R345 S.t20 S.n188 0.004
R346 S.t29 S.n81 0.004
R347 S.t20 S.n169 0.004
R348 S.t14 S.n220 0.004
R349 S.t16 S.n319 0.004
R350 S.t16 S.n323 0.004
R351 S.t4 S.n289 0.004
R352 S.n20 S.n215 0.003
R353 S.n15 S.n135 0.003
R354 S.n23 S.n102 0.003
R355 S.t22 S.n138 0.003
R356 S.t22 S.n60 0.003
R357 S.n18 S.n283 0.003
R358 S.t29 S.n99 0.003
R359 S.n17 S.n257 0.003
R360 S.t14 S.n240 0.003
R361 S.n347 S.n346 0.003
R362 S.n174 S.n171 0.003
R363 S.n55 S.n54 0.003
R364 S.t16 S.n321 0.003
R365 S.n42 S.n41 0.003
R366 S.t14 S.n196 0.002
R367 S.n17 S.n247 0.002
R368 S.n28 S.n205 0.002
R369 S.n1 S.n334 0.002
R370 S.n146 S.t22 0.002
R371 S.t20 S.n181 0.002
R372 S.t14 S.n246 0.002
R373 S.n276 S.n275 0.002
R374 S.n9 S.n177 0.002
R375 S.n343 S.n342 0.002
R376 S.n23 S.n66 0.002
R377 S.n28 S.n204 0.002
R378 S.n13 S.n43 0.002
R379 S.n16 S.n84 0.002
R380 S.n18 S.n259 0.002
R381 S.n1 S.n0 0.002
R382 S.n347 S.n336 0.002
R383 S.t20 S.n159 0.002
R384 S.n9 S.n175 0.002
R385 S.n1 S.n330 0.001
R386 S.n336 S.t16 0.001
R387 S.t22 S.n12 0.001
R388 S.n111 S.n110 0.001
R389 S.n266 S.n265 0.001
R390 S.n1 S.n332 0.001
R391 S.n0 S.n333 0.001
R392 S.n93 S.n92 0.001
R393 S.n112 S.n23 0.001
R394 S.n124 S.n123 0.001
R395 S.n76 S.n75 0.001
R396 S.n300 S.n299 0.001
R397 S.n234 S.n232 0.001
R398 S.n342 S.n341 0.001
R399 S.n190 S.t20 0.001
R400 S.n79 S.n78 0.001
R401 S.n238 S.n237 0.001
R402 S.n306 S.n290 0.001
R403 S.n9 S.n176 0.001
R404 S.n126 S.n125 0.001
R405 S.n302 S.n301 0.001
R406 S.n329 S.n1 0.001
R407 S.n212 S.n28 0.001
R408 S.t22 S.n24 0.001
R409 S.t4 S.n18 0.001
R410 S.n23 S.n22 0.001
R411 S.t4 S.n17 0.001
R412 S.t14 S.n21 0.001
R413 S.t22 S.n14 0.001
R414 S.t14 S.n20 0.001
R415 S.t4 S.n19 0.001
R416 S.t29 S.n16 0.001
R417 S.n23 S.t29 0.001
R418 S.t22 S.n13 0.001
R419 S.t22 S.n15 0.001
R420 S.t14 S.n213 0.001
R421 S.n213 S.n212 0.001
R422 S.n290 S.t4 0.001
R423 S.t29 S.n79 0.001
R424 S.t14 S.n238 0.001
R425 S.n307 S.n306 0.001
R426 S.n125 S.n124 0.001
R427 S.n75 S.n74 0.001
R428 S.n301 S.n300 0.001
R429 S.n232 S.n231 0.001
C0 D S 110.34fF
C1 G S 444.79fF
C2 D G 122.23fF
C3 D PW 369.09fF
C4 G PW -50.42fF
C5 S PW 191.15fF
C6 S.n0 PW 0.47fF
C7 S.n1 PW 25.80fF
C8 S.n2 PW 0.13fF
C9 S.n3 PW 0.13fF
C10 S.n4 PW 0.13fF
C11 S.n5 PW 0.13fF
C12 S.n6 PW 0.13fF
C13 S.n7 PW 0.13fF
C14 S.n8 PW 0.13fF
C15 S.n9 PW 22.54fF
C16 S.n10 PW 2.85fF
C17 S.n11 PW 2.95fF
C18 S.t20 PW 36.18fF
C19 S.n12 PW 1.53fF
C20 S.t22 PW 10.28fF
C21 S.n13 PW 1.66fF
C22 S.n14 PW 3.75fF
C23 S.n16 PW 1.90fF
C24 S.t29 PW 8.78fF
C25 S.n17 PW 5.00fF
C26 S.n18 PW 1.72fF
C27 S.n19 PW 0.05fF
C28 S.t4 PW 8.82fF
C29 S.t14 PW 13.07fF
C30 S.n21 PW 0.05fF
C31 S.n22 PW 0.05fF
C32 S.n23 PW 2.07fF
C33 S.n24 PW 0.05fF
C34 S.n25 PW 4.66fF
C35 S.n26 PW 5.05fF
C36 S.n27 PW 11.59fF
C37 S.n28 PW 1.19fF
C38 S.n29 PW 0.09fF
C39 S.n30 PW 0.09fF
C40 S.n31 PW 0.20fF
C41 S.n32 PW 0.06fF
C42 S.n33 PW 0.06fF
C43 S.n34 PW 0.05fF
C44 S.n35 PW 0.06fF
C45 S.n36 PW 0.11fF
C46 S.t45 PW 0.02fF
C47 S.n37 PW 0.18fF
C48 S.n38 PW 0.09fF
C49 S.n39 PW 0.64fF
C50 S.n40 PW 0.26fF
C51 S.n41 PW 1.39fF
C52 S.n42 PW 0.20fF
C53 S.n43 PW 1.74fF
C54 S.n44 PW 0.11fF
C55 S.t23 PW 0.02fF
C56 S.t56 PW 0.02fF
C57 S.n45 PW 0.23fF
C58 S.n46 PW 0.33fF
C59 S.n47 PW 0.57fF
C60 S.n48 PW 0.17fF
C61 S.n49 PW 0.71fF
C62 S.n50 PW 0.14fF
C63 S.n51 PW 0.34fF
C64 S.n52 PW 0.53fF
C65 S.n53 PW 0.20fF
C66 S.n54 PW 0.35fF
C67 S.n55 PW 0.44fF
C68 S.n56 PW 0.07fF
C69 S.t42 PW 0.02fF
C70 S.n57 PW 0.22fF
C71 S.n58 PW 0.86fF
C72 S.t24 PW 0.02fF
C73 S.n59 PW 0.11fF
C74 S.n60 PW 0.13fF
C75 S.n61 PW 1.58fF
C76 S.n62 PW 0.84fF
C77 S.n63 PW 0.15fF
C78 S.n64 PW 1.42fF
C79 S.n65 PW 0.33fF
C80 S.n66 PW 2.57fF
C81 S.n67 PW 0.11fF
C82 S.t40 PW 0.02fF
C83 S.t34 PW 0.02fF
C84 S.n68 PW 1.15fF
C85 S.n69 PW 0.57fF
C86 S.n70 PW 0.84fF
C87 S.n71 PW 0.83fF
C88 S.n72 PW 0.57fF
C89 S.n73 PW 0.90fF
C90 S.t0 PW 4.32fF
C91 S.n74 PW 6.52fF
C92 S.n76 PW 0.35fF
C93 S.n77 PW 2.28fF
C94 S.n78 PW 4.04fF
C95 S.n79 PW 0.24fF
C96 S.n80 PW 0.01fF
C97 S.t51 PW 0.02fF
C98 S.n81 PW 0.24fF
C99 S.t7 PW 0.02fF
C100 S.n82 PW 0.90fF
C101 S.n83 PW 0.66fF
C102 S.n84 PW 1.78fF
C103 S.n85 PW 0.77fF
C104 S.n86 PW 0.31fF
C105 S.t1 PW 0.02fF
C106 S.n87 PW 0.23fF
C107 S.n88 PW 0.33fF
C108 S.n89 PW 0.57fF
C109 S.n90 PW 0.11fF
C110 S.t30 PW 0.02fF
C111 S.n91 PW 0.21fF
C112 S.n92 PW 1.09fF
C113 S.n93 PW 0.21fF
C114 S.n94 PW 0.24fF
C115 S.n95 PW 0.08fF
C116 S.t53 PW 0.02fF
C117 S.n96 PW 0.22fF
C118 S.n97 PW 0.86fF
C119 S.t47 PW 0.02fF
C120 S.n98 PW 0.11fF
C121 S.n99 PW 0.13fF
C122 S.n100 PW 4.20fF
C123 S.t54 PW 0.02fF
C124 S.n101 PW 0.11fF
C125 S.n102 PW 0.13fF
C126 S.t28 PW 0.02fF
C127 S.n103 PW 0.22fF
C128 S.n104 PW 0.86fF
C129 S.t64 PW 0.02fF
C130 S.n105 PW 0.23fF
C131 S.n106 PW 0.33fF
C132 S.n107 PW 0.57fF
C133 S.n108 PW 0.28fF
C134 S.n109 PW 0.53fF
C135 S.n110 PW 0.44fF
C136 S.n111 PW 0.15fF
C137 S.n112 PW 1.84fF
C138 S.n113 PW 12.82fF
C139 S.n114 PW 19.19fF
C140 S.n115 PW 12.82fF
C141 S.n116 PW 19.19fF
C142 S.n117 PW 0.83fF
C143 S.n118 PW 0.25fF
C144 S.t6 PW 4.32fF
C145 S.n119 PW 0.83fF
C146 S.n120 PW 0.09fF
C147 S.n121 PW 1.55fF
C148 S.n122 PW 0.45fF
C149 S.n123 PW 1.09fF
C150 S.n125 PW 4.53fF
C151 S.n126 PW 1.32fF
C152 S.n127 PW 1.41fF
C153 S.n128 PW 1.23fF
C154 S.n129 PW 0.26fF
C155 S.n130 PW 0.23fF
C156 S.t58 PW 0.02fF
C157 S.n131 PW 0.60fF
C158 S.n132 PW 0.57fF
C159 S.t39 PW 0.02fF
C160 S.n133 PW 1.12fF
C161 S.t66 PW 0.02fF
C162 S.n134 PW 0.01fF
C163 S.n135 PW 0.24fF
C164 S.n136 PW 4.20fF
C165 S.t48 PW 0.02fF
C166 S.n137 PW 0.11fF
C167 S.n138 PW 0.13fF
C168 S.t38 PW 0.02fF
C169 S.n139 PW 0.22fF
C170 S.n140 PW 0.86fF
C171 S.t57 PW 0.02fF
C172 S.n141 PW 0.23fF
C173 S.n142 PW 0.33fF
C174 S.n143 PW 0.57fF
C175 S.n144 PW 1.83fF
C176 S.n145 PW 0.74fF
C177 S.n146 PW 1.90fF
C178 S.t52 PW 0.03fF
C179 S.t70 PW 0.02fF
C180 S.n147 PW 11.83fF
C181 S.n148 PW 1.97fF
C182 S.n149 PW 15.18fF
C183 S.n150 PW 0.88fF
C184 S.n151 PW 0.41fF
C185 S.t31 PW 4.85fF
C186 S.n152 PW 19.59fF
C187 S.n153 PW 19.59fF
C188 S.n154 PW 5.04fF
C189 S.n155 PW 0.99fF
C190 S.n156 PW 0.75fF
C191 S.n157 PW 0.43fF
C192 S.n158 PW 0.28fF
C193 S.n159 PW 3.08fF
C194 S.n160 PW 0.29fF
C195 S.n161 PW 0.21fF
C196 S.n162 PW 0.83fF
C197 S.n163 PW 0.64fF
C198 S.n164 PW 0.38fF
C199 S.n165 PW 0.32fF
C200 S.n166 PW 0.61fF
C201 S.t21 PW 0.02fF
C202 S.n167 PW 0.84fF
C203 S.n168 PW 0.02fF
C204 S.t41 PW 0.02fF
C205 S.n169 PW 0.35fF
C206 S.t68 PW 0.02fF
C207 S.n170 PW 0.84fF
C208 S.n171 PW 0.42fF
C209 S.n172 PW 0.17fF
C210 S.n173 PW 0.21fF
C211 S.n174 PW 1.38fF
C212 S.n175 PW 2.07fF
C213 S.n176 PW 4.03fF
C214 S.n177 PW 4.42fF
C215 S.n178 PW 12.82fF
C216 S.n179 PW 12.82fF
C217 S.n180 PW 5.23fF
C218 S.n181 PW 1.39fF
C219 S.n182 PW 0.83fF
C220 S.n183 PW 0.51fF
C221 S.n184 PW 0.41fF
C222 S.n185 PW 1.10fF
C223 S.t67 PW 0.02fF
C224 S.n186 PW 0.84fF
C225 S.n187 PW 0.02fF
C226 S.t32 PW 0.02fF
C227 S.n188 PW 0.35fF
C228 S.t50 PW 0.02fF
C229 S.n189 PW 0.84fF
C230 S.n190 PW 7.26fF
C231 S.n191 PW 17.94fF
C232 S.t11 PW 0.02fF
C233 S.n192 PW 1.15fF
C234 S.t69 PW 0.02fF
C235 S.n193 PW 0.22fF
C236 S.n194 PW 0.86fF
C237 S.n195 PW 1.72fF
C238 S.n196 PW 1.83fF
C239 S.n197 PW 0.11fF
C240 S.t65 PW 0.02fF
C241 S.t15 PW 0.02fF
C242 S.n198 PW 0.11fF
C243 S.n199 PW 0.13fF
C244 S.n200 PW 0.22fF
C245 S.t37 PW 0.02fF
C246 S.n201 PW 0.34fF
C247 S.n202 PW 0.34fF
C248 S.n203 PW 0.63fF
C249 S.n204 PW 1.48fF
C250 S.n205 PW 1.59fF
C251 S.n206 PW 0.29fF
C252 S.n207 PW 0.98fF
C253 S.n208 PW 0.46fF
C254 S.n209 PW 0.23fF
C255 S.t19 PW 0.02fF
C256 S.n210 PW 0.33fF
C257 S.n211 PW 0.59fF
C258 S.n212 PW 0.38fF
C259 S.n214 PW 0.11fF
C260 S.t59 PW 0.02fF
C261 S.n215 PW 0.13fF
C262 S.n216 PW 4.20fF
C263 S.t35 PW 0.02fF
C264 S.n217 PW 0.90fF
C265 S.n218 PW 0.66fF
C266 S.n219 PW 0.01fF
C267 S.t27 PW 0.02fF
C268 S.n220 PW 0.24fF
C269 S.t49 PW 0.02fF
C270 S.n221 PW 1.15fF
C271 S.n222 PW 0.34fF
C272 S.n223 PW 1.15fF
C273 S.n224 PW 0.09fF
C274 S.n225 PW 0.06fF
C275 S.n226 PW 0.57fF
C276 S.n227 PW 0.57fF
C277 S.n228 PW 0.90fF
C278 S.n229 PW 0.79fF
C279 S.n230 PW 0.02fF
C280 S.n231 PW 6.52fF
C281 S.t12 PW 4.32fF
C282 S.n233 PW 0.83fF
C283 S.n234 PW 0.35fF
C284 S.n235 PW 1.28fF
C285 S.n236 PW 2.28fF
C286 S.n237 PW 3.36fF
C287 S.n238 PW 0.24fF
C288 S.t26 PW 0.02fF
C289 S.n239 PW 0.11fF
C290 S.n240 PW 0.13fF
C291 S.t3 PW 0.02fF
C292 S.n241 PW 0.22fF
C293 S.n242 PW 0.86fF
C294 S.t25 PW 0.02fF
C295 S.n243 PW 0.23fF
C296 S.n244 PW 0.33fF
C297 S.n245 PW 0.57fF
C298 S.n246 PW 1.23fF
C299 S.n247 PW 1.77fF
C300 S.n248 PW 0.11fF
C301 S.t5 PW 0.02fF
C302 S.t43 PW 0.02fF
C303 S.n249 PW 0.23fF
C304 S.n250 PW 0.33fF
C305 S.n251 PW 0.57fF
C306 S.n252 PW 1.17fF
C307 S.n253 PW 0.66fF
C308 S.n254 PW 0.35fF
C309 S.n255 PW 0.33fF
C310 S.t44 PW 0.02fF
C311 S.n256 PW 0.11fF
C312 S.n257 PW 0.13fF
C313 S.n258 PW 4.20fF
C314 S.n259 PW 1.65fF
C315 S.n260 PW 0.16fF
C316 S.n261 PW 0.72fF
C317 S.n262 PW 0.30fF
C318 S.n263 PW 0.24fF
C319 S.n264 PW 0.28fF
C320 S.n265 PW 0.44fF
C321 S.n266 PW 0.15fF
C322 S.n267 PW 1.85fF
C323 S.t9 PW 0.02fF
C324 S.n268 PW 0.23fF
C325 S.n269 PW 0.33fF
C326 S.n270 PW 0.57fF
C327 S.n271 PW 0.11fF
C328 S.t62 PW 0.02fF
C329 S.n272 PW 0.17fF
C330 S.n273 PW 0.19fF
C331 S.n274 PW 0.62fF
C332 S.n275 PW 0.85fF
C333 S.n276 PW 0.21fF
C334 S.n277 PW 0.06fF
C335 S.n278 PW 0.05fF
C336 S.n279 PW 0.09fF
C337 S.n280 PW 0.20fF
C338 S.n281 PW 0.06fF
C339 S.t63 PW 0.02fF
C340 S.n282 PW 0.11fF
C341 S.n283 PW 0.13fF
C342 S.t8 PW 0.02fF
C343 S.n284 PW 0.22fF
C344 S.n285 PW 0.86fF
C345 S.t10 PW 0.02fF
C346 S.n286 PW 0.90fF
C347 S.n287 PW 0.66fF
C348 S.t55 PW 0.02fF
C349 S.n288 PW 0.01fF
C350 S.n289 PW 0.24fF
C351 S.n290 PW 0.24fF
C352 S.n291 PW 1.20fF
C353 S.n292 PW 0.18fF
C354 S.n293 PW 1.42fF
C355 S.n294 PW 0.32fF
C356 S.t2 PW 4.32fF
C357 S.n295 PW 0.56fF
C358 S.n296 PW 0.09fF
C359 S.n297 PW 1.55fF
C360 S.n298 PW 0.45fF
C361 S.n299 PW 1.09fF
C362 S.n301 PW 4.53fF
C363 S.n302 PW 1.32fF
C364 S.n303 PW 0.56fF
C365 S.n304 PW 0.19fF
C366 S.n305 PW 2.13fF
C367 S.n306 PW 1.02fF
C368 S.n307 PW 2.49fF
C369 S.t36 PW 0.02fF
C370 S.n308 PW 1.20fF
C371 S.n309 PW 1.21fF
C372 S.n310 PW 0.19fF
C373 S.n311 PW 2.06fF
C374 S.n312 PW 0.29fF
C375 S.n313 PW 0.29fF
C376 S.n314 PW 1.12fF
C377 S.n315 PW 0.31fF
C378 S.n316 PW 4.20fF
C379 S.t18 PW 0.02fF
C380 S.n317 PW 0.84fF
C381 S.t33 PW 0.02fF
C382 S.n318 PW 0.02fF
C383 S.n319 PW 0.35fF
C384 S.t17 PW 0.02fF
C385 S.n320 PW 0.84fF
C386 S.t46 PW 0.02fF
C387 S.n321 PW 0.42fF
C388 S.t13 PW 0.02fF
C389 S.n322 PW 0.02fF
C390 S.n323 PW 0.35fF
C391 S.t61 PW 0.02fF
C392 S.n324 PW 0.84fF
C393 S.t60 PW 0.02fF
C394 S.n325 PW 0.84fF
C395 S.n326 PW 0.96fF
C396 S.n327 PW 0.58fF
C397 S.n328 PW 0.83fF
C398 S.n329 PW 2.44fF
C399 S.n330 PW 1.45fF
C400 S.n331 PW 0.86fF
C401 S.n332 PW 0.37fF
C402 S.n333 PW 0.37fF
C403 S.n334 PW 1.47fF
C404 S.n335 PW 3.96fF
C405 S.t16 PW 30.14fF
C406 S.n336 PW 0.44fF
C407 S.n337 PW 2.00fF
C408 S.n338 PW 0.79fF
C409 S.n339 PW 0.12fF
C410 S.n340 PW 6.01fF
C411 S.n341 PW 2.31fF
C412 S.n342 PW 3.78fF
C413 S.n343 PW 5.74fF
C414 S.n344 PW 0.71fF
C415 S.n345 PW 4.44fF
C416 S.n346 PW 2.37fF
C417 S.n347 PW 6.81fF
C418 S.n348 PW 15.27fF
C419 S.n349 PW 16.74fF
C420 D.t1 PW 18.22fF
C421 D.t6 PW 70.07fF
C422 D.n0 PW 10.57fF
C423 D.t3 PW -0.05fF
C424 D.t7 PW 0.00fF
C425 D.t4 PW -0.00fF
C426 D.t5 PW -0.02fF
C427 D.t2 PW -0.02fF
C428 D.t0 PW -0.02fF
.ends

